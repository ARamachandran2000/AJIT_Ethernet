-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity AccessRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(3 downto 0);
    register_index : in  std_logic_vector(5 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity AccessRegister;
architecture AccessRegister_arch of AccessRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 43)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal register_index_buffer :  std_logic_vector(5 downto 0);
  signal register_index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal AccessRegister_CP_0_start: Boolean;
  signal AccessRegister_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "AccessRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 43) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(4 downto 1) <= bmask;
  bmask_buffer <= in_buffer_data_out(4 downto 1);
  in_buffer_data_in(10 downto 5) <= register_index;
  register_index_buffer <= in_buffer_data_out(10 downto 5);
  in_buffer_data_in(42 downto 11) <= wdata;
  wdata_buffer <= in_buffer_data_out(42 downto 11);
  in_buffer_data_in(tag_length + 42 downto 43) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 42 downto 43);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  AccessRegister_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "AccessRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  AccessRegister_CP_0: Block -- control-path 
    signal AccessRegister_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    AccessRegister_CP_0_elements(0) <= AccessRegister_CP_0_start;
    AccessRegister_CP_0_symbol <= AccessRegister_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_sample_start_
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/req
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_sample_start_
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/rr
      -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0); -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_sample_completed_
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_update_start_
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/ack
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/$entry
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0, ack => AccessRegister_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(1), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_update_completed_
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/$exit
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1, ack => AccessRegister_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_sample_completed_
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_update_start_
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/ra
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/$entry
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0, ack => AccessRegister_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(3), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_update_completed_
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/$exit
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1, ack => AccessRegister_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_77_to_assign_stmt_95/$exit
      -- 
    AccessRegister_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "AccessRegister_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= AccessRegister_CP_0_elements(4) & AccessRegister_CP_0_elements(2);
      gj_AccessRegister_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => AccessRegister_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u5_72_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u6_u38_75_wire : std_logic_vector(37 downto 0);
    signal request_77 : std_logic_vector(42 downto 0);
    signal response_89 : std_logic_vector(32 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_94_inst
    rdata_buffer <= response_89(31 downto 0);
    -- binary operator CONCAT_u1_u5_72_inst
    process(rwbar_buffer, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(rwbar_buffer, bmask_buffer, tmp_var);
      CONCAT_u1_u5_72_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u5_u43_76_inst
    process(CONCAT_u1_u5_72_wire, CONCAT_u6_u38_75_wire) -- 
      variable tmp_var : std_logic_vector(42 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_72_wire, CONCAT_u6_u38_75_wire, tmp_var);
      request_77 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u38_75_inst
    process(register_index_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(37 downto 0); -- 
    begin -- 
      ApConcat_proc(register_index_buffer, wdata_buffer, tmp_var);
      CONCAT_u6_u38_75_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_89 <= data_out(32 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_77;
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE", data_width => 43, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end AccessRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity NicRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity NicRegisterAccessDaemon;
architecture NicRegisterAccessDaemon_arch of NicRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal NicRegisterAccessDaemon_CP_116_start: Boolean;
  signal NicRegisterAccessDaemon_CP_116_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_179_branch_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1 : boolean;
  signal array_obj_ref_203_load_0_req_0 : boolean;
  signal array_obj_ref_203_load_0_ack_0 : boolean;
  signal array_obj_ref_203_load_0_req_1 : boolean;
  signal array_obj_ref_203_load_0_ack_1 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_req_0 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_ack_0 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_req_1 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_ack_1 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_req_0 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_ack_0 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_req_1 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_ack_1 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_req_0 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_ack_0 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_req_1 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_ack_1 : boolean;
  signal W_index_216_delayed_5_0_217_inst_req_0 : boolean;
  signal W_index_216_delayed_5_0_217_inst_ack_0 : boolean;
  signal W_index_216_delayed_5_0_217_inst_req_1 : boolean;
  signal W_index_216_delayed_5_0_217_inst_ack_1 : boolean;
  signal call_stmt_226_call_req_0 : boolean;
  signal call_stmt_226_call_ack_0 : boolean;
  signal call_stmt_226_call_req_1 : boolean;
  signal call_stmt_226_call_ack_1 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_req_0 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_ack_0 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_req_1 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_ack_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1 : boolean;
  signal do_while_stmt_179_branch_ack_0 : boolean;
  signal do_while_stmt_179_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  NicRegisterAccessDaemon_CP_116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  NicRegisterAccessDaemon_CP_116: Block -- control-path 
    signal NicRegisterAccessDaemon_CP_116_elements: BooleanArray(50 downto 0);
    -- 
  begin -- 
    NicRegisterAccessDaemon_CP_116_elements(0) <= NicRegisterAccessDaemon_CP_116_start;
    NicRegisterAccessDaemon_CP_116_symbol <= NicRegisterAccessDaemon_CP_116_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_178/$entry
      -- CP-element group 0: 	 branch_block_stmt_178/branch_block_stmt_178__entry__
      -- CP-element group 0: 	 branch_block_stmt_178/do_while_stmt_179__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	50 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_178/$exit
      -- CP-element group 1: 	 branch_block_stmt_178/branch_block_stmt_178__exit__
      -- CP-element group 1: 	 branch_block_stmt_178/do_while_stmt_179__exit__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(1) <= NicRegisterAccessDaemon_CP_116_elements(50);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_178/do_while_stmt_179/$entry
      -- CP-element group 2: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179__entry__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(2) <= NicRegisterAccessDaemon_CP_116_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	50 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179__exit__
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_178/do_while_stmt_179/loop_back
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	45 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	48 
    -- CP-element group 5: 	49 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/condition_done
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/$entry
      -- 
    NicRegisterAccessDaemon_CP_116_elements(5) <= NicRegisterAccessDaemon_CP_116_elements(45);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	47 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_178/do_while_stmt_179/loop_body_done
      -- 
    NicRegisterAccessDaemon_CP_116_elements(6) <= NicRegisterAccessDaemon_CP_116_elements(47);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/back_edge_to_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(7) <= NicRegisterAccessDaemon_CP_116_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/first_time_through_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(8) <= NicRegisterAccessDaemon_CP_116_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	45 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/loop_body_start
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/rr
      -- 
    rr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(10), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(9) & NicRegisterAccessDaemon_CP_116_elements(13);
      gj_NicRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	20 
    -- CP-element group 11: 	24 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	40 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_update_start_
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/cr
      -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(11), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(12) & NicRegisterAccessDaemon_CP_116_elements(20) & NicRegisterAccessDaemon_CP_116_elements(24) & NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(32) & NicRegisterAccessDaemon_CP_116_elements(40) & NicRegisterAccessDaemon_CP_116_elements(16);
      gj_NicRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/ra
      -- 
    ra_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	22 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	30 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (29) 
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/index_resize_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/index_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/scale_rename_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/scale_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resized_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scaled_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_computed_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/root_register_ack
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/rr
      -- 
    rr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(14), ack => array_obj_ref_203_load_0_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(37) & NicRegisterAccessDaemon_CP_116_elements(16);
      gj_NicRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	36 
    -- CP-element group 15: 	43 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_update_start_
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/cr
      -- 
    cr_212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => array_obj_ref_203_load_0_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(36) & NicRegisterAccessDaemon_CP_116_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	46 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/ra
      -- 
    ra_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_load_0_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17: 	42 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/merge_ack
      -- 
    ca_213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_load_0_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/req
      -- 
    req_226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(18), ack => W_rwbar_212_delayed_5_0_208_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(20);
      gj_NicRegisterAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	36 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_update_start_
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/req
      -- 
    req_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(19), ack => W_rwbar_212_delayed_5_0_208_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	11 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/ack
      -- 
    ack_227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_212_delayed_5_0_208_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/ack
      -- 
    ack_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_212_delayed_5_0_208_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/req
      -- 
    req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(22), ack => W_bmask_213_delayed_5_0_211_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(24);
      gj_NicRegisterAccessDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	36 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_update_start_
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/req
      -- 
    req_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(23), ack => W_bmask_213_delayed_5_0_211_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	11 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/ack
      -- 
    ack_241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_213_delayed_5_0_211_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/ack
      -- 
    ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_213_delayed_5_0_211_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/req
      -- 
    req_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(26), ack => W_wdata_215_delayed_5_0_214_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(28);
      gj_NicRegisterAccessDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	36 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_update_start_
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/req
      -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(27), ack => W_wdata_215_delayed_5_0_214_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: 	11 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/ack
      -- 
    ack_255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_215_delayed_5_0_214_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_215_delayed_5_0_214_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	13 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/req
      -- 
    req_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(30), ack => W_index_216_delayed_5_0_217_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(32);
      gj_NicRegisterAccessDaemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	36 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_update_start_
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/req
      -- 
    req_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(31), ack => W_index_216_delayed_5_0_217_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/ack
      -- 
    ack_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_216_delayed_5_0_217_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/ack
      -- 
    ack_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_216_delayed_5_0_217_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	46 
    -- CP-element group 34: 	17 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/crr
      -- 
    crr_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(34), ack => call_stmt_226_call_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 31,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(21) & NicRegisterAccessDaemon_CP_116_elements(25) & NicRegisterAccessDaemon_CP_116_elements(29) & NicRegisterAccessDaemon_CP_116_elements(33) & NicRegisterAccessDaemon_CP_116_elements(46) & NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_update_start_
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/ccr
      -- 
    ccr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(35), ack => call_stmt_226_call_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(37);
      gj_NicRegisterAccessDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	19 
    -- CP-element group 36: 	23 
    -- CP-element group 36: 	27 
    -- CP-element group 36: 	31 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	15 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/cra
      -- 
    cra_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_226_call_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	47 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/cca
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/ring_reenable_memory_space_0
      -- 
    cca_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_226_call_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/req
      -- 
    req_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(38), ack => W_rwbar_220_delayed_5_0_227_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(40);
      gj_NicRegisterAccessDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	43 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_update_start_
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/req
      -- 
    req_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(39), ack => W_rwbar_220_delayed_5_0_227_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: 	11 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/ack
      -- 
    ack_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_220_delayed_5_0_227_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/ack
      -- 
    ack_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_220_delayed_5_0_227_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	17 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/req
      -- 
    req_310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(42), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(41) & NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(44);
      gj_NicRegisterAccessDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	39 
    -- CP-element group 43: 	15 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_update_start_
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/req
      -- 
    ack_311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(43)); -- 
    req_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(43), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/ack
      -- 
    ack_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(44)); -- 
    -- CP-element group 45:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	9 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	5 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/condition_evaluated
      -- CP-element group 45: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(45), ack => do_while_stmt_179_branch_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(9), ack => NicRegisterAccessDaemon_CP_116_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	16 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	34 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_call_stmt_226_delay
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(16), ack => NicRegisterAccessDaemon_CP_116_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	37 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	6 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/$exit
      -- 
    NicRegisterAccessDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(37) & NicRegisterAccessDaemon_CP_116_elements(44);
      gj_NicRegisterAccessDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	5 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/$exit
      -- CP-element group 48: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/ack
      -- 
    ack_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_179_branch_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	5 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/$exit
      -- CP-element group 49: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/ack
      -- 
    ack_327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_179_branch_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(49)); -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	3 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	1 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_178/do_while_stmt_179/$exit
      -- 
    NicRegisterAccessDaemon_CP_116_elements(50) <= NicRegisterAccessDaemon_CP_116_elements(3);
    NicRegisterAccessDaemon_do_while_stmt_179_terminator_328: loop_terminator -- 
      generic map (name => " NicRegisterAccessDaemon_do_while_stmt_179_terminator_328", max_iterations_in_flight =>31) 
      port map(loop_body_exit => NicRegisterAccessDaemon_CP_116_elements(6),loop_continue => NicRegisterAccessDaemon_CP_116_elements(49),loop_terminate => NicRegisterAccessDaemon_CP_116_elements(48),loop_back => NicRegisterAccessDaemon_CP_116_elements(4),loop_exit => NicRegisterAccessDaemon_CP_116_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_141_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= NicRegisterAccessDaemon_CP_116_elements(7);
        preds(1)  <= NicRegisterAccessDaemon_CP_116_elements(8);
        entry_tmerge_141 : transition_merge -- 
          generic map(name => " entry_tmerge_141")
          port map (preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_index_202_resized : std_logic_vector(5 downto 0);
    signal R_index_202_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_203_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_192 : std_logic_vector(3 downto 0);
    signal bmask_213_delayed_5_0_213 : std_logic_vector(3 downto 0);
    signal index_196 : std_logic_vector(5 downto 0);
    signal index_216_delayed_5_0_219 : std_logic_vector(5 downto 0);
    signal konst_247_wire_constant : std_logic_vector(0 downto 0);
    signal rdata_236 : std_logic_vector(31 downto 0);
    signal req_183 : std_logic_vector(42 downto 0);
    signal resp_242 : std_logic_vector(32 downto 0);
    signal rval_204 : std_logic_vector(31 downto 0);
    signal rwbar_188 : std_logic_vector(0 downto 0);
    signal rwbar_212_delayed_5_0_210 : std_logic_vector(0 downto 0);
    signal rwbar_220_delayed_5_0_229 : std_logic_vector(0 downto 0);
    signal type_cast_234_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_200 : std_logic_vector(31 downto 0);
    signal wdata_215_delayed_5_0_216 : std_logic_vector(31 downto 0);
    signal wval_226 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_203_offset_scale_factor_0 <= "000001";
    array_obj_ref_203_resized_base_address <= "000000";
    array_obj_ref_203_word_offset_0 <= "000000";
    konst_247_wire_constant <= "1";
    type_cast_234_wire_constant <= "00000000000000000000000000000000";
    type_cast_239_wire_constant <= "0";
    -- flow-through select operator MUX_235_inst
    rdata_236 <= rval_204 when (rwbar_220_delayed_5_0_229(0) /=  '0') else type_cast_234_wire_constant;
    -- flow-through slice operator slice_187_inst
    rwbar_188 <= req_183(42 downto 42);
    -- flow-through slice operator slice_191_inst
    bmask_192 <= req_183(41 downto 38);
    -- flow-through slice operator slice_195_inst
    index_196 <= req_183(37 downto 32);
    -- flow-through slice operator slice_199_inst
    wdata_200 <= req_183(31 downto 0);
    W_bmask_213_delayed_5_0_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_213_delayed_5_0_211_inst_req_0;
      W_bmask_213_delayed_5_0_211_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_213_delayed_5_0_211_inst_req_1;
      W_bmask_213_delayed_5_0_211_inst_ack_1<= rack(0);
      W_bmask_213_delayed_5_0_211_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_213_delayed_5_0_211_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_213_delayed_5_0_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_216_delayed_5_0_217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_216_delayed_5_0_217_inst_req_0;
      W_index_216_delayed_5_0_217_inst_ack_0<= wack(0);
      rreq(0) <= W_index_216_delayed_5_0_217_inst_req_1;
      W_index_216_delayed_5_0_217_inst_ack_1<= rack(0);
      W_index_216_delayed_5_0_217_inst : InterlockBuffer generic map ( -- 
        name => "W_index_216_delayed_5_0_217_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_216_delayed_5_0_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_212_delayed_5_0_208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_212_delayed_5_0_208_inst_req_0;
      W_rwbar_212_delayed_5_0_208_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_212_delayed_5_0_208_inst_req_1;
      W_rwbar_212_delayed_5_0_208_inst_ack_1<= rack(0);
      W_rwbar_212_delayed_5_0_208_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_212_delayed_5_0_208_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_212_delayed_5_0_210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_220_delayed_5_0_227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_220_delayed_5_0_227_inst_req_0;
      W_rwbar_220_delayed_5_0_227_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_220_delayed_5_0_227_inst_req_1;
      W_rwbar_220_delayed_5_0_227_inst_ack_1<= rack(0);
      W_rwbar_220_delayed_5_0_227_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_220_delayed_5_0_227_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_220_delayed_5_0_229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_215_delayed_5_0_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_215_delayed_5_0_214_inst_req_0;
      W_wdata_215_delayed_5_0_214_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_215_delayed_5_0_214_inst_req_1;
      W_wdata_215_delayed_5_0_214_inst_ack_1<= rack(0);
      W_wdata_215_delayed_5_0_214_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_215_delayed_5_0_214_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_215_delayed_5_0_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_203_addr_0
    process(array_obj_ref_203_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_203_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_gather_scatter
    process(array_obj_ref_203_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_data_0;
      ov(31 downto 0) := iv;
      rval_204 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_0_rename
    process(R_index_202_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_202_resized;
      ov(5 downto 0) := iv;
      R_index_202_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_0_resize
    process(index_196) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_196;
      ov(5 downto 0) := iv;
      R_index_202_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_offset
    process(R_index_202_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_202_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_203_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_root_address_inst
    process(array_obj_ref_203_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_203_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_179_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_247_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_179_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_179_branch_req_0,
          ack0 => do_while_stmt_179_branch_ack_0,
          ack1 => do_while_stmt_179_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_241_inst
    process(type_cast_239_wire_constant, rdata_236) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_239_wire_constant, rdata_236, tmp_var);
      resp_242 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_203_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_203_load_0_req_0;
      array_obj_ref_203_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_203_load_0_req_1;
      array_obj_ref_203_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_203_word_address_0;
      array_obj_ref_203_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(42 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_183 <= data_out(42 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0", data_width => 43,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_242;
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_226_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_226_call_req_0;
      call_stmt_226_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_226_call_req_1;
      call_stmt_226_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_212_delayed_5_0_210(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_213_delayed_5_0_213 & rval_204 & wdata_215_delayed_5_0_216 & index_216_delayed_5_0_219;
      wval_226 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end NicRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ReceiveEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_call_data : out  std_logic_vector(35 downto 0);
    loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
    loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_return_data : in   std_logic_vector(0 downto 0);
    loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
    populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ReceiveEngineDaemon;
architecture ReceiveEngineDaemon_arch of ReceiveEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ReceiveEngineDaemon_CP_1868_start: Boolean;
  signal ReceiveEngineDaemon_CP_1868_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1523_call_ack_0 : boolean;
  signal W_pkt_cnt_1487_delayed_13_0_1491_inst_req_1 : boolean;
  signal W_pkt_cnt_1487_delayed_13_0_1491_inst_ack_0 : boolean;
  signal NOT_u1_u1_1466_inst_req_0 : boolean;
  signal W_pkt_cnt_1487_delayed_13_0_1491_inst_req_0 : boolean;
  signal call_stmt_1490_call_ack_0 : boolean;
  signal NOT_u1_u1_1456_inst_ack_1 : boolean;
  signal call_stmt_1510_call_ack_0 : boolean;
  signal NOT_u1_u1_1456_inst_ack_0 : boolean;
  signal call_stmt_1510_call_req_0 : boolean;
  signal call_stmt_1510_call_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_ack_1 : boolean;
  signal call_stmt_1510_call_ack_1 : boolean;
  signal call_stmt_1490_call_req_1 : boolean;
  signal call_stmt_1523_call_req_0 : boolean;
  signal NOT_u1_u1_1456_inst_req_1 : boolean;
  signal NOT_u1_u1_1466_inst_ack_1 : boolean;
  signal NOT_u1_u1_1466_inst_req_1 : boolean;
  signal call_stmt_1490_call_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_req_1 : boolean;
  signal NOT_u1_u1_1456_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_ack_1 : boolean;
  signal do_while_stmt_1411_branch_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_ack_1 : boolean;
  signal do_while_stmt_1411_branch_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_req_1 : boolean;
  signal if_stmt_1403_branch_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_ack_0 : boolean;
  signal if_stmt_1403_branch_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_req_0 : boolean;
  signal NOT_u1_u1_1466_inst_ack_0 : boolean;
  signal if_stmt_1403_branch_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_ack_0 : boolean;
  signal do_while_stmt_1411_branch_req_0 : boolean;
  signal phi_stmt_1413_req_0 : boolean;
  signal phi_stmt_1413_req_1 : boolean;
  signal phi_stmt_1413_ack_0 : boolean;
  signal npkt_cnt_1500_1415_buf_req_0 : boolean;
  signal npkt_cnt_1500_1415_buf_ack_0 : boolean;
  signal W_pkt_cnt_1482_delayed_13_0_1478_inst_ack_1 : boolean;
  signal W_pkt_cnt_1482_delayed_13_0_1478_inst_req_1 : boolean;
  signal npkt_cnt_1500_1415_buf_req_1 : boolean;
  signal npkt_cnt_1500_1415_buf_ack_1 : boolean;
  signal call_stmt_1490_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_req_0 : boolean;
  signal call_stmt_1425_call_req_0 : boolean;
  signal call_stmt_1523_call_ack_1 : boolean;
  signal call_stmt_1425_call_ack_0 : boolean;
  signal call_stmt_1425_call_req_1 : boolean;
  signal call_stmt_1523_call_req_1 : boolean;
  signal call_stmt_1425_call_ack_1 : boolean;
  signal call_stmt_1437_call_req_0 : boolean;
  signal call_stmt_1437_call_ack_0 : boolean;
  signal call_stmt_1437_call_req_1 : boolean;
  signal call_stmt_1437_call_ack_1 : boolean;
  signal W_pkt_cnt_1482_delayed_13_0_1478_inst_ack_0 : boolean;
  signal W_pkt_cnt_1482_delayed_13_0_1478_inst_req_0 : boolean;
  signal W_pkt_cnt_1487_delayed_13_0_1491_inst_ack_1 : boolean;
  signal call_stmt_1453_call_req_0 : boolean;
  signal call_stmt_1453_call_ack_0 : boolean;
  signal call_stmt_1453_call_req_1 : boolean;
  signal call_stmt_1453_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ReceiveEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ReceiveEngineDaemon_CP_1868_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ReceiveEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1868_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1868_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1868_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ReceiveEngineDaemon_CP_1868: Block -- control-path 
    signal ReceiveEngineDaemon_CP_1868_elements: BooleanArray(87 downto 0);
    -- 
  begin -- 
    ReceiveEngineDaemon_CP_1868_elements(0) <= ReceiveEngineDaemon_CP_1868_start;
    ReceiveEngineDaemon_CP_1868_symbol <= ReceiveEngineDaemon_CP_1868_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1399/$entry
      -- CP-element group 0: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_sample_start_
      -- CP-element group 0: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Sample/req
      -- 
    req_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(0), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_update_start_
      -- CP-element group 1: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Update/req
      -- 
    ack_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(1)); -- 
    req_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(1), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	87 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 branch_block_stmt_1400/merge_stmt_1402__entry___PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_1400/merge_stmt_1402__entry___PhiReq/$entry
      -- CP-element group 2: 	 assign_stmt_1399/$exit
      -- CP-element group 2: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1400/merge_stmt_1402_dead_link/$entry
      -- CP-element group 2: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1399/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_1400/$entry
      -- CP-element group 2: 	 branch_block_stmt_1400/branch_block_stmt_1400__entry__
      -- CP-element group 2: 	 branch_block_stmt_1400/merge_stmt_1402__entry__
      -- 
    ack_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_1400/$exit
      -- CP-element group 3: 	 branch_block_stmt_1400/branch_block_stmt_1400__exit__
      -- 
    ReceiveEngineDaemon_CP_1868_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	86 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	87 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1400/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1400/disable_loopback_PhiReq/$exit
      -- CP-element group 4: 	 branch_block_stmt_1400/do_while_stmt_1411__exit__
      -- CP-element group 4: 	 branch_block_stmt_1400/disable_loopback
      -- 
    ReceiveEngineDaemon_CP_1868_elements(4) <= ReceiveEngineDaemon_CP_1868_elements(86);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	87 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	87 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1400/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1400/not_enabled_yet_loopback_PhiReq/$exit
      -- CP-element group 5: 	 branch_block_stmt_1400/if_stmt_1403_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1400/if_stmt_1403_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1400/not_enabled_yet_loopback
      -- 
    if_choice_transition_1960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1403_branch_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	87 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_1400/if_stmt_1403__exit__
      -- CP-element group 6: 	 branch_block_stmt_1400/do_while_stmt_1411__entry__
      -- CP-element group 6: 	 branch_block_stmt_1400/if_stmt_1403_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1400/if_stmt_1403_else_link/else_choice_transition
      -- 
    else_choice_transition_1964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1403_branch_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1400/do_while_stmt_1411/$entry
      -- CP-element group 7: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411__entry__
      -- 
    ReceiveEngineDaemon_CP_1868_elements(7) <= ReceiveEngineDaemon_CP_1868_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	86 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411__exit__
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_back
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	84 
    -- CP-element group 10: 	85 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_taken/$entry
      -- CP-element group 10: 	 branch_block_stmt_1400/do_while_stmt_1411/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_exit/$entry
      -- 
    ReceiveEngineDaemon_CP_1868_elements(10) <= ReceiveEngineDaemon_CP_1868_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	83 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_body_done
      -- 
    ReceiveEngineDaemon_CP_1868_elements(11) <= ReceiveEngineDaemon_CP_1868_elements(83);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	21 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/back_edge_to_loop_body
      -- 
    ReceiveEngineDaemon_CP_1868_elements(12) <= ReceiveEngineDaemon_CP_1868_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	23 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/first_time_through_loop_body
      -- 
    ReceiveEngineDaemon_CP_1868_elements(13) <= ReceiveEngineDaemon_CP_1868_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	82 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	34 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/loop_body_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	82 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/condition_evaluated
      -- 
    condition_evaluated_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(15), ack => do_while_stmt_1411_branch_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(82) & ReceiveEngineDaemon_CP_1868_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	17 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_sample_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(17) & ReceiveEngineDaemon_CP_1868_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	65 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	16 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_sample_start_
      -- 
    ReceiveEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(14) & ReceiveEngineDaemon_CP_1868_elements(65) & ReceiveEngineDaemon_CP_1868_elements(19);
      gj_ReceiveEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	64 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_update_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(14) & ReceiveEngineDaemon_CP_1868_elements(56) & ReceiveEngineDaemon_CP_1868_elements(64);
      gj_ReceiveEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	63 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/aggregated_phi_sample_ack
      -- CP-element group 19: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_sample_completed__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	62 
    -- CP-element group 20: 	54 
    -- CP-element group 20: 	15 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/aggregated_phi_update_ack
      -- CP-element group 20: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_update_completed__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	12 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_loopback_trigger
      -- 
    ReceiveEngineDaemon_CP_1868_elements(21) <= ReceiveEngineDaemon_CP_1868_elements(12);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_loopback_sample_req_ps
      -- 
    phi_stmt_1413_loopback_sample_req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1413_loopback_sample_req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(22), ack => phi_stmt_1413_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	13 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_entry_trigger
      -- 
    ReceiveEngineDaemon_CP_1868_elements(23) <= ReceiveEngineDaemon_CP_1868_elements(13);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_entry_sample_req_ps
      -- 
    phi_stmt_1413_entry_sample_req_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1413_entry_sample_req_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(24), ack => phi_stmt_1413_req_1); -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/phi_stmt_1413_phi_mux_ack_ps
      -- 
    phi_stmt_1413_phi_mux_ack_2001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1413_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Sample/req
      -- 
    req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(26), ack => npkt_cnt_1500_1415_buf_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Update/req
      -- 
    req_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(27), ack => npkt_cnt_1500_1415_buf_req_1); -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Sample/ack
      -- 
    ack_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1500_1415_buf_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/R_npkt_cnt_1415_Update/ack
      -- 
    ack_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1500_1415_buf_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_sample_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_update_start_
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_update_completed__ps
      -- 
    ReceiveEngineDaemon_CP_1868_elements(32) <= ReceiveEngineDaemon_CP_1868_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/type_cast_1417_update_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_1868_elements(31), ack => ReceiveEngineDaemon_CP_1868_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	14 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	81 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Sample/crr
      -- 
    crr_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(34), ack => call_stmt_1425_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(14) & ReceiveEngineDaemon_CP_1868_elements(81) & ReceiveEngineDaemon_CP_1868_elements(36);
      gj_ReceiveEngineDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	52 
    -- CP-element group 35: 	48 
    -- CP-element group 35: 	44 
    -- CP-element group 35: 	81 
    -- CP-element group 35: 	76 
    -- CP-element group 35: 	68 
    -- CP-element group 35: 	40 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Update/ccr
      -- 
    ccr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(35), ack => call_stmt_1425_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(52) & ReceiveEngineDaemon_CP_1868_elements(48) & ReceiveEngineDaemon_CP_1868_elements(44) & ReceiveEngineDaemon_CP_1868_elements(81) & ReceiveEngineDaemon_CP_1868_elements(76) & ReceiveEngineDaemon_CP_1868_elements(68) & ReceiveEngineDaemon_CP_1868_elements(40);
      gj_ReceiveEngineDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Sample/cra
      -- 
    cra_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1425_call_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	50 
    -- CP-element group 37: 	46 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	74 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	42 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1425_Update/cca
      -- 
    cca_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1425_call_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	73 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Sample/crr
      -- 
    crr_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(38), ack => call_stmt_1437_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(37) & ReceiveEngineDaemon_CP_1868_elements(73) & ReceiveEngineDaemon_CP_1868_elements(40);
      gj_ReceiveEngineDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	73 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Update/ccr
      -- 
    ccr_2056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(39), ack => call_stmt_1437_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(73) & ReceiveEngineDaemon_CP_1868_elements(41);
      gj_ReceiveEngineDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	35 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Sample/cra
      -- 
    cra_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1437_call_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1437_Update/cca
      -- 
    cca_2057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1437_call_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	37 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Sample/crr
      -- 
    crr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(42), ack => call_stmt_1453_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(37) & ReceiveEngineDaemon_CP_1868_elements(44);
      gj_ReceiveEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	60 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	72 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Update/ccr
      -- 
    ccr_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(43), ack => call_stmt_1453_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(60) & ReceiveEngineDaemon_CP_1868_elements(80) & ReceiveEngineDaemon_CP_1868_elements(72);
      gj_ReceiveEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	35 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Sample/cra
      -- 
    cra_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1453_call_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45: 	78 
    -- CP-element group 45: 	70 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1453_Update/cca
      -- 
    cca_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1453_call_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	37 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_sample_start_
      -- 
    rr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(46), ack => NOT_u1_u1_1456_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(37) & ReceiveEngineDaemon_CP_1868_elements(48);
      gj_ReceiveEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	60 
    -- CP-element group 47: 	72 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Update/cr
      -- CP-element group 47: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_update_start_
      -- 
    cr_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(47), ack => NOT_u1_u1_1456_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(60) & ReceiveEngineDaemon_CP_1868_elements(72);
      gj_ReceiveEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: 	35 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_sample_completed_
      -- 
    ra_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1456_inst_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49: 	70 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1456_update_completed_
      -- 
    ca_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1456_inst_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	37 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Sample/rr
      -- 
    rr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(50), ack => NOT_u1_u1_1466_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(37) & ReceiveEngineDaemon_CP_1868_elements(52);
      gj_ReceiveEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	80 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Update/$entry
      -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(51), ack => NOT_u1_u1_1466_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1868_elements(80);
      gj_ReceiveEngineDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	35 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Sample/ra
      -- 
    ra_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1466_inst_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	78 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/NOT_u1_u1_1466_Update/$exit
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1466_inst_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	20 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Sample/req
      -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(54), ack => W_pkt_cnt_1482_delayed_13_0_1478_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(20) & ReceiveEngineDaemon_CP_1868_elements(56);
      gj_ReceiveEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	60 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Update/req
      -- CP-element group 55: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Update/$entry
      -- 
    req_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(55), ack => W_pkt_cnt_1482_delayed_13_0_1478_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1868_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	18 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Sample/ack
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1482_delayed_13_0_1478_inst_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Update/ack
      -- CP-element group 57: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1480_Update/$exit
      -- 
    ack_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1482_delayed_13_0_1478_inst_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	41 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Sample/crr
      -- CP-element group 58: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_sample_start_
      -- 
    crr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(58), ack => call_stmt_1490_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(45) & ReceiveEngineDaemon_CP_1868_elements(49) & ReceiveEngineDaemon_CP_1868_elements(57) & ReceiveEngineDaemon_CP_1868_elements(41) & ReceiveEngineDaemon_CP_1868_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Update/ccr
      -- CP-element group 59: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_update_start_
      -- 
    ccr_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(59), ack => call_stmt_1490_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1868_elements(61);
      gj_ReceiveEngineDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	47 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	55 
    -- CP-element group 60: 	43 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Sample/cra
      -- CP-element group 60: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_sample_completed_
      -- 
    cra_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1490_call_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	70 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1490_Update/cca
      -- 
    cca_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1490_call_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	20 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Sample/req
      -- CP-element group 62: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_sample_start_
      -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(62), ack => W_pkt_cnt_1487_delayed_13_0_1491_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(20) & ReceiveEngineDaemon_CP_1868_elements(64);
      gj_ReceiveEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Update/req
      -- CP-element group 63: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_update_start_
      -- 
    req_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(63), ack => W_pkt_cnt_1487_delayed_13_0_1491_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(19) & ReceiveEngineDaemon_CP_1868_elements(65);
      gj_ReceiveEngineDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	18 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_sample_completed_
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1487_delayed_13_0_1491_inst_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	83 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	17 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1493_Update/ack
      -- 
    ack_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1487_delayed_13_0_1491_inst_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Sample/req
      -- CP-element group 66: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_sample_start_
      -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(66), ack => W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(37) & ReceiveEngineDaemon_CP_1868_elements(68);
      gj_ReceiveEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	72 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Update/req
      -- CP-element group 67: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_update_start_
      -- 
    req_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(67), ack => W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1868_elements(72);
      gj_ReceiveEngineDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	35 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_sample_completed_
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Update/ack
      -- CP-element group 69: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1507_update_completed_
      -- 
    ack_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	45 
    -- CP-element group 70: 	49 
    -- CP-element group 70: 	61 
    -- CP-element group 70: 	69 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Sample/crr
      -- CP-element group 70: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_sample_start_
      -- 
    crr_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(70), ack => call_stmt_1510_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(45) & ReceiveEngineDaemon_CP_1868_elements(49) & ReceiveEngineDaemon_CP_1868_elements(61) & ReceiveEngineDaemon_CP_1868_elements(69) & ReceiveEngineDaemon_CP_1868_elements(72);
      gj_ReceiveEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Update/ccr
      -- CP-element group 71: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_update_start_
      -- 
    ccr_2168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(71), ack => call_stmt_1510_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1868_elements(73);
      gj_ReceiveEngineDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	47 
    -- CP-element group 72: 	67 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	43 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Sample/cra
      -- CP-element group 72: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_sample_completed_
      -- 
    cra_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1510_call_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	78 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	38 
    -- CP-element group 73: 	39 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_Update/cca
      -- CP-element group 73: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1510_update_completed_
      -- 
    cca_2169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1510_call_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	37 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Sample/req
      -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(74), ack => W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(37) & ReceiveEngineDaemon_CP_1868_elements(76);
      gj_ReceiveEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	80 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Update/req
      -- CP-element group 75: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Update/$entry
      -- 
    req_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(75), ack => W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1868_elements(80);
      gj_ReceiveEngineDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	35 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Sample/ack
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Update/ack
      -- CP-element group 77: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/assign_stmt_1515_Update/$exit
      -- 
    ack_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	45 
    -- CP-element group 78: 	53 
    -- CP-element group 78: 	77 
    -- CP-element group 78: 	73 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Sample/crr
      -- 
    crr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(78), ack => call_stmt_1523_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(45) & ReceiveEngineDaemon_CP_1868_elements(53) & ReceiveEngineDaemon_CP_1868_elements(77) & ReceiveEngineDaemon_CP_1868_elements(73) & ReceiveEngineDaemon_CP_1868_elements(80);
      gj_ReceiveEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_update_start_
      -- CP-element group 79: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Update/ccr
      -- CP-element group 79: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Update/$entry
      -- 
    ccr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(79), ack => call_stmt_1523_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1868_elements(81);
      gj_ReceiveEngineDaemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	51 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	75 
    -- CP-element group 80: 	43 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Sample/cra
      -- CP-element group 80: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Sample/$exit
      -- 
    cra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1523_call_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	34 
    -- CP-element group 81: 	35 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Update/cca
      -- CP-element group 81: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/call_stmt_1523_Update/$exit
      -- 
    cca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1523_call_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(81)); -- 
    -- CP-element group 82:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	14 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	15 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_1868_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_1868_elements(14), ack => ReceiveEngineDaemon_CP_1868_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	65 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	11 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1400/do_while_stmt_1411/do_while_stmt_1411_loop_body/$exit
      -- 
    ReceiveEngineDaemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1868_elements(65) & ReceiveEngineDaemon_CP_1868_elements(81);
      gj_ReceiveEngineDaemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	10 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_exit/ack
      -- CP-element group 84: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_exit/$exit
      -- 
    ack_2202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1411_branch_ack_0, ack => ReceiveEngineDaemon_CP_1868_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	10 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_taken/ack
      -- CP-element group 85: 	 branch_block_stmt_1400/do_while_stmt_1411/loop_taken/$exit
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1411_branch_ack_1, ack => ReceiveEngineDaemon_CP_1868_elements(85)); -- 
    -- CP-element group 86:  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	8 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	4 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1400/do_while_stmt_1411/$exit
      -- 
    ReceiveEngineDaemon_CP_1868_elements(86) <= ReceiveEngineDaemon_CP_1868_elements(8);
    -- CP-element group 87:  merge  branch  transition  place  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	2 
    -- CP-element group 87: 	4 
    -- CP-element group 87: 	5 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	5 
    -- CP-element group 87: 	6 
    -- CP-element group 87:  members (49) 
      -- CP-element group 87: 	 branch_block_stmt_1400/merge_stmt_1402_PhiAck/dummy
      -- CP-element group 87: 	 branch_block_stmt_1400/merge_stmt_1402_PhiAck/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/merge_stmt_1402_PhiAck/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/merge_stmt_1402__exit__
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403__entry__
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_dead_link/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Sample/req
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Update/req
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/BITSEL_u32_u1_1406_inputs/RPIPE_CONTROL_REGISTER_1404/Update/ack
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/BITSEL_u32_u1_1406/SplitProtocol/Update/ca
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Update/cr
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/NOT_u1_u1_1407/SplitProtocol/Update/ca
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_eval_test/branch_req
      -- CP-element group 87: 	 branch_block_stmt_1400/NOT_u1_u1_1407_place
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_if_link/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/if_stmt_1403_else_link/$entry
      -- CP-element group 87: 	 branch_block_stmt_1400/merge_stmt_1402_PhiReqMerge
      -- 
    branch_req_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1868_elements(87), ack => if_stmt_1403_branch_req_0); -- 
    ReceiveEngineDaemon_CP_1868_elements(87) <= OrReduce(ReceiveEngineDaemon_CP_1868_elements(2) & ReceiveEngineDaemon_CP_1868_elements(4) & ReceiveEngineDaemon_CP_1868_elements(5));
    ReceiveEngineDaemon_do_while_stmt_1411_terminator_2207: loop_terminator -- 
      generic map (name => " ReceiveEngineDaemon_do_while_stmt_1411_terminator_2207", max_iterations_in_flight =>31) 
      port map(loop_body_exit => ReceiveEngineDaemon_CP_1868_elements(11),loop_continue => ReceiveEngineDaemon_CP_1868_elements(85),loop_terminate => ReceiveEngineDaemon_CP_1868_elements(84),loop_back => ReceiveEngineDaemon_CP_1868_elements(9),loop_exit => ReceiveEngineDaemon_CP_1868_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1413_phi_seq_2029_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ReceiveEngineDaemon_CP_1868_elements(21);
      ReceiveEngineDaemon_CP_1868_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ReceiveEngineDaemon_CP_1868_elements(28);
      ReceiveEngineDaemon_CP_1868_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= ReceiveEngineDaemon_CP_1868_elements(29);
      ReceiveEngineDaemon_CP_1868_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= ReceiveEngineDaemon_CP_1868_elements(23);
      ReceiveEngineDaemon_CP_1868_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ReceiveEngineDaemon_CP_1868_elements(30);
      ReceiveEngineDaemon_CP_1868_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= ReceiveEngineDaemon_CP_1868_elements(32);
      ReceiveEngineDaemon_CP_1868_elements(24) <= phi_mux_reqs(1);
      phi_stmt_1413_phi_seq_2029 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1413_phi_seq_2029") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ReceiveEngineDaemon_CP_1868_elements(16), 
          phi_sample_ack => ReceiveEngineDaemon_CP_1868_elements(19), 
          phi_update_req => ReceiveEngineDaemon_CP_1868_elements(18), 
          phi_update_ack => ReceiveEngineDaemon_CP_1868_elements(20), 
          phi_mux_ack => ReceiveEngineDaemon_CP_1868_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1981_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ReceiveEngineDaemon_CP_1868_elements(12);
        preds(1)  <= ReceiveEngineDaemon_CP_1868_elements(13);
        entry_tmerge_1981 : transition_merge -- 
          generic map(name => " entry_tmerge_1981")
          port map (preds => preds, symbol_out => ReceiveEngineDaemon_CP_1868_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1406_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1528_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1407_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1459_1459_delayed_10_0_1457 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1461_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1466_1466_delayed_10_0_1467 : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1433_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_1486_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_1404_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1526_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1422_wire : std_logic_vector(35 downto 0);
    signal RPIPE_FREE_Q_1519_wire : std_logic_vector(35 downto 0);
    signal bad_packet_identifier_1453 : std_logic_vector(0 downto 0);
    signal cond_1477 : std_logic_vector(0 downto 0);
    signal free_flag_1472 : std_logic_vector(0 downto 0);
    signal ignore_resp0_1437 : std_logic_vector(31 downto 0);
    signal ignore_resp1_1490 : std_logic_vector(31 downto 0);
    signal konst_1398_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1405_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1434_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1475_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1487_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1527_wire_constant : std_logic_vector(31 downto 0);
    signal npkt_cnt_1500 : std_logic_vector(31 downto 0);
    signal npkt_cnt_1500_1415_buffered : std_logic_vector(31 downto 0);
    signal ok_flag_1463 : std_logic_vector(0 downto 0);
    signal pkt_cnt_1413 : std_logic_vector(31 downto 0);
    signal pkt_cnt_1482_delayed_13_0_1480 : std_logic_vector(31 downto 0);
    signal pkt_cnt_1487_delayed_13_0_1493 : std_logic_vector(31 downto 0);
    signal push_status_1523 : std_logic_vector(0 downto 0);
    signal rx_buffer_pointer_32_1425 : std_logic_vector(31 downto 0);
    signal rx_buffer_pointer_36_1443 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1497_delayed_10_0_1507 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1505_delayed_10_0_1515 : std_logic_vector(35 downto 0);
    signal slice_1521_wire : std_logic_vector(31 downto 0);
    signal status_1425 : std_logic_vector(0 downto 0);
    signal type_cast_1417_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1421_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1430_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1440_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1483_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1498_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1518_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1433_wire_constant <= "1111";
    NOT_u4_u4_1486_wire_constant <= "1111";
    konst_1398_wire_constant <= "000000";
    konst_1405_wire_constant <= "00000000000000000000000000000000";
    konst_1434_wire_constant <= "011000";
    konst_1475_wire_constant <= "1";
    konst_1487_wire_constant <= "011001";
    konst_1527_wire_constant <= "00000000000000000000000000000000";
    type_cast_1417_wire_constant <= "00000000000000000000000000000000";
    type_cast_1421_wire_constant <= "1";
    type_cast_1430_wire_constant <= "0";
    type_cast_1440_wire_constant <= "0000";
    type_cast_1483_wire_constant <= "0";
    type_cast_1498_wire_constant <= "00000000000000000000000000000001";
    type_cast_1518_wire_constant <= "1";
    phi_stmt_1413: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= npkt_cnt_1500_1415_buffered & type_cast_1417_wire_constant;
      req <= phi_stmt_1413_req_0 & phi_stmt_1413_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1413",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1413_ack_0,
          idata => idata,
          odata => pkt_cnt_1413,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1413
    -- flow-through slice operator slice_1521_inst
    slice_1521_wire <= rx_buffer_pointer_36_1505_delayed_10_0_1515(31 downto 0);
    W_pkt_cnt_1482_delayed_13_0_1478_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_cnt_1482_delayed_13_0_1478_inst_req_0;
      W_pkt_cnt_1482_delayed_13_0_1478_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_cnt_1482_delayed_13_0_1478_inst_req_1;
      W_pkt_cnt_1482_delayed_13_0_1478_inst_ack_1<= rack(0);
      W_pkt_cnt_1482_delayed_13_0_1478_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_cnt_1482_delayed_13_0_1478_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_cnt_1413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_cnt_1482_delayed_13_0_1480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pkt_cnt_1487_delayed_13_0_1491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_cnt_1487_delayed_13_0_1491_inst_req_0;
      W_pkt_cnt_1487_delayed_13_0_1491_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_cnt_1487_delayed_13_0_1491_inst_req_1;
      W_pkt_cnt_1487_delayed_13_0_1491_inst_ack_1<= rack(0);
      W_pkt_cnt_1487_delayed_13_0_1491_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_cnt_1487_delayed_13_0_1491_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_cnt_1413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_cnt_1487_delayed_13_0_1493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_req_0;
      W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_req_1;
      W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1497_delayed_10_0_1505_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_1443,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1497_delayed_10_0_1507,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_req_0;
      W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_req_1;
      W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1505_delayed_10_0_1513_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_1443,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1505_delayed_10_0_1515,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    npkt_cnt_1500_1415_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= npkt_cnt_1500_1415_buf_req_0;
      npkt_cnt_1500_1415_buf_ack_0<= wack(0);
      rreq(0) <= npkt_cnt_1500_1415_buf_req_1;
      npkt_cnt_1500_1415_buf_ack_1<= rack(0);
      npkt_cnt_1500_1415_buf : InterlockBuffer generic map ( -- 
        name => "npkt_cnt_1500_1415_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => npkt_cnt_1500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => npkt_cnt_1500_1415_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1411_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1528_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1411_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1411_branch_req_0,
          ack0 => do_while_stmt_1411_branch_ack_0,
          ack1 => do_while_stmt_1411_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1403_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1407_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1403_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1403_branch_req_0,
          ack0 => if_stmt_1403_branch_ack_0,
          ack1 => if_stmt_1403_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1499_inst
    process(pkt_cnt_1487_delayed_13_0_1493) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pkt_cnt_1487_delayed_13_0_1493, type_cast_1498_wire_constant, tmp_var);
      npkt_cnt_1500 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1462_inst
    process(NOT_u1_u1_1459_1459_delayed_10_0_1457, NOT_u1_u1_1461_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1459_1459_delayed_10_0_1457, NOT_u1_u1_1461_wire, tmp_var);
      ok_flag_1463 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1471_inst
    process(NOT_u1_u1_1466_1466_delayed_10_0_1467, bad_packet_identifier_1453) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1466_1466_delayed_10_0_1467, bad_packet_identifier_1453, tmp_var);
      free_flag_1472 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1406_inst
    process(RPIPE_CONTROL_REGISTER_1404_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1404_wire, konst_1405_wire_constant, tmp_var);
      BITSEL_u32_u1_1406_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1528_inst
    process(RPIPE_CONTROL_REGISTER_1526_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1526_wire, konst_1527_wire_constant, tmp_var);
      BITSEL_u32_u1_1528_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_1442_inst
    process(type_cast_1440_wire_constant, rx_buffer_pointer_32_1425) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1440_wire_constant, rx_buffer_pointer_32_1425, tmp_var);
      rx_buffer_pointer_36_1443 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1476_inst
    process(ok_flag_1463) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ok_flag_1463, konst_1475_wire_constant, tmp_var);
      cond_1477 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1407_inst
    process(BITSEL_u32_u1_1406_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1406_wire, tmp_var);
      NOT_u1_u1_1407_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (8) : NOT_u1_u1_1456_inst 
    ApIntNot_group_8: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1425;
      NOT_u1_u1_1459_1459_delayed_10_0_1457 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1456_inst_req_0;
      NOT_u1_u1_1456_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1456_inst_req_1;
      NOT_u1_u1_1456_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_8_gI: SplitGuardInterface generic map(name => "ApIntNot_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- unary operator NOT_u1_u1_1461_inst
    process(bad_packet_identifier_1453) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", bad_packet_identifier_1453, tmp_var);
      NOT_u1_u1_1461_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (10) : NOT_u1_u1_1466_inst 
    ApIntNot_group_10: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1425;
      NOT_u1_u1_1466_1466_delayed_10_0_1467 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1466_inst_req_0;
      NOT_u1_u1_1466_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1466_inst_req_1;
      NOT_u1_u1_1466_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_10_gI: SplitGuardInterface generic map(name => "ApIntNot_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1404_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1526_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1422_wire <= FREE_Q;
    RPIPE_FREE_Q_1519_wire <= FREE_Q;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1397_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_1398_wire_constant;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1425_call 
    popFromQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1425_call_req_0;
      call_stmt_1425_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1425_call_req_1;
      call_stmt_1425_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_0_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1421_wire_constant & RPIPE_FREE_Q_1422_wire;
      rx_buffer_pointer_32_1425 <= data_out(32 downto 1);
      status_1425 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1490_call call_stmt_1437_call 
    AccessRegister_call_group_1: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 4);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1490_call_req_0;
      reqL_unguarded(0) <= call_stmt_1437_call_req_0;
      call_stmt_1490_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1437_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1490_call_req_1;
      reqR_unguarded(0) <= call_stmt_1437_call_req_1;
      call_stmt_1490_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1437_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not status_1425(0);
      guard_vector(1)  <= ok_flag_1463(0);
      AccessRegister_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "AccessRegister_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "AccessRegister_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_1_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1483_wire_constant & NOT_u4_u4_1486_wire_constant & konst_1487_wire_constant & pkt_cnt_1482_delayed_13_0_1480 & type_cast_1430_wire_constant & NOT_u4_u4_1433_wire_constant & konst_1434_wire_constant & rx_buffer_pointer_32_1425;
      ignore_resp1_1490 <= data_out(63 downto 32);
      ignore_resp0_1437 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1453_call 
    loadBuffer_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1453_call_req_0;
      call_stmt_1453_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1453_call_req_1;
      call_stmt_1453_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not status_1425(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadBuffer_call_group_2_gI: SplitGuardInterface generic map(name => "loadBuffer_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1443;
      bad_packet_identifier_1453 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadBuffer_call_reqs(0),
          ackR => loadBuffer_call_acks(0),
          dataR => loadBuffer_call_data(35 downto 0),
          tagR => loadBuffer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => loadBuffer_return_acks(0), -- cross-over
          ackL => loadBuffer_return_reqs(0), -- cross-over
          dataL => loadBuffer_return_data(0 downto 0),
          tagL => loadBuffer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1510_call 
    populateRxQueue_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1510_call_req_0;
      call_stmt_1510_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1510_call_req_1;
      call_stmt_1510_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1463(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      populateRxQueue_call_group_3_gI: SplitGuardInterface generic map(name => "populateRxQueue_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1497_delayed_10_0_1507;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => populateRxQueue_call_reqs(0),
          ackR => populateRxQueue_call_acks(0),
          dataR => populateRxQueue_call_data(35 downto 0),
          tagR => populateRxQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => populateRxQueue_return_acks(0), -- cross-over
          ackL => populateRxQueue_return_reqs(0), -- cross-over
          tagL => populateRxQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1523_call 
    pushIntoQueue_call_group_4: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1523_call_req_0;
      call_stmt_1523_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1523_call_req_1;
      call_stmt_1523_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= free_flag_1472(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_4_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1518_wire_constant & RPIPE_FREE_Q_1519_wire & slice_1521_wire;
      push_status_1523 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end ReceiveEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity SoftwareRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
    CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
    AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
    NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity SoftwareRegisterAccessDaemon;
architecture SoftwareRegisterAccessDaemon_arch of SoftwareRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal SoftwareRegisterAccessDaemon_CP_2226_start: Boolean;
  signal SoftwareRegisterAccessDaemon_CP_2226_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_rwbar_1655_delayed_5_0_1678_inst_ack_1 : boolean;
  signal W_rwbar_1663_delayed_5_0_1688_inst_ack_0 : boolean;
  signal W_rwbar_1663_delayed_5_0_1688_inst_ack_1 : boolean;
  signal W_rwbar_1655_delayed_5_0_1678_inst_req_1 : boolean;
  signal W_rwbar_1663_delayed_5_0_1688_inst_req_0 : boolean;
  signal call_stmt_1687_call_req_0 : boolean;
  signal call_stmt_1687_call_ack_0 : boolean;
  signal phi_stmt_1537_req_1 : boolean;
  signal W_rwbar_1663_delayed_5_0_1688_inst_req_1 : boolean;
  signal do_while_stmt_1535_branch_req_0 : boolean;
  signal phi_stmt_1537_ack_0 : boolean;
  signal do_while_stmt_1535_branch_ack_1 : boolean;
  signal call_stmt_1687_call_ack_1 : boolean;
  signal phi_stmt_1537_req_0 : boolean;
  signal W_rwbar_1655_delayed_5_0_1678_inst_ack_0 : boolean;
  signal W_rwbar_1655_delayed_5_0_1678_inst_req_0 : boolean;
  signal call_stmt_1687_call_req_1 : boolean;
  signal do_while_stmt_1535_branch_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1704_inst_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1704_inst_req_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1704_inst_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1704_inst_req_0 : boolean;
  signal phi_stmt_1543_req_1 : boolean;
  signal phi_stmt_1543_req_0 : boolean;
  signal phi_stmt_1543_ack_0 : boolean;
  signal check_control_regsiter_1646_1547_buf_req_0 : boolean;
  signal check_control_regsiter_1646_1547_buf_ack_0 : boolean;
  signal check_control_regsiter_1646_1547_buf_req_1 : boolean;
  signal check_control_regsiter_1646_1547_buf_ack_1 : boolean;
  signal phi_stmt_1548_req_1 : boolean;
  signal phi_stmt_1548_req_0 : boolean;
  signal phi_stmt_1548_ack_0 : boolean;
  signal check_free_q_1655_1552_buf_req_0 : boolean;
  signal check_free_q_1655_1552_buf_ack_0 : boolean;
  signal check_free_q_1655_1552_buf_req_1 : boolean;
  signal check_free_q_1655_1552_buf_ack_1 : boolean;
  signal phi_stmt_1553_req_1 : boolean;
  signal phi_stmt_1553_req_0 : boolean;
  signal phi_stmt_1553_ack_0 : boolean;
  signal check_num_server_1664_1557_buf_req_0 : boolean;
  signal check_num_server_1664_1557_buf_ack_0 : boolean;
  signal check_num_server_1664_1557_buf_req_1 : boolean;
  signal check_num_server_1664_1557_buf_ack_1 : boolean;
  signal array_obj_ref_1562_load_0_req_0 : boolean;
  signal array_obj_ref_1562_load_0_ack_0 : boolean;
  signal array_obj_ref_1562_load_0_req_1 : boolean;
  signal array_obj_ref_1562_load_0_ack_1 : boolean;
  signal array_obj_ref_1593_load_0_req_0 : boolean;
  signal array_obj_ref_1593_load_0_ack_0 : boolean;
  signal array_obj_ref_1593_load_0_req_1 : boolean;
  signal array_obj_ref_1593_load_0_ack_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1591_inst_req_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1591_inst_ack_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1591_inst_req_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1591_inst_ack_1 : boolean;
  signal array_obj_ref_1598_load_0_req_0 : boolean;
  signal array_obj_ref_1598_load_0_ack_0 : boolean;
  signal array_obj_ref_1598_load_0_req_1 : boolean;
  signal array_obj_ref_1598_load_0_ack_1 : boolean;
  signal W_update_free_q_pipe_1585_delayed_5_0_1600_inst_req_0 : boolean;
  signal W_update_free_q_pipe_1585_delayed_5_0_1600_inst_ack_0 : boolean;
  signal W_update_free_q_pipe_1585_delayed_5_0_1600_inst_req_1 : boolean;
  signal W_update_free_q_pipe_1585_delayed_5_0_1600_inst_ack_1 : boolean;
  signal type_cast_1606_inst_req_0 : boolean;
  signal type_cast_1606_inst_ack_0 : boolean;
  signal type_cast_1606_inst_req_1 : boolean;
  signal type_cast_1606_inst_ack_1 : boolean;
  signal WPIPE_FREE_Q_1604_inst_req_0 : boolean;
  signal WPIPE_FREE_Q_1604_inst_ack_0 : boolean;
  signal WPIPE_FREE_Q_1604_inst_req_1 : boolean;
  signal WPIPE_FREE_Q_1604_inst_ack_1 : boolean;
  signal array_obj_ref_1611_load_0_req_0 : boolean;
  signal array_obj_ref_1611_load_0_ack_0 : boolean;
  signal array_obj_ref_1611_load_0_req_1 : boolean;
  signal array_obj_ref_1611_load_0_ack_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1609_inst_req_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1609_inst_ack_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1609_inst_req_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1609_inst_ack_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1614_inst_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1614_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1614_inst_req_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1614_inst_ack_1 : boolean;
  signal array_obj_ref_1667_load_0_req_0 : boolean;
  signal array_obj_ref_1667_load_0_ack_0 : boolean;
  signal array_obj_ref_1667_load_0_req_1 : boolean;
  signal array_obj_ref_1667_load_0_ack_1 : boolean;
  signal W_index_1659_delayed_5_0_1669_inst_req_0 : boolean;
  signal W_index_1659_delayed_5_0_1669_inst_ack_0 : boolean;
  signal W_index_1659_delayed_5_0_1669_inst_req_1 : boolean;
  signal W_index_1659_delayed_5_0_1669_inst_ack_1 : boolean;
  signal W_wdata_1658_delayed_5_0_1672_inst_req_0 : boolean;
  signal W_wdata_1658_delayed_5_0_1672_inst_ack_0 : boolean;
  signal W_wdata_1658_delayed_5_0_1672_inst_req_1 : boolean;
  signal W_wdata_1658_delayed_5_0_1672_inst_ack_1 : boolean;
  signal W_bmask_1656_delayed_5_0_1675_inst_req_0 : boolean;
  signal W_bmask_1656_delayed_5_0_1675_inst_ack_0 : boolean;
  signal W_bmask_1656_delayed_5_0_1675_inst_req_1 : boolean;
  signal W_bmask_1656_delayed_5_0_1675_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  SoftwareRegisterAccessDaemon_CP_2226_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2226_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2226_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2226_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  SoftwareRegisterAccessDaemon_CP_2226: Block -- control-path 
    signal SoftwareRegisterAccessDaemon_CP_2226_elements: BooleanArray(166 downto 0);
    -- 
  begin -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(0) <= SoftwareRegisterAccessDaemon_CP_2226_start;
    SoftwareRegisterAccessDaemon_CP_2226_symbol <= SoftwareRegisterAccessDaemon_CP_2226_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1534/do_while_stmt_1535__entry__
      -- CP-element group 0: 	 branch_block_stmt_1534/branch_block_stmt_1534__entry__
      -- CP-element group 0: 	 branch_block_stmt_1534/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	166 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1534/branch_block_stmt_1534__exit__
      -- CP-element group 1: 	 branch_block_stmt_1534/do_while_stmt_1535__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1534/$exit
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(166);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1534/do_while_stmt_1535/$entry
      -- CP-element group 2: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535__entry__
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(2) <= SoftwareRegisterAccessDaemon_CP_2226_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	166 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535__exit__
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_back
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	165 
    -- CP-element group 5: 	164 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1534/do_while_stmt_1535/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_exit/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(5) <= SoftwareRegisterAccessDaemon_CP_2226_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	163 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_body_done
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(6) <= SoftwareRegisterAccessDaemon_CP_2226_elements(163);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/back_edge_to_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(7) <= SoftwareRegisterAccessDaemon_CP_2226_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	78 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/first_time_through_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(8) <= SoftwareRegisterAccessDaemon_CP_2226_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	100 
    -- CP-element group 9: 	122 
    -- CP-element group 9: 	115 
    -- CP-element group 9: 	93 
    -- CP-element group 9: 	89 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_root_address_calculated
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	157 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/condition_evaluated
      -- 
    condition_evaluated_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(10), ack => do_while_stmt_1535_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(157) & SoftwareRegisterAccessDaemon_CP_2226_elements(14);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/aggregated_phi_sample_req
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(15) & SoftwareRegisterAccessDaemon_CP_2226_elements(32) & SoftwareRegisterAccessDaemon_CP_2226_elements(51) & SoftwareRegisterAccessDaemon_CP_2226_elements(70) & SoftwareRegisterAccessDaemon_CP_2226_elements(14);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	123 
    -- CP-element group 12: 	163 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_sample_completed_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(17) & SoftwareRegisterAccessDaemon_CP_2226_elements(35) & SoftwareRegisterAccessDaemon_CP_2226_elements(54) & SoftwareRegisterAccessDaemon_CP_2226_elements(73);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(16) & SoftwareRegisterAccessDaemon_CP_2226_elements(33) & SoftwareRegisterAccessDaemon_CP_2226_elements(52) & SoftwareRegisterAccessDaemon_CP_2226_elements(71);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/aggregated_phi_update_ack
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(18) & SoftwareRegisterAccessDaemon_CP_2226_elements(37) & SoftwareRegisterAccessDaemon_CP_2226_elements(56) & SoftwareRegisterAccessDaemon_CP_2226_elements(75);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	95 
    -- CP-element group 16: 	106 
    -- CP-element group 16: 	98 
    -- CP-element group 16: 	117 
    -- CP-element group 16: 	102 
    -- CP-element group 16: 	120 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(95) & SoftwareRegisterAccessDaemon_CP_2226_elements(106) & SoftwareRegisterAccessDaemon_CP_2226_elements(98) & SoftwareRegisterAccessDaemon_CP_2226_elements(117) & SoftwareRegisterAccessDaemon_CP_2226_elements(102) & SoftwareRegisterAccessDaemon_CP_2226_elements(120);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	104 
    -- CP-element group 18: 	119 
    -- CP-element group 18: 	100 
    -- CP-element group 18: 	115 
    -- CP-element group 18: 	97 
    -- CP-element group 18: 	93 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(19) <= SoftwareRegisterAccessDaemon_CP_2226_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_loopback_sample_req_ps
      -- 
    phi_stmt_1537_loopback_sample_req_2265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1537_loopback_sample_req_2265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(20), ack => phi_stmt_1537_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(21) <= SoftwareRegisterAccessDaemon_CP_2226_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_entry_sample_req
      -- 
    phi_stmt_1537_entry_sample_req_2268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1537_entry_sample_req_2268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(22), ack => phi_stmt_1537_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1537_phi_mux_ack_ps
      -- 
    phi_stmt_1537_phi_mux_ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1537_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_sample_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(26) <= SoftwareRegisterAccessDaemon_CP_2226_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1540_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(25), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_sample_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(30) <= SoftwareRegisterAccessDaemon_CP_2226_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1542_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(29), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	125 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	95 
    -- CP-element group 33: 	98 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(95) & SoftwareRegisterAccessDaemon_CP_2226_elements(98);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(34) <= SoftwareRegisterAccessDaemon_CP_2226_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(36) <= SoftwareRegisterAccessDaemon_CP_2226_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	97 
    -- CP-element group 37: 	93 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_update_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(38) <= SoftwareRegisterAccessDaemon_CP_2226_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_loopback_sample_req_ps
      -- 
    phi_stmt_1543_loopback_sample_req_2299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1543_loopback_sample_req_2299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(39), ack => phi_stmt_1543_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(40) <= SoftwareRegisterAccessDaemon_CP_2226_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_entry_sample_req_ps
      -- 
    phi_stmt_1543_entry_sample_req_2302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1543_entry_sample_req_2302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(41), ack => phi_stmt_1543_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1543_phi_mux_ack_ps
      -- 
    phi_stmt_1543_phi_mux_ack_2305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1543_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_sample_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(45) <= SoftwareRegisterAccessDaemon_CP_2226_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1546_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(44), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Sample/req
      -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(47), ack => check_control_regsiter_1646_1547_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Update/req
      -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(48), ack => check_control_regsiter_1646_1547_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Sample/ack
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1646_1547_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_control_regsiter_1547_Update/ack
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1646_1547_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	125 
    -- CP-element group 51: 	12 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	106 
    -- CP-element group 52: 	102 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(106) & SoftwareRegisterAccessDaemon_CP_2226_elements(102);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(53) <= SoftwareRegisterAccessDaemon_CP_2226_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(55) <= SoftwareRegisterAccessDaemon_CP_2226_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	104 
    -- CP-element group 56: 	100 
    -- CP-element group 56: 	14 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_update_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(57) <= SoftwareRegisterAccessDaemon_CP_2226_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_loopback_sample_req_ps
      -- 
    phi_stmt_1548_loopback_sample_req_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1548_loopback_sample_req_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(58), ack => phi_stmt_1548_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(59) <= SoftwareRegisterAccessDaemon_CP_2226_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_entry_sample_req_ps
      -- 
    phi_stmt_1548_entry_sample_req_2346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1548_entry_sample_req_2346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(60), ack => phi_stmt_1548_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1548_phi_mux_ack_ps
      -- 
    phi_stmt_1548_phi_mux_ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1548_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_sample_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(64) <= SoftwareRegisterAccessDaemon_CP_2226_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1551_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(63), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Sample/req
      -- 
    req_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(66), ack => check_free_q_1655_1552_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Update/req
      -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(67), ack => check_free_q_1655_1552_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Sample/ack
      -- 
    ack_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1655_1552_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_free_q_1552_Update/ack
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1655_1552_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	125 
    -- CP-element group 70: 	12 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	117 
    -- CP-element group 71: 	120 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(117) & SoftwareRegisterAccessDaemon_CP_2226_elements(120);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(72) <= SoftwareRegisterAccessDaemon_CP_2226_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(74) <= SoftwareRegisterAccessDaemon_CP_2226_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	119 
    -- CP-element group 75: 	115 
    -- CP-element group 75: 	14 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_update_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(76) <= SoftwareRegisterAccessDaemon_CP_2226_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_loopback_sample_req_ps
      -- 
    phi_stmt_1553_loopback_sample_req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1553_loopback_sample_req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(77), ack => phi_stmt_1553_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(78) <= SoftwareRegisterAccessDaemon_CP_2226_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_entry_sample_req_ps
      -- 
    phi_stmt_1553_entry_sample_req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1553_entry_sample_req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(79), ack => phi_stmt_1553_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/phi_stmt_1553_phi_mux_ack_ps
      -- 
    phi_stmt_1553_phi_mux_ack_2393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1553_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_sample_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_sample_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(83) <= SoftwareRegisterAccessDaemon_CP_2226_elements(84);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	83 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1556_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(82), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Sample/req
      -- 
    req_2414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(85), ack => check_num_server_1664_1557_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_update_start_
      -- CP-element group 86: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Update/req
      -- 
    req_2419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(86), ack => check_num_server_1664_1557_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Sample/ack
      -- 
    ack_2415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1664_1557_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_update_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/R_check_num_server_1557_Update/ack
      -- 
    ack_2420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1664_1557_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	9 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	149 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/word_access_start/$entry
      -- CP-element group 89: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/word_access_start/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/word_access_start/word_0/rr
      -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(89), ack => array_obj_ref_1562_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(91) & SoftwareRegisterAccessDaemon_CP_2226_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_update_start_
      -- CP-element group 90: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/word_access_complete/$entry
      -- CP-element group 90: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/word_access_complete/word_0/$entry
      -- CP-element group 90: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/word_access_complete/word_0/cr
      -- 
    cr_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(90), ack => array_obj_ref_1562_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(92);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	158 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/word_access_start/$exit
      -- CP-element group 91: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/word_access_start/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Sample/word_access_start/word_0/ra
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1562_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(91)); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	163 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/word_access_complete/$exit
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/word_access_complete/word_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/word_access_complete/word_0/ca
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/array_obj_ref_1562_Merge/$entry
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/array_obj_ref_1562_Merge/$exit
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/array_obj_ref_1562_Merge/merge_req
      -- CP-element group 92: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_Update/array_obj_ref_1562_Merge/merge_ack
      -- 
    ca_2450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1562_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: 	18 
    -- CP-element group 93: 	37 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	149 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/word_access_start/$entry
      -- CP-element group 93: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/word_access_start/word_0/$entry
      -- CP-element group 93: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/word_access_start/word_0/rr
      -- 
    rr_2472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(93), ack => array_obj_ref_1593_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(18) & SoftwareRegisterAccessDaemon_CP_2226_elements(37) & SoftwareRegisterAccessDaemon_CP_2226_elements(95) & SoftwareRegisterAccessDaemon_CP_2226_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	98 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/word_access_complete/word_0/cr
      -- 
    cr_2483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(94), ack => array_obj_ref_1593_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(98);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	159 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	16 
    -- CP-element group 95: 	33 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/word_access_start/$exit
      -- CP-element group 95: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Sample/word_access_start/word_0/ra
      -- 
    ra_2473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1593_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/word_access_complete/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/array_obj_ref_1593_Merge/$entry
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/array_obj_ref_1593_Merge/$exit
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/array_obj_ref_1593_Merge/merge_req
      -- CP-element group 96: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_Update/array_obj_ref_1593_Merge/merge_ack
      -- 
    ca_2484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1593_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: 	18 
    -- CP-element group 97: 	37 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Sample/req
      -- 
    req_2497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(97), ack => WPIPE_CONTROL_REGISTER_1591_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 31,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(96) & SoftwareRegisterAccessDaemon_CP_2226_elements(18) & SoftwareRegisterAccessDaemon_CP_2226_elements(37) & SoftwareRegisterAccessDaemon_CP_2226_elements(99);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	16 
    -- CP-element group 98: 	33 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Sample/ack
      -- CP-element group 98: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Update/req
      -- 
    ack_2498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1591_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(98)); -- 
    req_2502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(98), ack => WPIPE_CONTROL_REGISTER_1591_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	163 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_CONTROL_REGISTER_1591_Update/ack
      -- 
    ack_2503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1591_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	9 
    -- CP-element group 100: 	18 
    -- CP-element group 100: 	56 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: 	149 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/word_access_start/$entry
      -- CP-element group 100: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/word_access_start/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/word_access_start/word_0/rr
      -- 
    rr_2520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(100), ack => array_obj_ref_1598_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(18) & SoftwareRegisterAccessDaemon_CP_2226_elements(56) & SoftwareRegisterAccessDaemon_CP_2226_elements(102) & SoftwareRegisterAccessDaemon_CP_2226_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	110 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_update_start_
      -- CP-element group 101: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/word_access_complete/$entry
      -- CP-element group 101: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/word_access_complete/word_0/$entry
      -- CP-element group 101: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/word_access_complete/word_0/cr
      -- 
    cr_2531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(101), ack => array_obj_ref_1598_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	160 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	16 
    -- CP-element group 102: 	52 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/word_access_start/$exit
      -- CP-element group 102: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/word_access_start/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Sample/word_access_start/word_0/ra
      -- 
    ra_2521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1598_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	108 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/word_access_complete/$exit
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/word_access_complete/word_0/$exit
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/word_access_complete/word_0/ca
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/array_obj_ref_1598_Merge/$entry
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/array_obj_ref_1598_Merge/$exit
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/array_obj_ref_1598_Merge/merge_req
      -- CP-element group 103: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_Update/array_obj_ref_1598_Merge/merge_ack
      -- 
    ca_2532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1598_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	18 
    -- CP-element group 104: 	56 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Sample/req
      -- 
    req_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(104), ack => W_update_free_q_pipe_1585_delayed_5_0_1600_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(18) & SoftwareRegisterAccessDaemon_CP_2226_elements(56) & SoftwareRegisterAccessDaemon_CP_2226_elements(106);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	110 
    -- CP-element group 105: 	113 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_update_start_
      -- CP-element group 105: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Update/req
      -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(105), ack => W_update_free_q_pipe_1585_delayed_5_0_1600_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(110) & SoftwareRegisterAccessDaemon_CP_2226_elements(113);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	16 
    -- CP-element group 106: 	52 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Sample/ack
      -- 
    ack_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1585_delayed_5_0_1600_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1602_Update/ack
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1585_delayed_5_0_1600_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: 	103 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Sample/rr
      -- 
    rr_2559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(108), ack => type_cast_1606_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(107) & SoftwareRegisterAccessDaemon_CP_2226_elements(103) & SoftwareRegisterAccessDaemon_CP_2226_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	113 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Update/cr
      -- 
    cr_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(109), ack => type_cast_1606_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(113);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	101 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Sample/ra
      -- 
    ra_2560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/type_cast_1606_Update/ca
      -- 
    ca_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: 	107 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Sample/req
      -- 
    req_2573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(112), ack => WPIPE_FREE_Q_1604_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(111) & SoftwareRegisterAccessDaemon_CP_2226_elements(107) & SoftwareRegisterAccessDaemon_CP_2226_elements(114);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	109 
    -- CP-element group 113: 	105 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Update/req
      -- 
    ack_2574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1604_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(113)); -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(113), ack => WPIPE_FREE_Q_1604_inst_req_1); -- 
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	163 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_FREE_Q_1604_Update/ack
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1604_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	9 
    -- CP-element group 115: 	18 
    -- CP-element group 115: 	75 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: 	149 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/word_access_start/$entry
      -- CP-element group 115: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/word_access_start/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/word_access_start/word_0/rr
      -- 
    rr_2596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(115), ack => array_obj_ref_1611_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(18) & SoftwareRegisterAccessDaemon_CP_2226_elements(75) & SoftwareRegisterAccessDaemon_CP_2226_elements(117) & SoftwareRegisterAccessDaemon_CP_2226_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	120 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/word_access_complete/$entry
      -- CP-element group 116: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/word_access_complete/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/word_access_complete/word_0/cr
      -- 
    cr_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(116), ack => array_obj_ref_1611_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(120);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	161 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	16 
    -- CP-element group 117: 	71 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Sample/word_access_start/word_0/ra
      -- 
    ra_2597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1611_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/array_obj_ref_1611_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/array_obj_ref_1611_Merge/$exit
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/array_obj_ref_1611_Merge/merge_req
      -- CP-element group 118: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_Update/array_obj_ref_1611_Merge/merge_ack
      -- 
    ca_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1611_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: 	18 
    -- CP-element group 119: 	75 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Sample/req
      -- 
    req_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(119), ack => WPIPE_NUMBER_OF_SERVERS_1609_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 31,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(118) & SoftwareRegisterAccessDaemon_CP_2226_elements(18) & SoftwareRegisterAccessDaemon_CP_2226_elements(75) & SoftwareRegisterAccessDaemon_CP_2226_elements(121);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	16 
    -- CP-element group 120: 	71 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_update_start_
      -- CP-element group 120: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Update/req
      -- 
    ack_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1609_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(120)); -- 
    req_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(120), ack => WPIPE_NUMBER_OF_SERVERS_1609_inst_req_1); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	163 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_NUMBER_OF_SERVERS_1609_Update/ack
      -- 
    ack_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1609_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	9 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	125 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Sample/rr
      -- 
    rr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(122), ack => RPIPE_AFB_NIC_REQUEST_1614_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(9) & SoftwareRegisterAccessDaemon_CP_2226_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	12 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	132 
    -- CP-element group 123: 	128 
    -- CP-element group 123: 	140 
    -- CP-element group 123: 	144 
    -- CP-element group 123: 	136 
    -- CP-element group 123: 	152 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_update_start_
      -- CP-element group 123: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Update/cr
      -- 
    cr_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(123), ack => RPIPE_AFB_NIC_REQUEST_1614_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 31,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(124) & SoftwareRegisterAccessDaemon_CP_2226_elements(12) & SoftwareRegisterAccessDaemon_CP_2226_elements(132) & SoftwareRegisterAccessDaemon_CP_2226_elements(128) & SoftwareRegisterAccessDaemon_CP_2226_elements(140) & SoftwareRegisterAccessDaemon_CP_2226_elements(144) & SoftwareRegisterAccessDaemon_CP_2226_elements(136) & SoftwareRegisterAccessDaemon_CP_2226_elements(152);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Sample/ra
      -- 
    ra_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1614_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	130 
    -- CP-element group 125: 	134 
    -- CP-element group 125: 	138 
    -- CP-element group 125: 	126 
    -- CP-element group 125: 	142 
    -- CP-element group 125: 	150 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	32 
    -- CP-element group 125: 	51 
    -- CP-element group 125: 	70 
    -- CP-element group 125:  members (29) 
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/RPIPE_AFB_NIC_REQUEST_1614_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_word_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_root_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_offset_calculated
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_resized_0
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_scaled_0
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_computed_0
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_resize_0/$entry
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_resize_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_resize_0/index_resize_req
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_resize_0/index_resize_ack
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_scale_0/$entry
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_scale_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_scale_0/scale_rename_req
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_index_scale_0/scale_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_final_index_sum_regn/$entry
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_final_index_sum_regn/$exit
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_final_index_sum_regn/req
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_final_index_sum_regn/ack
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_base_plus_offset/$entry
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_base_plus_offset/$exit
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_base_plus_offset/sum_rename_req
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_base_plus_offset/sum_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_word_addrgen/$entry
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_word_addrgen/$exit
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_word_addrgen/root_register_req
      -- CP-element group 125: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_word_addrgen/root_register_ack
      -- 
    ca_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1614_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	128 
    -- CP-element group 126: 	149 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/word_access_start/$entry
      -- CP-element group 126: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/word_access_start/word_0/$entry
      -- CP-element group 126: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/word_access_start/word_0/rr
      -- 
    rr_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(126), ack => array_obj_ref_1667_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(128) & SoftwareRegisterAccessDaemon_CP_2226_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	155 
    -- CP-element group 127: 	148 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_update_start_
      -- CP-element group 127: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/word_access_complete/$entry
      -- CP-element group 127: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/word_access_complete/word_0/$entry
      -- CP-element group 127: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/word_access_complete/word_0/cr
      -- 
    cr_2698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(127), ack => array_obj_ref_1667_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(155) & SoftwareRegisterAccessDaemon_CP_2226_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	162 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	123 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/word_access_start/$exit
      -- CP-element group 128: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/word_access_start/word_0/$exit
      -- CP-element group 128: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Sample/word_access_start/word_0/ra
      -- 
    ra_2688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1667_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	146 
    -- CP-element group 129: 	154 
    -- CP-element group 129:  members (9) 
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/word_access_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/word_access_complete/word_0/$exit
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/word_access_complete/word_0/ca
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/array_obj_ref_1667_Merge/$entry
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/array_obj_ref_1667_Merge/$exit
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/array_obj_ref_1667_Merge/merge_req
      -- CP-element group 129: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_Update/array_obj_ref_1667_Merge/merge_ack
      -- 
    ca_2699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1667_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	125 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Sample/req
      -- 
    req_2712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(130), ack => W_index_1659_delayed_5_0_1669_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(132);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	148 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_update_start_
      -- CP-element group 131: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Update/req
      -- 
    req_2717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(131), ack => W_index_1659_delayed_5_0_1669_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	123 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Sample/ack
      -- 
    ack_2713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1659_delayed_5_0_1669_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	146 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1671_Update/ack
      -- 
    ack_2718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1659_delayed_5_0_1669_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	125 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	136 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Sample/req
      -- 
    req_2726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(134), ack => W_wdata_1658_delayed_5_0_1672_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(136);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	148 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_update_start_
      -- CP-element group 135: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Update/req
      -- 
    req_2731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(135), ack => W_wdata_1658_delayed_5_0_1672_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: 	123 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Sample/ack
      -- 
    ack_2727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1658_delayed_5_0_1672_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	146 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1674_Update/ack
      -- 
    ack_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1658_delayed_5_0_1672_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(137)); -- 
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	125 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Sample/req
      -- 
    req_2740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(138), ack => W_bmask_1656_delayed_5_0_1675_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(140);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	148 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_update_start_
      -- CP-element group 139: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Update/req
      -- 
    req_2745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(139), ack => W_bmask_1656_delayed_5_0_1675_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: 	123 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Sample/ack
      -- 
    ack_2741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1656_delayed_5_0_1675_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	146 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1677_Update/ack
      -- 
    ack_2746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1656_delayed_5_0_1675_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	125 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Sample/req
      -- CP-element group 142: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_sample_start_
      -- 
    req_2754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(142), ack => W_rwbar_1655_delayed_5_0_1678_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(144);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	148 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Update/req
      -- CP-element group 143: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_update_start_
      -- 
    req_2759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(143), ack => W_rwbar_1655_delayed_5_0_1678_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	123 
    -- CP-element group 144: 	142 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Sample/ack
      -- CP-element group 144: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_sample_completed_
      -- 
    ack_2755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1655_delayed_5_0_1678_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Update/ack
      -- CP-element group 145: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1680_Update/$exit
      -- 
    ack_2760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1655_delayed_5_0_1678_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	133 
    -- CP-element group 146: 	129 
    -- CP-element group 146: 	141 
    -- CP-element group 146: 	145 
    -- CP-element group 146: 	137 
    -- CP-element group 146: 	158 
    -- CP-element group 146: 	159 
    -- CP-element group 146: 	160 
    -- CP-element group 146: 	161 
    -- CP-element group 146: 	162 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Sample/crr
      -- CP-element group 146: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_sample_start_
      -- 
    crr_2768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(146), ack => call_stmt_1687_call_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 31,6 => 31,7 => 31,8 => 31,9 => 31,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(133) & SoftwareRegisterAccessDaemon_CP_2226_elements(129) & SoftwareRegisterAccessDaemon_CP_2226_elements(141) & SoftwareRegisterAccessDaemon_CP_2226_elements(145) & SoftwareRegisterAccessDaemon_CP_2226_elements(137) & SoftwareRegisterAccessDaemon_CP_2226_elements(158) & SoftwareRegisterAccessDaemon_CP_2226_elements(159) & SoftwareRegisterAccessDaemon_CP_2226_elements(160) & SoftwareRegisterAccessDaemon_CP_2226_elements(161) & SoftwareRegisterAccessDaemon_CP_2226_elements(162) & SoftwareRegisterAccessDaemon_CP_2226_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_update_start_
      -- CP-element group 147: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Update/ccr
      -- 
    ccr_2773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(147), ack => call_stmt_1687_call_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	131 
    -- CP-element group 148: 	139 
    -- CP-element group 148: 	127 
    -- CP-element group 148: 	143 
    -- CP-element group 148: 	146 
    -- CP-element group 148: 	135 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Sample/cra
      -- CP-element group 148: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Sample/$exit
      -- 
    cra_2769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1687_call_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	163 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	100 
    -- CP-element group 149: 	126 
    -- CP-element group 149: 	115 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	93 
    -- CP-element group 149: 	89 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_Update/cca
      -- CP-element group 149: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/call_stmt_1687_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/ring_reenable_memory_space_0
      -- 
    cca_2774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1687_call_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	125 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_sample_start_
      -- 
    req_2782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(150), ack => W_rwbar_1663_delayed_5_0_1688_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(125) & SoftwareRegisterAccessDaemon_CP_2226_elements(152);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	155 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Update/req
      -- CP-element group 151: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_update_start_
      -- 
    req_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(151), ack => W_rwbar_1663_delayed_5_0_1688_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2226_elements(155);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	123 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Sample/ack
      -- CP-element group 152: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_sample_completed_
      -- 
    ack_2783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1663_delayed_5_0_1688_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Update/ack
      -- CP-element group 153: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/assign_stmt_1690_Update/$exit
      -- 
    ack_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1663_delayed_5_0_1688_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	129 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Sample/req
      -- 
    req_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(154), ack => WPIPE_AFB_NIC_RESPONSE_1704_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(129) & SoftwareRegisterAccessDaemon_CP_2226_elements(153) & SoftwareRegisterAccessDaemon_CP_2226_elements(156);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	127 
    -- CP-element group 155: 	151 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Update/req
      -- CP-element group 155: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Sample/ack
      -- 
    ack_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1704_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(155)); -- 
    req_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2226_elements(155), ack => WPIPE_AFB_NIC_RESPONSE_1704_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	163 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Update/ack
      -- CP-element group 156: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/WPIPE_AFB_NIC_RESPONSE_1704_Update/$exit
      -- 
    ack_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1704_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(9), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	91 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	146 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1562_call_stmt_1687_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(158) is a control-delay.
    cp_element_158_delay: control_delay_element  generic map(name => " 158_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(91), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(158), clk => clk, reset =>reset);
    -- CP-element group 159:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	95 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	146 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1593_call_stmt_1687_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(159) is a control-delay.
    cp_element_159_delay: control_delay_element  generic map(name => " 159_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(95), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(159), clk => clk, reset =>reset);
    -- CP-element group 160:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	102 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	146 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1598_call_stmt_1687_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(160) is a control-delay.
    cp_element_160_delay: control_delay_element  generic map(name => " 160_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(102), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(160), clk => clk, reset =>reset);
    -- CP-element group 161:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	117 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	146 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1611_call_stmt_1687_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(161) is a control-delay.
    cp_element_161_delay: control_delay_element  generic map(name => " 161_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(117), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(161), clk => clk, reset =>reset);
    -- CP-element group 162:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	128 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	146 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/array_obj_ref_1667_call_stmt_1687_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2226_elements(162) is a control-delay.
    cp_element_162_delay: control_delay_element  generic map(name => " 162_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2226_elements(128), ack => SoftwareRegisterAccessDaemon_CP_2226_elements(162), clk => clk, reset =>reset);
    -- CP-element group 163:  join  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	156 
    -- CP-element group 163: 	99 
    -- CP-element group 163: 	121 
    -- CP-element group 163: 	114 
    -- CP-element group 163: 	92 
    -- CP-element group 163: 	149 
    -- CP-element group 163: 	12 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	6 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1534/do_while_stmt_1535/do_while_stmt_1535_loop_body/$exit
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31,6 => 31);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2226_elements(156) & SoftwareRegisterAccessDaemon_CP_2226_elements(99) & SoftwareRegisterAccessDaemon_CP_2226_elements(121) & SoftwareRegisterAccessDaemon_CP_2226_elements(114) & SoftwareRegisterAccessDaemon_CP_2226_elements(92) & SoftwareRegisterAccessDaemon_CP_2226_elements(149) & SoftwareRegisterAccessDaemon_CP_2226_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	5 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_exit/ack
      -- CP-element group 164: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_exit/$exit
      -- 
    ack_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1535_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	5 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_taken/$exit
      -- CP-element group 165: 	 branch_block_stmt_1534/do_while_stmt_1535/loop_taken/ack
      -- 
    ack_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1535_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2226_elements(165)); -- 
    -- CP-element group 166:  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	3 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	1 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_1534/do_while_stmt_1535/$exit
      -- 
    SoftwareRegisterAccessDaemon_CP_2226_elements(166) <= SoftwareRegisterAccessDaemon_CP_2226_elements(3);
    SoftwareRegisterAccessDaemon_do_while_stmt_1535_terminator_2818: loop_terminator -- 
      generic map (name => " SoftwareRegisterAccessDaemon_do_while_stmt_1535_terminator_2818", max_iterations_in_flight =>31) 
      port map(loop_body_exit => SoftwareRegisterAccessDaemon_CP_2226_elements(6),loop_continue => SoftwareRegisterAccessDaemon_CP_2226_elements(165),loop_terminate => SoftwareRegisterAccessDaemon_CP_2226_elements(164),loop_back => SoftwareRegisterAccessDaemon_CP_2226_elements(4),loop_exit => SoftwareRegisterAccessDaemon_CP_2226_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1537_phi_seq_2289_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(21);
      SoftwareRegisterAccessDaemon_CP_2226_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(24);
      SoftwareRegisterAccessDaemon_CP_2226_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(26);
      SoftwareRegisterAccessDaemon_CP_2226_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(19);
      SoftwareRegisterAccessDaemon_CP_2226_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(28);
      SoftwareRegisterAccessDaemon_CP_2226_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(30);
      SoftwareRegisterAccessDaemon_CP_2226_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1537_phi_seq_2289 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1537_phi_seq_2289") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2226_elements(11), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(17), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2226_elements(13), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(18), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1543_phi_seq_2333_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(40);
      SoftwareRegisterAccessDaemon_CP_2226_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(43);
      SoftwareRegisterAccessDaemon_CP_2226_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(45);
      SoftwareRegisterAccessDaemon_CP_2226_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(38);
      SoftwareRegisterAccessDaemon_CP_2226_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(49);
      SoftwareRegisterAccessDaemon_CP_2226_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(50);
      SoftwareRegisterAccessDaemon_CP_2226_elements(39) <= phi_mux_reqs(1);
      phi_stmt_1543_phi_seq_2333 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1543_phi_seq_2333") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2226_elements(34), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(35), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2226_elements(36), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(37), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1548_phi_seq_2377_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(59);
      SoftwareRegisterAccessDaemon_CP_2226_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(62);
      SoftwareRegisterAccessDaemon_CP_2226_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(64);
      SoftwareRegisterAccessDaemon_CP_2226_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(57);
      SoftwareRegisterAccessDaemon_CP_2226_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(68);
      SoftwareRegisterAccessDaemon_CP_2226_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(69);
      SoftwareRegisterAccessDaemon_CP_2226_elements(58) <= phi_mux_reqs(1);
      phi_stmt_1548_phi_seq_2377 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1548_phi_seq_2377") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2226_elements(53), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(54), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2226_elements(55), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(56), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1553_phi_seq_2421_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(78);
      SoftwareRegisterAccessDaemon_CP_2226_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(81);
      SoftwareRegisterAccessDaemon_CP_2226_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(83);
      SoftwareRegisterAccessDaemon_CP_2226_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(76);
      SoftwareRegisterAccessDaemon_CP_2226_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(87);
      SoftwareRegisterAccessDaemon_CP_2226_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(88);
      SoftwareRegisterAccessDaemon_CP_2226_elements(77) <= phi_mux_reqs(1);
      phi_stmt_1553_phi_seq_2421 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1553_phi_seq_2421") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2226_elements(72), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(73), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2226_elements(74), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(75), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2226_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2251_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(7);
        preds(1)  <= SoftwareRegisterAccessDaemon_CP_2226_elements(8);
        entry_tmerge_2251 : transition_merge -- 
          generic map(name => " entry_tmerge_2251")
          port map (preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2226_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1571_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1579_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1587_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1644_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1653_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1662_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1641_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1650_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1659_wire : std_logic_vector(0 downto 0);
    signal FREE_Q_32_1599 : std_logic_vector(31 downto 0);
    signal INIT_1537 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1568_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1576_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1584_wire : std_logic_vector(0 downto 0);
    signal R_index_1666_resized : std_logic_vector(5 downto 0);
    signal R_index_1666_scaled : std_logic_vector(5 downto 0);
    signal addr_1629 : std_logic_vector(35 downto 0);
    signal array_obj_ref_1562_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1562_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1593_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1593_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1593_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1598_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1598_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1611_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1611_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1611_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1667_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1667_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_1667_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1667_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1667_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1667_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1667_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_1625 : std_logic_vector(3 downto 0);
    signal bmask_1656_delayed_5_0_1677 : std_logic_vector(3 downto 0);
    signal check_control_regsiter_1646 : std_logic_vector(0 downto 0);
    signal check_control_regsiter_1646_1547_buffered : std_logic_vector(0 downto 0);
    signal check_free_q_1655 : std_logic_vector(0 downto 0);
    signal check_free_q_1655_1552_buffered : std_logic_vector(0 downto 0);
    signal check_num_server_1664 : std_logic_vector(0 downto 0);
    signal check_num_server_1664_1557_buffered : std_logic_vector(0 downto 0);
    signal control_data_1563 : std_logic_vector(31 downto 0);
    signal control_register_1543 : std_logic_vector(0 downto 0);
    signal free_q_1548 : std_logic_vector(0 downto 0);
    signal index_1637 : std_logic_vector(5 downto 0);
    signal index_1659_delayed_5_0_1671 : std_logic_vector(5 downto 0);
    signal konst_1640_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1643_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1649_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1652_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1658_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1661_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1708_wire_constant : std_logic_vector(0 downto 0);
    signal num_server_1553 : std_logic_vector(0 downto 0);
    signal rdata_1697 : std_logic_vector(31 downto 0);
    signal req_1615 : std_logic_vector(73 downto 0);
    signal resp_1703 : std_logic_vector(32 downto 0);
    signal rval_1668 : std_logic_vector(31 downto 0);
    signal rwbar_1621 : std_logic_vector(0 downto 0);
    signal rwbar_1655_delayed_5_0_1680 : std_logic_vector(0 downto 0);
    signal rwbar_1663_delayed_5_0_1690 : std_logic_vector(0 downto 0);
    signal type_cast_1540_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1542_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1546_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1551_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1556_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1606_wire : std_logic_vector(35 downto 0);
    signal type_cast_1695_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1700_wire_constant : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_1573 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1581 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1585_delayed_5_0_1602 : std_logic_vector(0 downto 0);
    signal update_server_num_1589 : std_logic_vector(0 downto 0);
    signal wdata_1633 : std_logic_vector(31 downto 0);
    signal wdata_1658_delayed_5_0_1674 : std_logic_vector(31 downto 0);
    signal wval_1687 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1562_word_address_0 <= "000000";
    array_obj_ref_1593_word_address_0 <= "000000";
    array_obj_ref_1598_word_address_0 <= "010010";
    array_obj_ref_1611_word_address_0 <= "000001";
    array_obj_ref_1667_offset_scale_factor_0 <= "000001";
    array_obj_ref_1667_resized_base_address <= "000000";
    array_obj_ref_1667_word_offset_0 <= "000000";
    konst_1640_wire_constant <= "000000";
    konst_1643_wire_constant <= "0";
    konst_1649_wire_constant <= "010010";
    konst_1652_wire_constant <= "0";
    konst_1658_wire_constant <= "000001";
    konst_1661_wire_constant <= "0";
    konst_1708_wire_constant <= "1";
    type_cast_1540_wire_constant <= "0";
    type_cast_1542_wire_constant <= "1";
    type_cast_1546_wire_constant <= "0";
    type_cast_1551_wire_constant <= "0";
    type_cast_1556_wire_constant <= "0";
    type_cast_1695_wire_constant <= "00000000000000000000000000000000";
    type_cast_1700_wire_constant <= "0";
    phi_stmt_1537: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1540_wire_constant & type_cast_1542_wire_constant;
      req <= phi_stmt_1537_req_0 & phi_stmt_1537_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1537",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1537_ack_0,
          idata => idata,
          odata => INIT_1537,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1537
    phi_stmt_1543: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1546_wire_constant & check_control_regsiter_1646_1547_buffered;
      req <= phi_stmt_1543_req_0 & phi_stmt_1543_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1543",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1543_ack_0,
          idata => idata,
          odata => control_register_1543,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1543
    phi_stmt_1548: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1551_wire_constant & check_free_q_1655_1552_buffered;
      req <= phi_stmt_1548_req_0 & phi_stmt_1548_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1548",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1548_ack_0,
          idata => idata,
          odata => free_q_1548,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1548
    phi_stmt_1553: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1556_wire_constant & check_num_server_1664_1557_buffered;
      req <= phi_stmt_1553_req_0 & phi_stmt_1553_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1553",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1553_ack_0,
          idata => idata,
          odata => num_server_1553,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1553
    -- flow-through select operator MUX_1696_inst
    rdata_1697 <= rval_1668 when (rwbar_1663_delayed_5_0_1690(0) /=  '0') else type_cast_1695_wire_constant;
    -- flow-through slice operator slice_1620_inst
    rwbar_1621 <= req_1615(72 downto 72);
    -- flow-through slice operator slice_1624_inst
    bmask_1625 <= req_1615(71 downto 68);
    -- flow-through slice operator slice_1628_inst
    addr_1629 <= req_1615(67 downto 32);
    -- flow-through slice operator slice_1632_inst
    wdata_1633 <= req_1615(31 downto 0);
    -- flow-through slice operator slice_1636_inst
    index_1637 <= addr_1629(7 downto 2);
    W_bmask_1656_delayed_5_0_1675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_1656_delayed_5_0_1675_inst_req_0;
      W_bmask_1656_delayed_5_0_1675_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_1656_delayed_5_0_1675_inst_req_1;
      W_bmask_1656_delayed_5_0_1675_inst_ack_1<= rack(0);
      W_bmask_1656_delayed_5_0_1675_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_1656_delayed_5_0_1675_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_1625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_1656_delayed_5_0_1677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_1659_delayed_5_0_1669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_1659_delayed_5_0_1669_inst_req_0;
      W_index_1659_delayed_5_0_1669_inst_ack_0<= wack(0);
      rreq(0) <= W_index_1659_delayed_5_0_1669_inst_req_1;
      W_index_1659_delayed_5_0_1669_inst_ack_1<= rack(0);
      W_index_1659_delayed_5_0_1669_inst : InterlockBuffer generic map ( -- 
        name => "W_index_1659_delayed_5_0_1669_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_1637,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_1659_delayed_5_0_1671,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1655_delayed_5_0_1678_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1655_delayed_5_0_1678_inst_req_0;
      W_rwbar_1655_delayed_5_0_1678_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1655_delayed_5_0_1678_inst_req_1;
      W_rwbar_1655_delayed_5_0_1678_inst_ack_1<= rack(0);
      W_rwbar_1655_delayed_5_0_1678_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1655_delayed_5_0_1678_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1655_delayed_5_0_1680,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1663_delayed_5_0_1688_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1663_delayed_5_0_1688_inst_req_0;
      W_rwbar_1663_delayed_5_0_1688_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1663_delayed_5_0_1688_inst_req_1;
      W_rwbar_1663_delayed_5_0_1688_inst_ack_1<= rack(0);
      W_rwbar_1663_delayed_5_0_1688_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1663_delayed_5_0_1688_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1663_delayed_5_0_1690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_update_free_q_pipe_1585_delayed_5_0_1600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_update_free_q_pipe_1585_delayed_5_0_1600_inst_req_0;
      W_update_free_q_pipe_1585_delayed_5_0_1600_inst_ack_0<= wack(0);
      rreq(0) <= W_update_free_q_pipe_1585_delayed_5_0_1600_inst_req_1;
      W_update_free_q_pipe_1585_delayed_5_0_1600_inst_ack_1<= rack(0);
      W_update_free_q_pipe_1585_delayed_5_0_1600_inst : InterlockBuffer generic map ( -- 
        name => "W_update_free_q_pipe_1585_delayed_5_0_1600_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => update_free_q_pipe_1581,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => update_free_q_pipe_1585_delayed_5_0_1602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_1658_delayed_5_0_1672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_1658_delayed_5_0_1672_inst_req_0;
      W_wdata_1658_delayed_5_0_1672_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_1658_delayed_5_0_1672_inst_req_1;
      W_wdata_1658_delayed_5_0_1672_inst_ack_1<= rack(0);
      W_wdata_1658_delayed_5_0_1672_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_1658_delayed_5_0_1672_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_1633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_1658_delayed_5_0_1674,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_control_regsiter_1646_1547_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_control_regsiter_1646_1547_buf_req_0;
      check_control_regsiter_1646_1547_buf_ack_0<= wack(0);
      rreq(0) <= check_control_regsiter_1646_1547_buf_req_1;
      check_control_regsiter_1646_1547_buf_ack_1<= rack(0);
      check_control_regsiter_1646_1547_buf : InterlockBuffer generic map ( -- 
        name => "check_control_regsiter_1646_1547_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_control_regsiter_1646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_control_regsiter_1646_1547_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_free_q_1655_1552_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_free_q_1655_1552_buf_req_0;
      check_free_q_1655_1552_buf_ack_0<= wack(0);
      rreq(0) <= check_free_q_1655_1552_buf_req_1;
      check_free_q_1655_1552_buf_ack_1<= rack(0);
      check_free_q_1655_1552_buf : InterlockBuffer generic map ( -- 
        name => "check_free_q_1655_1552_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_free_q_1655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_free_q_1655_1552_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_num_server_1664_1557_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_num_server_1664_1557_buf_req_0;
      check_num_server_1664_1557_buf_ack_0<= wack(0);
      rreq(0) <= check_num_server_1664_1557_buf_req_1;
      check_num_server_1664_1557_buf_ack_1<= rack(0);
      check_num_server_1664_1557_buf : InterlockBuffer generic map ( -- 
        name => "check_num_server_1664_1557_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_num_server_1664,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_num_server_1664_1557_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1606_inst_req_0;
      type_cast_1606_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1606_inst_req_1;
      type_cast_1606_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  update_free_q_pipe_1585_delayed_5_0_1602(0);
      type_cast_1606_inst_gI: SplitGuardInterface generic map(name => "type_cast_1606_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => FREE_Q_32_1599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1606_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1562_gather_scatter
    process(array_obj_ref_1562_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1562_data_0;
      ov(31 downto 0) := iv;
      control_data_1563 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1593_gather_scatter
    process(array_obj_ref_1593_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1593_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1593_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1598_gather_scatter
    process(array_obj_ref_1598_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1598_data_0;
      ov(31 downto 0) := iv;
      FREE_Q_32_1599 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1611_gather_scatter
    process(array_obj_ref_1611_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1611_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1611_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1667_addr_0
    process(array_obj_ref_1667_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1667_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_1667_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1667_gather_scatter
    process(array_obj_ref_1667_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1667_data_0;
      ov(31 downto 0) := iv;
      rval_1668 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1667_index_0_rename
    process(R_index_1666_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1666_resized;
      ov(5 downto 0) := iv;
      R_index_1666_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1667_index_0_resize
    process(index_1637) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_1637;
      ov(5 downto 0) := iv;
      R_index_1666_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1667_index_offset
    process(R_index_1666_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1666_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_1667_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1667_root_address_inst
    process(array_obj_ref_1667_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1667_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_1667_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_1535_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1708_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1535_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1535_branch_req_0,
          ack0 => do_while_stmt_1535_branch_ack_0,
          ack1 => do_while_stmt_1535_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1571_inst
    process(INIT_1537, control_register_1543) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1537, control_register_1543, tmp_var);
      AND_u1_u1_1571_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1579_inst
    process(INIT_1537, free_q_1548) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1537, free_q_1548, tmp_var);
      AND_u1_u1_1579_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1587_inst
    process(INIT_1537, num_server_1553) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1537, num_server_1553, tmp_var);
      AND_u1_u1_1587_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1645_inst
    process(EQ_u6_u1_1641_wire, EQ_u1_u1_1644_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1641_wire, EQ_u1_u1_1644_wire, tmp_var);
      check_control_regsiter_1646 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1654_inst
    process(EQ_u6_u1_1650_wire, EQ_u1_u1_1653_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1650_wire, EQ_u1_u1_1653_wire, tmp_var);
      check_free_q_1655 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1663_inst
    process(EQ_u6_u1_1659_wire, EQ_u1_u1_1662_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1659_wire, EQ_u1_u1_1662_wire, tmp_var);
      check_num_server_1664 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_1702_inst
    process(type_cast_1700_wire_constant, rdata_1697) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1700_wire_constant, rdata_1697, tmp_var);
      resp_1703 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1644_inst
    process(rwbar_1621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1621, konst_1643_wire_constant, tmp_var);
      EQ_u1_u1_1644_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1653_inst
    process(rwbar_1621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1621, konst_1652_wire_constant, tmp_var);
      EQ_u1_u1_1653_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1662_inst
    process(rwbar_1621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1621, konst_1661_wire_constant, tmp_var);
      EQ_u1_u1_1662_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1641_inst
    process(index_1637) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1637, konst_1640_wire_constant, tmp_var);
      EQ_u6_u1_1641_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1650_inst
    process(index_1637) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1637, konst_1649_wire_constant, tmp_var);
      EQ_u6_u1_1650_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1659_inst
    process(index_1637) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1637, konst_1658_wire_constant, tmp_var);
      EQ_u6_u1_1659_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1568_inst
    process(INIT_1537) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1537, tmp_var);
      NOT_u1_u1_1568_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1576_inst
    process(INIT_1537) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1537, tmp_var);
      NOT_u1_u1_1576_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1584_inst
    process(INIT_1537) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1537, tmp_var);
      NOT_u1_u1_1584_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1572_inst
    process(NOT_u1_u1_1568_wire, AND_u1_u1_1571_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1568_wire, AND_u1_u1_1571_wire, tmp_var);
      update_control_register_pipe_1573 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1580_inst
    process(NOT_u1_u1_1576_wire, AND_u1_u1_1579_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1576_wire, AND_u1_u1_1579_wire, tmp_var);
      update_free_q_pipe_1581 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1588_inst
    process(NOT_u1_u1_1584_wire, AND_u1_u1_1587_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1584_wire, AND_u1_u1_1587_wire, tmp_var);
      update_server_num_1589 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_1562_load_0 array_obj_ref_1667_load_0 array_obj_ref_1611_load_0 array_obj_ref_1593_load_0 array_obj_ref_1598_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => true, 1 => true, 2 => true, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5, 4 => 5);
      -- 
    begin -- 
      reqL_unguarded(4) <= array_obj_ref_1562_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_1667_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1611_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1593_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1598_load_0_req_0;
      array_obj_ref_1562_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_1667_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1611_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1593_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1598_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= array_obj_ref_1562_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_1667_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1611_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1593_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1598_load_0_req_1;
      array_obj_ref_1562_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_1667_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1611_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1593_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1598_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= update_free_q_pipe_1581(0);
      guard_vector(1)  <= update_control_register_pipe_1573(0);
      guard_vector(2)  <= update_server_num_1589(0);
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1562_word_address_0 & array_obj_ref_1667_word_address_0 & array_obj_ref_1611_word_address_0 & array_obj_ref_1593_word_address_0 & array_obj_ref_1598_word_address_0;
      array_obj_ref_1562_data_0 <= data_out(159 downto 128);
      array_obj_ref_1667_data_0 <= data_out(127 downto 96);
      array_obj_ref_1611_data_0 <= data_out(95 downto 64);
      array_obj_ref_1593_data_0 <= data_out(63 downto 32);
      array_obj_ref_1598_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_AFB_NIC_REQUEST_1614_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(73 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1614_inst_req_0;
      RPIPE_AFB_NIC_REQUEST_1614_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1614_inst_req_1;
      RPIPE_AFB_NIC_REQUEST_1614_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_1615 <= data_out(73 downto 0);
      AFB_NIC_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST_read_0", data_width => 74,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_REQUEST_pipe_read_req(0),
          oack => AFB_NIC_REQUEST_pipe_read_ack(0),
          odata => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_AFB_NIC_RESPONSE_1704_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1704_inst_req_0;
      WPIPE_AFB_NIC_RESPONSE_1704_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1704_inst_req_1;
      WPIPE_AFB_NIC_RESPONSE_1704_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_1703;
      AFB_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_RESPONSE_pipe_write_req(0),
          oack => AFB_NIC_RESPONSE_pipe_write_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_CONTROL_REGISTER_1591_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1591_inst_req_0;
      WPIPE_CONTROL_REGISTER_1591_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1591_inst_req_1;
      WPIPE_CONTROL_REGISTER_1591_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_1573(0);
      data_in <= array_obj_ref_1593_wire;
      CONTROL_REGISTER_write_1_gI: SplitGuardInterface generic map(name => "CONTROL_REGISTER_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      CONTROL_REGISTER_write_1: OutputPortRevised -- 
        generic map ( name => "CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => CONTROL_REGISTER_pipe_write_req(0),
          oack => CONTROL_REGISTER_pipe_write_ack(0),
          odata => CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_FREE_Q_1604_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_FREE_Q_1604_inst_req_0;
      WPIPE_FREE_Q_1604_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_FREE_Q_1604_inst_req_1;
      WPIPE_FREE_Q_1604_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_free_q_pipe_1585_delayed_5_0_1602(0);
      data_in <= type_cast_1606_wire;
      FREE_Q_write_2_gI: SplitGuardInterface generic map(name => "FREE_Q_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      FREE_Q_write_2: OutputPortRevised -- 
        generic map ( name => "FREE_Q", data_width => 36, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => FREE_Q_pipe_write_req(0),
          oack => FREE_Q_pipe_write_ack(0),
          odata => FREE_Q_pipe_write_data(35 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_NUMBER_OF_SERVERS_1609_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1609_inst_req_0;
      WPIPE_NUMBER_OF_SERVERS_1609_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1609_inst_req_1;
      WPIPE_NUMBER_OF_SERVERS_1609_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_server_num_1589(0);
      data_in <= array_obj_ref_1611_wire;
      NUMBER_OF_SERVERS_write_3_gI: SplitGuardInterface generic map(name => "NUMBER_OF_SERVERS_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NUMBER_OF_SERVERS_write_3: OutputPortRevised -- 
        generic map ( name => "NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1687_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1687_call_req_0;
      call_stmt_1687_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1687_call_req_1;
      call_stmt_1687_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_1655_delayed_5_0_1680(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_1656_delayed_5_0_1677 & rval_1668 & wdata_1658_delayed_5_0_1674 & index_1659_delayed_5_0_1671;
      wval_1687 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end SoftwareRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity UpdateRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    bmask : in  std_logic_vector(3 downto 0);
    rval : in  std_logic_vector(31 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    index : in  std_logic_vector(5 downto 0);
    wval : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity UpdateRegister;
architecture UpdateRegister_arch of UpdateRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 74)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal rval_buffer :  std_logic_vector(31 downto 0);
  signal rval_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(5 downto 0);
  signal index_update_enable: Boolean;
  -- output port buffer signals
  signal wval_buffer :  std_logic_vector(31 downto 0);
  signal wval_update_enable: Boolean;
  signal UpdateRegister_CP_34_start: Boolean;
  signal UpdateRegister_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u16_u32_170_inst_req_0 : boolean;
  signal CONCAT_u16_u32_170_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_170_inst_req_1 : boolean;
  signal CONCAT_u16_u32_170_inst_ack_1 : boolean;
  signal array_obj_ref_173_store_0_req_0 : boolean;
  signal array_obj_ref_173_store_0_ack_0 : boolean;
  signal array_obj_ref_173_store_0_req_1 : boolean;
  signal array_obj_ref_173_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "UpdateRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 74) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(3 downto 0) <= bmask;
  bmask_buffer <= in_buffer_data_out(3 downto 0);
  in_buffer_data_in(35 downto 4) <= rval;
  rval_buffer <= in_buffer_data_out(35 downto 4);
  in_buffer_data_in(67 downto 36) <= wdata;
  wdata_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(73 downto 68) <= index;
  index_buffer <= in_buffer_data_out(73 downto 68);
  in_buffer_data_in(tag_length + 73 downto 74) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 73 downto 74);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  UpdateRegister_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "UpdateRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wval_buffer;
  wval <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  UpdateRegister_CP_34: Block -- control-path 
    signal UpdateRegister_CP_34_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    UpdateRegister_CP_34_elements(0) <= UpdateRegister_CP_34_start;
    UpdateRegister_CP_34_symbol <= UpdateRegister_CP_34_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0:  members (39) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_sample_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_update_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/rr
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/cr
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_update_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_offset_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resized_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_computed_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/root_register_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/cr
      -- 
    cr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => array_obj_ref_173_store_0_req_1); -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_170_inst_req_0); -- 
    cr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_170_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_sample_completed_
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_170_inst_ack_0, ack => UpdateRegister_CP_34_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_update_completed_
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/$exit
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/ca
      -- 
    ca_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_170_inst_ack_1, ack => UpdateRegister_CP_34_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_sample_start_
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/$exit
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/split_req
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/split_ack
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/rr
      -- 
    rr_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(3), ack => array_obj_ref_173_store_0_req_0); -- 
    UpdateRegister_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "UpdateRegister_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= UpdateRegister_CP_34_elements(0) & UpdateRegister_CP_34_elements(2);
      gj_UpdateRegister_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => UpdateRegister_CP_34_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_sample_completed_
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/ra
      -- 
    ra_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_store_0_ack_0, ack => UpdateRegister_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_update_completed_
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/ca
      -- 
    ca_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_store_0_ack_1, ack => UpdateRegister_CP_34_elements(5)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_160_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_169_wire : std_logic_vector(15 downto 0);
    signal MUX_155_wire : std_logic_vector(7 downto 0);
    signal MUX_159_wire : std_logic_vector(7 downto 0);
    signal MUX_164_wire : std_logic_vector(7 downto 0);
    signal MUX_168_wire : std_logic_vector(7 downto 0);
    signal R_index_172_resized : std_logic_vector(5 downto 0);
    signal R_index_172_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_173_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_word_offset_0 : std_logic_vector(5 downto 0);
    signal b0_106 : std_logic_vector(0 downto 0);
    signal b1_110 : std_logic_vector(0 downto 0);
    signal b2_114 : std_logic_vector(0 downto 0);
    signal b3_118 : std_logic_vector(0 downto 0);
    signal r0_122 : std_logic_vector(7 downto 0);
    signal r1_126 : std_logic_vector(7 downto 0);
    signal r2_130 : std_logic_vector(7 downto 0);
    signal r3_134 : std_logic_vector(7 downto 0);
    signal w0_138 : std_logic_vector(7 downto 0);
    signal w1_142 : std_logic_vector(7 downto 0);
    signal w2_146 : std_logic_vector(7 downto 0);
    signal w3_150 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_173_offset_scale_factor_0 <= "000001";
    array_obj_ref_173_resized_base_address <= "000000";
    array_obj_ref_173_word_offset_0 <= "000000";
    -- flow-through select operator MUX_155_inst
    MUX_155_wire <= w0_138 when (b0_106(0) /=  '0') else r0_122;
    -- flow-through select operator MUX_159_inst
    MUX_159_wire <= w1_142 when (b1_110(0) /=  '0') else r1_126;
    -- flow-through select operator MUX_164_inst
    MUX_164_wire <= w2_146 when (b2_114(0) /=  '0') else r2_130;
    -- flow-through select operator MUX_168_inst
    MUX_168_wire <= w3_150 when (b3_118(0) /=  '0') else r3_134;
    -- flow-through slice operator slice_105_inst
    b0_106 <= bmask_buffer(3 downto 3);
    -- flow-through slice operator slice_109_inst
    b1_110 <= bmask_buffer(2 downto 2);
    -- flow-through slice operator slice_113_inst
    b2_114 <= bmask_buffer(1 downto 1);
    -- flow-through slice operator slice_117_inst
    b3_118 <= bmask_buffer(0 downto 0);
    -- flow-through slice operator slice_121_inst
    r0_122 <= rval_buffer(31 downto 24);
    -- flow-through slice operator slice_125_inst
    r1_126 <= rval_buffer(23 downto 16);
    -- flow-through slice operator slice_129_inst
    r2_130 <= rval_buffer(15 downto 8);
    -- flow-through slice operator slice_133_inst
    r3_134 <= rval_buffer(7 downto 0);
    -- flow-through slice operator slice_137_inst
    w0_138 <= wdata_buffer(31 downto 24);
    -- flow-through slice operator slice_141_inst
    w1_142 <= wdata_buffer(23 downto 16);
    -- flow-through slice operator slice_145_inst
    w2_146 <= wdata_buffer(15 downto 8);
    -- flow-through slice operator slice_149_inst
    w3_150 <= wdata_buffer(7 downto 0);
    -- equivalence array_obj_ref_173_addr_0
    process(array_obj_ref_173_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_173_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_173_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_gather_scatter
    process(wval_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := wval_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_173_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_0_rename
    process(R_index_172_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_172_resized;
      ov(5 downto 0) := iv;
      R_index_172_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(5 downto 0) := iv;
      R_index_172_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_offset
    process(R_index_172_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_172_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_173_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_root_address_inst
    process(array_obj_ref_173_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_173_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_173_root_address <= ov(5 downto 0);
      --
    end process;
    -- shared split operator group (0) : CONCAT_u16_u32_170_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_160_wire & CONCAT_u8_u16_169_wire;
      wval_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_170_inst_req_0;
      CONCAT_u16_u32_170_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_170_inst_req_1;
      CONCAT_u16_u32_170_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator CONCAT_u8_u16_160_inst
    process(MUX_155_wire, MUX_159_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_155_wire, MUX_159_wire, tmp_var);
      CONCAT_u8_u16_160_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_169_inst
    process(MUX_164_wire, MUX_168_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_164_wire, MUX_168_wire, tmp_var);
      CONCAT_u8_u16_169_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_173_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_173_store_0_req_0;
      array_obj_ref_173_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_173_store_0_req_1;
      array_obj_ref_173_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_173_word_address_0;
      data_in <= array_obj_ref_173_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(5 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end UpdateRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity accessMemory is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(7 downto 0);
    addr : in  std_logic_vector(35 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemory;
architecture accessMemory_arch of accessMemory is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 110)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(7 downto 0);
  signal bmask_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemory_CP_329_start: Boolean;
  signal accessMemory_CP_329_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemory_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 110) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(9 downto 2) <= bmask;
  bmask_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(45 downto 10) <= addr;
  addr_buffer <= in_buffer_data_out(45 downto 10);
  in_buffer_data_in(109 downto 46) <= wdata;
  wdata_buffer <= in_buffer_data_out(109 downto 46);
  in_buffer_data_in(tag_length + 109 downto 110) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 109 downto 110);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= lock_update_enable & rwbar_update_enable & bmask_update_enable & addr_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemory_CP_329_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemory_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_329_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemory_CP_329_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_329_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemory_CP_329: Block -- control-path 
    signal accessMemory_CP_329_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    accessMemory_CP_329_elements(0) <= accessMemory_CP_329_start;
    accessMemory_CP_329_symbol <= accessMemory_CP_329_elements(22);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	11 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_267_to_stmt_287/$entry
      -- 
    accessMemory_CP_329_elements(1) <= accessMemory_CP_329_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_267_to_stmt_287/lock_update_enable
      -- CP-element group 2: 	 assign_stmt_267_to_stmt_287/lock_update_enable_out
      -- 
    accessMemory_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	9 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_267_to_stmt_287/rwbar_update_enable
      -- CP-element group 3: 	 assign_stmt_267_to_stmt_287/rwbar_update_enable_out
      -- 
    accessMemory_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	9 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	18 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_267_to_stmt_287/bmask_update_enable
      -- CP-element group 4: 	 assign_stmt_267_to_stmt_287/bmask_update_enable_out
      -- 
    accessMemory_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	9 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_267_to_stmt_287/addr_update_enable
      -- CP-element group 5: 	 assign_stmt_267_to_stmt_287/addr_update_enable_out
      -- 
    accessMemory_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	20 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_267_to_stmt_287/wdata_update_enable
      -- CP-element group 6: 	 assign_stmt_267_to_stmt_287/wdata_update_enable_out
      -- 
    accessMemory_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	21 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_267_to_stmt_287/rdata_update_enable
      -- CP-element group 7: 	 assign_stmt_267_to_stmt_287/rdata_update_enable_in
      -- 
    accessMemory_CP_329_elements(7) <= accessMemory_CP_329_elements(21);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_sample_start_
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/req
      -- 
    req_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(8), ack => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0); -- 
    accessMemory_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(1) & accessMemory_CP_329_elements(10);
      gj_accessMemory_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	5 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	2 
    -- CP-element group 9: 	3 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_sample_completed_
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_update_start_
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/ack
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/$entry
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/req
      -- 
    ack_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0, ack => accessMemory_CP_329_elements(9)); -- 
    req_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(9), ack => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_update_completed_
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/$exit
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/ack
      -- 
    ack_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1, ack => accessMemory_CP_329_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_sample_start_
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/rr
      -- 
    rr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(11), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0); -- 
    accessMemory_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(1) & accessMemory_CP_329_elements(14);
      gj_accessMemory_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	7 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_update_start_
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/$entry
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/cr
      -- 
    cr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(12), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1); -- 
    accessMemory_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(13) & accessMemory_CP_329_elements(7);
      gj_accessMemory_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	12 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_sample_completed_
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/ra
      -- 
    ra_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0, ack => accessMemory_CP_329_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_update_completed_
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/$exit
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/ca
      -- 
    ca_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1, ack => accessMemory_CP_329_elements(14)); -- 
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 assign_stmt_267_to_stmt_287/$exit
      -- 
    accessMemory_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(14) & accessMemory_CP_329_elements(10);
      gj_accessMemory_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 lock_update_enable
      -- 
    accessMemory_CP_329_elements(16) <= accessMemory_CP_329_elements(2);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 rwbar_update_enable
      -- 
    accessMemory_CP_329_elements(17) <= accessMemory_CP_329_elements(3);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	4 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 bmask_update_enable
      -- 
    accessMemory_CP_329_elements(18) <= accessMemory_CP_329_elements(4);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 addr_update_enable
      -- 
    accessMemory_CP_329_elements(19) <= accessMemory_CP_329_elements(5);
    -- CP-element group 20:  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 wdata_update_enable
      -- 
    accessMemory_CP_329_elements(20) <= accessMemory_CP_329_elements(6);
    -- CP-element group 21:  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	7 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 rdata_update_enable
      -- 
    -- CP-element group 22:  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 $exit
      -- 
    accessMemory_CP_329_elements(22) <= accessMemory_CP_329_elements(15);
    --  hookup: inputs to control-path 
    accessMemory_CP_329_elements(21) <= rdata_update_enable;
    -- hookup: output from control-path 
    lock_update_enable <= accessMemory_CP_329_elements(16);
    rwbar_update_enable <= accessMemory_CP_329_elements(17);
    bmask_update_enable <= accessMemory_CP_329_elements(18);
    addr_update_enable <= accessMemory_CP_329_elements(19);
    wdata_update_enable <= accessMemory_CP_329_elements(20);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_260_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_262_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_265_wire : std_logic_vector(99 downto 0);
    signal err_277 : std_logic_vector(0 downto 0);
    signal request_267 : std_logic_vector(109 downto 0);
    signal response_273 : std_logic_vector(64 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_276_inst
    err_277 <= response_273(64 downto 64);
    -- flow-through slice operator slice_280_inst
    rdata_buffer <= response_273(63 downto 0);
    -- binary operator CONCAT_u10_u110_266_inst
    process(CONCAT_u2_u10_262_wire, CONCAT_u36_u100_265_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_262_wire, CONCAT_u36_u100_265_wire, tmp_var);
      request_267 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_260_inst
    process(lock_buffer, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(lock_buffer, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_260_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u10_262_inst
    process(CONCAT_u1_u2_260_wire, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_260_wire, bmask_buffer, tmp_var);
      CONCAT_u2_u10_262_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_265_inst
    process(addr_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_buffer, wdata_buffer, tmp_var);
      CONCAT_u36_u100_265_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0;
      RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1;
      RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_273 <= data_out(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE_read_0", data_width => 65,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_TO_MEMORY_REQUEST_268_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0;
      WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1;
      WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_267;
      NIC_TO_MEMORY_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_write_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemory_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity acquireLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    m_ok : out  std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity acquireLock;
architecture acquireLock_arch of acquireLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal m_ok_buffer :  std_logic_vector(0 downto 0);
  signal acquireLock_CP_381_start: Boolean;
  signal acquireLock_CP_381_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_311_call_req_1 : boolean;
  signal call_stmt_539_call_ack_1 : boolean;
  signal call_stmt_539_call_req_1 : boolean;
  signal if_stmt_449_branch_ack_0 : boolean;
  signal call_stmt_335_call_ack_1 : boolean;
  signal if_stmt_449_branch_ack_1 : boolean;
  signal call_stmt_335_call_req_1 : boolean;
  signal call_stmt_539_call_ack_0 : boolean;
  signal call_stmt_335_call_ack_0 : boolean;
  signal call_stmt_539_call_req_0 : boolean;
  signal call_stmt_335_call_req_0 : boolean;
  signal call_stmt_466_call_ack_1 : boolean;
  signal call_stmt_466_call_req_1 : boolean;
  signal call_stmt_311_call_ack_0 : boolean;
  signal if_stmt_449_branch_req_0 : boolean;
  signal call_stmt_466_call_ack_0 : boolean;
  signal call_stmt_311_call_req_0 : boolean;
  signal call_stmt_466_call_req_0 : boolean;
  signal call_stmt_311_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "acquireLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  acquireLock_CP_381_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "acquireLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  m_ok_buffer <= "1";
  out_buffer_data_in(0 downto 0) <= m_ok_buffer;
  m_ok <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_381_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= acquireLock_CP_381_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_381_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  acquireLock_CP_381: Block -- control-path 
    signal acquireLock_CP_381_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    acquireLock_CP_381_elements(0) <= acquireLock_CP_381_start;
    acquireLock_CP_381_symbol <= acquireLock_CP_381_elements(10);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_292/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_299__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_299__entry__
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_298__exit__
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_298__entry__
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_299__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_292/branch_block_stmt_292__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_298/$exit
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_298/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_299_dead_link/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	11 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Sample/$exit
      -- 
    cra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_311_call_ack_0, ack => acquireLock_CP_381_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Sample/crr
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Update/cca
      -- 
    cca_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_311_call_ack_1, ack => acquireLock_CP_381_elements(2)); -- 
    crr_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(2), ack => call_stmt_335_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_sample_completed_
      -- 
    cra_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_335_call_ack_0, ack => acquireLock_CP_381_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	11 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448__exit__
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_else_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/EQ_u8_u1_454_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/EQ_u8_u1_454_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/EQ_u8_u1_454_place
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449__entry__
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_449_eval_test/EQ_u8_u1_454/SplitProtocol/Sample/rr
      -- 
    cca_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_335_call_ack_1, ack => acquireLock_CP_381_elements(4)); -- 
    branch_req_459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(4), ack => if_stmt_449_branch_req_0); -- 
    -- CP-element group 5:  fork  transition  place  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (10) 
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466__entry__
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466/$entry
      -- CP-element group 5: 	 branch_block_stmt_292/if_stmt_449_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_292/if_stmt_449_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Update/ccr
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Sample/crr
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_update_start_
      -- 
    if_choice_transition_464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_449_branch_ack_1, ack => acquireLock_CP_381_elements(5)); -- 
    ccr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(5), ack => call_stmt_466_call_req_1); -- 
    crr_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(5), ack => call_stmt_466_call_req_0); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: 	10 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/$entry
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Update/ccr
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_292/if_stmt_449_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_292/if_stmt_449_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_update_start_
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539__entry__
      -- CP-element group 6: 	 branch_block_stmt_292/if_stmt_449__exit__
      -- 
    else_choice_transition_468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_449_branch_ack_0, ack => acquireLock_CP_381_elements(6)); -- 
    ccr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(6), ack => call_stmt_539_call_req_1); -- 
    crr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(6), ack => call_stmt_539_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Sample/cra
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_sample_completed_
      -- 
    cra_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_466_call_ack_0, ack => acquireLock_CP_381_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (8) 
      -- CP-element group 8: 	 branch_block_stmt_292/call_stmt_466__exit__
      -- CP-element group 8: 	 branch_block_stmt_292/call_stmt_466/$exit
      -- CP-element group 8: 	 branch_block_stmt_292/loopback
      -- CP-element group 8: 	 branch_block_stmt_292/loopback_PhiReq/$exit
      -- CP-element group 8: 	 branch_block_stmt_292/loopback_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Update/cca
      -- CP-element group 8: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_292/call_stmt_466/call_stmt_466_update_completed_
      -- 
    cca_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_466_call_ack_1, ack => acquireLock_CP_381_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Sample/cra
      -- CP-element group 9: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_sample_completed_
      -- 
    cra_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_539_call_ack_0, ack => acquireLock_CP_381_elements(9)); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	6 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 branch_block_stmt_292/$exit
      -- CP-element group 10: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Update/cca
      -- CP-element group 10: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/call_stmt_539_update_completed_
      -- CP-element group 10: 	 $exit
      -- CP-element group 10: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539/$exit
      -- CP-element group 10: 	 branch_block_stmt_292/branch_block_stmt_292__exit__
      -- CP-element group 10: 	 assign_stmt_544/$exit
      -- CP-element group 10: 	 assign_stmt_544/$entry
      -- CP-element group 10: 	 branch_block_stmt_292/assign_stmt_525_to_call_stmt_539__exit__
      -- 
    cca_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_539_call_ack_1, ack => acquireLock_CP_381_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: 	4 
    -- CP-element group 11: 	1 
    -- CP-element group 11:  members (16) 
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Update/ccr
      -- CP-element group 11: 	 branch_block_stmt_292/merge_stmt_299_PhiAck/dummy
      -- CP-element group 11: 	 branch_block_stmt_292/merge_stmt_299_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_292/merge_stmt_299_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Update/ccr
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448__entry__
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_292/merge_stmt_299_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/$entry
      -- CP-element group 11: 	 branch_block_stmt_292/merge_stmt_299__exit__
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Sample/crr
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_311_update_start_
      -- CP-element group 11: 	 branch_block_stmt_292/call_stmt_311_to_assign_stmt_448/call_stmt_335_update_start_
      -- 
    ccr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(11), ack => call_stmt_311_call_req_1); -- 
    ccr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(11), ack => call_stmt_335_call_req_1); -- 
    crr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_381_elements(11), ack => call_stmt_311_call_req_0); -- 
    acquireLock_CP_381_elements(11) <= OrReduce(acquireLock_CP_381_elements(8) & acquireLock_CP_381_elements(0));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_482_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_495_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_509_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_522_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_496_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_523_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u4_u36_331_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u4_u36_534_wire : std_logic_vector(35 downto 0);
    signal EQ_u8_u1_454_wire : std_logic_vector(0 downto 0);
    signal MUX_412_wire : std_logic_vector(7 downto 0);
    signal MUX_416_wire : std_logic_vector(7 downto 0);
    signal MUX_421_wire : std_logic_vector(7 downto 0);
    signal MUX_425_wire : std_logic_vector(7 downto 0);
    signal MUX_431_wire : std_logic_vector(7 downto 0);
    signal MUX_435_wire : std_logic_vector(7 downto 0);
    signal MUX_440_wire : std_logic_vector(7 downto 0);
    signal MUX_444_wire : std_logic_vector(7 downto 0);
    signal MUX_475_wire : std_logic_vector(0 downto 0);
    signal MUX_481_wire : std_logic_vector(0 downto 0);
    signal MUX_488_wire : std_logic_vector(0 downto 0);
    signal MUX_494_wire : std_logic_vector(0 downto 0);
    signal MUX_502_wire : std_logic_vector(0 downto 0);
    signal MUX_508_wire : std_logic_vector(0 downto 0);
    signal MUX_515_wire : std_logic_vector(0 downto 0);
    signal MUX_521_wire : std_logic_vector(0 downto 0);
    signal NOT_u64_u64_537_wire_constant : std_logic_vector(63 downto 0);
    signal NOT_u8_u8_306_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_327_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_453_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_461_wire_constant : std_logic_vector(7 downto 0);
    signal OR_u8_u8_417_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_426_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_427_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_436_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_445_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_446_wire : std_logic_vector(7 downto 0);
    signal err_466 : std_logic_vector(63 downto 0);
    signal ignore_539 : std_logic_vector(63 downto 0);
    signal konst_370_wire_constant : std_logic_vector(2 downto 0);
    signal konst_375_wire_constant : std_logic_vector(2 downto 0);
    signal konst_380_wire_constant : std_logic_vector(2 downto 0);
    signal konst_385_wire_constant : std_logic_vector(2 downto 0);
    signal konst_390_wire_constant : std_logic_vector(2 downto 0);
    signal konst_395_wire_constant : std_logic_vector(2 downto 0);
    signal konst_400_wire_constant : std_logic_vector(2 downto 0);
    signal konst_405_wire_constant : std_logic_vector(2 downto 0);
    signal konst_411_wire_constant : std_logic_vector(7 downto 0);
    signal konst_415_wire_constant : std_logic_vector(7 downto 0);
    signal konst_420_wire_constant : std_logic_vector(7 downto 0);
    signal konst_424_wire_constant : std_logic_vector(7 downto 0);
    signal konst_430_wire_constant : std_logic_vector(7 downto 0);
    signal konst_434_wire_constant : std_logic_vector(7 downto 0);
    signal konst_439_wire_constant : std_logic_vector(7 downto 0);
    signal konst_443_wire_constant : std_logic_vector(7 downto 0);
    signal l0_339 : std_logic_vector(7 downto 0);
    signal l1_343 : std_logic_vector(7 downto 0);
    signal l2_347 : std_logic_vector(7 downto 0);
    signal l3_351 : std_logic_vector(7 downto 0);
    signal l4_355 : std_logic_vector(7 downto 0);
    signal l5_359 : std_logic_vector(7 downto 0);
    signal l6_363 : std_logic_vector(7 downto 0);
    signal l7_367 : std_logic_vector(7 downto 0);
    signal lock_addr_32_315 : std_logic_vector(31 downto 0);
    signal lock_address_pointer_298 : std_logic_vector(35 downto 0);
    signal lock_val_448 : std_logic_vector(7 downto 0);
    signal lock_values_335 : std_logic_vector(63 downto 0);
    signal msg_size_plus_lock_311 : std_logic_vector(63 downto 0);
    signal new_bmask_525 : std_logic_vector(7 downto 0);
    signal s0_372 : std_logic_vector(0 downto 0);
    signal s1_377 : std_logic_vector(0 downto 0);
    signal s2_382 : std_logic_vector(0 downto 0);
    signal s3_387 : std_logic_vector(0 downto 0);
    signal s4_392 : std_logic_vector(0 downto 0);
    signal s5_397 : std_logic_vector(0 downto 0);
    signal s6_402 : std_logic_vector(0 downto 0);
    signal s7_407 : std_logic_vector(0 downto 0);
    signal sel_320 : std_logic_vector(2 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_301_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_303_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_309_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_322_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_324_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_329_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_333_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_456_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_464_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_472_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_474_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_480_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_485_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_487_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_491_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_493_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_501_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_505_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_507_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_514_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_518_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_527_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_529_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_532_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    NOT_u64_u64_537_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    NOT_u8_u8_306_wire_constant <= "11111111";
    NOT_u8_u8_327_wire_constant <= "11111111";
    NOT_u8_u8_453_wire_constant <= "11111111";
    NOT_u8_u8_461_wire_constant <= "11111111";
    konst_370_wire_constant <= "000";
    konst_375_wire_constant <= "001";
    konst_380_wire_constant <= "010";
    konst_385_wire_constant <= "011";
    konst_390_wire_constant <= "100";
    konst_395_wire_constant <= "101";
    konst_400_wire_constant <= "110";
    konst_405_wire_constant <= "111";
    konst_411_wire_constant <= "00000000";
    konst_415_wire_constant <= "00000000";
    konst_420_wire_constant <= "00000000";
    konst_424_wire_constant <= "00000000";
    konst_430_wire_constant <= "00000000";
    konst_434_wire_constant <= "00000000";
    konst_439_wire_constant <= "00000000";
    konst_443_wire_constant <= "00000000";
    type_cast_296_wire_constant <= "000000000000000000000000000000010000";
    type_cast_301_wire_constant <= "1";
    type_cast_303_wire_constant <= "1";
    type_cast_309_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_322_wire_constant <= "1";
    type_cast_324_wire_constant <= "1";
    type_cast_329_wire_constant <= "0000";
    type_cast_333_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_456_wire_constant <= "0";
    type_cast_458_wire_constant <= "1";
    type_cast_464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_472_wire_constant <= "1";
    type_cast_474_wire_constant <= "0";
    type_cast_478_wire_constant <= "1";
    type_cast_480_wire_constant <= "0";
    type_cast_485_wire_constant <= "1";
    type_cast_487_wire_constant <= "0";
    type_cast_491_wire_constant <= "1";
    type_cast_493_wire_constant <= "0";
    type_cast_499_wire_constant <= "1";
    type_cast_501_wire_constant <= "0";
    type_cast_505_wire_constant <= "1";
    type_cast_507_wire_constant <= "0";
    type_cast_512_wire_constant <= "1";
    type_cast_514_wire_constant <= "0";
    type_cast_518_wire_constant <= "1";
    type_cast_520_wire_constant <= "0";
    type_cast_527_wire_constant <= "0";
    type_cast_529_wire_constant <= "0";
    type_cast_532_wire_constant <= "0000";
    -- flow-through select operator MUX_412_inst
    MUX_412_wire <= l0_339 when (s0_372(0) /=  '0') else konst_411_wire_constant;
    -- flow-through select operator MUX_416_inst
    MUX_416_wire <= l1_343 when (s1_377(0) /=  '0') else konst_415_wire_constant;
    -- flow-through select operator MUX_421_inst
    MUX_421_wire <= l2_347 when (s2_382(0) /=  '0') else konst_420_wire_constant;
    -- flow-through select operator MUX_425_inst
    MUX_425_wire <= l3_351 when (s3_387(0) /=  '0') else konst_424_wire_constant;
    -- flow-through select operator MUX_431_inst
    MUX_431_wire <= l4_355 when (s4_392(0) /=  '0') else konst_430_wire_constant;
    -- flow-through select operator MUX_435_inst
    MUX_435_wire <= l5_359 when (s5_397(0) /=  '0') else konst_434_wire_constant;
    -- flow-through select operator MUX_440_inst
    MUX_440_wire <= l6_363 when (s6_402(0) /=  '0') else konst_439_wire_constant;
    -- flow-through select operator MUX_444_inst
    MUX_444_wire <= l7_367 when (s7_407(0) /=  '0') else konst_443_wire_constant;
    -- flow-through select operator MUX_475_inst
    MUX_475_wire <= type_cast_472_wire_constant when (s0_372(0) /=  '0') else type_cast_474_wire_constant;
    -- flow-through select operator MUX_481_inst
    MUX_481_wire <= type_cast_478_wire_constant when (s1_377(0) /=  '0') else type_cast_480_wire_constant;
    -- flow-through select operator MUX_488_inst
    MUX_488_wire <= type_cast_485_wire_constant when (s2_382(0) /=  '0') else type_cast_487_wire_constant;
    -- flow-through select operator MUX_494_inst
    MUX_494_wire <= type_cast_491_wire_constant when (s3_387(0) /=  '0') else type_cast_493_wire_constant;
    -- flow-through select operator MUX_502_inst
    MUX_502_wire <= type_cast_499_wire_constant when (s4_392(0) /=  '0') else type_cast_501_wire_constant;
    -- flow-through select operator MUX_508_inst
    MUX_508_wire <= type_cast_505_wire_constant when (s5_397(0) /=  '0') else type_cast_507_wire_constant;
    -- flow-through select operator MUX_515_inst
    MUX_515_wire <= type_cast_512_wire_constant when (s6_402(0) /=  '0') else type_cast_514_wire_constant;
    -- flow-through select operator MUX_521_inst
    MUX_521_wire <= type_cast_518_wire_constant when (s7_407(0) /=  '0') else type_cast_520_wire_constant;
    -- flow-through slice operator slice_314_inst
    lock_addr_32_315 <= msg_size_plus_lock_311(31 downto 0);
    -- flow-through slice operator slice_319_inst
    sel_320 <= lock_addr_32_315(2 downto 0);
    -- flow-through slice operator slice_338_inst
    l0_339 <= lock_values_335(63 downto 56);
    -- flow-through slice operator slice_342_inst
    l1_343 <= lock_values_335(55 downto 48);
    -- flow-through slice operator slice_346_inst
    l2_347 <= lock_values_335(47 downto 40);
    -- flow-through slice operator slice_350_inst
    l3_351 <= lock_values_335(39 downto 32);
    -- flow-through slice operator slice_354_inst
    l4_355 <= lock_values_335(31 downto 24);
    -- flow-through slice operator slice_358_inst
    l5_359 <= lock_values_335(23 downto 16);
    -- flow-through slice operator slice_362_inst
    l6_363 <= lock_values_335(15 downto 8);
    -- flow-through slice operator slice_366_inst
    l7_367 <= lock_values_335(7 downto 0);
    if_stmt_449_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u8_u1_454_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_449_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_449_branch_req_0,
          ack0 => if_stmt_449_branch_ack_0,
          ack1 => if_stmt_449_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u36_u36_297_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_296_wire_constant, tmp_var);
      lock_address_pointer_298 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_482_inst
    process(MUX_475_wire, MUX_481_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_475_wire, MUX_481_wire, tmp_var);
      CONCAT_u1_u2_482_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_495_inst
    process(MUX_488_wire, MUX_494_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_488_wire, MUX_494_wire, tmp_var);
      CONCAT_u1_u2_495_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_509_inst
    process(MUX_502_wire, MUX_508_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_502_wire, MUX_508_wire, tmp_var);
      CONCAT_u1_u2_509_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_522_inst
    process(MUX_515_wire, MUX_521_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_515_wire, MUX_521_wire, tmp_var);
      CONCAT_u1_u2_522_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_496_inst
    process(CONCAT_u1_u2_482_wire, CONCAT_u1_u2_495_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_482_wire, CONCAT_u1_u2_495_wire, tmp_var);
      CONCAT_u2_u4_496_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_523_inst
    process(CONCAT_u1_u2_509_wire, CONCAT_u1_u2_522_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_509_wire, CONCAT_u1_u2_522_wire, tmp_var);
      CONCAT_u2_u4_523_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_331_inst
    process(type_cast_329_wire_constant, lock_addr_32_315) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_329_wire_constant, lock_addr_32_315, tmp_var);
      CONCAT_u4_u36_331_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_534_inst
    process(type_cast_532_wire_constant, lock_addr_32_315) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_532_wire_constant, lock_addr_32_315, tmp_var);
      CONCAT_u4_u36_534_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_524_inst
    process(CONCAT_u2_u4_496_wire, CONCAT_u2_u4_523_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_496_wire, CONCAT_u2_u4_523_wire, tmp_var);
      new_bmask_525 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_371_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_370_wire_constant, tmp_var);
      s0_372 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_376_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_375_wire_constant, tmp_var);
      s1_377 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_381_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_380_wire_constant, tmp_var);
      s2_382 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_386_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_385_wire_constant, tmp_var);
      s3_387 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_391_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_390_wire_constant, tmp_var);
      s4_392 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_396_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_395_wire_constant, tmp_var);
      s5_397 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_401_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_400_wire_constant, tmp_var);
      s6_402 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_406_inst
    process(sel_320) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_320, konst_405_wire_constant, tmp_var);
      s7_407 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_454_inst
    process(lock_val_448) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(lock_val_448, NOT_u8_u8_453_wire_constant, tmp_var);
      EQ_u8_u1_454_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_417_inst
    process(MUX_412_wire, MUX_416_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_412_wire, MUX_416_wire, tmp_var);
      OR_u8_u8_417_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_426_inst
    process(MUX_421_wire, MUX_425_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_421_wire, MUX_425_wire, tmp_var);
      OR_u8_u8_426_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_427_inst
    process(OR_u8_u8_417_wire, OR_u8_u8_426_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_417_wire, OR_u8_u8_426_wire, tmp_var);
      OR_u8_u8_427_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_436_inst
    process(MUX_431_wire, MUX_435_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_431_wire, MUX_435_wire, tmp_var);
      OR_u8_u8_436_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_445_inst
    process(MUX_440_wire, MUX_444_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_440_wire, MUX_444_wire, tmp_var);
      OR_u8_u8_445_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_446_inst
    process(OR_u8_u8_436_wire, OR_u8_u8_445_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_436_wire, OR_u8_u8_445_wire, tmp_var);
      OR_u8_u8_446_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_447_inst
    process(OR_u8_u8_427_wire, OR_u8_u8_446_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_427_wire, OR_u8_u8_446_wire, tmp_var);
      lock_val_448 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_311_call call_stmt_539_call call_stmt_466_call call_stmt_335_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(439 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= call_stmt_311_call_req_0;
      reqL_unguarded(2) <= call_stmt_539_call_req_0;
      reqL_unguarded(1) <= call_stmt_466_call_req_0;
      reqL_unguarded(0) <= call_stmt_335_call_req_0;
      call_stmt_311_call_ack_0 <= ackL_unguarded(3);
      call_stmt_539_call_ack_0 <= ackL_unguarded(2);
      call_stmt_466_call_ack_0 <= ackL_unguarded(1);
      call_stmt_335_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= call_stmt_311_call_req_1;
      reqR_unguarded(2) <= call_stmt_539_call_req_1;
      reqR_unguarded(1) <= call_stmt_466_call_req_1;
      reqR_unguarded(0) <= call_stmt_335_call_req_1;
      call_stmt_311_call_ack_1 <= ackR_unguarded(3);
      call_stmt_539_call_ack_1 <= ackR_unguarded(2);
      call_stmt_466_call_ack_1 <= ackR_unguarded(1);
      call_stmt_335_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_3: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_301_wire_constant & type_cast_303_wire_constant & NOT_u8_u8_306_wire_constant & lock_address_pointer_298 & type_cast_309_wire_constant & type_cast_527_wire_constant & type_cast_529_wire_constant & new_bmask_525 & CONCAT_u4_u36_534_wire & NOT_u64_u64_537_wire_constant & type_cast_456_wire_constant & type_cast_458_wire_constant & NOT_u8_u8_461_wire_constant & lock_address_pointer_298 & type_cast_464_wire_constant & type_cast_322_wire_constant & type_cast_324_wire_constant & NOT_u8_u8_327_wire_constant & CONCAT_u4_u36_331_wire & type_cast_333_wire_constant;
      msg_size_plus_lock_311 <= data_out(255 downto 192);
      ignore_539 <= data_out(191 downto 128);
      err_466 <= data_out(127 downto 64);
      lock_values_335 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 440,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 4,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 256,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 4) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end acquireLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity delay_time_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    T : in  std_logic_vector(31 downto 0);
    delay_done : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity delay_time_Operator;
architecture delay_time_Operator_arch of delay_time_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal T_buffer :  std_logic_vector(31 downto 0);
  signal T_update_enable: Boolean;
  signal T_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal delay_done_buffer :  std_logic_vector(0 downto 0);
  signal delay_time_CP_1459_start: Boolean;
  signal delay_time_CP_1459_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1288_branch_ack_1 : boolean;
  signal nR_1299_1292_buf_ack_1 : boolean;
  signal nR_1299_1292_buf_req_1 : boolean;
  signal phi_stmt_1290_req_1 : boolean;
  signal do_while_stmt_1288_branch_ack_0 : boolean;
  signal nR_1299_1292_buf_req_0 : boolean;
  signal nR_1299_1292_buf_ack_0 : boolean;
  signal do_while_stmt_1288_branch_req_0 : boolean;
  signal T_1293_buf_ack_1 : boolean;
  signal T_1293_buf_req_1 : boolean;
  signal phi_stmt_1290_ack_0 : boolean;
  signal phi_stmt_1290_req_0 : boolean;
  signal T_1293_buf_ack_0 : boolean;
  signal T_1293_buf_req_0 : boolean;
  -- 
begin --  
  sample_ack <= delay_time_CP_1459_symbol;
  -- input handling ------------------------------------------------
  T_buffer <= T;
  delay_time_CP_1459_start <= sample_req;
  -- output handling  -------------------------------------------------------
  delay_done_buffer <= "1";
  delay_done <= delay_done_buffer;
  update_ack_symbol <= delay_time_CP_1459_symbol;
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  delay_time_CP_1459: Block -- control-path 
    signal delay_time_CP_1459_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    delay_time_CP_1459_elements(0) <= delay_time_CP_1459_start;
    delay_time_CP_1459_symbol <= delay_time_CP_1459_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1287/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1287/do_while_stmt_1288__entry__
      -- CP-element group 0: 	 branch_block_stmt_1287/branch_block_stmt_1287__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	32 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (8) 
      -- CP-element group 1: 	 branch_block_stmt_1287/assign_stmt_1306/$entry
      -- CP-element group 1: 	 branch_block_stmt_1287/assign_stmt_1306/$exit
      -- CP-element group 1: 	 branch_block_stmt_1287/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1287/assign_stmt_1306__exit__
      -- CP-element group 1: 	 branch_block_stmt_1287/assign_stmt_1306__entry__
      -- CP-element group 1: 	 branch_block_stmt_1287/do_while_stmt_1288__exit__
      -- CP-element group 1: 	 branch_block_stmt_1287/branch_block_stmt_1287__exit__
      -- 
    delay_time_CP_1459_elements(1) <= delay_time_CP_1459_elements(32);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1287/do_while_stmt_1288/$entry
      -- CP-element group 2: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288__entry__
      -- 
    delay_time_CP_1459_elements(2) <= delay_time_CP_1459_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	32 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288__exit__
      -- 
    -- Element group delay_time_CP_1459_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_back
      -- 
    -- Element group delay_time_CP_1459_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	31 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1287/do_while_stmt_1288/condition_done
      -- 
    delay_time_CP_1459_elements(5) <= delay_time_CP_1459_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	14 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_body_done
      -- 
    delay_time_CP_1459_elements(6) <= delay_time_CP_1459_elements(14);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/back_edge_to_loop_body
      -- 
    delay_time_CP_1459_elements(7) <= delay_time_CP_1459_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/first_time_through_loop_body
      -- 
    delay_time_CP_1459_elements(8) <= delay_time_CP_1459_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	29 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/$entry
      -- 
    -- Element group delay_time_CP_1459_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	29 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/condition_evaluated
      -- 
    condition_evaluated_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1459_elements(10), ack => do_while_stmt_1288_branch_req_0); -- 
    delay_time_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1459_elements(15) & delay_time_CP_1459_elements(29);
      gj_delay_time_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1459_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/aggregated_phi_sample_req
      -- 
    delay_time_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1459_elements(12) & delay_time_CP_1459_elements(15);
      gj_delay_time_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1459_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_sample_start_
      -- 
    delay_time_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1459_elements(9) & delay_time_CP_1459_elements(14);
      gj_delay_time_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1459_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_update_start_
      -- 
    delay_time_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1459_elements(9) & delay_time_CP_1459_elements(15);
      gj_delay_time_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1459_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_sample_completed__ps
      -- CP-element group 14: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/$exit
      -- 
    -- Element group delay_time_CP_1459_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_update_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_update_completed_
      -- 
    -- Element group delay_time_CP_1459_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_loopback_trigger
      -- 
    delay_time_CP_1459_elements(16) <= delay_time_CP_1459_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_loopback_sample_req_ps
      -- CP-element group 17: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_loopback_sample_req
      -- 
    phi_stmt_1290_loopback_sample_req_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1290_loopback_sample_req_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1459_elements(17), ack => phi_stmt_1290_req_0); -- 
    -- Element group delay_time_CP_1459_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_entry_trigger
      -- 
    delay_time_CP_1459_elements(18) <= delay_time_CP_1459_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_entry_sample_req_ps
      -- 
    phi_stmt_1290_entry_sample_req_1503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1290_entry_sample_req_1503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1459_elements(19), ack => phi_stmt_1290_req_1); -- 
    -- Element group delay_time_CP_1459_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/phi_stmt_1290_phi_mux_ack_ps
      -- 
    phi_stmt_1290_phi_mux_ack_1506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1290_ack_0, ack => delay_time_CP_1459_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Sample/req
      -- CP-element group 21: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_sample_start__ps
      -- 
    req_1519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1459_elements(21), ack => nR_1299_1292_buf_req_0); -- 
    -- Element group delay_time_CP_1459_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Update/req
      -- CP-element group 22: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_update_start__ps
      -- 
    req_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1459_elements(22), ack => nR_1299_1292_buf_req_1); -- 
    -- Element group delay_time_CP_1459_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Sample/ack
      -- CP-element group 23: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_sample_completed__ps
      -- 
    ack_1520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1299_1292_buf_ack_0, ack => delay_time_CP_1459_elements(23)); -- 
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Update/ack
      -- CP-element group 24: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_nR_1292_update_completed__ps
      -- 
    ack_1525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1299_1292_buf_ack_1, ack => delay_time_CP_1459_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Sample/req
      -- CP-element group 25: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Sample/$entry
      -- 
    req_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1459_elements(25), ack => T_1293_buf_req_0); -- 
    -- Element group delay_time_CP_1459_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Update/req
      -- CP-element group 26: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_update_start_
      -- 
    req_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1459_elements(26), ack => T_1293_buf_req_1); -- 
    -- Element group delay_time_CP_1459_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Sample/$exit
      -- 
    ack_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1293_buf_ack_0, ack => delay_time_CP_1459_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Update/ack
      -- CP-element group 28: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/R_T_1293_Update/$exit
      -- 
    ack_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1293_buf_ack_1, ack => delay_time_CP_1459_elements(28)); -- 
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	9 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	10 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1287/do_while_stmt_1288/do_while_stmt_1288_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group delay_time_CP_1459_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => delay_time_CP_1459_elements(9), ack => delay_time_CP_1459_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_exit/ack
      -- CP-element group 30: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_exit/$exit
      -- 
    ack_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1288_branch_ack_0, ack => delay_time_CP_1459_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_taken/$exit
      -- CP-element group 31: 	 branch_block_stmt_1287/do_while_stmt_1288/loop_taken/ack
      -- 
    ack_1553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1288_branch_ack_1, ack => delay_time_CP_1459_elements(31)); -- 
    -- CP-element group 32:  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	3 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	1 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1287/do_while_stmt_1288/$exit
      -- 
    delay_time_CP_1459_elements(32) <= delay_time_CP_1459_elements(3);
    delay_time_do_while_stmt_1288_terminator_1554: loop_terminator -- 
      generic map (name => " delay_time_do_while_stmt_1288_terminator_1554", max_iterations_in_flight =>7) 
      port map(loop_body_exit => delay_time_CP_1459_elements(6),loop_continue => delay_time_CP_1459_elements(31),loop_terminate => delay_time_CP_1459_elements(30),loop_back => delay_time_CP_1459_elements(4),loop_exit => delay_time_CP_1459_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1290_phi_seq_1544_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= delay_time_CP_1459_elements(16);
      delay_time_CP_1459_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= delay_time_CP_1459_elements(23);
      delay_time_CP_1459_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= delay_time_CP_1459_elements(24);
      delay_time_CP_1459_elements(17) <= phi_mux_reqs(0);
      triggers(1)  <= delay_time_CP_1459_elements(18);
      delay_time_CP_1459_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= delay_time_CP_1459_elements(27);
      delay_time_CP_1459_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= delay_time_CP_1459_elements(28);
      delay_time_CP_1459_elements(19) <= phi_mux_reqs(1);
      phi_stmt_1290_phi_seq_1544 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1290_phi_seq_1544") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => delay_time_CP_1459_elements(11), 
          phi_sample_ack => delay_time_CP_1459_elements(14), 
          phi_update_req => delay_time_CP_1459_elements(13), 
          phi_update_ack => delay_time_CP_1459_elements(15), 
          phi_mux_ack => delay_time_CP_1459_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1486_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= delay_time_CP_1459_elements(7);
        preds(1)  <= delay_time_CP_1459_elements(8);
        entry_tmerge_1486 : transition_merge -- 
          generic map(name => " entry_tmerge_1486")
          port map (preds => preds, symbol_out => delay_time_CP_1459_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_1290 : std_logic_vector(31 downto 0);
    signal T_1293_buffered : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_1303_wire : std_logic_vector(0 downto 0);
    signal konst_1297_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1302_wire_constant : std_logic_vector(31 downto 0);
    signal nR_1299 : std_logic_vector(31 downto 0);
    signal nR_1299_1292_buffered : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_1297_wire_constant <= "00000000000000000000000000000001";
    konst_1302_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_1290: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nR_1299_1292_buffered & T_1293_buffered;
      req <= phi_stmt_1290_req_0 & phi_stmt_1290_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1290",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1290_ack_0,
          idata => idata,
          odata => R_1290,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1290
    T_1293_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= T_1293_buf_req_0;
      T_1293_buf_ack_0<= wack(0);
      rreq(0) <= T_1293_buf_req_1;
      T_1293_buf_ack_1<= rack(0);
      T_1293_buf : InterlockBuffer generic map ( -- 
        name => "T_1293_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_1293_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nR_1299_1292_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_1299_1292_buf_req_0;
      nR_1299_1292_buf_ack_0<= wack(0);
      rreq(0) <= nR_1299_1292_buf_req_1;
      nR_1299_1292_buf_ack_1<= rack(0);
      nR_1299_1292_buf : InterlockBuffer generic map ( -- 
        name => "nR_1299_1292_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_1299,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_1299_1292_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1288_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u32_u1_1303_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1288_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1288_branch_req_0,
          ack0 => do_while_stmt_1288_branch_ack_0,
          ack1 => do_while_stmt_1288_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator SUB_u32_u32_1298_inst
    process(R_1290) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_1290, konst_1297_wire_constant, tmp_var);
      nR_1299 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1303_inst
    process(R_1290) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(R_1290, konst_1302_wire_constant, tmp_var);
      UGT_u32_u1_1303_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end delay_time_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    read_index : in  std_logic_vector(31 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueElement;
architecture getQueueElement_arch of getQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal read_index_buffer :  std_logic_vector(31 downto 0);
  signal read_index_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal getQueueElement_CP_626_start: Boolean;
  signal getQueueElement_CP_626_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_664_call_req_0 : boolean;
  signal call_stmt_664_call_ack_0 : boolean;
  signal call_stmt_664_call_req_1 : boolean;
  signal call_stmt_664_call_ack_1 : boolean;
  signal MUX_679_inst_req_0 : boolean;
  signal MUX_679_inst_ack_0 : boolean;
  signal MUX_679_inst_req_1 : boolean;
  signal MUX_679_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= read_index;
  read_index_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueElement_CP_626_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_626_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueElement_CP_626_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_626_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueElement_CP_626: Block -- control-path 
    signal getQueueElement_CP_626_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueElement_CP_626_elements(0) <= getQueueElement_CP_626_start;
    getQueueElement_CP_626_symbol <= getQueueElement_CP_626_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/$entry
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_sample_start_
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_update_start_
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Sample/crr
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Update/$entry
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Update/ccr
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_update_start_
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_complete/$entry
      -- CP-element group 0: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_complete/req
      -- 
    ccr_644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_626_elements(0), ack => call_stmt_664_call_req_1); -- 
    req_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_626_elements(0), ack => MUX_679_inst_req_1); -- 
    crr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_626_elements(0), ack => call_stmt_664_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_sample_completed_
      -- CP-element group 1: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Sample/cra
      -- 
    cra_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_664_call_ack_0, ack => getQueueElement_CP_626_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_update_completed_
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Update/$exit
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_680/call_stmt_664_Update/cca
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_sample_start_
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_start/$entry
      -- CP-element group 2: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_start/req
      -- 
    cca_645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_664_call_ack_1, ack => getQueueElement_CP_626_elements(2)); -- 
    req_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_626_elements(2), ack => MUX_679_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_sample_completed_
      -- CP-element group 3: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_start/$exit
      -- CP-element group 3: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_start/ack
      -- 
    ack_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_679_inst_ack_0, ack => getQueueElement_CP_626_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 assign_stmt_640_to_assign_stmt_680/$exit
      -- CP-element group 4: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_update_completed_
      -- CP-element group 4: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_complete/$exit
      -- CP-element group 4: 	 assign_stmt_640_to_assign_stmt_680/MUX_679_complete/ack
      -- 
    ack_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_679_inst_ack_1, ack => getQueueElement_CP_626_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_676_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_648_wire : std_logic_vector(33 downto 0);
    signal NOT_u8_u8_659_wire_constant : std_logic_vector(7 downto 0);
    signal buffer_address_640 : std_logic_vector(35 downto 0);
    signal e0_668 : std_logic_vector(31 downto 0);
    signal e1_672 : std_logic_vector(31 downto 0);
    signal element_pair_664 : std_logic_vector(63 downto 0);
    signal element_pair_address_652 : std_logic_vector(35 downto 0);
    signal konst_675_wire_constant : std_logic_vector(31 downto 0);
    signal slice_645_wire : std_logic_vector(30 downto 0);
    signal type_cast_638_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_650_wire : std_logic_vector(35 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_656_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_662_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_659_wire_constant <= "11111111";
    konst_675_wire_constant <= "00000000000000000000000000000000";
    type_cast_638_wire_constant <= "000000000000000000000000000000011000";
    type_cast_647_wire_constant <= "000";
    type_cast_654_wire_constant <= "0";
    type_cast_656_wire_constant <= "1";
    type_cast_662_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    MUX_679_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_679_inst_req_0;
      MUX_679_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_679_inst_req_1;
      MUX_679_inst_ack_1<= update_ack(0);
      MUX_679_inst: SelectSplitProtocol generic map(name => "MUX_679_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => e1_672, y => e0_668, sel => BITSEL_u32_u1_676_wire, z => q_r_data_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_645_inst
    slice_645_wire <= read_index_buffer(31 downto 1);
    -- flow-through slice operator slice_667_inst
    e0_668 <= element_pair_664(63 downto 32);
    -- flow-through slice operator slice_671_inst
    e1_672 <= element_pair_664(31 downto 0);
    -- interlock type_cast_650_inst
    process(CONCAT_u31_u34_648_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_648_wire(33 downto 0);
      type_cast_650_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_639_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_638_wire_constant, tmp_var);
      buffer_address_640 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_651_inst
    process(buffer_address_640, type_cast_650_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_640, type_cast_650_wire, tmp_var);
      element_pair_address_652 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_676_inst
    process(read_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(read_index_buffer, konst_675_wire_constant, tmp_var);
      BITSEL_u32_u1_676_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_648_inst
    process(slice_645_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_645_wire, type_cast_647_wire_constant, tmp_var);
      CONCAT_u31_u34_648_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_664_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_664_call_req_0;
      call_stmt_664_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_664_call_req_1;
      call_stmt_664_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_654_wire_constant & type_cast_656_wire_constant & NOT_u8_u8_659_wire_constant & element_pair_address_652 & type_cast_662_wire_constant;
      element_pair_664 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueueLength is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    Queue_Length : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueLength;
architecture getQueueLength_arch of getQueueLength is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal Queue_Length_buffer :  std_logic_vector(31 downto 0);
  signal Queue_Length_update_enable: Boolean;
  signal getQueueLength_CP_558_start: Boolean;
  signal getQueueLength_CP_558_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_605_call_req_0 : boolean;
  signal call_stmt_605_call_ack_0 : boolean;
  signal call_stmt_605_call_req_1 : boolean;
  signal call_stmt_605_call_ack_1 : boolean;
  signal slice_608_inst_req_0 : boolean;
  signal slice_608_inst_ack_0 : boolean;
  signal slice_608_inst_req_1 : boolean;
  signal slice_608_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueLength_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueLength_CP_558_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueLength_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= Queue_Length_buffer;
  Queue_Length <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_558_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueLength_CP_558_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_558_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueLength_CP_558: Block -- control-path 
    signal getQueueLength_CP_558_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueLength_CP_558_elements(0) <= getQueueLength_CP_558_start;
    getQueueLength_CP_558_symbol <= getQueueLength_CP_558_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/$entry
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_sample_start_
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_update_start_
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Sample/$entry
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Sample/crr
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Update/$entry
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Update/ccr
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/slice_608_update_start_
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/slice_608_Update/$entry
      -- CP-element group 0: 	 call_stmt_605_to_assign_stmt_609/slice_608_Update/cr
      -- 
    crr_571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_558_elements(0), ack => call_stmt_605_call_req_0); -- 
    ccr_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_558_elements(0), ack => call_stmt_605_call_req_1); -- 
    cr_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_558_elements(0), ack => slice_608_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_sample_completed_
      -- CP-element group 1: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Sample/$exit
      -- CP-element group 1: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Sample/cra
      -- 
    cra_572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_605_call_ack_0, ack => getQueueLength_CP_558_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_update_completed_
      -- CP-element group 2: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Update/$exit
      -- CP-element group 2: 	 call_stmt_605_to_assign_stmt_609/call_stmt_605_Update/cca
      -- CP-element group 2: 	 call_stmt_605_to_assign_stmt_609/slice_608_sample_start_
      -- CP-element group 2: 	 call_stmt_605_to_assign_stmt_609/slice_608_Sample/$entry
      -- CP-element group 2: 	 call_stmt_605_to_assign_stmt_609/slice_608_Sample/rr
      -- 
    cca_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_605_call_ack_1, ack => getQueueLength_CP_558_elements(2)); -- 
    rr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_558_elements(2), ack => slice_608_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_605_to_assign_stmt_609/slice_608_sample_completed_
      -- CP-element group 3: 	 call_stmt_605_to_assign_stmt_609/slice_608_Sample/$exit
      -- CP-element group 3: 	 call_stmt_605_to_assign_stmt_609/slice_608_Sample/ra
      -- 
    ra_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_608_inst_ack_0, ack => getQueueLength_CP_558_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_605_to_assign_stmt_609/$exit
      -- CP-element group 4: 	 call_stmt_605_to_assign_stmt_609/slice_608_update_completed_
      -- CP-element group 4: 	 call_stmt_605_to_assign_stmt_609/slice_608_Update/$exit
      -- CP-element group 4: 	 call_stmt_605_to_assign_stmt_609/slice_608_Update/ca
      -- 
    ca_591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_608_inst_ack_1, ack => getQueueLength_CP_558_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_601_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_598_wire_constant : std_logic_vector(7 downto 0);
    signal konst_600_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_593_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_595_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_603_wire_constant : std_logic_vector(63 downto 0);
    signal wi_and_len_605 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_598_wire_constant <= "11111111";
    konst_600_wire_constant <= "000000000000000000000000000000001000";
    type_cast_593_wire_constant <= "0";
    type_cast_595_wire_constant <= "1";
    type_cast_603_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    slice_608_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_608_inst_req_0;
      slice_608_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_608_inst_req_1;
      slice_608_inst_ack_1<= update_ack(0);
      slice_608_inst: SliceSplitProtocol generic map(name => "slice_608_inst", in_data_width => 64, high_index => 31, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => wi_and_len_605, dout => Queue_Length_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- binary operator ADD_u36_u36_601_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_600_wire_constant, tmp_var);
      ADD_u36_u36_601_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_605_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_605_call_req_0;
      call_stmt_605_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_605_call_req_1;
      call_stmt_605_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_593_wire_constant & type_cast_595_wire_constant & NOT_u8_u8_598_wire_constant & ADD_u36_u36_601_wire & type_cast_603_wire_constant;
      wi_and_len_605 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueLength_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : out  std_logic_vector(31 downto 0);
    rp : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointers;
architecture getQueuePointers_arch of getQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  signal getQueuePointers_CP_524_start: Boolean;
  signal getQueuePointers_CP_524_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_575_call_req_0 : boolean;
  signal call_stmt_575_call_ack_0 : boolean;
  signal call_stmt_575_call_req_1 : boolean;
  signal call_stmt_575_call_ack_1 : boolean;
  signal call_stmt_561_call_req_0 : boolean;
  signal call_stmt_561_call_ack_0 : boolean;
  signal call_stmt_561_call_req_1 : boolean;
  signal call_stmt_561_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointers_CP_524_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wp_buffer;
  wp <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= rp_buffer;
  rp <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_524_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointers_CP_524_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_524_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointers_CP_524: Block -- control-path 
    signal getQueuePointers_CP_524_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueuePointers_CP_524_elements(0) <= getQueuePointers_CP_524_start;
    getQueuePointers_CP_524_symbol <= getQueuePointers_CP_524_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Update/$entry
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Update/ccr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Sample/$entry
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Sample/crr
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Update/$entry
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_update_start_
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/$entry
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_sample_start_
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Update/ccr
      -- CP-element group 0: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_update_start_
      -- 
    crr_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_524_elements(0), ack => call_stmt_561_call_req_0); -- 
    ccr_542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_524_elements(0), ack => call_stmt_561_call_req_1); -- 
    ccr_556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_524_elements(0), ack => call_stmt_575_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Sample/$exit
      -- CP-element group 1: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Sample/cra
      -- CP-element group 1: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_sample_completed_
      -- 
    cra_538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_561_call_ack_0, ack => getQueuePointers_CP_524_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Sample/$entry
      -- CP-element group 2: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Sample/crr
      -- CP-element group 2: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Update/$exit
      -- CP-element group 2: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_update_completed_
      -- CP-element group 2: 	 call_stmt_561_to_assign_stmt_583/call_stmt_561_Update/cca
      -- CP-element group 2: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_sample_start_
      -- 
    cca_543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_561_call_ack_1, ack => getQueuePointers_CP_524_elements(2)); -- 
    crr_551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_524_elements(2), ack => call_stmt_575_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Sample/$exit
      -- CP-element group 3: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Sample/cra
      -- CP-element group 3: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_sample_completed_
      -- 
    cra_552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_575_call_ack_0, ack => getQueuePointers_CP_524_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Update/$exit
      -- CP-element group 4: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_Update/cca
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_561_to_assign_stmt_583/$exit
      -- CP-element group 4: 	 call_stmt_561_to_assign_stmt_583/call_stmt_575_update_completed_
      -- 
    cca_557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_575_call_ack_1, ack => getQueuePointers_CP_524_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_571_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_556_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_568_wire_constant : std_logic_vector(7 downto 0);
    signal konst_570_wire_constant : std_logic_vector(35 downto 0);
    signal msgs_rp_561 : std_logic_vector(63 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_559_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_563_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_565_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_573_wire_constant : std_logic_vector(63 downto 0);
    signal wp_len_575 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_556_wire_constant <= "11111111";
    NOT_u8_u8_568_wire_constant <= "11111111";
    konst_570_wire_constant <= "000000000000000000000000000000001000";
    type_cast_551_wire_constant <= "0";
    type_cast_553_wire_constant <= "1";
    type_cast_559_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_563_wire_constant <= "0";
    type_cast_565_wire_constant <= "1";
    type_cast_573_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through slice operator slice_578_inst
    rp_buffer <= msgs_rp_561(31 downto 0);
    -- flow-through slice operator slice_582_inst
    wp_buffer <= wp_len_575(63 downto 32);
    -- binary operator ADD_u36_u36_571_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_570_wire_constant, tmp_var);
      ADD_u36_u36_571_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_561_call call_stmt_575_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_561_call_req_0;
      reqL_unguarded(0) <= call_stmt_575_call_req_0;
      call_stmt_561_call_ack_0 <= ackL_unguarded(1);
      call_stmt_575_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_561_call_req_1;
      reqR_unguarded(0) <= call_stmt_575_call_req_1;
      call_stmt_561_call_ack_1 <= ackR_unguarded(1);
      call_stmt_575_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_551_wire_constant & type_cast_553_wire_constant & NOT_u8_u8_556_wire_constant & q_base_address_buffer & type_cast_559_wire_constant & type_cast_563_wire_constant & type_cast_565_wire_constant & NOT_u8_u8_568_wire_constant & ADD_u36_u36_571_wire & type_cast_573_wire_constant;
      msgs_rp_561 <= data_out(127 downto 64);
      wp_len_575 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    total_msgs : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTotalMessages;
architecture getTotalMessages_arch of getTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal total_msgs_update_enable: Boolean;
  signal getTotalMessages_CP_592_start: Boolean;
  signal getTotalMessages_CP_592_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_625_call_req_0 : boolean;
  signal call_stmt_625_call_ack_0 : boolean;
  signal call_stmt_625_call_req_1 : boolean;
  signal call_stmt_625_call_ack_1 : boolean;
  signal slice_628_inst_req_0 : boolean;
  signal slice_628_inst_ack_0 : boolean;
  signal slice_628_inst_req_1 : boolean;
  signal slice_628_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTotalMessages_CP_592_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= total_msgs_buffer;
  total_msgs <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_592_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTotalMessages_CP_592_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_592_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTotalMessages_CP_592: Block -- control-path 
    signal getTotalMessages_CP_592_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getTotalMessages_CP_592_elements(0) <= getTotalMessages_CP_592_start;
    getTotalMessages_CP_592_symbol <= getTotalMessages_CP_592_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/$entry
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_sample_start_
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_update_start_
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Sample/$entry
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Sample/crr
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Update/$entry
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Update/ccr
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/slice_628_update_start_
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/slice_628_Update/$entry
      -- CP-element group 0: 	 call_stmt_625_to_assign_stmt_629/slice_628_Update/cr
      -- 
    crr_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_592_elements(0), ack => call_stmt_625_call_req_0); -- 
    ccr_610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_592_elements(0), ack => call_stmt_625_call_req_1); -- 
    cr_624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_592_elements(0), ack => slice_628_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_sample_completed_
      -- CP-element group 1: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Sample/$exit
      -- CP-element group 1: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Sample/cra
      -- 
    cra_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_625_call_ack_0, ack => getTotalMessages_CP_592_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_update_completed_
      -- CP-element group 2: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Update/$exit
      -- CP-element group 2: 	 call_stmt_625_to_assign_stmt_629/call_stmt_625_Update/cca
      -- CP-element group 2: 	 call_stmt_625_to_assign_stmt_629/slice_628_sample_start_
      -- CP-element group 2: 	 call_stmt_625_to_assign_stmt_629/slice_628_Sample/$entry
      -- CP-element group 2: 	 call_stmt_625_to_assign_stmt_629/slice_628_Sample/rr
      -- 
    cca_611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_625_call_ack_1, ack => getTotalMessages_CP_592_elements(2)); -- 
    rr_619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_592_elements(2), ack => slice_628_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_625_to_assign_stmt_629/slice_628_sample_completed_
      -- CP-element group 3: 	 call_stmt_625_to_assign_stmt_629/slice_628_Sample/$exit
      -- CP-element group 3: 	 call_stmt_625_to_assign_stmt_629/slice_628_Sample/ra
      -- 
    ra_620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_628_inst_ack_0, ack => getTotalMessages_CP_592_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_625_to_assign_stmt_629/$exit
      -- CP-element group 4: 	 call_stmt_625_to_assign_stmt_629/slice_628_update_completed_
      -- CP-element group 4: 	 call_stmt_625_to_assign_stmt_629/slice_628_Update/$exit
      -- CP-element group 4: 	 call_stmt_625_to_assign_stmt_629/slice_628_Update/ca
      -- 
    ca_625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_628_inst_ack_1, ack => getTotalMessages_CP_592_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u8_u8_620_wire_constant : std_logic_vector(7 downto 0);
    signal rdata_625 : std_logic_vector(63 downto 0);
    signal type_cast_615_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_617_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_623_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_620_wire_constant <= "11111111";
    type_cast_615_wire_constant <= "0";
    type_cast_617_wire_constant <= "1";
    type_cast_623_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    slice_628_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_628_inst_req_0;
      slice_628_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_628_inst_req_1;
      slice_628_inst_ack_1<= update_ack(0);
      slice_628_inst: SliceSplitProtocol generic map(name => "slice_628_inst", in_data_width => 64, high_index => 63, low_index => 32, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdata_625, dout => total_msgs_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- shared call operator group (0) : call_stmt_625_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_625_call_req_0;
      call_stmt_625_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_625_call_req_1;
      call_stmt_625_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_615_wire_constant & type_cast_617_wire_constant & NOT_u8_u8_620_wire_constant & q_base_address_buffer & type_cast_623_wire_constant;
      rdata_625 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getTxPacketPointerFromServer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_index : in  std_logic_vector(5 downto 0);
    pkt_pointer : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTxPacketPointerFromServer;
architecture getTxPacketPointerFromServer_arch of getTxPacketPointerFromServer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 6)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_index_buffer :  std_logic_vector(5 downto 0);
  signal queue_index_update_enable: Boolean;
  -- output port buffer signals
  signal pkt_pointer_buffer :  std_logic_vector(31 downto 0);
  signal pkt_pointer_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal getTxPacketPointerFromServer_CP_2819_start: Boolean;
  signal getTxPacketPointerFromServer_CP_2819_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1742_call_req_1 : boolean;
  signal call_stmt_1742_call_ack_0 : boolean;
  signal call_stmt_1742_call_ack_1 : boolean;
  signal call_stmt_1730_call_req_0 : boolean;
  signal call_stmt_1730_call_ack_0 : boolean;
  signal call_stmt_1730_call_ack_1 : boolean;
  signal call_stmt_1730_call_req_1 : boolean;
  signal call_stmt_1742_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 6) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= queue_index;
  queue_index_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(tag_length + 5 downto 6) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 5 downto 6);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 7);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= queue_index_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTxPacketPointerFromServer_CP_2819_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= pkt_pointer_buffer;
  pkt_pointer <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2819_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  pkt_pointer_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "pkt_pointer_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_pkt_pointer_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => pkt_pointer_update_enable, clk => clk, reset => reset); --
  end block;
  status_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "status_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_status_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => status_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2819_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2819_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTxPacketPointerFromServer_CP_2819: Block -- control-path 
    signal getTxPacketPointerFromServer_CP_2819_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    getTxPacketPointerFromServer_CP_2819_elements(0) <= getTxPacketPointerFromServer_CP_2819_start;
    getTxPacketPointerFromServer_CP_2819_symbol <= getTxPacketPointerFromServer_CP_2819_elements(16);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_1720_to_stmt_1747/$entry
      -- 
    getTxPacketPointerFromServer_CP_2819_elements(1) <= getTxPacketPointerFromServer_CP_2819_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_1720_to_stmt_1747/queue_index_update_enable_out
      -- CP-element group 2: 	 assign_stmt_1720_to_stmt_1747/queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_2819_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2819_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	14 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_1720_to_stmt_1747/pkt_pointer_update_enable
      -- CP-element group 3: 	 assign_stmt_1720_to_stmt_1747/pkt_pointer_update_enable_in
      -- 
    getTxPacketPointerFromServer_CP_2819_elements(3) <= getTxPacketPointerFromServer_CP_2819_elements(14);
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_1720_to_stmt_1747/status_update_enable
      -- CP-element group 4: 	 assign_stmt_1720_to_stmt_1747/status_update_enable_in
      -- 
    getTxPacketPointerFromServer_CP_2819_elements(4) <= getTxPacketPointerFromServer_CP_2819_elements(15);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_sample_start_
      -- CP-element group 5: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Sample/crr
      -- 
    crr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2819_elements(5), ack => call_stmt_1730_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2819_elements(1) & getTxPacketPointerFromServer_CP_2819_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2819_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_update_start_
      -- CP-element group 6: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Update/ccr
      -- CP-element group 6: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Update/$entry
      -- 
    ccr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2819_elements(6), ack => call_stmt_1730_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2819_elements(8) & getTxPacketPointerFromServer_CP_2819_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2819_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_sample_completed_
      -- CP-element group 7: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Sample/cra
      -- 
    cra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1730_call_ack_0, ack => getTxPacketPointerFromServer_CP_2819_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_update_completed_
      -- CP-element group 8: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Update/cca
      -- CP-element group 8: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1730_Update/$exit
      -- 
    cca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1730_call_ack_1, ack => getTxPacketPointerFromServer_CP_2819_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_sample_start_
      -- CP-element group 9: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Sample/crr
      -- 
    crr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2819_elements(9), ack => call_stmt_1742_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2819_elements(8) & getTxPacketPointerFromServer_CP_2819_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2819_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Update/$entry
      -- CP-element group 10: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_update_start_
      -- CP-element group 10: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Update/ccr
      -- 
    ccr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2819_elements(10), ack => call_stmt_1742_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "getTxPacketPointerFromServer_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2819_elements(3) & getTxPacketPointerFromServer_CP_2819_elements(4) & getTxPacketPointerFromServer_CP_2819_elements(12);
      gj_getTxPacketPointerFromServer_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2819_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_sample_completed_
      -- CP-element group 11: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Sample/cra
      -- CP-element group 11: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Sample/$exit
      -- 
    cra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1742_call_ack_0, ack => getTxPacketPointerFromServer_CP_2819_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Update/$exit
      -- CP-element group 12: 	 assign_stmt_1720_to_stmt_1747/$exit
      -- CP-element group 12: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_Update/cca
      -- CP-element group 12: 	 assign_stmt_1720_to_stmt_1747/call_stmt_1742_update_completed_
      -- 
    cca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1742_call_ack_1, ack => getTxPacketPointerFromServer_CP_2819_elements(12)); -- 
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_CP_2819_elements(13) <= getTxPacketPointerFromServer_CP_2819_elements(2);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 pkt_pointer_update_enable
      -- 
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 status_update_enable
      -- 
    -- CP-element group 16:  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 $exit
      -- 
    getTxPacketPointerFromServer_CP_2819_elements(16) <= getTxPacketPointerFromServer_CP_2819_elements(12);
    --  hookup: inputs to control-path 
    getTxPacketPointerFromServer_CP_2819_elements(14) <= pkt_pointer_update_enable;
    getTxPacketPointerFromServer_CP_2819_elements(15) <= status_update_enable;
    -- hookup: output from control-path 
    queue_index_update_enable <= getTxPacketPointerFromServer_CP_2819_elements(13);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1718_wire : std_logic_vector(5 downto 0);
    signal NOT_u4_u4_1725_wire_constant : std_logic_vector(3 downto 0);
    signal R_TX_QUEUES_REG_START_OFFSET_1717_wire_constant : std_logic_vector(5 downto 0);
    signal register_index_1720 : std_logic_vector(5 downto 0);
    signal tx_queue_pointer_32_1730 : std_logic_vector(31 downto 0);
    signal tx_queue_pointer_36_1736 : std_logic_vector(35 downto 0);
    signal type_cast_1722_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1728_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1733_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1738_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1725_wire_constant <= "1111";
    R_TX_QUEUES_REG_START_OFFSET_1717_wire_constant <= "001010";
    type_cast_1722_wire_constant <= "1";
    type_cast_1728_wire_constant <= "00000000000000000000000000000000";
    type_cast_1733_wire_constant <= "0000";
    type_cast_1738_wire_constant <= "1";
    -- interlock type_cast_1719_inst
    process(ADD_u6_u6_1718_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1718_wire(5 downto 0);
      register_index_1720 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u6_u6_1718_inst
    process(queue_index_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(queue_index_buffer, R_TX_QUEUES_REG_START_OFFSET_1717_wire_constant, tmp_var);
      ADD_u6_u6_1718_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_1735_inst
    process(type_cast_1733_wire_constant, tx_queue_pointer_32_1730) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1733_wire_constant, tx_queue_pointer_32_1730, tmp_var);
      tx_queue_pointer_36_1736 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1730_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1730_call_req_0;
      call_stmt_1730_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1730_call_req_1;
      call_stmt_1730_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1722_wire_constant & NOT_u4_u4_1725_wire_constant & register_index_1720 & type_cast_1728_wire_constant;
      tx_queue_pointer_32_1730 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1742_call 
    popFromQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1742_call_req_0;
      call_stmt_1742_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1742_call_req_1;
      call_stmt_1742_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_1_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1738_wire_constant & tx_queue_pointer_36_1736;
      pkt_pointer_buffer <= data_out(32 downto 1);
      status_buffer <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getTxPacketPointerFromServer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity loadBuffer is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
    writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
    writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
    writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadBuffer;
architecture loadBuffer_arch of loadBuffer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal loadBuffer_CP_1205_start: Boolean;
  signal loadBuffer_CP_1205_symbol: Boolean;
  -- volatile/operator module components. 
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1120_call_ack_1 : boolean;
  signal W_bad_packet_identifier_1136_delayed_8_0_1130_inst_ack_0 : boolean;
  signal call_stmt_1120_call_req_1 : boolean;
  signal W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_ack_0 : boolean;
  signal W_bad_packet_identifier_1136_delayed_8_0_1130_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_req_0 : boolean;
  signal W_bad_packet_identifier_1136_delayed_8_0_1130_inst_req_1 : boolean;
  signal call_stmt_1129_call_req_0 : boolean;
  signal call_stmt_1120_call_ack_0 : boolean;
  signal W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_req_1 : boolean;
  signal call_stmt_1129_call_ack_0 : boolean;
  signal call_stmt_1120_call_req_0 : boolean;
  signal call_stmt_1140_call_req_1 : boolean;
  signal call_stmt_1140_call_req_0 : boolean;
  signal call_stmt_1140_call_ack_0 : boolean;
  signal call_stmt_1129_call_ack_1 : boolean;
  signal call_stmt_1129_call_req_1 : boolean;
  signal W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_req_0 : boolean;
  signal W_bad_packet_identifier_1136_delayed_8_0_1130_inst_req_0 : boolean;
  signal call_stmt_1140_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadBuffer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 31);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_buffer_pointer_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadBuffer_CP_1205_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadBuffer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1205_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  bad_packet_identifier_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 40) := "bad_packet_identifier_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_bad_packet_identifier_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => bad_packet_identifier_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 31,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadBuffer_CP_1205_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1205_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadBuffer_CP_1205: Block -- control-path 
    signal loadBuffer_CP_1205_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    loadBuffer_CP_1205_elements(0) <= loadBuffer_CP_1205_start;
    loadBuffer_CP_1205_symbol <= loadBuffer_CP_1205_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	20 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_1120_to_call_stmt_1140/$entry
      -- 
    loadBuffer_CP_1205_elements(1) <= loadBuffer_CP_1205_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	6 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	28 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_1120_to_call_stmt_1140/rx_buffer_pointer_update_enable
      -- CP-element group 2: 	 call_stmt_1120_to_call_stmt_1140/rx_buffer_pointer_update_enable_out
      -- 
    loadBuffer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(22) & loadBuffer_CP_1205_elements(10) & loadBuffer_CP_1205_elements(6);
      gj_loadBuffer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	29 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_1120_to_call_stmt_1140/bad_packet_identifier_update_enable_in
      -- CP-element group 3: 	 call_stmt_1120_to_call_stmt_1140/bad_packet_identifier_update_enable
      -- 
    loadBuffer_CP_1205_elements(3) <= loadBuffer_CP_1205_elements(29);
    -- CP-element group 4:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	27 
    -- CP-element group 4: 	6 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_sample_start_
      -- CP-element group 4: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Sample/crr
      -- CP-element group 4: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Sample/$entry
      -- 
    crr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(4), ack => call_stmt_1120_call_req_0); -- 
    loadBuffer_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(1) & loadBuffer_CP_1205_elements(27) & loadBuffer_CP_1205_elements(6);
      gj_loadBuffer_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	27 
    -- CP-element group 5: 	7 
    -- CP-element group 5: 	14 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_update_start_
      -- CP-element group 5: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Update/$entry
      -- CP-element group 5: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Update/ccr
      -- 
    ccr_1227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(5), ack => call_stmt_1120_call_req_1); -- 
    loadBuffer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(27) & loadBuffer_CP_1205_elements(7) & loadBuffer_CP_1205_elements(14);
      gj_loadBuffer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: marked-successors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: 	4 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_sample_completed_
      -- CP-element group 6: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Sample/cra
      -- CP-element group 6: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Sample/$exit
      -- 
    cra_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1120_call_ack_0, ack => loadBuffer_CP_1205_elements(6)); -- 
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Update/cca
      -- CP-element group 7: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_Update/$exit
      -- CP-element group 7: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1120_update_completed_
      -- 
    cca_1228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1120_call_ack_1, ack => loadBuffer_CP_1205_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_sample_start_
      -- CP-element group 8: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Sample/req
      -- 
    req_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(8), ack => W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_req_0); -- 
    loadBuffer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(1) & loadBuffer_CP_1205_elements(10);
      gj_loadBuffer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_update_start_
      -- CP-element group 9: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Update/req
      -- CP-element group 9: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Update/$entry
      -- 
    req_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(9), ack => W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_req_1); -- 
    loadBuffer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(11) & loadBuffer_CP_1205_elements(14);
      gj_loadBuffer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: 	2 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_sample_completed_
      -- CP-element group 10: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Sample/ack
      -- CP-element group 10: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Sample/$exit
      -- 
    ack_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_ack_0, ack => loadBuffer_CP_1205_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_update_completed_
      -- CP-element group 11: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Update/ack
      -- CP-element group 11: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1123_Update/$exit
      -- 
    ack_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_ack_1, ack => loadBuffer_CP_1205_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_sample_start_
      -- CP-element group 12: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Sample/crr
      -- CP-element group 12: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Sample/$entry
      -- 
    crr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(12), ack => call_stmt_1129_call_req_0); -- 
    loadBuffer_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(7) & loadBuffer_CP_1205_elements(11) & loadBuffer_CP_1205_elements(14);
      gj_loadBuffer_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	26 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Update/ccr
      -- CP-element group 13: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Update/$entry
      -- CP-element group 13: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_update_start_
      -- 
    ccr_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(13), ack => call_stmt_1129_call_req_1); -- 
    loadBuffer_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(3) & loadBuffer_CP_1205_elements(15) & loadBuffer_CP_1205_elements(18) & loadBuffer_CP_1205_elements(26);
      gj_loadBuffer_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	5 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_sample_completed_
      -- CP-element group 14: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Sample/$exit
      -- CP-element group 14: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Sample/cra
      -- 
    cra_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1129_call_ack_0, ack => loadBuffer_CP_1205_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	24 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Update/cca
      -- CP-element group 15: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_Update/$exit
      -- CP-element group 15: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1129_update_completed_
      -- 
    cca_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1129_call_ack_1, ack => loadBuffer_CP_1205_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Sample/$entry
      -- CP-element group 16: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_sample_start_
      -- CP-element group 16: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Sample/req
      -- 
    req_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(16), ack => W_bad_packet_identifier_1136_delayed_8_0_1130_inst_req_0); -- 
    loadBuffer_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(15) & loadBuffer_CP_1205_elements(18);
      gj_loadBuffer_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	26 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Update/$entry
      -- CP-element group 17: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_update_start_
      -- CP-element group 17: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Update/req
      -- 
    req_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(17), ack => W_bad_packet_identifier_1136_delayed_8_0_1130_inst_req_1); -- 
    loadBuffer_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(19) & loadBuffer_CP_1205_elements(26);
      gj_loadBuffer_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	13 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Sample/ack
      -- CP-element group 18: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Sample/$exit
      -- CP-element group 18: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_sample_completed_
      -- 
    ack_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1136_delayed_8_0_1130_inst_ack_0, ack => loadBuffer_CP_1205_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Update/$exit
      -- CP-element group 19: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_Update/ack
      -- CP-element group 19: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1132_update_completed_
      -- 
    ack_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1136_delayed_8_0_1130_inst_ack_1, ack => loadBuffer_CP_1205_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	1 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_sample_start_
      -- CP-element group 20: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Sample/req
      -- CP-element group 20: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Sample/$entry
      -- 
    req_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(20), ack => W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_req_0); -- 
    loadBuffer_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(1) & loadBuffer_CP_1205_elements(22);
      gj_loadBuffer_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	26 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Update/req
      -- CP-element group 21: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Update/$entry
      -- CP-element group 21: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_update_start_
      -- 
    req_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(21), ack => W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_req_1); -- 
    loadBuffer_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(23) & loadBuffer_CP_1205_elements(26);
      gj_loadBuffer_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	2 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Sample/ack
      -- CP-element group 22: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_sample_completed_
      -- CP-element group 22: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Sample/$exit
      -- 
    ack_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_ack_0, ack => loadBuffer_CP_1205_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Update/$exit
      -- CP-element group 23: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_update_completed_
      -- CP-element group 23: 	 call_stmt_1120_to_call_stmt_1140/assign_stmt_1135_Update/ack
      -- 
    ack_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_ack_1, ack => loadBuffer_CP_1205_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_sample_start_
      -- CP-element group 24: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Sample/crr
      -- CP-element group 24: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Sample/$entry
      -- 
    crr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(24), ack => call_stmt_1140_call_req_0); -- 
    loadBuffer_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1205_elements(15) & loadBuffer_CP_1205_elements(19) & loadBuffer_CP_1205_elements(23) & loadBuffer_CP_1205_elements(26);
      gj_loadBuffer_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_update_start_
      -- CP-element group 25: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Update/ccr
      -- CP-element group 25: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Update/$entry
      -- 
    ccr_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1205_elements(25), ack => call_stmt_1140_call_req_1); -- 
    loadBuffer_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadBuffer_CP_1205_elements(27);
      gj_loadBuffer_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1205_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	17 
    -- CP-element group 26: 	21 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	13 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_sample_completed_
      -- CP-element group 26: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Sample/cra
      -- CP-element group 26: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Sample/$exit
      -- 
    cra_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1140_call_ack_0, ack => loadBuffer_CP_1205_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: 	4 
    -- CP-element group 27: 	5 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_update_completed_
      -- CP-element group 27: 	 call_stmt_1120_to_call_stmt_1140/$exit
      -- CP-element group 27: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Update/$exit
      -- CP-element group 27: 	 call_stmt_1120_to_call_stmt_1140/call_stmt_1140_Update/cca
      -- 
    cca_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1140_call_ack_1, ack => loadBuffer_CP_1205_elements(27)); -- 
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 rx_buffer_pointer_update_enable
      -- 
    loadBuffer_CP_1205_elements(28) <= loadBuffer_CP_1205_elements(2);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	3 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 bad_packet_identifier_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    loadBuffer_CP_1205_elements(30) <= loadBuffer_CP_1205_elements(27);
    --  hookup: inputs to control-path 
    loadBuffer_CP_1205_elements(29) <= bad_packet_identifier_update_enable;
    -- hookup: output from control-path 
    rx_buffer_pointer_update_enable <= loadBuffer_CP_1205_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal bad_packet_identifier_1136_delayed_8_0_1132 : std_logic_vector(0 downto 0);
    signal last_keep_1129 : std_logic_vector(7 downto 0);
    signal new_buf_pointer_1120 : std_logic_vector(35 downto 0);
    signal packet_size_1129 : std_logic_vector(7 downto 0);
    signal rx_buffer_pointer_1130_delayed_4_0_1123 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_1137_delayed_8_0_1135 : std_logic_vector(35 downto 0);
    -- 
  begin -- 
    W_bad_packet_identifier_1136_delayed_8_0_1130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bad_packet_identifier_1136_delayed_8_0_1130_inst_req_0;
      W_bad_packet_identifier_1136_delayed_8_0_1130_inst_ack_0<= wack(0);
      rreq(0) <= W_bad_packet_identifier_1136_delayed_8_0_1130_inst_req_1;
      W_bad_packet_identifier_1136_delayed_8_0_1130_inst_ack_1<= rack(0);
      W_bad_packet_identifier_1136_delayed_8_0_1130_inst : InterlockBuffer generic map ( -- 
        name => "W_bad_packet_identifier_1136_delayed_8_0_1130_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bad_packet_identifier_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bad_packet_identifier_1136_delayed_8_0_1132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_req_0;
      W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_req_1;
      W_rx_buffer_pointer_1130_delayed_4_0_1121_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1130_delayed_4_0_1121_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1130_delayed_4_0_1121_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1130_delayed_4_0_1123,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_req_0;
      W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_req_1;
      W_rx_buffer_pointer_1137_delayed_8_0_1133_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1137_delayed_8_0_1133_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1137_delayed_8_0_1133_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1137_delayed_8_0_1135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared call operator group (0) : call_stmt_1120_call 
    writeEthernetHeaderToMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1120_call_req_0;
      call_stmt_1120_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1120_call_req_1;
      call_stmt_1120_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeEthernetHeaderToMem_call_group_0_gI: SplitGuardInterface generic map(name => "writeEthernetHeaderToMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer;
      new_buf_pointer_1120 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeEthernetHeaderToMem_call_reqs(0),
          ackR => writeEthernetHeaderToMem_call_acks(0),
          dataR => writeEthernetHeaderToMem_call_data(35 downto 0),
          tagR => writeEthernetHeaderToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeEthernetHeaderToMem_return_acks(0), -- cross-over
          ackL => writeEthernetHeaderToMem_return_reqs(0), -- cross-over
          dataL => writeEthernetHeaderToMem_return_data(35 downto 0),
          tagL => writeEthernetHeaderToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1129_call 
    writePayloadToMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(16 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1129_call_req_0;
      call_stmt_1129_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1129_call_req_1;
      call_stmt_1129_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writePayloadToMem_call_group_1_gI: SplitGuardInterface generic map(name => "writePayloadToMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_1130_delayed_4_0_1123 & new_buf_pointer_1120;
      packet_size_1129 <= data_out(16 downto 9);
      bad_packet_identifier_buffer <= data_out(8 downto 8);
      last_keep_1129 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writePayloadToMem_call_reqs(0),
          ackR => writePayloadToMem_call_acks(0),
          dataR => writePayloadToMem_call_data(71 downto 0),
          tagR => writePayloadToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 17,
          owidth => 17,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writePayloadToMem_return_acks(0), -- cross-over
          ackL => writePayloadToMem_return_reqs(0), -- cross-over
          dataL => writePayloadToMem_return_data(16 downto 0),
          tagL => writePayloadToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1140_call 
    writeControlInformationToMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(51 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1140_call_req_0;
      call_stmt_1140_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1140_call_req_1;
      call_stmt_1140_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not bad_packet_identifier_1136_delayed_8_0_1132(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeControlInformationToMem_call_group_2_gI: SplitGuardInterface generic map(name => "writeControlInformationToMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_1137_delayed_8_0_1135 & packet_size_1129 & last_keep_1129;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 52,
        owidth => 52,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeControlInformationToMem_call_reqs(0),
          ackR => writeControlInformationToMem_call_acks(0),
          dataR => writeControlInformationToMem_call_data(51 downto 0),
          tagR => writeControlInformationToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeControlInformationToMem_return_acks(0), -- cross-over
          ackL => writeControlInformationToMem_return_reqs(0), -- cross-over
          tagL => writeControlInformationToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end loadBuffer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nextLSTATE_Volatile is -- 
  port ( -- 
    RX : in  std_logic_vector(72 downto 0);
    LSTATE : in  std_logic_vector(1 downto 0);
    nLSTATE : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity nextLSTATE_Volatile;
architecture nextLSTATE_Volatile_arch of nextLSTATE_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal RX_buffer :  std_logic_vector(72 downto 0);
  signal LSTATE_buffer :  std_logic_vector(1 downto 0);
  -- output port buffer signals
  signal nLSTATE_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  RX_buffer <= RX;
  LSTATE_buffer <= LSTATE;
  -- output handling  -------------------------------------------------------
  nLSTATE <= nLSTATE_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1784_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1792_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1768_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1774_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1781_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1790_wire : std_logic_vector(0 downto 0);
    signal MUX_1771_wire : std_logic_vector(1 downto 0);
    signal MUX_1777_wire : std_logic_vector(1 downto 0);
    signal MUX_1787_wire : std_logic_vector(1 downto 0);
    signal MUX_1795_wire : std_logic_vector(1 downto 0);
    signal NOT_u1_u1_1783_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_1778_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_1796_wire : std_logic_vector(1 downto 0);
    signal R_S0_1767_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1793_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1769_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1773_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1775_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1780_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1785_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1789_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1762_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1770_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1776_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1786_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1794_wire_constant : std_logic_vector(1 downto 0);
    signal last_word_1764 : std_logic_vector(0 downto 0);
    signal tlast_1759 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_S0_1767_wire_constant <= "00";
    R_S0_1793_wire_constant <= "00";
    R_S1_1769_wire_constant <= "01";
    R_S1_1773_wire_constant <= "01";
    R_S2_1775_wire_constant <= "10";
    R_S2_1780_wire_constant <= "10";
    R_S2_1785_wire_constant <= "10";
    R_S2_1789_wire_constant <= "10";
    konst_1762_wire_constant <= "1";
    konst_1770_wire_constant <= "00";
    konst_1776_wire_constant <= "00";
    konst_1786_wire_constant <= "00";
    konst_1794_wire_constant <= "00";
    -- flow-through select operator MUX_1771_inst
    MUX_1771_wire <= R_S1_1769_wire_constant when (EQ_u2_u1_1768_wire(0) /=  '0') else konst_1770_wire_constant;
    -- flow-through select operator MUX_1777_inst
    MUX_1777_wire <= R_S2_1775_wire_constant when (EQ_u2_u1_1774_wire(0) /=  '0') else konst_1776_wire_constant;
    -- flow-through select operator MUX_1787_inst
    MUX_1787_wire <= R_S2_1785_wire_constant when (AND_u1_u1_1784_wire(0) /=  '0') else konst_1786_wire_constant;
    -- flow-through select operator MUX_1795_inst
    MUX_1795_wire <= R_S0_1793_wire_constant when (AND_u1_u1_1792_wire(0) /=  '0') else konst_1794_wire_constant;
    -- flow-through slice operator slice_1758_inst
    tlast_1759 <= RX_buffer(72 downto 72);
    -- binary operator AND_u1_u1_1784_inst
    process(EQ_u2_u1_1781_wire, NOT_u1_u1_1783_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1781_wire, NOT_u1_u1_1783_wire, tmp_var);
      AND_u1_u1_1784_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1792_inst
    process(EQ_u2_u1_1790_wire, last_word_1764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1790_wire, last_word_1764, tmp_var);
      AND_u1_u1_1792_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1763_inst
    process(tlast_1759) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tlast_1759, konst_1762_wire_constant, tmp_var);
      last_word_1764 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1768_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S0_1767_wire_constant, tmp_var);
      EQ_u2_u1_1768_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1774_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S1_1773_wire_constant, tmp_var);
      EQ_u2_u1_1774_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1781_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1780_wire_constant, tmp_var);
      EQ_u2_u1_1781_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1790_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1789_wire_constant, tmp_var);
      EQ_u2_u1_1790_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1783_inst
    process(last_word_1764) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_word_1764, tmp_var);
      NOT_u1_u1_1783_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u2_u2_1778_inst
    process(MUX_1771_wire, MUX_1777_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1771_wire, MUX_1777_wire, tmp_var);
      OR_u2_u2_1778_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1796_inst
    process(MUX_1787_wire, MUX_1795_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1787_wire, MUX_1795_wire, tmp_var);
      OR_u2_u2_1796_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1797_inst
    process(OR_u2_u2_1778_wire, OR_u2_u2_1796_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_1778_wire, OR_u2_u2_1796_wire, tmp_var);
      nLSTATE_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end nextLSTATE_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nicRxFromMacDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
    nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(1 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(1 downto 0);
    AccessRegister_call_data : out  std_logic_vector(85 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(1 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(1 downto 0);
    AccessRegister_return_data : in   std_logic_vector(63 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicRxFromMacDaemon;
architecture nicRxFromMacDaemon_arch of nicRxFromMacDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicRxFromMacDaemon_CP_2868_start: Boolean;
  signal nicRxFromMacDaemon_CP_2868_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component nextLSTATE_Volatile is -- 
    port ( -- 
      RX : in  std_logic_vector(72 downto 0);
      LSTATE : in  std_logic_vector(1 downto 0);
      nLSTATE : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal call_stmt_1813_call_ack_0 : boolean;
  signal nLSTATE_1853_1837_buf_req_1 : boolean;
  signal call_stmt_1831_call_req_0 : boolean;
  signal call_stmt_1831_call_ack_0 : boolean;
  signal nLSTATE_1853_1837_buf_ack_1 : boolean;
  signal phi_stmt_1834_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_1840_inst_ack_0 : boolean;
  signal phi_stmt_1834_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_1840_inst_req_1 : boolean;
  signal phi_stmt_1834_ack_0 : boolean;
  signal do_while_stmt_1832_branch_req_0 : boolean;
  signal nLSTATE_1853_1837_buf_req_0 : boolean;
  signal if_stmt_1814_branch_req_0 : boolean;
  signal call_stmt_1813_call_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_1840_inst_req_0 : boolean;
  signal call_stmt_1813_call_ack_1 : boolean;
  signal if_stmt_1814_branch_ack_1 : boolean;
  signal nLSTATE_1853_1837_buf_ack_0 : boolean;
  signal if_stmt_1814_branch_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_1840_inst_ack_1 : boolean;
  signal call_stmt_1813_call_req_0 : boolean;
  signal phi_stmt_1841_req_1 : boolean;
  signal phi_stmt_1841_ack_0 : boolean;
  signal npkt_cnt_1891_1845_buf_req_1 : boolean;
  signal npkt_cnt_1891_1845_buf_ack_1 : boolean;
  signal call_stmt_1831_call_ack_1 : boolean;
  signal call_stmt_1831_call_req_1 : boolean;
  signal phi_stmt_1841_req_0 : boolean;
  signal npkt_cnt_1891_1845_buf_req_0 : boolean;
  signal npkt_cnt_1891_1845_buf_ack_0 : boolean;
  signal MUX_1873_inst_req_0 : boolean;
  signal MUX_1873_inst_ack_0 : boolean;
  signal MUX_1873_inst_req_1 : boolean;
  signal MUX_1873_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_1864_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_header_1864_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_header_1864_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_header_1864_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_packet_1875_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1875_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1875_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_packet_1875_inst_ack_1 : boolean;
  signal call_stmt_1901_call_req_0 : boolean;
  signal call_stmt_1901_call_ack_0 : boolean;
  signal call_stmt_1901_call_req_1 : boolean;
  signal call_stmt_1901_call_ack_1 : boolean;
  signal do_while_stmt_1832_branch_ack_0 : boolean;
  signal do_while_stmt_1832_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicRxFromMacDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicRxFromMacDaemon_CP_2868_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicRxFromMacDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2868_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2868_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2868_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicRxFromMacDaemon_CP_2868: Block -- control-path 
    signal nicRxFromMacDaemon_CP_2868_elements: BooleanArray(82 downto 0);
    -- 
  begin -- 
    nicRxFromMacDaemon_CP_2868_elements(0) <= nicRxFromMacDaemon_CP_2868_start;
    nicRxFromMacDaemon_CP_2868_symbol <= nicRxFromMacDaemon_CP_2868_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	82 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_1801/branch_block_stmt_1801__entry__
      -- CP-element group 0: 	 branch_block_stmt_1801/merge_stmt_1803__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1801/$entry
      -- CP-element group 0: 	 branch_block_stmt_1801/merge_stmt_1803_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1801/merge_stmt_1803__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1801/merge_stmt_1803__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1801/branch_block_stmt_1801__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1801/$exit
      -- 
    nicRxFromMacDaemon_CP_2868_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	81 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	82 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_1801/do_while_stmt_1832__exit__
      -- CP-element group 2: 	 branch_block_stmt_1801/disable_loopback
      -- CP-element group 2: 	 branch_block_stmt_1801/disable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1801/disable_loopback_PhiReq/$exit
      -- 
    nicRxFromMacDaemon_CP_2868_elements(2) <= nicRxFromMacDaemon_CP_2868_elements(81);
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	82 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Sample/$exit
      -- 
    cra_2898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1813_call_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	82 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (49) 
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814__entry__
      -- CP-element group 4: 	 branch_block_stmt_1801/call_stmt_1813__exit__
      -- CP-element group 4: 	 branch_block_stmt_1801/NOT_u1_u1_1818_place
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Sample/req
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Sample/ack
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Update/req
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/BITSEL_u32_u1_1817_inputs/RPIPE_CONTROL_REGISTER_1815/Update/ack
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/BITSEL_u32_u1_1817/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1801/call_stmt_1813/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/NOT_u1_u1_1818/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1801/if_stmt_1814_else_link/$entry
      -- 
    cca_2903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1813_call_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(4)); -- 
    branch_req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(4), ack => if_stmt_1814_branch_req_0); -- 
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	82 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1801/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1801/if_stmt_1814_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1801/if_stmt_1814_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1801/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1801/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_2964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1814_branch_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(5)); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831__entry__
      -- CP-element group 6: 	 branch_block_stmt_1801/if_stmt_1814__exit__
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1801/if_stmt_1814_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1801/if_stmt_1814_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831/$entry
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Update/ccr
      -- CP-element group 6: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Update/$entry
      -- 
    else_choice_transition_2968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1814_branch_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(6)); -- 
    crr_2980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(6), ack => call_stmt_1831_call_req_0); -- 
    ccr_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(6), ack => call_stmt_1831_call_req_1); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Sample/cra
      -- CP-element group 7: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Sample/$exit
      -- 
    cra_2981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1831_call_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1801/call_stmt_1831__exit__
      -- CP-element group 8: 	 branch_block_stmt_1801/do_while_stmt_1832__entry__
      -- CP-element group 8: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1801/call_stmt_1831/$exit
      -- CP-element group 8: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Update/cca
      -- CP-element group 8: 	 branch_block_stmt_1801/call_stmt_1831/call_stmt_1831_Update/$exit
      -- 
    cca_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1831_call_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(8)); -- 
    -- CP-element group 9:  transition  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832__entry__
      -- CP-element group 9: 	 branch_block_stmt_1801/do_while_stmt_1832/$entry
      -- 
    nicRxFromMacDaemon_CP_2868_elements(9) <= nicRxFromMacDaemon_CP_2868_elements(8);
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	81 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832__exit__
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(10) is bound as output of CP function.
    -- CP-element group 11:  merge  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_back
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(11) is bound as output of CP function.
    -- CP-element group 12:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	80 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1801/do_while_stmt_1832/condition_done
      -- CP-element group 12: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_exit/$entry
      -- CP-element group 12: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_taken/$entry
      -- 
    nicRxFromMacDaemon_CP_2868_elements(12) <= nicRxFromMacDaemon_CP_2868_elements(17);
    -- CP-element group 13:  branch  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	78 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_body_done
      -- 
    nicRxFromMacDaemon_CP_2868_elements(13) <= nicRxFromMacDaemon_CP_2868_elements(78);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	50 
    -- CP-element group 14: 	28 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/back_edge_to_loop_body
      -- 
    nicRxFromMacDaemon_CP_2868_elements(14) <= nicRxFromMacDaemon_CP_2868_elements(11);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	52 
    -- CP-element group 15: 	30 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/first_time_through_loop_body
      -- 
    nicRxFromMacDaemon_CP_2868_elements(15) <= nicRxFromMacDaemon_CP_2868_elements(9);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	46 
    -- CP-element group 16: 	47 
    -- CP-element group 16: 	77 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	22 
    -- CP-element group 16: 	23 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1838_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/$entry
      -- CP-element group 16: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/loop_body_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(16) is bound as output of CP function.
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	77 
    -- CP-element group 17: 	21 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/condition_evaluated
      -- 
    condition_evaluated_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(17), ack => do_while_stmt_1832_branch_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(77) & nicRxFromMacDaemon_CP_2868_elements(21);
      gj_nicRxFromMacDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	46 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	22 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	24 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/aggregated_phi_sample_req
      -- CP-element group 18: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_sample_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(46) & nicRxFromMacDaemon_CP_2868_elements(16) & nicRxFromMacDaemon_CP_2868_elements(22) & nicRxFromMacDaemon_CP_2868_elements(21);
      gj_nicRxFromMacDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	48 
    -- CP-element group 19: 	25 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	78 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	46 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1838_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/aggregated_phi_sample_ack
      -- CP-element group 19: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_sample_completed_
      -- 
    nicRxFromMacDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(44) & nicRxFromMacDaemon_CP_2868_elements(48) & nicRxFromMacDaemon_CP_2868_elements(25);
      gj_nicRxFromMacDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	41 
    -- CP-element group 20: 	47 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	26 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_update_start__ps
      -- CP-element group 20: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/aggregated_phi_update_req
      -- 
    nicRxFromMacDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(41) & nicRxFromMacDaemon_CP_2868_elements(47) & nicRxFromMacDaemon_CP_2868_elements(23);
      gj_nicRxFromMacDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	45 
    -- CP-element group 21: 	49 
    -- CP-element group 21: 	27 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/aggregated_phi_update_ack
      -- 
    nicRxFromMacDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(45) & nicRxFromMacDaemon_CP_2868_elements(49) & nicRxFromMacDaemon_CP_2868_elements(27);
      gj_nicRxFromMacDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(16) & nicRxFromMacDaemon_CP_2868_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	65 
    -- CP-element group 23: 	68 
    -- CP-element group 23: 	75 
    -- CP-element group 23: 	27 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(16) & nicRxFromMacDaemon_CP_2868_elements(65) & nicRxFromMacDaemon_CP_2868_elements(68) & nicRxFromMacDaemon_CP_2868_elements(75) & nicRxFromMacDaemon_CP_2868_elements(27);
      gj_nicRxFromMacDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_sample_start__ps
      -- 
    nicRxFromMacDaemon_CP_2868_elements(24) <= nicRxFromMacDaemon_CP_2868_elements(18);
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	19 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_update_start__ps
      -- 
    nicRxFromMacDaemon_CP_2868_elements(26) <= nicRxFromMacDaemon_CP_2868_elements(20);
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	63 
    -- CP-element group 27: 	67 
    -- CP-element group 27: 	73 
    -- CP-element group 27: 	21 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	23 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	14 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_2868_elements(28) <= nicRxFromMacDaemon_CP_2868_elements(14);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_loopback_sample_req_ps
      -- CP-element group 29: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_loopback_sample_req
      -- 
    phi_stmt_1834_loopback_sample_req_3016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1834_loopback_sample_req_3016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(29), ack => phi_stmt_1834_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_2868_elements(30) <= nicRxFromMacDaemon_CP_2868_elements(15);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_entry_sample_req
      -- CP-element group 31: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_entry_sample_req_ps
      -- 
    phi_stmt_1834_entry_sample_req_3019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1834_entry_sample_req_3019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(31), ack => phi_stmt_1834_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_phi_mux_ack
      -- CP-element group 32: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1834_phi_mux_ack_ps
      -- 
    phi_stmt_1834_phi_mux_ack_3022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1834_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_sample_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_update_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_2868_elements(35) <= nicRxFromMacDaemon_CP_2868_elements(36);
    -- CP-element group 36:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	35 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_S0_1836_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(36) is a control-delay.
    cp_element_36_delay: control_delay_element  generic map(name => " 36_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2868_elements(34), ack => nicRxFromMacDaemon_CP_2868_elements(36), clk => clk, reset =>reset);
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_sample_start__ps
      -- 
    req_3043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(37), ack => nLSTATE_1853_1837_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Update/req
      -- CP-element group 38: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Update/$entry
      -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(38), ack => nLSTATE_1853_1837_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Sample/ack
      -- 
    ack_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1853_1837_buf_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_nLSTATE_1837_update_completed_
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1853_1837_buf_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	65 
    -- CP-element group 41: 	71 
    -- CP-element group 41: 	75 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1838_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(16) & nicRxFromMacDaemon_CP_2868_elements(65) & nicRxFromMacDaemon_CP_2868_elements(71) & nicRxFromMacDaemon_CP_2868_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Sample/rr
      -- 
    rr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(42), ack => RPIPE_mac_to_nic_data_1840_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(18) & nicRxFromMacDaemon_CP_2868_elements(45);
      gj_nicRxFromMacDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Update/cr
      -- 
    cr_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(43), ack => RPIPE_mac_to_nic_data_1840_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(44) & nicRxFromMacDaemon_CP_2868_elements(20);
      gj_nicRxFromMacDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	19 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Sample/$exit
      -- 
    ra_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1840_inst_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	63 
    -- CP-element group 45: 	70 
    -- CP-element group 45: 	73 
    -- CP-element group 45: 	21 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	42 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1838_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/RPIPE_mac_to_nic_data_1840_Update/ca
      -- 
    ca_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1840_inst_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(45)); -- 
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	16 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	19 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	18 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(16) & nicRxFromMacDaemon_CP_2868_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: 	75 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	20 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(16) & nicRxFromMacDaemon_CP_2868_elements(49) & nicRxFromMacDaemon_CP_2868_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	19 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	73 
    -- CP-element group 49: 	21 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_update_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	14 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_2868_elements(50) <= nicRxFromMacDaemon_CP_2868_elements(14);
    -- CP-element group 51:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_loopback_sample_req_ps
      -- CP-element group 51: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_loopback_sample_req
      -- 
    phi_stmt_1841_loopback_sample_req_3078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1841_loopback_sample_req_3078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(51), ack => phi_stmt_1841_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	15 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_2868_elements(52) <= nicRxFromMacDaemon_CP_2868_elements(15);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_entry_sample_req_ps
      -- CP-element group 53: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_entry_sample_req
      -- 
    phi_stmt_1841_entry_sample_req_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1841_entry_sample_req_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(53), ack => phi_stmt_1841_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_phi_mux_ack
      -- CP-element group 54: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/phi_stmt_1841_phi_mux_ack_ps
      -- 
    phi_stmt_1841_phi_mux_ack_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1841_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_sample_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_update_start__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_2868_elements(57) <= nicRxFromMacDaemon_CP_2868_elements(58);
    -- CP-element group 58:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	57 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/type_cast_1844_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2868_elements(56), ack => nicRxFromMacDaemon_CP_2868_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_sample_start__ps
      -- CP-element group 59: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Sample/req
      -- 
    req_3105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(59), ack => npkt_cnt_1891_1845_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(59) is bound as output of CP function.
    -- CP-element group 60:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (4) 
      -- CP-element group 60: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Update/req
      -- CP-element group 60: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_update_start__ps
      -- CP-element group 60: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Update/$entry
      -- 
    req_3110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(60), ack => npkt_cnt_1891_1845_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_sample_completed__ps
      -- CP-element group 61: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Sample/ack
      -- 
    ack_3106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1891_1845_buf_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(61)); -- 
    -- CP-element group 62:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_update_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/R_npkt_cnt_1845_Update/$exit
      -- 
    ack_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1891_1845_buf_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	45 
    -- CP-element group 63: 	27 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_start/req
      -- 
    req_3120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(63), ack => MUX_1873_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(45) & nicRxFromMacDaemon_CP_2868_elements(27) & nicRxFromMacDaemon_CP_2868_elements(65);
      gj_nicRxFromMacDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: 	68 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_update_start_
      -- CP-element group 64: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_complete/req
      -- 
    req_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(64), ack => MUX_1873_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(66) & nicRxFromMacDaemon_CP_2868_elements(68);
      gj_nicRxFromMacDaemon_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	41 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	23 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_start/ack
      -- 
    ack_3121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1873_inst_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(65)); -- 
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/MUX_1873_complete/ack
      -- 
    ack_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1873_inst_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: 	27 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Sample/req
      -- 
    req_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(67), ack => WPIPE_nic_rx_to_header_1864_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(66) & nicRxFromMacDaemon_CP_2868_elements(27) & nicRxFromMacDaemon_CP_2868_elements(69);
      gj_nicRxFromMacDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: 	23 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_update_start_
      -- CP-element group 68: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Update/req
      -- 
    ack_3135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1864_inst_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(68)); -- 
    req_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(68), ack => WPIPE_nic_rx_to_header_1864_inst_req_1); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	78 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_header_1864_Update/ack
      -- 
    ack_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1864_inst_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	45 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Sample/req
      -- 
    req_3148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(70), ack => WPIPE_nic_rx_to_packet_1875_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(45) & nicRxFromMacDaemon_CP_2868_elements(72);
      gj_nicRxFromMacDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	41 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Update/req
      -- 
    ack_3149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1875_inst_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(71)); -- 
    req_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(71), ack => WPIPE_nic_rx_to_packet_1875_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	78 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/WPIPE_nic_rx_to_packet_1875_Update/ack
      -- 
    ack_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1875_inst_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	45 
    -- CP-element group 73: 	49 
    -- CP-element group 73: 	27 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Sample/crr
      -- 
    crr_3162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(73), ack => call_stmt_1901_call_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 7,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(45) & nicRxFromMacDaemon_CP_2868_elements(49) & nicRxFromMacDaemon_CP_2868_elements(27) & nicRxFromMacDaemon_CP_2868_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_update_start_
      -- CP-element group 74: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Update/ccr
      -- 
    ccr_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(74), ack => call_stmt_1901_call_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicRxFromMacDaemon_CP_2868_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: 	47 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	23 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Sample/cra
      -- 
    cra_3163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1901_call_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(75)); -- 
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/call_stmt_1901_Update/cca
      -- 
    cca_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1901_call_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(76)); -- 
    -- CP-element group 77:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	16 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	17 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_2868_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2868_elements(16), ack => nicRxFromMacDaemon_CP_2868_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	69 
    -- CP-element group 78: 	72 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	19 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	13 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1801/do_while_stmt_1832/do_while_stmt_1832_loop_body/$exit
      -- 
    nicRxFromMacDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2868_elements(69) & nicRxFromMacDaemon_CP_2868_elements(72) & nicRxFromMacDaemon_CP_2868_elements(76) & nicRxFromMacDaemon_CP_2868_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	12 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_exit/$exit
      -- CP-element group 79: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_exit/ack
      -- 
    ack_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1832_branch_ack_0, ack => nicRxFromMacDaemon_CP_2868_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	12 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_taken/$exit
      -- CP-element group 80: 	 branch_block_stmt_1801/do_while_stmt_1832/loop_taken/ack
      -- 
    ack_3177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1832_branch_ack_1, ack => nicRxFromMacDaemon_CP_2868_elements(80)); -- 
    -- CP-element group 81:  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	10 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	2 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1801/do_while_stmt_1832/$exit
      -- 
    nicRxFromMacDaemon_CP_2868_elements(81) <= nicRxFromMacDaemon_CP_2868_elements(10);
    -- CP-element group 82:  merge  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	0 
    -- CP-element group 82: 	2 
    -- CP-element group 82: 	5 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	3 
    -- CP-element group 82: 	4 
    -- CP-element group 82:  members (13) 
      -- CP-element group 82: 	 branch_block_stmt_1801/merge_stmt_1803__exit__
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813__entry__
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813/$entry
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Update/ccr
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1801/call_stmt_1813/call_stmt_1813_Sample/crr
      -- CP-element group 82: 	 branch_block_stmt_1801/merge_stmt_1803_PhiReqMerge
      -- CP-element group 82: 	 branch_block_stmt_1801/merge_stmt_1803_PhiAck/$entry
      -- CP-element group 82: 	 branch_block_stmt_1801/merge_stmt_1803_PhiAck/$exit
      -- CP-element group 82: 	 branch_block_stmt_1801/merge_stmt_1803_PhiAck/dummy
      -- 
    ccr_2902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(82), ack => call_stmt_1813_call_req_1); -- 
    crr_2897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2868_elements(82), ack => call_stmt_1813_call_req_0); -- 
    nicRxFromMacDaemon_CP_2868_elements(82) <= OrReduce(nicRxFromMacDaemon_CP_2868_elements(0) & nicRxFromMacDaemon_CP_2868_elements(2) & nicRxFromMacDaemon_CP_2868_elements(5));
    nicRxFromMacDaemon_do_while_stmt_1832_terminator_3178: loop_terminator -- 
      generic map (name => " nicRxFromMacDaemon_do_while_stmt_1832_terminator_3178", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicRxFromMacDaemon_CP_2868_elements(13),loop_continue => nicRxFromMacDaemon_CP_2868_elements(80),loop_terminate => nicRxFromMacDaemon_CP_2868_elements(79),loop_back => nicRxFromMacDaemon_CP_2868_elements(11),loop_exit => nicRxFromMacDaemon_CP_2868_elements(10),clk => clk, reset => reset); -- 
    phi_stmt_1834_phi_seq_3050_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_2868_elements(30);
      nicRxFromMacDaemon_CP_2868_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_2868_elements(33);
      nicRxFromMacDaemon_CP_2868_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_2868_elements(35);
      nicRxFromMacDaemon_CP_2868_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_2868_elements(28);
      nicRxFromMacDaemon_CP_2868_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_2868_elements(39);
      nicRxFromMacDaemon_CP_2868_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_2868_elements(40);
      nicRxFromMacDaemon_CP_2868_elements(29) <= phi_mux_reqs(1);
      phi_stmt_1834_phi_seq_3050 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1834_phi_seq_3050") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_2868_elements(24), 
          phi_sample_ack => nicRxFromMacDaemon_CP_2868_elements(25), 
          phi_update_req => nicRxFromMacDaemon_CP_2868_elements(26), 
          phi_update_ack => nicRxFromMacDaemon_CP_2868_elements(27), 
          phi_mux_ack => nicRxFromMacDaemon_CP_2868_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1841_phi_seq_3112_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_2868_elements(52);
      nicRxFromMacDaemon_CP_2868_elements(55)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_2868_elements(55);
      nicRxFromMacDaemon_CP_2868_elements(56)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_2868_elements(57);
      nicRxFromMacDaemon_CP_2868_elements(53) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_2868_elements(50);
      nicRxFromMacDaemon_CP_2868_elements(59)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_2868_elements(61);
      nicRxFromMacDaemon_CP_2868_elements(60)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_2868_elements(62);
      nicRxFromMacDaemon_CP_2868_elements(51) <= phi_mux_reqs(1);
      phi_stmt_1841_phi_seq_3112 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1841_phi_seq_3112") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_2868_elements(18), 
          phi_sample_ack => nicRxFromMacDaemon_CP_2868_elements(48), 
          phi_update_req => nicRxFromMacDaemon_CP_2868_elements(20), 
          phi_update_ack => nicRxFromMacDaemon_CP_2868_elements(49), 
          phi_mux_ack => nicRxFromMacDaemon_CP_2868_elements(54), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3002_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicRxFromMacDaemon_CP_2868_elements(14);
        preds(1)  <= nicRxFromMacDaemon_CP_2868_elements(15);
        entry_tmerge_3002 : transition_merge -- 
          generic map(name => " entry_tmerge_3002")
          port map (preds => preds, symbol_out => nicRxFromMacDaemon_CP_2868_elements(16));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1888_wire : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_1817_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1908_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u65_u73_1871_wire : std_logic_vector(72 downto 0);
    signal EQ_u2_u1_1857_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1860_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1867_wire : std_logic_vector(0 downto 0);
    signal LSTATE_1834 : std_logic_vector(1 downto 0);
    signal MUX_1873_wire : std_logic_vector(72 downto 0);
    signal NOT_u1_u1_1818_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1808_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_1826_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_1897_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_1815_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1906_wire : std_logic_vector(31 downto 0);
    signal RPIPE_mac_to_nic_data_1840_wire : std_logic_vector(72 downto 0);
    signal RX_1838 : std_logic_vector(72 downto 0);
    signal R_HEADER_TKEEP_1870_wire_constant : std_logic_vector(7 downto 0);
    signal R_S0_1836_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1856_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1880_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1859_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1866_wire_constant : std_logic_vector(1 downto 0);
    signal ignore_resp0_1813 : std_logic_vector(31 downto 0);
    signal ignore_resp1_1831 : std_logic_vector(31 downto 0);
    signal ignore_resp2_1901 : std_logic_vector(31 downto 0);
    signal konst_1809_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1816_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1827_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1898_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1907_wire_constant : std_logic_vector(31 downto 0);
    signal nLSTATE_1853 : std_logic_vector(1 downto 0);
    signal nLSTATE_1853_1837_buffered : std_logic_vector(1 downto 0);
    signal npkt_cnt_1891 : std_logic_vector(31 downto 0);
    signal npkt_cnt_1891_1845_buffered : std_logic_vector(31 downto 0);
    signal pkt_cnt_1841 : std_logic_vector(31 downto 0);
    signal pkt_complete_1882 : std_logic_vector(0 downto 0);
    signal slice_1869_wire : std_logic_vector(64 downto 0);
    signal type_cast_1805_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1811_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1823_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1829_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1844_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1887_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1894_wire_constant : std_logic_vector(0 downto 0);
    signal write_to_header_1862 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1808_wire_constant <= "1111";
    NOT_u4_u4_1826_wire_constant <= "1111";
    NOT_u4_u4_1897_wire_constant <= "1111";
    R_HEADER_TKEEP_1870_wire_constant <= "00111111";
    R_S0_1836_wire_constant <= "00";
    R_S0_1856_wire_constant <= "00";
    R_S0_1880_wire_constant <= "00";
    R_S1_1859_wire_constant <= "01";
    R_S1_1866_wire_constant <= "01";
    konst_1809_wire_constant <= "010110";
    konst_1816_wire_constant <= "00000000000000000000000000000000";
    konst_1827_wire_constant <= "010110";
    konst_1898_wire_constant <= "010111";
    konst_1907_wire_constant <= "00000000000000000000000000000000";
    type_cast_1805_wire_constant <= "0";
    type_cast_1811_wire_constant <= "00000000000000000000000000000000";
    type_cast_1823_wire_constant <= "0";
    type_cast_1829_wire_constant <= "00000000000000000000000000000001";
    type_cast_1844_wire_constant <= "00000000000000000000000000000000";
    type_cast_1887_wire_constant <= "00000000000000000000000000000001";
    type_cast_1894_wire_constant <= "0";
    phi_stmt_1834: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_S0_1836_wire_constant & nLSTATE_1853_1837_buffered;
      req <= phi_stmt_1834_req_0 & phi_stmt_1834_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1834",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1834_ack_0,
          idata => idata,
          odata => LSTATE_1834,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1834
    phi_stmt_1841: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1844_wire_constant & npkt_cnt_1891_1845_buffered;
      req <= phi_stmt_1841_req_0 & phi_stmt_1841_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1841",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1841_ack_0,
          idata => idata,
          odata => pkt_cnt_1841,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1841
    MUX_1873_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= MUX_1873_inst_req_0;
      MUX_1873_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= MUX_1873_inst_req_1;
      MUX_1873_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  write_to_header_1862(0);
      MUX_1873_inst_gI: SplitGuardInterface generic map(name => "MUX_1873_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      MUX_1873_inst: SelectSplitProtocol generic map(name => "MUX_1873_inst", data_width => 73, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u65_u73_1871_wire, y => RX_1838, sel => EQ_u2_u1_1867_wire, z => MUX_1873_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1890_inst
    npkt_cnt_1891 <= ADD_u32_u32_1888_wire when (pkt_complete_1882(0) /=  '0') else pkt_cnt_1841;
    -- flow-through slice operator slice_1869_inst
    slice_1869_wire <= RX_1838(72 downto 8);
    nLSTATE_1853_1837_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nLSTATE_1853_1837_buf_req_0;
      nLSTATE_1853_1837_buf_ack_0<= wack(0);
      rreq(0) <= nLSTATE_1853_1837_buf_req_1;
      nLSTATE_1853_1837_buf_ack_1<= rack(0);
      nLSTATE_1853_1837_buf : InterlockBuffer generic map ( -- 
        name => "nLSTATE_1853_1837_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nLSTATE_1853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nLSTATE_1853_1837_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    npkt_cnt_1891_1845_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= npkt_cnt_1891_1845_buf_req_0;
      npkt_cnt_1891_1845_buf_ack_0<= wack(0);
      rreq(0) <= npkt_cnt_1891_1845_buf_req_1;
      npkt_cnt_1891_1845_buf_ack_1<= rack(0);
      npkt_cnt_1891_1845_buf : InterlockBuffer generic map ( -- 
        name => "npkt_cnt_1891_1845_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => npkt_cnt_1891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => npkt_cnt_1891_1845_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1838
    process(RPIPE_mac_to_nic_data_1840_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_mac_to_nic_data_1840_wire(72 downto 0);
      RX_1838 <= tmp_var; -- 
    end process;
    do_while_stmt_1832_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1908_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1832_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1832_branch_req_0,
          ack0 => do_while_stmt_1832_branch_ack_0,
          ack1 => do_while_stmt_1832_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1814_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1818_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1814_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1814_branch_req_0,
          ack0 => if_stmt_1814_branch_ack_0,
          ack1 => if_stmt_1814_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1888_inst
    process(pkt_cnt_1841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pkt_cnt_1841, type_cast_1887_wire_constant, tmp_var);
      ADD_u32_u32_1888_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1817_inst
    process(RPIPE_CONTROL_REGISTER_1815_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1815_wire, konst_1816_wire_constant, tmp_var);
      BITSEL_u32_u1_1817_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1908_inst
    process(RPIPE_CONTROL_REGISTER_1906_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1906_wire, konst_1907_wire_constant, tmp_var);
      BITSEL_u32_u1_1908_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u65_u73_1871_inst
    process(slice_1869_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1869_wire, R_HEADER_TKEEP_1870_wire_constant, tmp_var);
      CONCAT_u65_u73_1871_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1857_inst
    process(LSTATE_1834) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1834, R_S0_1856_wire_constant, tmp_var);
      EQ_u2_u1_1857_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1860_inst
    process(LSTATE_1834) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1834, R_S1_1859_wire_constant, tmp_var);
      EQ_u2_u1_1860_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1867_inst
    process(LSTATE_1834) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1834, R_S1_1866_wire_constant, tmp_var);
      EQ_u2_u1_1867_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1881_inst
    process(nLSTATE_1853) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(nLSTATE_1853, R_S0_1880_wire_constant, tmp_var);
      pkt_complete_1882 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1818_inst
    process(BITSEL_u32_u1_1817_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1817_wire, tmp_var);
      NOT_u1_u1_1818_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1861_inst
    process(EQ_u2_u1_1857_wire, EQ_u2_u1_1860_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_1857_wire, EQ_u2_u1_1860_wire, tmp_var);
      write_to_header_1862 <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1815_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1906_wire <= CONTROL_REGISTER;
    -- shared inport operator group (2) : RPIPE_mac_to_nic_data_1840_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_1840_inst_req_0;
      RPIPE_mac_to_nic_data_1840_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_1840_inst_req_1;
      RPIPE_mac_to_nic_data_1840_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_1840_wire <= data_out(72 downto 0);
      mac_to_nic_data_read_2_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_read_2: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_read_2", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_pipe_read_req(0),
          oack => mac_to_nic_data_pipe_read_ack(0),
          odata => mac_to_nic_data_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_nic_rx_to_header_1864_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_header_1864_inst_req_0;
      WPIPE_nic_rx_to_header_1864_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_header_1864_inst_req_1;
      WPIPE_nic_rx_to_header_1864_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_to_header_1862(0);
      data_in <= MUX_1873_wire;
      nic_rx_to_header_write_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_write_0: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_header", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_header_pipe_write_req(0),
          oack => nic_rx_to_header_pipe_write_ack(0),
          odata => nic_rx_to_header_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_rx_to_packet_1875_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1875_inst_req_0;
      WPIPE_nic_rx_to_packet_1875_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1875_inst_req_1;
      WPIPE_nic_rx_to_packet_1875_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= RX_1838;
      nic_rx_to_packet_write_1_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_write_1: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_packet", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_packet_pipe_write_req(0),
          oack => nic_rx_to_packet_pipe_write_ack(0),
          odata => nic_rx_to_packet_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1813_call call_stmt_1831_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1813_call_req_0;
      reqL_unguarded(0) <= call_stmt_1831_call_req_0;
      call_stmt_1813_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1831_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1813_call_req_1;
      reqR_unguarded(0) <= call_stmt_1831_call_req_1;
      call_stmt_1813_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1831_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      AccessRegister_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1805_wire_constant & NOT_u4_u4_1808_wire_constant & konst_1809_wire_constant & type_cast_1811_wire_constant & type_cast_1823_wire_constant & NOT_u4_u4_1826_wire_constant & konst_1827_wire_constant & type_cast_1829_wire_constant;
      ignore_resp0_1813 <= data_out(63 downto 32);
      ignore_resp1_1831 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(1),
          ackR => AccessRegister_call_acks(1),
          dataR => AccessRegister_call_data(85 downto 43),
          tagR => AccessRegister_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(1), -- cross-over
          ackL => AccessRegister_return_reqs(1), -- cross-over
          dataL => AccessRegister_return_data(63 downto 32),
          tagL => AccessRegister_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_nextLSTATE_4691: nextLSTATE_Volatile port map(RX => RX_1838, LSTATE => LSTATE_1834, nLSTATE => nLSTATE_1853); 
    -- shared call operator group (2) : call_stmt_1901_call 
    AccessRegister_call_group_2: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1901_call_req_0;
      call_stmt_1901_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1901_call_req_1;
      call_stmt_1901_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= pkt_complete_1882(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_2_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1894_wire_constant & NOT_u4_u4_1897_wire_constant & konst_1898_wire_constant & pkt_cnt_1841;
      ignore_resp2_1901 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end nicRxFromMacDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity popFromQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(35 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(35 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_call_data : out  std_logic_vector(67 downto 0);
    getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_return_data : in   std_logic_vector(31 downto 0);
    getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(35 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
    updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity popFromQueue;
architecture popFromQueue_arch of popFromQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 37)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal popFromQueue_CP_748_start: Boolean;
  signal popFromQueue_CP_748_symbol: Boolean;
  -- volatile/operator module components. 
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_911_call_req_0 : boolean;
  signal call_stmt_957_call_req_0 : boolean;
  signal call_stmt_911_call_ack_0 : boolean;
  signal call_stmt_939_call_ack_0 : boolean;
  signal call_stmt_934_call_req_0 : boolean;
  signal call_stmt_898_call_ack_1 : boolean;
  signal call_stmt_957_call_req_1 : boolean;
  signal call_stmt_946_call_ack_1 : boolean;
  signal call_stmt_939_call_req_0 : boolean;
  signal call_stmt_939_call_req_1 : boolean;
  signal call_stmt_957_call_ack_0 : boolean;
  signal call_stmt_903_call_req_0 : boolean;
  signal call_stmt_898_call_req_0 : boolean;
  signal call_stmt_914_call_req_0 : boolean;
  signal call_stmt_911_call_ack_1 : boolean;
  signal call_stmt_911_call_req_1 : boolean;
  signal call_stmt_903_call_ack_1 : boolean;
  signal W_status_958_inst_ack_1 : boolean;
  signal W_status_958_inst_req_1 : boolean;
  signal call_stmt_903_call_ack_0 : boolean;
  signal call_stmt_934_call_ack_0 : boolean;
  signal call_stmt_939_call_ack_1 : boolean;
  signal call_stmt_914_call_ack_0 : boolean;
  signal call_stmt_946_call_req_0 : boolean;
  signal call_stmt_898_call_ack_0 : boolean;
  signal call_stmt_898_call_req_1 : boolean;
  signal call_stmt_903_call_req_1 : boolean;
  signal call_stmt_957_call_ack_1 : boolean;
  signal call_stmt_934_call_ack_1 : boolean;
  signal call_stmt_934_call_req_1 : boolean;
  signal call_stmt_914_call_ack_1 : boolean;
  signal W_status_958_inst_req_0 : boolean;
  signal W_status_958_inst_ack_0 : boolean;
  signal call_stmt_946_call_req_1 : boolean;
  signal call_stmt_914_call_req_1 : boolean;
  signal call_stmt_946_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "popFromQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 37) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(tag_length + 36 downto 37) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 36 downto 37);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  popFromQueue_CP_748_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "popFromQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_748_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= popFromQueue_CP_748_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_748_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  popFromQueue_CP_748: Block -- control-path 
    signal popFromQueue_CP_748_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    popFromQueue_CP_748_elements(0) <= popFromQueue_CP_748_start;
    popFromQueue_CP_748_symbol <= popFromQueue_CP_748_elements(22);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_898/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_898/call_stmt_898_sample_start_
      -- CP-element group 0: 	 call_stmt_898/call_stmt_898_Sample/crr
      -- CP-element group 0: 	 call_stmt_898/call_stmt_898_update_start_
      -- CP-element group 0: 	 call_stmt_898/call_stmt_898_Update/$entry
      -- CP-element group 0: 	 call_stmt_898/call_stmt_898_Update/ccr
      -- CP-element group 0: 	 call_stmt_898/call_stmt_898_Sample/$entry
      -- 
    crr_761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(0), ack => call_stmt_898_call_req_0); -- 
    ccr_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(0), ack => call_stmt_898_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_898/call_stmt_898_sample_completed_
      -- CP-element group 1: 	 call_stmt_898/call_stmt_898_Sample/cra
      -- CP-element group 1: 	 call_stmt_898/call_stmt_898_Sample/$exit
      -- 
    cra_762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_898_call_ack_0, ack => popFromQueue_CP_748_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (26) 
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_update_start_
      -- CP-element group 2: 	 call_stmt_898/$exit
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Update/$entry
      -- CP-element group 2: 	 call_stmt_898/call_stmt_898_Update/$exit
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_update_start_
      -- CP-element group 2: 	 call_stmt_898/call_stmt_898_Update/cca
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Update/$entry
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Update/ccr
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Sample/crr
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Sample/$entry
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_update_start_
      -- CP-element group 2: 	 call_stmt_898/call_stmt_898_update_completed_
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Update/ccr
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_update_start_
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Update/$entry
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Update/$entry
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Update/ccr
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Update/ccr
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_sample_start_
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Update/$entry
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_update_start_
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_update_start_
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/$entry
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Update/ccr
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Update/ccr
      -- CP-element group 2: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Update/$entry
      -- 
    cca_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_898_call_ack_1, ack => popFromQueue_CP_748_elements(2)); -- 
    crr_778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(2), ack => call_stmt_903_call_req_0); -- 
    ccr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(2), ack => call_stmt_903_call_req_1); -- 
    ccr_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(2), ack => call_stmt_911_call_req_1); -- 
    ccr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(2), ack => call_stmt_914_call_req_1); -- 
    ccr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(2), ack => call_stmt_934_call_req_1); -- 
    ccr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(2), ack => call_stmt_939_call_req_1); -- 
    ccr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(2), ack => call_stmt_946_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Sample/$exit
      -- CP-element group 3: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_sample_completed_
      -- CP-element group 3: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Sample/cra
      -- 
    cra_779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_903_call_ack_0, ack => popFromQueue_CP_748_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	9 
    -- CP-element group 4: 	12 
    -- CP-element group 4: 	15 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Sample/crr
      -- CP-element group 4: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_sample_start_
      -- CP-element group 4: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_update_completed_
      -- CP-element group 4: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Update/cca
      -- CP-element group 4: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Sample/$entry
      -- CP-element group 4: 	 call_stmt_903_to_call_stmt_946/call_stmt_903_Update/$exit
      -- 
    cca_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_903_call_ack_1, ack => popFromQueue_CP_748_elements(4)); -- 
    crr_792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(4), ack => call_stmt_911_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Sample/cra
      -- CP-element group 5: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_sample_completed_
      -- CP-element group 5: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Sample/$exit
      -- 
    cra_793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_911_call_ack_0, ack => popFromQueue_CP_748_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	12 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Sample/$entry
      -- CP-element group 6: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Sample/crr
      -- CP-element group 6: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Update/cca
      -- CP-element group 6: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_Update/$exit
      -- CP-element group 6: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_sample_start_
      -- CP-element group 6: 	 call_stmt_903_to_call_stmt_946/call_stmt_911_update_completed_
      -- 
    cca_798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_911_call_ack_1, ack => popFromQueue_CP_748_elements(6)); -- 
    crr_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(6), ack => call_stmt_914_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_sample_completed_
      -- CP-element group 7: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Sample/$exit
      -- CP-element group 7: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Sample/cra
      -- 
    cra_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_914_call_ack_0, ack => popFromQueue_CP_748_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	15 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Update/$exit
      -- CP-element group 8: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_Update/cca
      -- CP-element group 8: 	 call_stmt_903_to_call_stmt_946/call_stmt_914_update_completed_
      -- 
    cca_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_914_call_ack_1, ack => popFromQueue_CP_748_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Sample/crr
      -- CP-element group 9: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Sample/$entry
      -- CP-element group 9: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_sample_start_
      -- 
    crr_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(9), ack => call_stmt_934_call_req_0); -- 
    popFromQueue_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "popFromQueue_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_748_elements(4) & popFromQueue_CP_748_elements(8);
      gj_popFromQueue_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_748_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Sample/$exit
      -- CP-element group 10: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Sample/cra
      -- CP-element group 10: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_sample_completed_
      -- 
    cra_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_934_call_ack_0, ack => popFromQueue_CP_748_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_update_completed_
      -- CP-element group 11: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Update/cca
      -- CP-element group 11: 	 call_stmt_903_to_call_stmt_946/call_stmt_934_Update/$exit
      -- 
    cca_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_934_call_ack_1, ack => popFromQueue_CP_748_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	4 
    -- CP-element group 12: 	6 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Sample/crr
      -- CP-element group 12: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Sample/$entry
      -- CP-element group 12: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_sample_start_
      -- 
    crr_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(12), ack => call_stmt_939_call_req_0); -- 
    popFromQueue_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= popFromQueue_CP_748_elements(4) & popFromQueue_CP_748_elements(6) & popFromQueue_CP_748_elements(11);
      gj_popFromQueue_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_748_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Sample/$exit
      -- CP-element group 13: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Sample/cra
      -- CP-element group 13: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_sample_completed_
      -- 
    cra_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_939_call_ack_0, ack => popFromQueue_CP_748_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_update_completed_
      -- CP-element group 14: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Update/$exit
      -- CP-element group 14: 	 call_stmt_903_to_call_stmt_946/call_stmt_939_Update/cca
      -- 
    cca_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_939_call_ack_1, ack => popFromQueue_CP_748_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	8 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_sample_start_
      -- CP-element group 15: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Sample/$entry
      -- CP-element group 15: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Sample/crr
      -- 
    crr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(15), ack => call_stmt_946_call_req_0); -- 
    popFromQueue_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= popFromQueue_CP_748_elements(4) & popFromQueue_CP_748_elements(8) & popFromQueue_CP_748_elements(14);
      gj_popFromQueue_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_748_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Sample/$exit
      -- CP-element group 16: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_sample_completed_
      -- CP-element group 16: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Sample/cra
      -- 
    cra_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_946_call_ack_0, ack => popFromQueue_CP_748_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (17) 
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Sample/crr
      -- CP-element group 17: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Update/$exit
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Update/ccr
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_update_start_
      -- CP-element group 17: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_Update/cca
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Sample/$entry
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_sample_start_
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Update/req
      -- CP-element group 17: 	 call_stmt_903_to_call_stmt_946/call_stmt_946_update_completed_
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_update_start_
      -- CP-element group 17: 	 call_stmt_903_to_call_stmt_946/$exit
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_sample_start_
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/$entry
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Update/$entry
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Update/$entry
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Sample/req
      -- CP-element group 17: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Sample/$entry
      -- 
    cca_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_946_call_ack_1, ack => popFromQueue_CP_748_elements(17)); -- 
    crr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(17), ack => call_stmt_957_call_req_0); -- 
    ccr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(17), ack => call_stmt_957_call_req_1); -- 
    req_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(17), ack => W_status_958_inst_req_0); -- 
    req_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_748_elements(17), ack => W_status_958_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Sample/$exit
      -- CP-element group 18: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Sample/cra
      -- CP-element group 18: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_sample_completed_
      -- 
    cra_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_957_call_ack_0, ack => popFromQueue_CP_748_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Update/$exit
      -- CP-element group 19: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_update_completed_
      -- CP-element group 19: 	 call_stmt_957_to_assign_stmt_960/call_stmt_957_Update/cca
      -- 
    cca_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_957_call_ack_1, ack => popFromQueue_CP_748_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_sample_completed_
      -- CP-element group 20: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Sample/$exit
      -- CP-element group 20: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Sample/ack
      -- 
    ack_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_958_inst_ack_0, ack => popFromQueue_CP_748_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_update_completed_
      -- CP-element group 21: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Update/ack
      -- CP-element group 21: 	 call_stmt_957_to_assign_stmt_960/assign_stmt_960_Update/$exit
      -- 
    ack_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_958_inst_ack_1, ack => popFromQueue_CP_748_elements(21)); -- 
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 $exit
      -- CP-element group 22: 	 call_stmt_957_to_assign_stmt_960/$exit
      -- 
    popFromQueue_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_748_elements(19) & popFromQueue_CP_748_elements(21);
      gj_popFromQueue_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_748_elements(22), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_927_wire : std_logic_vector(31 downto 0);
    signal Queue_Length_911 : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_919_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_945_wire : std_logic_vector(31 downto 0);
    signal konst_918_wire_constant : std_logic_vector(31 downto 0);
    signal konst_924_wire_constant : std_logic_vector(31 downto 0);
    signal konst_926_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_898 : std_logic_vector(0 downto 0);
    signal next_ri_929 : std_logic_vector(31 downto 0);
    signal q_empty_908 : std_logic_vector(0 downto 0);
    signal read_index_903 : std_logic_vector(31 downto 0);
    signal round_off_921 : std_logic_vector(0 downto 0);
    signal total_msgs_914 : std_logic_vector(31 downto 0);
    signal type_cast_944_wire_constant : std_logic_vector(31 downto 0);
    signal write_index_903 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_918_wire_constant <= "00000000000000000000000000000001";
    konst_924_wire_constant <= "00000000000000000000000000000000";
    konst_926_wire_constant <= "00000000000000000000000000000001";
    type_cast_944_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_928_inst
    next_ri_929 <= konst_924_wire_constant when (round_off_921(0) /=  '0') else ADD_u32_u32_927_wire;
    W_status_958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_958_inst_req_0;
      W_status_958_inst_ack_0<= wack(0);
      rreq(0) <= W_status_958_inst_req_1;
      W_status_958_inst_ack_1<= rack(0);
      W_status_958_inst : InterlockBuffer generic map ( -- 
        name => "W_status_958_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_empty_908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator ADD_u32_u32_927_inst
    process(read_index_903) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(read_index_903, konst_926_wire_constant, tmp_var);
      ADD_u32_u32_927_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_907_inst
    process(write_index_903, read_index_903) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_index_903, read_index_903, tmp_var);
      q_empty_908 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_920_inst
    process(read_index_903, SUB_u32_u32_919_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(read_index_903, SUB_u32_u32_919_wire, tmp_var);
      round_off_921 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_919_inst
    process(Queue_Length_911) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(Queue_Length_911, konst_918_wire_constant, tmp_var);
      SUB_u32_u32_919_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_945_inst
    process(total_msgs_914) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(total_msgs_914, type_cast_944_wire_constant, tmp_var);
      SUB_u32_u32_945_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_898_call 
    acquireLock_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_898_call_req_0;
      call_stmt_898_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_898_call_req_1;
      call_stmt_898_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_0_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_898 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(35 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_903_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_903_call_req_0;
      call_stmt_903_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_903_call_req_1;
      call_stmt_903_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_index_903 <= data_out(63 downto 32);
      read_index_903 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_911_call 
    getQueueLength_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_911_call_req_0;
      call_stmt_911_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_911_call_req_1;
      call_stmt_911_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_2_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      Queue_Length_911 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(35 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_914_call 
    getTotalMessages_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_914_call_req_0;
      call_stmt_914_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_914_call_req_1;
      call_stmt_914_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_3_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      total_msgs_914 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(35 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_934_call 
    getQueueElement_call_group_4: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_934_call_req_0;
      call_stmt_934_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_934_call_req_1;
      call_stmt_934_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_908(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueElement_call_group_4_gI: SplitGuardInterface generic map(name => "getQueueElement_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & read_index_903;
      q_r_data_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueElement_call_reqs(0),
          ackR => getQueueElement_call_acks(0),
          dataR => getQueueElement_call_data(67 downto 0),
          tagR => getQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueElement_return_acks(0), -- cross-over
          ackL => getQueueElement_return_reqs(0), -- cross-over
          dataL => getQueueElement_return_data(31 downto 0),
          tagL => getQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_939_call 
    setQueuePointers_call_group_5: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_939_call_req_0;
      call_stmt_939_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_939_call_req_1;
      call_stmt_939_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_908(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_5_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_index_903 & next_ri_929;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_946_call 
    updateTotalMessages_call_group_6: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_946_call_req_0;
      call_stmt_946_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_946_call_req_1;
      call_stmt_946_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_908(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateTotalMessages_call_group_6_gI: SplitGuardInterface generic map(name => "updateTotalMessages_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & SUB_u32_u32_945_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateTotalMessages_call_reqs(0),
          ackR => updateTotalMessages_call_acks(0),
          dataR => updateTotalMessages_call_data(67 downto 0),
          tagR => updateTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => updateTotalMessages_return_acks(0), -- cross-over
          ackL => updateTotalMessages_return_reqs(0), -- cross-over
          tagL => updateTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_957_call 
    releaseLock_call_group_7: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_957_call_req_0;
      call_stmt_957_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_957_call_req_1;
      call_stmt_957_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_7_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(35 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- 
  end Block; -- data_path
  -- 
end popFromQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity populateRxQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity populateRxQueue;
architecture populateRxQueue_arch of populateRxQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal populateRxQueue_CP_1558_start: Boolean;
  signal populateRxQueue_CP_1558_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component delay_time_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      T : in  std_logic_vector(31 downto 0);
      delay_done : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1346_call_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_ack_1 : boolean;
  signal if_stmt_1377_branch_ack_1 : boolean;
  signal if_stmt_1377_branch_req_0 : boolean;
  signal call_stmt_1363_call_ack_0 : boolean;
  signal AND_u6_u6_1372_inst_req_1 : boolean;
  signal AND_u6_u6_1372_inst_req_0 : boolean;
  signal call_stmt_1382_call_ack_1 : boolean;
  signal AND_u6_u6_1372_inst_ack_0 : boolean;
  signal AND_u6_u6_1372_inst_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_req_1 : boolean;
  signal if_stmt_1377_branch_ack_0 : boolean;
  signal call_stmt_1363_call_req_0 : boolean;
  signal if_stmt_1383_branch_req_0 : boolean;
  signal phi_stmt_1315_ack_0 : boolean;
  signal AND_u6_u6_1324_inst_req_0 : boolean;
  signal AND_u6_u6_1324_inst_ack_0 : boolean;
  signal call_stmt_1382_call_req_1 : boolean;
  signal n_q_index_1373_1325_buf_req_1 : boolean;
  signal phi_stmt_1315_req_0 : boolean;
  signal AND_u6_u6_1324_inst_ack_1 : boolean;
  signal AND_u6_u6_1324_inst_req_1 : boolean;
  signal n_q_index_1373_1325_buf_req_0 : boolean;
  signal phi_stmt_1315_req_1 : boolean;
  signal n_q_index_1373_1325_buf_ack_1 : boolean;
  signal n_q_index_1373_1325_buf_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_req_0 : boolean;
  signal call_stmt_1382_call_ack_0 : boolean;
  signal call_stmt_1382_call_req_0 : boolean;
  signal call_stmt_1346_call_ack_1 : boolean;
  signal if_stmt_1383_branch_ack_0 : boolean;
  signal call_stmt_1346_call_req_1 : boolean;
  signal if_stmt_1383_branch_ack_1 : boolean;
  signal call_stmt_1363_call_ack_1 : boolean;
  signal call_stmt_1363_call_req_1 : boolean;
  signal call_stmt_1346_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "populateRxQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  populateRxQueue_CP_1558_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "populateRxQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1558_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= populateRxQueue_CP_1558_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1558_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  populateRxQueue_CP_1558: Block -- control-path 
    signal populateRxQueue_CP_1558_elements: BooleanArray(25 downto 0);
    -- 
  begin -- 
    populateRxQueue_CP_1558_elements(0) <= populateRxQueue_CP_1558_start;
    populateRxQueue_CP_1558_symbol <= populateRxQueue_CP_1558_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1313/merge_stmt_1314__entry__
      -- CP-element group 0: 	 branch_block_stmt_1313/$entry
      -- CP-element group 0: 	 branch_block_stmt_1313/branch_block_stmt_1313__entry__
      -- CP-element group 0: 	 branch_block_stmt_1313/merge_stmt_1314_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	16 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1313/$exit
      -- CP-element group 1: 	 branch_block_stmt_1313/if_stmt_1377__exit__
      -- CP-element group 1: 	 branch_block_stmt_1313/branch_block_stmt_1313__exit__
      -- 
    populateRxQueue_CP_1558_elements(1) <= OrReduce(populateRxQueue_CP_1558_elements(14) & populateRxQueue_CP_1558_elements(16));
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	25 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Sample/cra
      -- 
    cra_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1346_call_ack_0, ack => populateRxQueue_CP_1558_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	25 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Update/$exit
      -- 
    cca_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1346_call_ack_1, ack => populateRxQueue_CP_1558_elements(3)); -- 
    crr_1596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(3), ack => call_stmt_1363_call_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Sample/cra
      -- CP-element group 4: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Sample/$exit
      -- 
    cra_1597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1363_call_ack_0, ack => populateRxQueue_CP_1558_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Update/cca
      -- 
    cca_1602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1363_call_ack_1, ack => populateRxQueue_CP_1558_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	25 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_sample_completed_
      -- 
    ra_1611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1372_inst_ack_0, ack => populateRxQueue_CP_1558_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	25 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_update_completed_
      -- 
    ca_1616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1372_inst_ack_1, ack => populateRxQueue_CP_1558_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (22) 
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/branch_req
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/$exit
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_else_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/$exit
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377_eval_test/NOT_u1_u1_1379/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1313/NOT_u1_u1_1379_place
      -- CP-element group 8: 	 branch_block_stmt_1313/if_stmt_1377__entry__
      -- CP-element group 8: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373__exit__
      -- 
    branch_req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(8), ack => if_stmt_1377_branch_req_0); -- 
    populateRxQueue_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "populateRxQueue_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1558_elements(5) & populateRxQueue_CP_1558_elements(7);
      gj_populateRxQueue_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1558_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_1313/if_stmt_1377_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_1313/if_stmt_1377_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Update/ccr
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382__entry__
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Sample/crr
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1313/call_stmt_1382/$entry
      -- 
    if_choice_transition_1645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1377_branch_ack_1, ack => populateRxQueue_CP_1558_elements(9)); -- 
    ccr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(9), ack => call_stmt_1382_call_req_1); -- 
    crr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(9), ack => call_stmt_1382_call_req_0); -- 
    -- CP-element group 10:  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_1313/assign_stmt_1392/$entry
      -- CP-element group 10: 	 branch_block_stmt_1313/assign_stmt_1392__entry__
      -- CP-element group 10: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1313/if_stmt_1377_else_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_1313/if_stmt_1377_else_link/else_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Sample/req
      -- CP-element group 10: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Sample/$entry
      -- 
    else_choice_transition_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1377_branch_ack_0, ack => populateRxQueue_CP_1558_elements(10)); -- 
    req_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(10), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Sample/cra
      -- CP-element group 11: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_sample_completed_
      -- 
    cra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1382_call_ack_0, ack => populateRxQueue_CP_1558_elements(11)); -- 
    -- CP-element group 12:  branch  transition  place  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (27) 
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Update/cca
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/EQ_u1_u1_1386_place
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/SplitProtocol/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/EQ_u1_u1_1386_inputs/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/EQ_u1_u1_1386_inputs/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_eval_test/EQ_u1_u1_1386/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/call_stmt_1382/call_stmt_1382_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_else_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/call_stmt_1382/$exit
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383__entry__
      -- CP-element group 12: 	 branch_block_stmt_1313/if_stmt_1383_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_1313/call_stmt_1382__exit__
      -- 
    cca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1382_call_ack_1, ack => populateRxQueue_CP_1558_elements(12)); -- 
    branch_req_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(12), ack => if_stmt_1383_branch_req_0); -- 
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	21 
    -- CP-element group 13: 	22 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Update/req
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/$entry
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Sample/req
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/$entry
      -- CP-element group 13: 	 branch_block_stmt_1313/loopback
      -- CP-element group 13: 	 branch_block_stmt_1313/if_stmt_1383_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_1313/if_stmt_1383_if_link/$exit
      -- 
    if_choice_transition_1702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_1, ack => populateRxQueue_CP_1558_elements(13)); -- 
    req_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(13), ack => n_q_index_1373_1325_buf_req_1); -- 
    req_1855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(13), ack => n_q_index_1373_1325_buf_req_0); -- 
    -- CP-element group 14:  merge  transition  place  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	1 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1313/if_stmt_1383_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_1313/if_stmt_1383_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_1313/if_stmt_1383__exit__
      -- 
    else_choice_transition_1706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_0, ack => populateRxQueue_CP_1558_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Update/req
      -- CP-element group 15: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Sample/ack
      -- CP-element group 15: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Sample/$exit
      -- 
    ack_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_ack_0, ack => populateRxQueue_CP_1558_elements(15)); -- 
    req_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(15), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_req_1); -- 
    -- CP-element group 16:  transition  place  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	1 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Update/ack
      -- CP-element group 16: 	 branch_block_stmt_1313/assign_stmt_1392__exit__
      -- CP-element group 16: 	 branch_block_stmt_1313/assign_stmt_1392/$exit
      -- CP-element group 16: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1313/assign_stmt_1392/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_Update/$exit
      -- 
    ack_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_ack_1, ack => populateRxQueue_CP_1558_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (71) 
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Update/req
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Update/req
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/ADD_u6_u6_1319_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/ADD_u6_u6_1319/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SUB_u32_u32_1322/SUB_u32_u32_1322_inputs/RPIPE_NUMBER_OF_SERVERS_1320/$exit
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/AND_u6_u6_1324_inputs/type_cast_1323/SplitProtocol/$exit
      -- 
    rr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(17), ack => AND_u6_u6_1324_inst_req_0); -- 
    cr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(17), ack => AND_u6_u6_1324_inst_req_1); -- 
    populateRxQueue_CP_1558_elements(17) <= populateRxQueue_CP_1558_elements(0);
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Sample/$exit
      -- 
    ra_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1324_inst_ack_0, ack => populateRxQueue_CP_1558_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/Update/$exit
      -- 
    ca_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1324_inst_ack_1, ack => populateRxQueue_CP_1558_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	24 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/$exit
      -- CP-element group 20: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/$exit
      -- CP-element group 20: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_req
      -- CP-element group 20: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/SplitProtocol/$exit
      -- CP-element group 20: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/AND_u6_u6_1324/$exit
      -- CP-element group 20: 	 branch_block_stmt_1313/merge_stmt_1314__entry___PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$exit
      -- 
    phi_stmt_1315_req_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1315_req_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(20), ack => phi_stmt_1315_req_0); -- 
    populateRxQueue_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1558_elements(18) & populateRxQueue_CP_1558_elements(19);
      gj_populateRxQueue_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1558_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	13 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Sample/ack
      -- 
    ack_1856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1373_1325_buf_ack_0, ack => populateRxQueue_CP_1558_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/Update/ack
      -- 
    ack_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1373_1325_buf_ack_1, ack => populateRxQueue_CP_1558_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/$exit
      -- CP-element group 23: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/$exit
      -- CP-element group 23: 	 branch_block_stmt_1313/loopback_PhiReq/$exit
      -- CP-element group 23: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_req
      -- CP-element group 23: 	 branch_block_stmt_1313/loopback_PhiReq/phi_stmt_1315/phi_stmt_1315_sources/Interlock/$exit
      -- 
    phi_stmt_1315_req_1862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1315_req_1862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(23), ack => phi_stmt_1315_req_1); -- 
    populateRxQueue_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1558_elements(21) & populateRxQueue_CP_1558_elements(22);
      gj_populateRxQueue_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1558_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  merge  transition  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1313/merge_stmt_1314_PhiAck/$entry
      -- CP-element group 24: 	 branch_block_stmt_1313/merge_stmt_1314_PhiReqMerge
      -- 
    populateRxQueue_CP_1558_elements(24) <= OrReduce(populateRxQueue_CP_1558_elements(20) & populateRxQueue_CP_1558_elements(23));
    -- CP-element group 25:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: 	3 
    -- CP-element group 25: 	5 
    -- CP-element group 25: 	6 
    -- CP-element group 25: 	7 
    -- CP-element group 25:  members (20) 
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/$entry
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Sample/crr
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1313/merge_stmt_1314__exit__
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373__entry__
      -- CP-element group 25: 	 branch_block_stmt_1313/merge_stmt_1314_PhiAck/$exit
      -- CP-element group 25: 	 branch_block_stmt_1313/merge_stmt_1314_PhiAck/phi_stmt_1315_ack
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/AND_u6_u6_1372_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Update/ccr
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1346_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1313/assign_stmt_1334_to_assign_stmt_1373/call_stmt_1363_Update/ccr
      -- 
    phi_stmt_1315_ack_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1315_ack_0, ack => populateRxQueue_CP_1558_elements(25)); -- 
    crr_1582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(25), ack => call_stmt_1346_call_req_0); -- 
    cr_1615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(25), ack => AND_u6_u6_1372_inst_req_1); -- 
    rr_1610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(25), ack => AND_u6_u6_1372_inst_req_0); -- 
    ccr_1587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(25), ack => call_stmt_1346_call_req_1); -- 
    ccr_1601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1558_elements(25), ack => call_stmt_1363_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1319_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_1332_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_1367_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_1324_wire : std_logic_vector(5 downto 0);
    signal EQ_u1_u1_1386_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1379_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1341_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1320_wire : std_logic_vector(31 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1368_wire : std_logic_vector(31 downto 0);
    signal R_RX_QUEUES_REG_START_OFFSET_1331_wire_constant : std_logic_vector(5 downto 0);
    signal SUB_u32_u32_1322_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1370_wire : std_logic_vector(31 downto 0);
    signal konst_1318_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1321_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1366_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1369_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1380_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1385_wire_constant : std_logic_vector(0 downto 0);
    signal n_q_index_1373 : std_logic_vector(5 downto 0);
    signal n_q_index_1373_1325_buffered : std_logic_vector(5 downto 0);
    signal push_status_1363 : std_logic_vector(0 downto 0);
    signal q_index_1315 : std_logic_vector(5 downto 0);
    signal register_index_1334 : std_logic_vector(5 downto 0);
    signal rx_queue_pointer_32_1346 : std_logic_vector(31 downto 0);
    signal rx_queue_pointer_36_1352 : std_logic_vector(35 downto 0);
    signal slice_1361_wire : std_logic_vector(31 downto 0);
    signal status_1382 : std_logic_vector(0 downto 0);
    signal type_cast_1323_wire : std_logic_vector(5 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1349_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1358_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1371_wire : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1341_wire_constant <= "1111";
    R_RX_QUEUES_REG_START_OFFSET_1331_wire_constant <= "000010";
    konst_1318_wire_constant <= "000001";
    konst_1321_wire_constant <= "00000000000000000000000000000001";
    konst_1366_wire_constant <= "000001";
    konst_1369_wire_constant <= "00000000000000000000000000000001";
    konst_1380_wire_constant <= "00000000000000000000000000100000";
    konst_1385_wire_constant <= "0";
    type_cast_1338_wire_constant <= "1";
    type_cast_1344_wire_constant <= "00000000000000000000000000000000";
    type_cast_1349_wire_constant <= "0000";
    type_cast_1358_wire_constant <= "0";
    phi_stmt_1315: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= AND_u6_u6_1324_wire & n_q_index_1373_1325_buffered;
      req <= phi_stmt_1315_req_0 & phi_stmt_1315_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1315",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1315_ack_0,
          idata => idata,
          odata => q_index_1315,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1315
    -- flow-through slice operator slice_1361_inst
    slice_1361_wire <= rx_buffer_pointer_buffer(31 downto 0);
    n_q_index_1373_1325_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_q_index_1373_1325_buf_req_0;
      n_q_index_1373_1325_buf_ack_0<= wack(0);
      rreq(0) <= n_q_index_1373_1325_buf_req_1;
      n_q_index_1373_1325_buf_ack_1<= rack(0);
      n_q_index_1373_1325_buf : InterlockBuffer generic map ( -- 
        name => "n_q_index_1373_1325_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_q_index_1373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_q_index_1373_1325_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1323_inst
    process(SUB_u32_u32_1322_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1322_wire(5 downto 0);
      type_cast_1323_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1333_inst
    process(ADD_u6_u6_1332_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1332_wire(5 downto 0);
      register_index_1334 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1371_inst
    process(SUB_u32_u32_1370_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1370_wire(5 downto 0);
      type_cast_1371_wire <= tmp_var; -- 
    end process;
    if_stmt_1377_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1379_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1377_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1377_branch_req_0,
          ack0 => if_stmt_1377_branch_ack_0,
          ack1 => if_stmt_1377_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1383_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_1386_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1383_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1383_branch_req_0,
          ack0 => if_stmt_1383_branch_ack_0,
          ack1 => if_stmt_1383_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u6_u6_1319_inst
    process(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317_wire, konst_1318_wire_constant, tmp_var);
      ADD_u6_u6_1319_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_1332_inst
    process(q_index_1315) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_1315, R_RX_QUEUES_REG_START_OFFSET_1331_wire_constant, tmp_var);
      ADD_u6_u6_1332_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_1367_inst
    process(q_index_1315) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_1315, konst_1366_wire_constant, tmp_var);
      ADD_u6_u6_1367_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_1324_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1319_wire & type_cast_1323_wire;
      AND_u6_u6_1324_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1324_inst_req_0;
      AND_u6_u6_1324_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1324_inst_req_1;
      AND_u6_u6_1324_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : AND_u6_u6_1372_inst 
    ApIntAnd_group_4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1367_wire & type_cast_1371_wire;
      n_q_index_1373 <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1372_inst_req_0;
      AND_u6_u6_1372_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1372_inst_req_1;
      AND_u6_u6_1372_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator CONCAT_u4_u36_1351_inst
    process(type_cast_1349_wire_constant, rx_queue_pointer_32_1346) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1349_wire_constant, rx_queue_pointer_32_1346, tmp_var);
      rx_queue_pointer_36_1352 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1386_inst
    process(status_1382) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(status_1382, konst_1385_wire_constant, tmp_var);
      EQ_u1_u1_1386_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1379_inst
    process(push_status_1363) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", push_status_1363, tmp_var);
      NOT_u1_u1_1379_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u32_u32_1322_inst
    process(RPIPE_NUMBER_OF_SERVERS_1320_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1320_wire, konst_1321_wire_constant, tmp_var);
      SUB_u32_u32_1322_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1370_inst
    process(RPIPE_NUMBER_OF_SERVERS_1368_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1368_wire, konst_1369_wire_constant, tmp_var);
      SUB_u32_u32_1370_wire <= tmp_var; --
    end process;
    -- read from input-signal LAST_WRITTEN_RX_QUEUE_INDEX
    RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1317_wire <= LAST_WRITTEN_RX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_1320_wire <= NUMBER_OF_SERVERS;
    RPIPE_NUMBER_OF_SERVERS_1368_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1390_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= q_index_1315;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1346_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1346_call_req_0;
      call_stmt_1346_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1346_call_req_1;
      call_stmt_1346_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1338_wire_constant & NOT_u4_u4_1341_wire_constant & register_index_1334 & type_cast_1344_wire_constant;
      rx_queue_pointer_32_1346 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1363_call 
    pushIntoQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1363_call_req_0;
      call_stmt_1363_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1363_call_req_1;
      call_stmt_1363_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_1_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1358_wire_constant & rx_queue_pointer_36_1352 & slice_1361_wire;
      push_status_1363 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    operator_delay_time_2931_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_1382_call_req_0;
      call_stmt_1382_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_1382_call_req_1;
      call_stmt_1382_call_ack_1<= update_ack(0);
      call_stmt_1382_call: delay_time_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        T => konst_1380_wire_constant,
        delay_done => status_1382,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end populateRxQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity pushIntoQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(35 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(35 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(35 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
    updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_call_data : out  std_logic_vector(99 downto 0);
    setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity pushIntoQueue;
architecture pushIntoQueue_arch of pushIntoQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 69)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal pushIntoQueue_CP_1321_start: Boolean;
  signal pushIntoQueue_CP_1321_symbol: Boolean;
  -- volatile/operator module components. 
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1217_call_req_0 : boolean;
  signal call_stmt_1217_call_ack_0 : boolean;
  signal call_stmt_1217_call_req_1 : boolean;
  signal call_stmt_1217_call_ack_1 : boolean;
  signal call_stmt_1225_call_req_0 : boolean;
  signal call_stmt_1225_call_ack_0 : boolean;
  signal call_stmt_1225_call_req_1 : boolean;
  signal call_stmt_1225_call_ack_1 : boolean;
  signal call_stmt_1228_call_req_0 : boolean;
  signal call_stmt_1228_call_ack_0 : boolean;
  signal call_stmt_1228_call_req_1 : boolean;
  signal call_stmt_1228_call_ack_1 : boolean;
  signal call_stmt_1231_call_req_0 : boolean;
  signal call_stmt_1231_call_ack_0 : boolean;
  signal call_stmt_1231_call_req_1 : boolean;
  signal call_stmt_1231_call_ack_1 : boolean;
  signal call_stmt_1262_call_req_0 : boolean;
  signal call_stmt_1262_call_ack_0 : boolean;
  signal call_stmt_1262_call_req_1 : boolean;
  signal call_stmt_1262_call_ack_1 : boolean;
  signal call_stmt_1267_call_req_0 : boolean;
  signal call_stmt_1267_call_ack_0 : boolean;
  signal call_stmt_1267_call_req_1 : boolean;
  signal call_stmt_1267_call_ack_1 : boolean;
  signal call_stmt_1274_call_req_0 : boolean;
  signal call_stmt_1274_call_ack_0 : boolean;
  signal call_stmt_1274_call_req_1 : boolean;
  signal call_stmt_1274_call_ack_1 : boolean;
  signal call_stmt_1278_call_req_0 : boolean;
  signal call_stmt_1278_call_ack_0 : boolean;
  signal call_stmt_1278_call_req_1 : boolean;
  signal call_stmt_1278_call_ack_1 : boolean;
  signal NOT_u1_u1_1281_inst_req_0 : boolean;
  signal NOT_u1_u1_1281_inst_ack_0 : boolean;
  signal NOT_u1_u1_1281_inst_req_1 : boolean;
  signal NOT_u1_u1_1281_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "pushIntoQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 69) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(68 downto 37) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(68 downto 37);
  in_buffer_data_in(tag_length + 68 downto 69) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 68 downto 69);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  pushIntoQueue_CP_1321_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "pushIntoQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1321_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1321_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1321_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  pushIntoQueue_CP_1321: Block -- control-path 
    signal pushIntoQueue_CP_1321_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    pushIntoQueue_CP_1321_elements(0) <= pushIntoQueue_CP_1321_start;
    pushIntoQueue_CP_1321_symbol <= pushIntoQueue_CP_1321_elements(22);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1217/$entry
      -- CP-element group 0: 	 call_stmt_1217/call_stmt_1217_sample_start_
      -- CP-element group 0: 	 call_stmt_1217/call_stmt_1217_update_start_
      -- CP-element group 0: 	 call_stmt_1217/call_stmt_1217_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1217/call_stmt_1217_Sample/crr
      -- CP-element group 0: 	 call_stmt_1217/call_stmt_1217_Update/$entry
      -- CP-element group 0: 	 call_stmt_1217/call_stmt_1217_Update/ccr
      -- 
    ccr_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(0), ack => call_stmt_1217_call_req_1); -- 
    crr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(0), ack => call_stmt_1217_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1217/call_stmt_1217_sample_completed_
      -- CP-element group 1: 	 call_stmt_1217/call_stmt_1217_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1217/call_stmt_1217_Sample/cra
      -- 
    cra_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1217_call_ack_0, ack => pushIntoQueue_CP_1321_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (26) 
      -- CP-element group 2: 	 call_stmt_1217/$exit
      -- CP-element group 2: 	 call_stmt_1217/call_stmt_1217_update_completed_
      -- CP-element group 2: 	 call_stmt_1217/call_stmt_1217_Update/$exit
      -- CP-element group 2: 	 call_stmt_1217/call_stmt_1217_Update/cca
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_sample_start_
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_update_start_
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Sample/crr
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Update/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Update/ccr
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_update_start_
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Update/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Update/ccr
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_update_start_
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Update/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Update/ccr
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_update_start_
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Update/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Update/ccr
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_update_start_
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Update/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Update/ccr
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_update_start_
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Update/$entry
      -- CP-element group 2: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Update/ccr
      -- 
    cca_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1217_call_ack_1, ack => pushIntoQueue_CP_1321_elements(2)); -- 
    crr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(2), ack => call_stmt_1225_call_req_0); -- 
    ccr_1356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(2), ack => call_stmt_1225_call_req_1); -- 
    ccr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(2), ack => call_stmt_1228_call_req_1); -- 
    ccr_1384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(2), ack => call_stmt_1231_call_req_1); -- 
    ccr_1398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(2), ack => call_stmt_1262_call_req_1); -- 
    ccr_1412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(2), ack => call_stmt_1267_call_req_1); -- 
    ccr_1426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(2), ack => call_stmt_1274_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_sample_completed_
      -- CP-element group 3: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Sample/$exit
      -- CP-element group 3: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Sample/cra
      -- 
    cra_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1225_call_ack_0, ack => pushIntoQueue_CP_1321_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	9 
    -- CP-element group 4: 	12 
    -- CP-element group 4: 	15 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_update_completed_
      -- CP-element group 4: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Update/$exit
      -- CP-element group 4: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1225_Update/cca
      -- CP-element group 4: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_sample_start_
      -- CP-element group 4: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Sample/crr
      -- 
    cca_1357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1225_call_ack_1, ack => pushIntoQueue_CP_1321_elements(4)); -- 
    crr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(4), ack => call_stmt_1228_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_sample_completed_
      -- CP-element group 5: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Sample/$exit
      -- CP-element group 5: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Sample/cra
      -- 
    cra_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1228_call_ack_0, ack => pushIntoQueue_CP_1321_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6: 	12 
    -- CP-element group 6: 	15 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_update_completed_
      -- CP-element group 6: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Update/$exit
      -- CP-element group 6: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1228_Update/cca
      -- CP-element group 6: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_sample_start_
      -- CP-element group 6: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Sample/crr
      -- 
    cca_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1228_call_ack_1, ack => pushIntoQueue_CP_1321_elements(6)); -- 
    crr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(6), ack => call_stmt_1231_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_sample_completed_
      -- CP-element group 7: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Sample/$exit
      -- CP-element group 7: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Sample/cra
      -- 
    cra_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1231_call_ack_0, ack => pushIntoQueue_CP_1321_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	15 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_update_completed_
      -- CP-element group 8: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Update/$exit
      -- CP-element group 8: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1231_Update/cca
      -- 
    cca_1385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1231_call_ack_1, ack => pushIntoQueue_CP_1321_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_sample_start_
      -- CP-element group 9: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Sample/$entry
      -- CP-element group 9: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Sample/crr
      -- 
    crr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(9), ack => call_stmt_1262_call_req_0); -- 
    pushIntoQueue_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "pushIntoQueue_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1321_elements(4) & pushIntoQueue_CP_1321_elements(6) & pushIntoQueue_CP_1321_elements(8);
      gj_pushIntoQueue_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1321_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_sample_completed_
      -- CP-element group 10: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Sample/$exit
      -- CP-element group 10: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Sample/cra
      -- 
    cra_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1262_call_ack_0, ack => pushIntoQueue_CP_1321_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_update_completed_
      -- CP-element group 11: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Update/$exit
      -- CP-element group 11: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1262_Update/cca
      -- 
    cca_1399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1262_call_ack_1, ack => pushIntoQueue_CP_1321_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	4 
    -- CP-element group 12: 	6 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_sample_start_
      -- CP-element group 12: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Sample/$entry
      -- CP-element group 12: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Sample/crr
      -- 
    crr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(12), ack => call_stmt_1267_call_req_0); -- 
    pushIntoQueue_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1321_elements(4) & pushIntoQueue_CP_1321_elements(6) & pushIntoQueue_CP_1321_elements(11);
      gj_pushIntoQueue_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1321_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_sample_completed_
      -- CP-element group 13: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Sample/$exit
      -- CP-element group 13: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Sample/cra
      -- 
    cra_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1267_call_ack_0, ack => pushIntoQueue_CP_1321_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_update_completed_
      -- CP-element group 14: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Update/$exit
      -- CP-element group 14: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1267_Update/cca
      -- 
    cca_1413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1267_call_ack_1, ack => pushIntoQueue_CP_1321_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	6 
    -- CP-element group 15: 	8 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_sample_start_
      -- CP-element group 15: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Sample/$entry
      -- CP-element group 15: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Sample/crr
      -- 
    crr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(15), ack => call_stmt_1274_call_req_0); -- 
    pushIntoQueue_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1321_elements(4) & pushIntoQueue_CP_1321_elements(6) & pushIntoQueue_CP_1321_elements(8) & pushIntoQueue_CP_1321_elements(14);
      gj_pushIntoQueue_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1321_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_sample_completed_
      -- CP-element group 16: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Sample/$exit
      -- CP-element group 16: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Sample/cra
      -- 
    cra_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1274_call_ack_0, ack => pushIntoQueue_CP_1321_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (17) 
      -- CP-element group 17: 	 call_stmt_1225_to_call_stmt_1274/$exit
      -- CP-element group 17: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_update_completed_
      -- CP-element group 17: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Update/$exit
      -- CP-element group 17: 	 call_stmt_1225_to_call_stmt_1274/call_stmt_1274_Update/cca
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/$entry
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_sample_start_
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_update_start_
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Sample/$entry
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Sample/crr
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Update/$entry
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Update/ccr
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_sample_start_
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_update_start_
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Sample/$entry
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Sample/rr
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Update/$entry
      -- CP-element group 17: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Update/cr
      -- 
    cca_1427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1274_call_ack_1, ack => pushIntoQueue_CP_1321_elements(17)); -- 
    crr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(17), ack => call_stmt_1278_call_req_0); -- 
    ccr_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(17), ack => call_stmt_1278_call_req_1); -- 
    rr_1452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(17), ack => NOT_u1_u1_1281_inst_req_0); -- 
    cr_1457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1321_elements(17), ack => NOT_u1_u1_1281_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_sample_completed_
      -- CP-element group 18: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Sample/$exit
      -- CP-element group 18: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Sample/cra
      -- 
    cra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1278_call_ack_0, ack => pushIntoQueue_CP_1321_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_update_completed_
      -- CP-element group 19: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Update/$exit
      -- CP-element group 19: 	 call_stmt_1278_to_assign_stmt_1282/call_stmt_1278_Update/cca
      -- 
    cca_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1278_call_ack_1, ack => pushIntoQueue_CP_1321_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_sample_completed_
      -- CP-element group 20: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Sample/$exit
      -- CP-element group 20: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Sample/ra
      -- 
    ra_1453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1281_inst_ack_0, ack => pushIntoQueue_CP_1321_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_update_completed_
      -- CP-element group 21: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Update/$exit
      -- CP-element group 21: 	 call_stmt_1278_to_assign_stmt_1282/NOT_u1_u1_1281_Update/ca
      -- 
    ca_1458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1281_inst_ack_1, ack => pushIntoQueue_CP_1321_elements(21)); -- 
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 $exit
      -- CP-element group 22: 	 call_stmt_1278_to_assign_stmt_1282/$exit
      -- 
    pushIntoQueue_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1321_elements(19) & pushIntoQueue_CP_1321_elements(21);
      gj_pushIntoQueue_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1321_elements(22), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1244_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1273_wire : std_logic_vector(31 downto 0);
    signal Queue_Length_1228 : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1236_wire : std_logic_vector(31 downto 0);
    signal konst_1235_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1241_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1243_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_1217 : std_logic_vector(0 downto 0);
    signal next_wi_1246 : std_logic_vector(31 downto 0);
    signal q_full_1251 : std_logic_vector(0 downto 0);
    signal read_index_1225 : std_logic_vector(31 downto 0);
    signal round_off_1238 : std_logic_vector(0 downto 0);
    signal total_msgs_1231 : std_logic_vector(31 downto 0);
    signal type_cast_1272_wire_constant : std_logic_vector(31 downto 0);
    signal write_index_1225 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_1235_wire_constant <= "00000000000000000000000000000001";
    konst_1241_wire_constant <= "00000000000000000000000000000000";
    konst_1243_wire_constant <= "00000000000000000000000000000001";
    type_cast_1272_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_1245_inst
    next_wi_1246 <= konst_1241_wire_constant when (round_off_1238(0) /=  '0') else ADD_u32_u32_1244_wire;
    -- binary operator ADD_u32_u32_1244_inst
    process(write_index_1225) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(write_index_1225, konst_1243_wire_constant, tmp_var);
      ADD_u32_u32_1244_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1273_inst
    process(total_msgs_1231) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(total_msgs_1231, type_cast_1272_wire_constant, tmp_var);
      ADD_u32_u32_1273_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1237_inst
    process(write_index_1225, SUB_u32_u32_1236_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_index_1225, SUB_u32_u32_1236_wire, tmp_var);
      round_off_1238 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1250_inst
    process(next_wi_1246, read_index_1225) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_wi_1246, read_index_1225, tmp_var);
      q_full_1251 <= tmp_var; --
    end process;
    -- shared split operator group (4) : NOT_u1_u1_1281_inst 
    ApIntNot_group_4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= q_full_1251;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1281_inst_req_0;
      NOT_u1_u1_1281_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1281_inst_req_1;
      NOT_u1_u1_1281_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_4_gI: SplitGuardInterface generic map(name => "ApIntNot_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator SUB_u32_u32_1236_inst
    process(Queue_Length_1228) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(Queue_Length_1228, konst_1235_wire_constant, tmp_var);
      SUB_u32_u32_1236_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1217_call 
    acquireLock_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1217_call_req_0;
      call_stmt_1217_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1217_call_req_1;
      call_stmt_1217_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_0_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_1217 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(35 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1225_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1225_call_req_0;
      call_stmt_1225_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1225_call_req_1;
      call_stmt_1225_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_index_1225 <= data_out(63 downto 32);
      read_index_1225 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1228_call 
    getQueueLength_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1228_call_req_0;
      call_stmt_1228_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1228_call_req_1;
      call_stmt_1228_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_2_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      Queue_Length_1228 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(35 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1231_call 
    getTotalMessages_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1231_call_req_0;
      call_stmt_1231_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1231_call_req_1;
      call_stmt_1231_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_3_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      total_msgs_1231 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(35 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1262_call 
    setQueueElement_call_group_4: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1262_call_req_0;
      call_stmt_1262_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1262_call_req_1;
      call_stmt_1262_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1251(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueueElement_call_group_4_gI: SplitGuardInterface generic map(name => "setQueueElement_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_index_1225 & q_w_data_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueueElement_call_reqs(0),
          ackR => setQueueElement_call_acks(0),
          dataR => setQueueElement_call_data(99 downto 0),
          tagR => setQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueueElement_return_acks(0), -- cross-over
          ackL => setQueueElement_return_reqs(0), -- cross-over
          tagL => setQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1267_call 
    setQueuePointers_call_group_5: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1267_call_req_0;
      call_stmt_1267_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1267_call_req_1;
      call_stmt_1267_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1251(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_5_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & next_wi_1246 & read_index_1225;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_1274_call 
    updateTotalMessages_call_group_6: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1274_call_req_0;
      call_stmt_1274_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1274_call_req_1;
      call_stmt_1274_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1251(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateTotalMessages_call_group_6_gI: SplitGuardInterface generic map(name => "updateTotalMessages_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & ADD_u32_u32_1273_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateTotalMessages_call_reqs(0),
          ackR => updateTotalMessages_call_acks(0),
          dataR => updateTotalMessages_call_data(67 downto 0),
          tagR => updateTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => updateTotalMessages_return_acks(0), -- cross-over
          ackL => updateTotalMessages_return_reqs(0), -- cross-over
          tagL => updateTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_1278_call 
    releaseLock_call_group_7: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1278_call_req_0;
      call_stmt_1278_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1278_call_req_1;
      call_stmt_1278_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_7_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(35 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- 
  end Block; -- data_path
  -- 
end pushIntoQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity releaseLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity releaseLock;
architecture releaseLock_arch of releaseLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal releaseLock_CP_714_start: Boolean;
  signal releaseLock_CP_714_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_888_call_ack_0 : boolean;
  signal call_stmt_888_call_ack_1 : boolean;
  signal call_stmt_888_call_req_1 : boolean;
  signal call_stmt_888_call_req_0 : boolean;
  signal call_stmt_770_call_ack_1 : boolean;
  signal call_stmt_770_call_req_1 : boolean;
  signal call_stmt_770_call_ack_0 : boolean;
  signal call_stmt_770_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "releaseLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  releaseLock_CP_714_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "releaseLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_714_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= releaseLock_CP_714_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_714_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  releaseLock_CP_714: Block -- control-path 
    signal releaseLock_CP_714_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    releaseLock_CP_714_elements(0) <= releaseLock_CP_714_start;
    releaseLock_CP_714_symbol <= releaseLock_CP_714_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Update/ccr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_update_start_
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/$entry
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_update_start_
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_sample_start_
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Update/$entry
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Update/ccr
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Update/$entry
      -- CP-element group 0: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Sample/crr
      -- 
    crr_727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_714_elements(0), ack => call_stmt_770_call_req_0); -- 
    ccr_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_714_elements(0), ack => call_stmt_770_call_req_1); -- 
    ccr_746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_714_elements(0), ack => call_stmt_888_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_sample_completed_
      -- CP-element group 1: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Sample/cra
      -- CP-element group 1: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Sample/$exit
      -- 
    cra_728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_770_call_ack_0, ack => releaseLock_CP_714_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_sample_start_
      -- CP-element group 2: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_update_completed_
      -- CP-element group 2: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Sample/crr
      -- CP-element group 2: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Update/cca
      -- CP-element group 2: 	 assign_stmt_758_to_call_stmt_888/call_stmt_770_Update/$exit
      -- 
    cca_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_770_call_ack_1, ack => releaseLock_CP_714_elements(2)); -- 
    crr_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_714_elements(2), ack => call_stmt_888_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Sample/cra
      -- CP-element group 3: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_sample_completed_
      -- CP-element group 3: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Sample/$exit
      -- 
    cra_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_888_call_ack_0, ack => releaseLock_CP_714_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Update/cca
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 assign_stmt_758_to_call_stmt_888/$exit
      -- CP-element group 4: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_update_completed_
      -- CP-element group 4: 	 assign_stmt_758_to_call_stmt_888/call_stmt_888_Update/$exit
      -- 
    cca_747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_888_call_ack_1, ack => releaseLock_CP_714_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_832_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_845_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_859_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_872_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_846_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_873_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u4_u36_884_wire : std_logic_vector(35 downto 0);
    signal MUX_825_wire : std_logic_vector(0 downto 0);
    signal MUX_831_wire : std_logic_vector(0 downto 0);
    signal MUX_838_wire : std_logic_vector(0 downto 0);
    signal MUX_844_wire : std_logic_vector(0 downto 0);
    signal MUX_852_wire : std_logic_vector(0 downto 0);
    signal MUX_858_wire : std_logic_vector(0 downto 0);
    signal MUX_865_wire : std_logic_vector(0 downto 0);
    signal MUX_871_wire : std_logic_vector(0 downto 0);
    signal NOT_u8_u8_765_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_888 : std_logic_vector(63 downto 0);
    signal konst_781_wire_constant : std_logic_vector(2 downto 0);
    signal konst_786_wire_constant : std_logic_vector(2 downto 0);
    signal konst_791_wire_constant : std_logic_vector(2 downto 0);
    signal konst_796_wire_constant : std_logic_vector(2 downto 0);
    signal konst_801_wire_constant : std_logic_vector(2 downto 0);
    signal konst_806_wire_constant : std_logic_vector(2 downto 0);
    signal konst_811_wire_constant : std_logic_vector(2 downto 0);
    signal konst_816_wire_constant : std_logic_vector(2 downto 0);
    signal lock_addr_32_774 : std_logic_vector(31 downto 0);
    signal lock_address_pointer_758 : std_logic_vector(35 downto 0);
    signal msg_size_plus_lock_770 : std_logic_vector(63 downto 0);
    signal new_bmask_875 : std_logic_vector(7 downto 0);
    signal s0_783 : std_logic_vector(0 downto 0);
    signal s1_788 : std_logic_vector(0 downto 0);
    signal s2_793 : std_logic_vector(0 downto 0);
    signal s3_798 : std_logic_vector(0 downto 0);
    signal s4_803 : std_logic_vector(0 downto 0);
    signal s5_808 : std_logic_vector(0 downto 0);
    signal s6_813 : std_logic_vector(0 downto 0);
    signal s7_818 : std_logic_vector(0 downto 0);
    signal sel_778 : std_logic_vector(2 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_762_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_768_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_822_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_828_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_830_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_835_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_837_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_841_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_843_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_849_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_851_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_855_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_857_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_862_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_864_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_868_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_877_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_879_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_882_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_765_wire_constant <= "11111111";
    konst_781_wire_constant <= "000";
    konst_786_wire_constant <= "001";
    konst_791_wire_constant <= "010";
    konst_796_wire_constant <= "011";
    konst_801_wire_constant <= "100";
    konst_806_wire_constant <= "101";
    konst_811_wire_constant <= "110";
    konst_816_wire_constant <= "111";
    type_cast_756_wire_constant <= "000000000000000000000000000000010000";
    type_cast_760_wire_constant <= "0";
    type_cast_762_wire_constant <= "1";
    type_cast_768_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_822_wire_constant <= "1";
    type_cast_824_wire_constant <= "0";
    type_cast_828_wire_constant <= "1";
    type_cast_830_wire_constant <= "0";
    type_cast_835_wire_constant <= "1";
    type_cast_837_wire_constant <= "0";
    type_cast_841_wire_constant <= "1";
    type_cast_843_wire_constant <= "0";
    type_cast_849_wire_constant <= "1";
    type_cast_851_wire_constant <= "0";
    type_cast_855_wire_constant <= "1";
    type_cast_857_wire_constant <= "0";
    type_cast_862_wire_constant <= "1";
    type_cast_864_wire_constant <= "0";
    type_cast_868_wire_constant <= "1";
    type_cast_870_wire_constant <= "0";
    type_cast_877_wire_constant <= "1";
    type_cast_879_wire_constant <= "0";
    type_cast_882_wire_constant <= "0000";
    type_cast_886_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_825_inst
    MUX_825_wire <= type_cast_822_wire_constant when (s0_783(0) /=  '0') else type_cast_824_wire_constant;
    -- flow-through select operator MUX_831_inst
    MUX_831_wire <= type_cast_828_wire_constant when (s1_788(0) /=  '0') else type_cast_830_wire_constant;
    -- flow-through select operator MUX_838_inst
    MUX_838_wire <= type_cast_835_wire_constant when (s2_793(0) /=  '0') else type_cast_837_wire_constant;
    -- flow-through select operator MUX_844_inst
    MUX_844_wire <= type_cast_841_wire_constant when (s3_798(0) /=  '0') else type_cast_843_wire_constant;
    -- flow-through select operator MUX_852_inst
    MUX_852_wire <= type_cast_849_wire_constant when (s4_803(0) /=  '0') else type_cast_851_wire_constant;
    -- flow-through select operator MUX_858_inst
    MUX_858_wire <= type_cast_855_wire_constant when (s5_808(0) /=  '0') else type_cast_857_wire_constant;
    -- flow-through select operator MUX_865_inst
    MUX_865_wire <= type_cast_862_wire_constant when (s6_813(0) /=  '0') else type_cast_864_wire_constant;
    -- flow-through select operator MUX_871_inst
    MUX_871_wire <= type_cast_868_wire_constant when (s7_818(0) /=  '0') else type_cast_870_wire_constant;
    -- flow-through slice operator slice_773_inst
    lock_addr_32_774 <= msg_size_plus_lock_770(31 downto 0);
    -- flow-through slice operator slice_777_inst
    sel_778 <= lock_addr_32_774(2 downto 0);
    -- binary operator ADD_u36_u36_757_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_756_wire_constant, tmp_var);
      lock_address_pointer_758 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_832_inst
    process(MUX_825_wire, MUX_831_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_825_wire, MUX_831_wire, tmp_var);
      CONCAT_u1_u2_832_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_845_inst
    process(MUX_838_wire, MUX_844_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_838_wire, MUX_844_wire, tmp_var);
      CONCAT_u1_u2_845_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_859_inst
    process(MUX_852_wire, MUX_858_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_852_wire, MUX_858_wire, tmp_var);
      CONCAT_u1_u2_859_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_872_inst
    process(MUX_865_wire, MUX_871_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_865_wire, MUX_871_wire, tmp_var);
      CONCAT_u1_u2_872_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_846_inst
    process(CONCAT_u1_u2_832_wire, CONCAT_u1_u2_845_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_832_wire, CONCAT_u1_u2_845_wire, tmp_var);
      CONCAT_u2_u4_846_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_873_inst
    process(CONCAT_u1_u2_859_wire, CONCAT_u1_u2_872_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_859_wire, CONCAT_u1_u2_872_wire, tmp_var);
      CONCAT_u2_u4_873_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_884_inst
    process(type_cast_882_wire_constant, lock_addr_32_774) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_882_wire_constant, lock_addr_32_774, tmp_var);
      CONCAT_u4_u36_884_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_874_inst
    process(CONCAT_u2_u4_846_wire, CONCAT_u2_u4_873_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_846_wire, CONCAT_u2_u4_873_wire, tmp_var);
      new_bmask_875 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_782_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_781_wire_constant, tmp_var);
      s0_783 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_787_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_786_wire_constant, tmp_var);
      s1_788 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_792_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_791_wire_constant, tmp_var);
      s2_793 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_797_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_796_wire_constant, tmp_var);
      s3_798 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_802_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_801_wire_constant, tmp_var);
      s4_803 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_807_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_806_wire_constant, tmp_var);
      s5_808 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_812_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_811_wire_constant, tmp_var);
      s6_813 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_817_inst
    process(sel_778) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_778, konst_816_wire_constant, tmp_var);
      s7_818 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_888_call call_stmt_770_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_888_call_req_0;
      reqL_unguarded(0) <= call_stmt_770_call_req_0;
      call_stmt_888_call_ack_0 <= ackL_unguarded(1);
      call_stmt_770_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_888_call_req_1;
      reqR_unguarded(0) <= call_stmt_770_call_req_1;
      call_stmt_888_call_ack_1 <= ackR_unguarded(1);
      call_stmt_770_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_877_wire_constant & type_cast_879_wire_constant & new_bmask_875 & CONCAT_u4_u36_884_wire & type_cast_886_wire_constant & type_cast_760_wire_constant & type_cast_762_wire_constant & NOT_u8_u8_765_wire_constant & lock_address_pointer_758 & type_cast_768_wire_constant;
      ignore_888 <= data_out(127 downto 64);
      msg_size_plus_lock_770 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end releaseLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    write_index : in  std_logic_vector(31 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueueElement;
architecture setQueueElement_arch of setQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal write_index_buffer :  std_logic_vector(31 downto 0);
  signal write_index_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal setQueueElement_CP_1301_start: Boolean;
  signal setQueueElement_CP_1301_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1207_call_req_0 : boolean;
  signal call_stmt_1207_call_ack_0 : boolean;
  signal call_stmt_1207_call_req_1 : boolean;
  signal call_stmt_1207_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= write_index;
  write_index_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueueElement_CP_1301_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1301_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueueElement_CP_1301_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1301_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueueElement_CP_1301: Block -- control-path 
    signal setQueueElement_CP_1301_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueueElement_CP_1301_elements(0) <= setQueueElement_CP_1301_start;
    setQueueElement_CP_1301_symbol <= setQueueElement_CP_1301_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1151_to_call_stmt_1207/$entry
      -- CP-element group 0: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_sample_start_
      -- CP-element group 0: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_update_start_
      -- CP-element group 0: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Update/ccr
      -- 
    crr_1314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1301_elements(0), ack => call_stmt_1207_call_req_0); -- 
    ccr_1319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1301_elements(0), ack => call_stmt_1207_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Sample/cra
      -- 
    cra_1315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1207_call_ack_0, ack => setQueueElement_CP_1301_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1151_to_call_stmt_1207/$exit
      -- CP-element group 2: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_update_completed_
      -- CP-element group 2: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1151_to_call_stmt_1207/call_stmt_1207_Update/cca
      -- 
    cca_1320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1207_call_ack_1, ack => setQueueElement_CP_1301_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1165_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1183_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_1158_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u32_u64_1187_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1191_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_1171_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_1177_wire_constant : std_logic_vector(7 downto 0);
    signal bmask_1179 : std_logic_vector(7 downto 0);
    signal buffer_address_1151 : std_logic_vector(35 downto 0);
    signal element_pair_address_1161 : std_logic_vector(35 downto 0);
    signal ignore_1207 : std_logic_vector(63 downto 0);
    signal konst_1164_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1182_wire_constant : std_logic_vector(31 downto 0);
    signal slice_1155_wire : std_logic_vector(30 downto 0);
    signal type_cast_1149_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_1157_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_1159_wire : std_logic_vector(35 downto 0);
    signal type_cast_1185_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1190_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1200_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1202_wire_constant : std_logic_vector(0 downto 0);
    signal wval_1193 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_1171_wire_constant <= "00001111";
    CONCAT_u4_u8_1177_wire_constant <= "11110000";
    konst_1164_wire_constant <= "00000000000000000000000000000000";
    konst_1182_wire_constant <= "00000000000000000000000000000000";
    type_cast_1149_wire_constant <= "000000000000000000000000000000011000";
    type_cast_1157_wire_constant <= "000";
    type_cast_1185_wire_constant <= "00000000000000000000000000000000";
    type_cast_1190_wire_constant <= "00000000000000000000000000000000";
    type_cast_1200_wire_constant <= "0";
    type_cast_1202_wire_constant <= "0";
    -- flow-through select operator MUX_1178_inst
    bmask_1179 <= CONCAT_u4_u8_1171_wire_constant when (BITSEL_u32_u1_1165_wire(0) /=  '0') else CONCAT_u4_u8_1177_wire_constant;
    -- flow-through select operator MUX_1192_inst
    wval_1193 <= CONCAT_u32_u64_1187_wire when (BITSEL_u32_u1_1183_wire(0) /=  '0') else CONCAT_u32_u64_1191_wire;
    -- flow-through slice operator slice_1155_inst
    slice_1155_wire <= write_index_buffer(31 downto 1);
    -- interlock type_cast_1159_inst
    process(CONCAT_u31_u34_1158_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_1158_wire(33 downto 0);
      type_cast_1159_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_1150_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_1149_wire_constant, tmp_var);
      buffer_address_1151 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_1160_inst
    process(buffer_address_1151, type_cast_1159_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_1151, type_cast_1159_wire, tmp_var);
      element_pair_address_1161 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1165_inst
    process(write_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_index_buffer, konst_1164_wire_constant, tmp_var);
      BITSEL_u32_u1_1165_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1183_inst
    process(write_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_index_buffer, konst_1182_wire_constant, tmp_var);
      BITSEL_u32_u1_1183_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_1158_inst
    process(slice_1155_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1155_wire, type_cast_1157_wire_constant, tmp_var);
      CONCAT_u31_u34_1158_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_1187_inst
    process(type_cast_1185_wire_constant, q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1185_wire_constant, q_w_data_buffer, tmp_var);
      CONCAT_u32_u64_1187_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_1191_inst
    process(q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(q_w_data_buffer, type_cast_1190_wire_constant, tmp_var);
      CONCAT_u32_u64_1191_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1207_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1207_call_req_0;
      call_stmt_1207_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1207_call_req_1;
      call_stmt_1207_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1200_wire_constant & type_cast_1202_wire_constant & bmask_1179 & element_pair_address_1161 & wval_1193;
      ignore_1207 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : in  std_logic_vector(31 downto 0);
    rp : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueuePointers;
architecture setQueuePointers_arch of setQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  -- output port buffer signals
  signal setQueuePointers_CP_660_start: Boolean;
  signal setQueuePointers_CP_660_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_710_call_req_0 : boolean;
  signal call_stmt_710_call_ack_0 : boolean;
  signal call_stmt_710_call_req_1 : boolean;
  signal call_stmt_710_call_ack_1 : boolean;
  signal call_stmt_728_call_req_0 : boolean;
  signal call_stmt_728_call_ack_0 : boolean;
  signal call_stmt_728_call_req_1 : boolean;
  signal call_stmt_728_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= wp;
  wp_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= rp;
  rp_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueuePointers_CP_660_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_660_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueuePointers_CP_660_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_660_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueuePointers_CP_660: Block -- control-path 
    signal setQueuePointers_CP_660_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    setQueuePointers_CP_660_elements(0) <= setQueuePointers_CP_660_start;
    setQueuePointers_CP_660_symbol <= setQueuePointers_CP_660_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/$entry
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_sample_start_
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_update_start_
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Sample/$entry
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Sample/crr
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Update/$entry
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Update/ccr
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_update_start_
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Update/$entry
      -- CP-element group 0: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Update/ccr
      -- 
    crr_673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_660_elements(0), ack => call_stmt_710_call_req_0); -- 
    ccr_678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_660_elements(0), ack => call_stmt_710_call_req_1); -- 
    ccr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_660_elements(0), ack => call_stmt_728_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_sample_completed_
      -- CP-element group 1: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Sample/$exit
      -- CP-element group 1: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Sample/cra
      -- 
    cra_674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_0, ack => setQueuePointers_CP_660_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_update_completed_
      -- CP-element group 2: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Update/$exit
      -- CP-element group 2: 	 call_stmt_710_to_call_stmt_728/call_stmt_710_Update/cca
      -- CP-element group 2: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_sample_start_
      -- CP-element group 2: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Sample/$entry
      -- CP-element group 2: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Sample/crr
      -- 
    cca_679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_1, ack => setQueuePointers_CP_660_elements(2)); -- 
    crr_687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_660_elements(2), ack => call_stmt_728_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_sample_completed_
      -- CP-element group 3: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Sample/$exit
      -- CP-element group 3: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Sample/cra
      -- 
    cra_688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_728_call_ack_0, ack => setQueuePointers_CP_660_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_710_to_call_stmt_728/$exit
      -- CP-element group 4: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_update_completed_
      -- CP-element group 4: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Update/$exit
      -- CP-element group 4: 	 call_stmt_710_to_call_stmt_728/call_stmt_728_Update/cca
      -- 
    cca_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_728_call_ack_1, ack => setQueuePointers_CP_660_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_723_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u32_u64_708_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_726_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_704_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_720_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_1_728 : std_logic_vector(63 downto 0);
    signal ignore_710 : std_logic_vector(63 downto 0);
    signal konst_722_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_696_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_712_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_714_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_704_wire_constant <= "00001111";
    CONCAT_u4_u8_720_wire_constant <= "11110000";
    konst_722_wire_constant <= "000000000000000000000000000000001000";
    type_cast_696_wire_constant <= "0";
    type_cast_698_wire_constant <= "0";
    type_cast_712_wire_constant <= "0";
    type_cast_714_wire_constant <= "0";
    -- binary operator ADD_u36_u36_723_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_722_wire_constant, tmp_var);
      ADD_u36_u36_723_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_708_inst
    process(rp_buffer, rp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(rp_buffer, rp_buffer, tmp_var);
      CONCAT_u32_u64_708_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_726_inst
    process(wp_buffer, wp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(wp_buffer, wp_buffer, tmp_var);
      CONCAT_u32_u64_726_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_728_call call_stmt_710_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_728_call_req_0;
      reqL_unguarded(0) <= call_stmt_710_call_req_0;
      call_stmt_728_call_ack_0 <= ackL_unguarded(1);
      call_stmt_710_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_728_call_req_1;
      reqR_unguarded(0) <= call_stmt_710_call_req_1;
      call_stmt_728_call_ack_1 <= ackR_unguarded(1);
      call_stmt_710_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_712_wire_constant & type_cast_714_wire_constant & CONCAT_u4_u8_720_wire_constant & ADD_u36_u36_723_wire & CONCAT_u32_u64_726_wire & type_cast_696_wire_constant & type_cast_698_wire_constant & CONCAT_u4_u8_704_wire_constant & q_base_address_buffer & CONCAT_u32_u64_708_wire;
      ignore_1_728 <= data_out(127 downto 64);
      ignore_710 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
    getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
    getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
    transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_call_data : out  std_logic_vector(31 downto 0);
    transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
    transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_return_data : in   std_logic_vector(0 downto 0);
    transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitEngineDaemon;
architecture transmitEngineDaemon_arch of transmitEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal transmitEngineDaemon_CP_3465_start: Boolean;
  signal transmitEngineDaemon_CP_3465_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_req_1 : boolean;
  signal if_stmt_2038_branch_req_0 : boolean;
  signal if_stmt_2038_branch_ack_1 : boolean;
  signal if_stmt_2038_branch_ack_0 : boolean;
  signal do_while_stmt_2046_branch_req_0 : boolean;
  signal AND_u6_u6_2057_inst_req_0 : boolean;
  signal AND_u6_u6_2057_inst_ack_0 : boolean;
  signal AND_u6_u6_2057_inst_req_1 : boolean;
  signal AND_u6_u6_2057_inst_ack_1 : boolean;
  signal phi_stmt_2058_req_0 : boolean;
  signal phi_stmt_2058_req_1 : boolean;
  signal phi_stmt_2058_ack_0 : boolean;
  signal ncount_2132_2060_buf_req_0 : boolean;
  signal ncount_2132_2060_buf_ack_0 : boolean;
  signal ncount_2132_2060_buf_req_1 : boolean;
  signal ncount_2132_2060_buf_ack_1 : boolean;
  signal call_stmt_2069_call_req_0 : boolean;
  signal call_stmt_2069_call_ack_0 : boolean;
  signal call_stmt_2069_call_req_1 : boolean;
  signal call_stmt_2069_call_ack_1 : boolean;
  signal call_stmt_2073_call_req_0 : boolean;
  signal call_stmt_2073_call_ack_0 : boolean;
  signal call_stmt_2073_call_req_1 : boolean;
  signal call_stmt_2073_call_ack_1 : boolean;
  signal NOT_u1_u1_2083_inst_req_0 : boolean;
  signal NOT_u1_u1_2083_inst_ack_0 : boolean;
  signal NOT_u1_u1_2083_inst_req_1 : boolean;
  signal NOT_u1_u1_2083_inst_ack_1 : boolean;
  signal W_pkt_pointer_2078_delayed_4_0_2093_inst_req_0 : boolean;
  signal W_pkt_pointer_2078_delayed_4_0_2093_inst_ack_0 : boolean;
  signal W_pkt_pointer_2078_delayed_4_0_2093_inst_req_1 : boolean;
  signal W_pkt_pointer_2078_delayed_4_0_2093_inst_ack_1 : boolean;
  signal call_stmt_2102_call_req_0 : boolean;
  signal call_stmt_2102_call_ack_0 : boolean;
  signal call_stmt_2102_call_req_1 : boolean;
  signal call_stmt_2102_call_ack_1 : boolean;
  signal W_count_2091_delayed_14_0_2106_inst_req_0 : boolean;
  signal W_count_2091_delayed_14_0_2106_inst_ack_0 : boolean;
  signal W_count_2091_delayed_14_0_2106_inst_req_1 : boolean;
  signal W_count_2091_delayed_14_0_2106_inst_ack_1 : boolean;
  signal call_stmt_2118_call_req_0 : boolean;
  signal call_stmt_2118_call_ack_0 : boolean;
  signal call_stmt_2118_call_req_1 : boolean;
  signal call_stmt_2118_call_ack_1 : boolean;
  signal W_count_2099_delayed_14_0_2119_inst_req_0 : boolean;
  signal W_count_2099_delayed_14_0_2119_inst_ack_0 : boolean;
  signal W_count_2099_delayed_14_0_2119_inst_req_1 : boolean;
  signal W_count_2099_delayed_14_0_2119_inst_ack_1 : boolean;
  signal ADD_u32_u32_2125_inst_req_0 : boolean;
  signal ADD_u32_u32_2125_inst_ack_0 : boolean;
  signal ADD_u32_u32_2125_inst_req_1 : boolean;
  signal ADD_u32_u32_2125_inst_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_ack_1 : boolean;
  signal do_while_stmt_2046_branch_ack_0 : boolean;
  signal do_while_stmt_2046_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitEngineDaemon_CP_3465_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3465_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3465_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3465_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitEngineDaemon_CP_3465: Block -- control-path 
    signal transmitEngineDaemon_CP_3465_elements: BooleanArray(86 downto 0);
    -- 
  begin -- 
    transmitEngineDaemon_CP_3465_elements(0) <= transmitEngineDaemon_CP_3465_start;
    transmitEngineDaemon_CP_3465_symbol <= transmitEngineDaemon_CP_3465_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_sample_start_
      -- CP-element group 0: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Sample/req
      -- CP-element group 0: 	 assign_stmt_2035/$entry
      -- 
    req_3478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(0), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Sample/ack
      -- CP-element group 1: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_update_start_
      -- CP-element group 1: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_sample_completed_
      -- CP-element group 1: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Update/$entry
      -- CP-element group 1: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Update/req
      -- 
    ack_3479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(1)); -- 
    req_3483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(1), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	86 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 branch_block_stmt_2036/merge_stmt_2037__entry__
      -- CP-element group 2: 	 branch_block_stmt_2036/branch_block_stmt_2036__entry__
      -- CP-element group 2: 	 branch_block_stmt_2036/$entry
      -- CP-element group 2: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Update/ack
      -- CP-element group 2: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_update_completed_
      -- CP-element group 2: 	 assign_stmt_2035/WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_Update/$exit
      -- CP-element group 2: 	 assign_stmt_2035/$exit
      -- CP-element group 2: 	 branch_block_stmt_2036/merge_stmt_2037_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_2036/merge_stmt_2037__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_2036/merge_stmt_2037__entry___PhiReq/$exit
      -- 
    ack_3484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_2036/branch_block_stmt_2036__exit__
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_2036/$exit
      -- 
    transmitEngineDaemon_CP_3465_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	85 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	86 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_2036/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_2036/do_while_stmt_2046__exit__
      -- CP-element group 4: 	 branch_block_stmt_2036/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_2036/disable_loopback_PhiReq/$exit
      -- 
    transmitEngineDaemon_CP_3465_elements(4) <= transmitEngineDaemon_CP_3465_elements(85);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	86 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	86 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_2036/if_stmt_2038_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_2036/if_stmt_2038_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_2036/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_2036/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_2036/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_3557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2038_branch_ack_1, ack => transmitEngineDaemon_CP_3465_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	86 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_2036/do_while_stmt_2046__entry__
      -- CP-element group 6: 	 branch_block_stmt_2036/if_stmt_2038__exit__
      -- CP-element group 6: 	 branch_block_stmt_2036/if_stmt_2038_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_2036/if_stmt_2038_else_link/else_choice_transition
      -- 
    else_choice_transition_3561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2038_branch_ack_0, ack => transmitEngineDaemon_CP_3465_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_2036/do_while_stmt_2046/$entry
      -- CP-element group 7: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046__entry__
      -- 
    transmitEngineDaemon_CP_3465_elements(7) <= transmitEngineDaemon_CP_3465_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	85 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046__exit__
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_back
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	83 
    -- CP-element group 10: 	84 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2036/do_while_stmt_2046/condition_done
      -- CP-element group 10: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_taken/$entry
      -- 
    transmitEngineDaemon_CP_3465_elements(10) <= transmitEngineDaemon_CP_3465_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	82 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_body_done
      -- 
    transmitEngineDaemon_CP_3465_elements(11) <= transmitEngineDaemon_CP_3465_elements(82);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/back_edge_to_loop_body
      -- 
    transmitEngineDaemon_CP_3465_elements(12) <= transmitEngineDaemon_CP_3465_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	31 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/first_time_through_loop_body
      -- 
    transmitEngineDaemon_CP_3465_elements(13) <= transmitEngineDaemon_CP_3465_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	25 
    -- CP-element group 14: 	26 
    -- CP-element group 14: 	81 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2048_sample_start_
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	81 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/condition_evaluated
      -- 
    condition_evaluated_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(15), ack => do_while_stmt_2046_branch_req_0); -- 
    transmitEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(19) & transmitEngineDaemon_CP_3465_elements(81);
      gj_transmitEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	25 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_sample_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(14) & transmitEngineDaemon_CP_3465_elements(25) & transmitEngineDaemon_CP_3465_elements(19);
      gj_transmitEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	23 
    -- CP-element group 17: 	27 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	47 
    -- CP-element group 17: 	51 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	75 
    -- CP-element group 17: 	82 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	25 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2048_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_sample_completed_
      -- 
    transmitEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(23) & transmitEngineDaemon_CP_3465_elements(27);
      gj_transmitEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	26 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_update_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(20) & transmitEngineDaemon_CP_3465_elements(26);
      gj_transmitEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	28 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/aggregated_phi_update_ack
      -- 
    transmitEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(24) & transmitEngineDaemon_CP_3465_elements(28);
      gj_transmitEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	44 
    -- CP-element group 20: 	79 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2048_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(14) & transmitEngineDaemon_CP_3465_elements(44) & transmitEngineDaemon_CP_3465_elements(79);
      gj_transmitEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Sample/rr
      -- 
    rr_3594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(21), ack => AND_u6_u6_2057_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(16) & transmitEngineDaemon_CP_3465_elements(23);
      gj_transmitEngineDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_update_start_
      -- CP-element group 22: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Update/cr
      -- 
    cr_3599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(22), ack => AND_u6_u6_2057_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(18) & transmitEngineDaemon_CP_3465_elements(24);
      gj_transmitEngineDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Sample/ra
      -- 
    ra_3595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_2057_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	42 
    -- CP-element group 24: 	78 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2048_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/AND_u6_u6_2057_Update/ca
      -- 
    ca_3600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_2057_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(24)); -- 
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	14 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	17 
    -- CP-element group 25: 	49 
    -- CP-element group 25: 	53 
    -- CP-element group 25: 	73 
    -- CP-element group 25: 	77 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	16 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_sample_start_
      -- 
    transmitEngineDaemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(14) & transmitEngineDaemon_CP_3465_elements(17) & transmitEngineDaemon_CP_3465_elements(49) & transmitEngineDaemon_CP_3465_elements(53) & transmitEngineDaemon_CP_3465_elements(73) & transmitEngineDaemon_CP_3465_elements(77);
      gj_transmitEngineDaemon_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	64 
    -- CP-element group 26: 	72 
    -- CP-element group 26: 	76 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	18 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(14) & transmitEngineDaemon_CP_3465_elements(64) & transmitEngineDaemon_CP_3465_elements(72) & transmitEngineDaemon_CP_3465_elements(76);
      gj_transmitEngineDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	17 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_sample_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	19 
    -- CP-element group 28: 	62 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_update_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	12 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_loopback_trigger
      -- 
    transmitEngineDaemon_CP_3465_elements(29) <= transmitEngineDaemon_CP_3465_elements(12);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_loopback_sample_req
      -- CP-element group 30: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_loopback_sample_req_ps
      -- 
    phi_stmt_2058_loopback_sample_req_3610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2058_loopback_sample_req_3610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(30), ack => phi_stmt_2058_req_0); -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(30) is bound as output of CP function.
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	13 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_entry_trigger
      -- 
    transmitEngineDaemon_CP_3465_elements(31) <= transmitEngineDaemon_CP_3465_elements(13);
    -- CP-element group 32:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_entry_sample_req
      -- CP-element group 32: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_entry_sample_req_ps
      -- 
    phi_stmt_2058_entry_sample_req_3613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2058_entry_sample_req_3613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(32), ack => phi_stmt_2058_req_1); -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_phi_mux_ack
      -- CP-element group 33: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/phi_stmt_2058_phi_mux_ack_ps
      -- 
    phi_stmt_2058_phi_mux_ack_3616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2058_ack_0, ack => transmitEngineDaemon_CP_3465_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Sample/req
      -- 
    req_3629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(34), ack => ncount_2132_2060_buf_req_0); -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_update_start_
      -- CP-element group 35: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Update/req
      -- 
    req_3634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(35), ack => ncount_2132_2060_buf_req_1); -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Sample/ack
      -- 
    ack_3630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_2132_2060_buf_ack_0, ack => transmitEngineDaemon_CP_3465_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/R_ncount_2060_Update/ack
      -- 
    ack_3635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_2132_2060_buf_ack_1, ack => transmitEngineDaemon_CP_3465_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_sample_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_update_start_
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_update_completed__ps
      -- 
    transmitEngineDaemon_CP_3465_elements(40) <= transmitEngineDaemon_CP_3465_elements(41);
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	40 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/type_cast_2062_update_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3465_elements(39), ack => transmitEngineDaemon_CP_3465_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	24 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	69 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Sample/crr
      -- 
    crr_3652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(42), ack => call_stmt_2069_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(24) & transmitEngineDaemon_CP_3465_elements(44) & transmitEngineDaemon_CP_3465_elements(61) & transmitEngineDaemon_CP_3465_elements(69);
      gj_transmitEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	48 
    -- CP-element group 43: 	52 
    -- CP-element group 43: 	56 
    -- CP-element group 43: 	61 
    -- CP-element group 43: 	69 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_update_start_
      -- CP-element group 43: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Update/ccr
      -- 
    ccr_3657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(43), ack => call_stmt_2069_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(48) & transmitEngineDaemon_CP_3465_elements(52) & transmitEngineDaemon_CP_3465_elements(56) & transmitEngineDaemon_CP_3465_elements(61) & transmitEngineDaemon_CP_3465_elements(69);
      gj_transmitEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	20 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Sample/cra
      -- 
    cra_3653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2069_call_ack_0, ack => transmitEngineDaemon_CP_3465_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	50 
    -- CP-element group 45: 	54 
    -- CP-element group 45: 	66 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2069_Update/cca
      -- 
    cca_3658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2069_call_ack_1, ack => transmitEngineDaemon_CP_3465_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Sample/crr
      -- 
    crr_3666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(46), ack => call_stmt_2073_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(45) & transmitEngineDaemon_CP_3465_elements(48);
      gj_transmitEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	17 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	60 
    -- CP-element group 47: 	68 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_update_start_
      -- CP-element group 47: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Update/ccr
      -- 
    ccr_3671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(47), ack => call_stmt_2073_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(17) & transmitEngineDaemon_CP_3465_elements(60) & transmitEngineDaemon_CP_3465_elements(68);
      gj_transmitEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Sample/cra
      -- 
    cra_3667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2073_call_ack_0, ack => transmitEngineDaemon_CP_3465_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49: 	66 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	25 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2073_Update/cca
      -- 
    cca_3672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2073_call_ack_1, ack => transmitEngineDaemon_CP_3465_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Sample/rr
      -- 
    rr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(50), ack => NOT_u1_u1_2083_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(45) & transmitEngineDaemon_CP_3465_elements(52);
      gj_transmitEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	17 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	60 
    -- CP-element group 51: 	68 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_update_start_
      -- CP-element group 51: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Update/cr
      -- 
    cr_3685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(51), ack => NOT_u1_u1_2083_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(17) & transmitEngineDaemon_CP_3465_elements(60) & transmitEngineDaemon_CP_3465_elements(68);
      gj_transmitEngineDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	43 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Sample/ra
      -- 
    ra_3681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_2083_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	58 
    -- CP-element group 53: 	66 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	25 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/NOT_u1_u1_2083_Update/ca
      -- 
    ca_3686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_2083_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	45 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Sample/req
      -- 
    req_3694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(54), ack => W_pkt_pointer_2078_delayed_4_0_2093_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(45) & transmitEngineDaemon_CP_3465_elements(56);
      gj_transmitEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	60 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_update_start_
      -- CP-element group 55: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Update/req
      -- 
    req_3699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(55), ack => W_pkt_pointer_2078_delayed_4_0_2093_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3465_elements(60);
      gj_transmitEngineDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Sample/ack
      -- 
    ack_3695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_2078_delayed_4_0_2093_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2095_Update/ack
      -- 
    ack_3700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_2078_delayed_4_0_2093_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	57 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Sample/crr
      -- 
    crr_3708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(58), ack => call_stmt_2102_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(49) & transmitEngineDaemon_CP_3465_elements(53) & transmitEngineDaemon_CP_3465_elements(57) & transmitEngineDaemon_CP_3465_elements(60);
      gj_transmitEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_update_start_
      -- CP-element group 59: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Update/ccr
      -- 
    ccr_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(59), ack => call_stmt_2102_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3465_elements(61);
      gj_transmitEngineDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	47 
    -- CP-element group 60: 	51 
    -- CP-element group 60: 	55 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Sample/cra
      -- 
    cra_3709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2102_call_ack_0, ack => transmitEngineDaemon_CP_3465_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	82 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	42 
    -- CP-element group 61: 	43 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2102_Update/cca
      -- 
    cca_3714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2102_call_ack_1, ack => transmitEngineDaemon_CP_3465_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	28 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Sample/req
      -- 
    req_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(62), ack => W_count_2091_delayed_14_0_2106_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(28) & transmitEngineDaemon_CP_3465_elements(64);
      gj_transmitEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_update_start_
      -- CP-element group 63: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Update/req
      -- 
    req_3727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(63), ack => W_count_2091_delayed_14_0_2106_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3465_elements(68);
      gj_transmitEngineDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	26 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Sample/ack
      -- 
    ack_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2091_delayed_14_0_2106_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2108_Update/ack
      -- 
    ack_3728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2091_delayed_14_0_2106_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	45 
    -- CP-element group 66: 	49 
    -- CP-element group 66: 	53 
    -- CP-element group 66: 	65 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Sample/crr
      -- 
    crr_3736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(66), ack => call_stmt_2118_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(45) & transmitEngineDaemon_CP_3465_elements(49) & transmitEngineDaemon_CP_3465_elements(53) & transmitEngineDaemon_CP_3465_elements(65) & transmitEngineDaemon_CP_3465_elements(68);
      gj_transmitEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_update_start_
      -- CP-element group 67: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Update/ccr
      -- 
    ccr_3741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(67), ack => call_stmt_2118_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3465_elements(69);
      gj_transmitEngineDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	47 
    -- CP-element group 68: 	51 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Sample/cra
      -- 
    cra_3737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2118_call_ack_0, ack => transmitEngineDaemon_CP_3465_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	82 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	42 
    -- CP-element group 69: 	43 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/call_stmt_2118_Update/cca
      -- 
    cca_3742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2118_call_ack_1, ack => transmitEngineDaemon_CP_3465_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	28 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Sample/req
      -- 
    req_3750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(70), ack => W_count_2099_delayed_14_0_2119_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(28) & transmitEngineDaemon_CP_3465_elements(72);
      gj_transmitEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	17 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_update_start_
      -- CP-element group 71: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Update/req
      -- 
    req_3755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(71), ack => W_count_2099_delayed_14_0_2119_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(17) & transmitEngineDaemon_CP_3465_elements(73);
      gj_transmitEngineDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	26 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Sample/ack
      -- 
    ack_3751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2099_delayed_14_0_2119_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	82 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	25 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/assign_stmt_2121_Update/ack
      -- 
    ack_3756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_2099_delayed_14_0_2119_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Sample/rr
      -- 
    rr_3764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(74), ack => ADD_u32_u32_2125_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(28) & transmitEngineDaemon_CP_3465_elements(76);
      gj_transmitEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_update_start_
      -- CP-element group 75: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Update/cr
      -- 
    cr_3769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(75), ack => ADD_u32_u32_2125_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(17) & transmitEngineDaemon_CP_3465_elements(77);
      gj_transmitEngineDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	26 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Sample/ra
      -- 
    ra_3765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2125_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	82 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	25 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/ADD_u32_u32_2125_Update/ca
      -- 
    ca_3770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_2125_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	24 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Sample/req
      -- 
    req_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(78), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(24) & transmitEngineDaemon_CP_3465_elements(80);
      gj_transmitEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	20 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_update_start_
      -- CP-element group 79: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Sample/ack
      -- CP-element group 79: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Update/req
      -- 
    ack_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_ack_0, ack => transmitEngineDaemon_CP_3465_elements(79)); -- 
    req_3783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(79), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_Update/ack
      -- 
    ack_3784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_ack_1, ack => transmitEngineDaemon_CP_3465_elements(80)); -- 
    -- CP-element group 81:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	15 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitEngineDaemon_CP_3465_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3465_elements(14), ack => transmitEngineDaemon_CP_3465_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  join  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	17 
    -- CP-element group 82: 	61 
    -- CP-element group 82: 	69 
    -- CP-element group 82: 	73 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	11 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2036/do_while_stmt_2046/do_while_stmt_2046_loop_body/$exit
      -- 
    transmitEngineDaemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3465_elements(17) & transmitEngineDaemon_CP_3465_elements(61) & transmitEngineDaemon_CP_3465_elements(69) & transmitEngineDaemon_CP_3465_elements(73) & transmitEngineDaemon_CP_3465_elements(77) & transmitEngineDaemon_CP_3465_elements(80);
      gj_transmitEngineDaemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	10 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_exit/$exit
      -- CP-element group 83: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_exit/ack
      -- 
    ack_3789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2046_branch_ack_0, ack => transmitEngineDaemon_CP_3465_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	10 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_taken/$exit
      -- CP-element group 84: 	 branch_block_stmt_2036/do_while_stmt_2046/loop_taken/ack
      -- 
    ack_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2046_branch_ack_1, ack => transmitEngineDaemon_CP_3465_elements(84)); -- 
    -- CP-element group 85:  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	4 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2036/do_while_stmt_2046/$exit
      -- 
    transmitEngineDaemon_CP_3465_elements(85) <= transmitEngineDaemon_CP_3465_elements(8);
    -- CP-element group 86:  merge  branch  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	2 
    -- CP-element group 86: 	5 
    -- CP-element group 86: 	4 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	5 
    -- CP-element group 86: 	6 
    -- CP-element group 86:  members (49) 
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038__entry__
      -- CP-element group 86: 	 branch_block_stmt_2036/merge_stmt_2037__exit__
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Sample/req
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Sample/ack
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Update/req
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/BITSEL_u32_u1_2041_inputs/RPIPE_CONTROL_REGISTER_2039/Update/ack
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/BITSEL_u32_u1_2041/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/NOT_u1_u1_2042/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_2036/NOT_u1_u1_2042_place
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/if_stmt_2038_else_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/merge_stmt_2037_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_2036/merge_stmt_2037_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_2036/merge_stmt_2037_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_2036/merge_stmt_2037_PhiAck/dummy
      -- 
    branch_req_3552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3465_elements(86), ack => if_stmt_2038_branch_req_0); -- 
    transmitEngineDaemon_CP_3465_elements(86) <= OrReduce(transmitEngineDaemon_CP_3465_elements(2) & transmitEngineDaemon_CP_3465_elements(5) & transmitEngineDaemon_CP_3465_elements(4));
    transmitEngineDaemon_do_while_stmt_2046_terminator_3794: loop_terminator -- 
      generic map (name => " transmitEngineDaemon_do_while_stmt_2046_terminator_3794", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitEngineDaemon_CP_3465_elements(11),loop_continue => transmitEngineDaemon_CP_3465_elements(84),loop_terminate => transmitEngineDaemon_CP_3465_elements(83),loop_back => transmitEngineDaemon_CP_3465_elements(9),loop_exit => transmitEngineDaemon_CP_3465_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_2058_phi_seq_3644_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitEngineDaemon_CP_3465_elements(29);
      transmitEngineDaemon_CP_3465_elements(34)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitEngineDaemon_CP_3465_elements(36);
      transmitEngineDaemon_CP_3465_elements(35)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitEngineDaemon_CP_3465_elements(37);
      transmitEngineDaemon_CP_3465_elements(30) <= phi_mux_reqs(0);
      triggers(1)  <= transmitEngineDaemon_CP_3465_elements(31);
      transmitEngineDaemon_CP_3465_elements(38)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitEngineDaemon_CP_3465_elements(38);
      transmitEngineDaemon_CP_3465_elements(39)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitEngineDaemon_CP_3465_elements(40);
      transmitEngineDaemon_CP_3465_elements(32) <= phi_mux_reqs(1);
      phi_stmt_2058_phi_seq_3644 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_2058_phi_seq_3644") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitEngineDaemon_CP_3465_elements(16), 
          phi_sample_ack => transmitEngineDaemon_CP_3465_elements(27), 
          phi_update_req => transmitEngineDaemon_CP_3465_elements(18), 
          phi_update_ack => transmitEngineDaemon_CP_3465_elements(28), 
          phi_mux_ack => transmitEngineDaemon_CP_3465_elements(33), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3578_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitEngineDaemon_CP_3465_elements(12);
        preds(1)  <= transmitEngineDaemon_CP_3465_elements(13);
        entry_tmerge_3578 : transition_merge -- 
          generic map(name => " entry_tmerge_3578")
          port map (preds => preds, symbol_out => transmitEngineDaemon_CP_3465_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_2098_2098_delayed_14_0_2126 : std_logic_vector(31 downto 0);
    signal ADD_u6_u6_2052_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_2057_wire : std_logic_vector(5 downto 0);
    signal BITSEL_u32_u1_2041_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_2141_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2042_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2067_2067_delayed_4_0_2084 : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_2114_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_2039_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_2139_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_2099_wire : std_logic_vector(35 downto 0);
    signal RPIPE_LAST_READ_TX_QUEUE_INDEX_2050_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_2053_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_2055_wire : std_logic_vector(31 downto 0);
    signal count_2058 : std_logic_vector(31 downto 0);
    signal count_2091_delayed_14_0_2108 : std_logic_vector(31 downto 0);
    signal count_2099_delayed_14_0_2121 : std_logic_vector(31 downto 0);
    signal ignore_resp_2118 : std_logic_vector(31 downto 0);
    signal konst_2034_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2040_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2051_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2054_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2115_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2124_wire_constant : std_logic_vector(31 downto 0);
    signal konst_2140_wire_constant : std_logic_vector(31 downto 0);
    signal ncount_2132 : std_logic_vector(31 downto 0);
    signal ncount_2132_2060_buffered : std_logic_vector(31 downto 0);
    signal pkt_pointer_2069 : std_logic_vector(31 downto 0);
    signal pkt_pointer_2078_delayed_4_0_2095 : std_logic_vector(31 downto 0);
    signal push_pointer_back_to_free_Q_2089 : std_logic_vector(0 downto 0);
    signal push_status_2102 : std_logic_vector(0 downto 0);
    signal transmitted_flag_2073 : std_logic_vector(0 downto 0);
    signal tx_flag_2069 : std_logic_vector(0 downto 0);
    signal tx_q_index_2048 : std_logic_vector(5 downto 0);
    signal type_cast_2056_wire : std_logic_vector(5 downto 0);
    signal type_cast_2062_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2098_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2111_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_2114_wire_constant <= "1111";
    konst_2034_wire_constant <= "000000";
    konst_2040_wire_constant <= "00000000000000000000000000000000";
    konst_2051_wire_constant <= "000001";
    konst_2054_wire_constant <= "00000000000000000000000000000001";
    konst_2115_wire_constant <= "010101";
    konst_2124_wire_constant <= "00000000000000000000000000000001";
    konst_2140_wire_constant <= "00000000000000000000000000000000";
    type_cast_2062_wire_constant <= "00000000000000000000000000000001";
    type_cast_2098_wire_constant <= "1";
    type_cast_2111_wire_constant <= "0";
    phi_stmt_2058: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ncount_2132_2060_buffered & type_cast_2062_wire_constant;
      req <= phi_stmt_2058_req_0 & phi_stmt_2058_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2058",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2058_ack_0,
          idata => idata,
          odata => count_2058,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2058
    -- flow-through select operator MUX_2131_inst
    ncount_2132 <= ADD_u32_u32_2098_2098_delayed_14_0_2126 when (push_pointer_back_to_free_Q_2089(0) /=  '0') else count_2099_delayed_14_0_2121;
    W_count_2091_delayed_14_0_2106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_2091_delayed_14_0_2106_inst_req_0;
      W_count_2091_delayed_14_0_2106_inst_ack_0<= wack(0);
      rreq(0) <= W_count_2091_delayed_14_0_2106_inst_req_1;
      W_count_2091_delayed_14_0_2106_inst_ack_1<= rack(0);
      W_count_2091_delayed_14_0_2106_inst : InterlockBuffer generic map ( -- 
        name => "W_count_2091_delayed_14_0_2106_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_2058,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_2091_delayed_14_0_2108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_2099_delayed_14_0_2119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_2099_delayed_14_0_2119_inst_req_0;
      W_count_2099_delayed_14_0_2119_inst_ack_0<= wack(0);
      rreq(0) <= W_count_2099_delayed_14_0_2119_inst_req_1;
      W_count_2099_delayed_14_0_2119_inst_ack_1<= rack(0);
      W_count_2099_delayed_14_0_2119_inst : InterlockBuffer generic map ( -- 
        name => "W_count_2099_delayed_14_0_2119_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_2058,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_2099_delayed_14_0_2121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pkt_pointer_2078_delayed_4_0_2093_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_pointer_2078_delayed_4_0_2093_inst_req_0;
      W_pkt_pointer_2078_delayed_4_0_2093_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_pointer_2078_delayed_4_0_2093_inst_req_1;
      W_pkt_pointer_2078_delayed_4_0_2093_inst_ack_1<= rack(0);
      W_pkt_pointer_2078_delayed_4_0_2093_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_pointer_2078_delayed_4_0_2093_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_pointer_2069,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_pointer_2078_delayed_4_0_2095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ncount_2132_2060_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_2132_2060_buf_req_0;
      ncount_2132_2060_buf_ack_0<= wack(0);
      rreq(0) <= ncount_2132_2060_buf_req_1;
      ncount_2132_2060_buf_ack_1<= rack(0);
      ncount_2132_2060_buf : InterlockBuffer generic map ( -- 
        name => "ncount_2132_2060_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_2132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_2132_2060_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2048
    process(AND_u6_u6_2057_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := AND_u6_u6_2057_wire(5 downto 0);
      tx_q_index_2048 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2056_inst
    process(SUB_u32_u32_2055_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_2055_wire(5 downto 0);
      type_cast_2056_wire <= tmp_var; -- 
    end process;
    do_while_stmt_2046_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_2141_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2046_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2046_branch_req_0,
          ack0 => do_while_stmt_2046_branch_ack_0,
          ack1 => do_while_stmt_2046_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2038_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2042_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2038_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2038_branch_req_0,
          ack0 => if_stmt_2038_branch_ack_0,
          ack1 => if_stmt_2038_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_2125_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= count_2058;
      ADD_u32_u32_2098_2098_delayed_14_0_2126 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_2125_inst_req_0;
      ADD_u32_u32_2125_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_2125_inst_req_1;
      ADD_u32_u32_2125_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u6_u6_2052_inst
    process(RPIPE_LAST_READ_TX_QUEUE_INDEX_2050_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_READ_TX_QUEUE_INDEX_2050_wire, konst_2051_wire_constant, tmp_var);
      ADD_u6_u6_2052_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2088_inst
    process(NOT_u1_u1_2067_2067_delayed_4_0_2084, transmitted_flag_2073) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_2067_2067_delayed_4_0_2084, transmitted_flag_2073, tmp_var);
      push_pointer_back_to_free_Q_2089 <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_2057_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_2052_wire & type_cast_2056_wire;
      AND_u6_u6_2057_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_2057_inst_req_0;
      AND_u6_u6_2057_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_2057_inst_req_1;
      AND_u6_u6_2057_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator BITSEL_u32_u1_2041_inst
    process(RPIPE_CONTROL_REGISTER_2039_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_2039_wire, konst_2040_wire_constant, tmp_var);
      BITSEL_u32_u1_2041_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_2141_inst
    process(RPIPE_CONTROL_REGISTER_2139_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_2139_wire, konst_2140_wire_constant, tmp_var);
      BITSEL_u32_u1_2141_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2042_inst
    process(BITSEL_u32_u1_2041_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_2041_wire, tmp_var);
      NOT_u1_u1_2042_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (7) : NOT_u1_u1_2083_inst 
    ApIntNot_group_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tx_flag_2069;
      NOT_u1_u1_2067_2067_delayed_4_0_2084 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_2083_inst_req_0;
      NOT_u1_u1_2083_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_2083_inst_req_1;
      NOT_u1_u1_2083_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_7_gI: SplitGuardInterface generic map(name => "ApIntNot_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u32_u32_2055_inst
    process(RPIPE_NUMBER_OF_SERVERS_2053_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_2053_wire, konst_2054_wire_constant, tmp_var);
      SUB_u32_u32_2055_wire <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_2039_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_2139_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_2099_wire <= FREE_Q;
    -- read from input-signal LAST_READ_TX_QUEUE_INDEX
    RPIPE_LAST_READ_TX_QUEUE_INDEX_2050_wire <= LAST_READ_TX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_2053_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2033_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2034_wire_constant;
      LAST_READ_TX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 6),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_2135_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= tx_q_index_2048;
      LAST_READ_TX_QUEUE_INDEX_write_1_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_1: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2069_call 
    getTxPacketPointerFromServer_call_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2069_call_req_0;
      call_stmt_2069_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2069_call_req_1;
      call_stmt_2069_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTxPacketPointerFromServer_call_group_0_gI: SplitGuardInterface generic map(name => "getTxPacketPointerFromServer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_q_index_2048;
      pkt_pointer_2069 <= data_out(32 downto 1);
      tx_flag_2069 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 6,
        owidth => 6,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTxPacketPointerFromServer_call_reqs(0),
          ackR => getTxPacketPointerFromServer_call_acks(0),
          dataR => getTxPacketPointerFromServer_call_data(5 downto 0),
          tagR => getTxPacketPointerFromServer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTxPacketPointerFromServer_return_acks(0), -- cross-over
          ackL => getTxPacketPointerFromServer_return_reqs(0), -- cross-over
          dataL => getTxPacketPointerFromServer_return_data(32 downto 0),
          tagL => getTxPacketPointerFromServer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_2073_call 
    transmitPacket_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2073_call_req_0;
      call_stmt_2073_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2073_call_req_1;
      call_stmt_2073_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not tx_flag_2069(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      transmitPacket_call_group_1_gI: SplitGuardInterface generic map(name => "transmitPacket_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pkt_pointer_2069;
      transmitted_flag_2073 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => transmitPacket_call_reqs(0),
          ackR => transmitPacket_call_acks(0),
          dataR => transmitPacket_call_data(31 downto 0),
          tagR => transmitPacket_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => transmitPacket_return_acks(0), -- cross-over
          ackL => transmitPacket_return_reqs(0), -- cross-over
          dataL => transmitPacket_return_data(0 downto 0),
          tagL => transmitPacket_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_2102_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2102_call_req_0;
      call_stmt_2102_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2102_call_req_1;
      call_stmt_2102_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_2089(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2098_wire_constant & RPIPE_FREE_Q_2099_wire & pkt_pointer_2078_delayed_4_0_2095;
      push_status_2102 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_2118_call 
    AccessRegister_call_group_3: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2118_call_req_0;
      call_stmt_2118_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2118_call_req_1;
      call_stmt_2118_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_2089(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_3_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2111_wire_constant & NOT_u4_u4_2114_wire_constant & konst_2115_wire_constant & count_2091_delayed_14_0_2108;
      ignore_resp_2118 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end transmitEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitPacket is -- 
  generic (tag_length : integer); 
  port ( -- 
    packet_pointer : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_call_acks : in   std_logic_vector(1 downto 0);
    accessMemory_call_data : out  std_logic_vector(219 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_return_acks : in   std_logic_vector(1 downto 0);
    accessMemory_return_data : in   std_logic_vector(127 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitPacket;
architecture transmitPacket_arch of transmitPacket is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal packet_pointer_buffer :  std_logic_vector(31 downto 0);
  signal packet_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal transmitPacket_CP_3197_start: Boolean;
  signal transmitPacket_CP_3197_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal nmem_addr_1986_1954_buf_ack_0 : boolean;
  signal call_stmt_2011_call_req_1 : boolean;
  signal EQ_u8_u1_2028_inst_req_1 : boolean;
  signal EQ_u8_u1_2028_inst_ack_1 : boolean;
  signal CONCAT_u65_u73_2020_inst_ack_1 : boolean;
  signal CONCAT_u65_u73_2020_inst_req_1 : boolean;
  signal call_stmt_1968_call_ack_1 : boolean;
  signal nmem_addr_1986_1954_buf_req_0 : boolean;
  signal EQ_u8_u1_2028_inst_req_0 : boolean;
  signal CONCAT_u65_u73_2020_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2014_inst_ack_1 : boolean;
  signal call_stmt_1968_call_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2014_inst_req_1 : boolean;
  signal do_while_stmt_1944_branch_ack_1 : boolean;
  signal EQ_u8_u1_2028_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_1975_inst_req_0 : boolean;
  signal CONCAT_u65_u73_2020_inst_req_0 : boolean;
  signal nmem_addr_1986_1954_buf_ack_1 : boolean;
  signal nmem_addr_1986_1954_buf_req_1 : boolean;
  signal CONCAT_u65_u73_1975_inst_ack_0 : boolean;
  signal do_while_stmt_1944_branch_ack_0 : boolean;
  signal call_stmt_1968_call_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1969_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1969_inst_req_1 : boolean;
  signal call_stmt_1968_call_req_0 : boolean;
  signal call_stmt_2011_call_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1969_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1969_inst_req_0 : boolean;
  signal call_stmt_2011_call_ack_0 : boolean;
  signal call_stmt_2011_call_req_0 : boolean;
  signal ADD_u36_u36_1957_inst_ack_1 : boolean;
  signal ADD_u36_u36_1957_inst_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2014_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_2014_inst_req_0 : boolean;
  signal ADD_u36_u36_1957_inst_ack_0 : boolean;
  signal ADD_u36_u36_1957_inst_req_0 : boolean;
  signal CONCAT_u65_u73_1975_inst_ack_1 : boolean;
  signal CONCAT_u65_u73_1975_inst_req_1 : boolean;
  signal call_stmt_1931_call_req_0 : boolean;
  signal call_stmt_1931_call_ack_0 : boolean;
  signal call_stmt_1931_call_req_1 : boolean;
  signal call_stmt_1931_call_ack_1 : boolean;
  signal do_while_stmt_1944_branch_req_0 : boolean;
  signal phi_stmt_1946_req_1 : boolean;
  signal phi_stmt_1946_req_0 : boolean;
  signal phi_stmt_1946_ack_0 : boolean;
  signal SUB_u8_u8_1950_inst_req_0 : boolean;
  signal SUB_u8_u8_1950_inst_ack_0 : boolean;
  signal SUB_u8_u8_1950_inst_req_1 : boolean;
  signal SUB_u8_u8_1950_inst_ack_1 : boolean;
  signal ncount_down_1981_1951_buf_req_0 : boolean;
  signal ncount_down_1981_1951_buf_ack_0 : boolean;
  signal ncount_down_1981_1951_buf_req_1 : boolean;
  signal ncount_down_1981_1951_buf_ack_1 : boolean;
  signal phi_stmt_1952_req_0 : boolean;
  signal phi_stmt_1952_req_1 : boolean;
  signal phi_stmt_1952_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitPacket_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= packet_pointer;
  packet_pointer_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitPacket_CP_3197_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitPacket_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_3197_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitPacket_CP_3197_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_3197_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitPacket_CP_3197: Block -- control-path 
    signal transmitPacket_CP_3197_elements: BooleanArray(81 downto 0);
    -- 
  begin -- 
    transmitPacket_CP_3197_elements(0) <= transmitPacket_CP_3197_start;
    transmitPacket_CP_3197_symbol <= transmitPacket_CP_3197_elements(81);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1918_to_assign_stmt_1939/$entry
      -- CP-element group 0: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_sample_start_
      -- CP-element group 0: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_update_start_
      -- CP-element group 0: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Update/ccr
      -- 
    ccr_3215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(0), ack => call_stmt_1931_call_req_1); -- 
    crr_3210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(0), ack => call_stmt_1931_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Sample/cra
      -- 
    cra_3211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1931_call_ack_0, ack => transmitPacket_CP_3197_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_1918_to_assign_stmt_1939/$exit
      -- CP-element group 2: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_update_completed_
      -- CP-element group 2: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1918_to_assign_stmt_1939/call_stmt_1931_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1943/$entry
      -- CP-element group 2: 	 branch_block_stmt_1943/branch_block_stmt_1943__entry__
      -- CP-element group 2: 	 branch_block_stmt_1943/do_while_stmt_1944__entry__
      -- 
    cca_3216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1931_call_ack_1, ack => transmitPacket_CP_3197_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	72 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	79 
    -- CP-element group 3: 	80 
    -- CP-element group 3: 	76 
    -- CP-element group 3: 	73 
    -- CP-element group 3: 	74 
    -- CP-element group 3:  members (18) 
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/$entry
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1943/do_while_stmt_1944__exit__
      -- CP-element group 3: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029__entry__
      -- 
    ccr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(3), ack => call_stmt_2011_call_req_1); -- 
    cr_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(3), ack => EQ_u8_u1_2028_inst_req_1); -- 
    cr_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(3), ack => CONCAT_u65_u73_2020_inst_req_1); -- 
    rr_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(3), ack => EQ_u8_u1_2028_inst_req_0); -- 
    crr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(3), ack => call_stmt_2011_call_req_0); -- 
    transmitPacket_CP_3197_elements(3) <= transmitPacket_CP_3197_elements(72);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_1943/do_while_stmt_1944/$entry
      -- CP-element group 4: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944__entry__
      -- 
    transmitPacket_CP_3197_elements(4) <= transmitPacket_CP_3197_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	72 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944__exit__
      -- 
    -- Element group transmitPacket_CP_3197_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_back
      -- 
    -- Element group transmitPacket_CP_3197_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	70 
    -- CP-element group 7: 	71 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_taken/$entry
      -- CP-element group 7: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_1943/do_while_stmt_1944/condition_done
      -- 
    transmitPacket_CP_3197_elements(7) <= transmitPacket_CP_3197_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	69 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_body_done
      -- 
    transmitPacket_CP_3197_elements(8) <= transmitPacket_CP_3197_elements(69);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	42 
    -- CP-element group 9: 	23 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/back_edge_to_loop_body
      -- 
    transmitPacket_CP_3197_elements(9) <= transmitPacket_CP_3197_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	44 
    -- CP-element group 10: 	25 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/first_time_through_loop_body
      -- 
    transmitPacket_CP_3197_elements(10) <= transmitPacket_CP_3197_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	68 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	38 
    -- CP-element group 11: 	39 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/loop_body_start
      -- 
    -- Element group transmitPacket_CP_3197_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	68 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	22 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/condition_evaluated
      -- 
    condition_evaluated_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(12), ack => do_while_stmt_1944_branch_req_0); -- 
    transmitPacket_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(68) & transmitPacket_CP_3197_elements(16) & transmitPacket_CP_3197_elements(22);
      gj_transmitPacket_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: 	38 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/aggregated_phi_sample_req
      -- CP-element group 13: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_sample_start__ps
      -- 
    transmitPacket_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(17) & transmitPacket_CP_3197_elements(38) & transmitPacket_CP_3197_elements(16);
      gj_transmitPacket_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	40 
    -- CP-element group 14: 	20 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	69 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	38 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_sample_completed_
      -- 
    transmitPacket_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(40) & transmitPacket_CP_3197_elements(20);
      gj_transmitPacket_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	39 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	21 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/aggregated_phi_update_req
      -- CP-element group 15: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_update_start__ps
      -- 
    transmitPacket_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(18) & transmitPacket_CP_3197_elements(39);
      gj_transmitPacket_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	22 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/aggregated_phi_update_ack
      -- 
    transmitPacket_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(41) & transmitPacket_CP_3197_elements(22);
      gj_transmitPacket_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_sample_start_
      -- 
    transmitPacket_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(11) & transmitPacket_CP_3197_elements(14);
      gj_transmitPacket_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_update_start_
      -- 
    transmitPacket_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(11) & transmitPacket_CP_3197_elements(22);
      gj_transmitPacket_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_sample_start__ps
      -- 
    transmitPacket_CP_3197_elements(19) <= transmitPacket_CP_3197_elements(13);
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_update_start__ps
      -- 
    transmitPacket_CP_3197_elements(21) <= transmitPacket_CP_3197_elements(15);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: 	12 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	9 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_loopback_trigger
      -- 
    transmitPacket_CP_3197_elements(23) <= transmitPacket_CP_3197_elements(9);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_loopback_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_loopback_sample_req_ps
      -- 
    phi_stmt_1946_loopback_sample_req_3255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1946_loopback_sample_req_3255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(24), ack => phi_stmt_1946_req_1); -- 
    -- Element group transmitPacket_CP_3197_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_entry_trigger
      -- 
    transmitPacket_CP_3197_elements(25) <= transmitPacket_CP_3197_elements(10);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_entry_sample_req
      -- CP-element group 26: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_entry_sample_req_ps
      -- 
    phi_stmt_1946_entry_sample_req_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1946_entry_sample_req_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(26), ack => phi_stmt_1946_req_0); -- 
    -- Element group transmitPacket_CP_3197_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_phi_mux_ack
      -- CP-element group 27: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1946_phi_mux_ack_ps
      -- 
    phi_stmt_1946_phi_mux_ack_3261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1946_ack_0, ack => transmitPacket_CP_3197_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_update_start__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Sample/rr
      -- 
    rr_3274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(30), ack => SUB_u8_u8_1950_inst_req_0); -- 
    transmitPacket_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(28) & transmitPacket_CP_3197_elements(32);
      gj_transmitPacket_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Update/cr
      -- 
    cr_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(31), ack => SUB_u8_u8_1950_inst_req_1); -- 
    transmitPacket_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(29) & transmitPacket_CP_3197_elements(33);
      gj_transmitPacket_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Sample/ra
      -- 
    ra_3275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u8_u8_1950_inst_ack_0, ack => transmitPacket_CP_3197_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/SUB_u8_u8_1950_Update/ca
      -- 
    ca_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u8_u8_1950_inst_ack_1, ack => transmitPacket_CP_3197_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Sample/req
      -- 
    req_3292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(34), ack => ncount_down_1981_1951_buf_req_0); -- 
    -- Element group transmitPacket_CP_3197_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Update/req
      -- 
    req_3297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(35), ack => ncount_down_1981_1951_buf_req_1); -- 
    -- Element group transmitPacket_CP_3197_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_sample_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Sample/ack
      -- 
    ack_3293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1981_1951_buf_ack_0, ack => transmitPacket_CP_3197_elements(36)); -- 
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_update_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_ncount_down_1951_Update/ack
      -- 
    ack_3298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1981_1951_buf_ack_1, ack => transmitPacket_CP_3197_elements(37)); -- 
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	13 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_sample_start_
      -- 
    transmitPacket_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(11) & transmitPacket_CP_3197_elements(14);
      gj_transmitPacket_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	11 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	59 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	15 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_update_start_
      -- 
    transmitPacket_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(11) & transmitPacket_CP_3197_elements(59) & transmitPacket_CP_3197_elements(41);
      gj_transmitPacket_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	14 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	16 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	9 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_loopback_trigger
      -- 
    transmitPacket_CP_3197_elements(42) <= transmitPacket_CP_3197_elements(9);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_loopback_sample_req_ps
      -- 
    phi_stmt_1952_loopback_sample_req_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1952_loopback_sample_req_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(43), ack => phi_stmt_1952_req_0); -- 
    -- Element group transmitPacket_CP_3197_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	10 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_entry_trigger
      -- 
    transmitPacket_CP_3197_elements(44) <= transmitPacket_CP_3197_elements(10);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_entry_sample_req
      -- CP-element group 45: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_entry_sample_req_ps
      -- 
    phi_stmt_1952_entry_sample_req_3312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1952_entry_sample_req_3312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(45), ack => phi_stmt_1952_req_1); -- 
    -- Element group transmitPacket_CP_3197_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/phi_stmt_1952_phi_mux_ack_ps
      -- 
    phi_stmt_1952_phi_mux_ack_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1952_ack_0, ack => transmitPacket_CP_3197_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_sample_start__ps
      -- 
    req_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(47), ack => nmem_addr_1986_1954_buf_req_0); -- 
    -- Element group transmitPacket_CP_3197_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Update/req
      -- CP-element group 48: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_update_start__ps
      -- 
    req_3333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(48), ack => nmem_addr_1986_1954_buf_req_1); -- 
    -- Element group transmitPacket_CP_3197_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_sample_completed__ps
      -- 
    ack_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1986_1954_buf_ack_0, ack => transmitPacket_CP_3197_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/R_nmem_addr_1954_update_completed__ps
      -- 
    ack_3334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1986_1954_buf_ack_1, ack => transmitPacket_CP_3197_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_update_start__ps
      -- 
    -- Element group transmitPacket_CP_3197_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_sample_start_
      -- 
    rr_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(53), ack => ADD_u36_u36_1957_inst_req_0); -- 
    transmitPacket_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(51) & transmitPacket_CP_3197_elements(55);
      gj_transmitPacket_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Update/cr
      -- CP-element group 54: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_update_start_
      -- 
    cr_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(54), ack => ADD_u36_u36_1957_inst_req_1); -- 
    transmitPacket_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(52) & transmitPacket_CP_3197_elements(56);
      gj_transmitPacket_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_sample_completed_
      -- 
    ra_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1957_inst_ack_0, ack => transmitPacket_CP_3197_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/ADD_u36_u36_1957_update_completed_
      -- 
    ca_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1957_inst_ack_1, ack => transmitPacket_CP_3197_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Sample/crr
      -- CP-element group 57: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_sample_start_
      -- 
    crr_3361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(57), ack => call_stmt_1968_call_req_0); -- 
    transmitPacket_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(41) & transmitPacket_CP_3197_elements(59);
      gj_transmitPacket_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	63 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Update/ccr
      -- CP-element group 58: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_update_start_
      -- 
    ccr_3366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(58), ack => call_stmt_1968_call_req_1); -- 
    transmitPacket_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(60) & transmitPacket_CP_3197_elements(63);
      gj_transmitPacket_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: 	39 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Sample/cra
      -- CP-element group 59: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_sample_completed_
      -- 
    cra_3362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1968_call_ack_0, ack => transmitPacket_CP_3197_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Update/cca
      -- CP-element group 60: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/call_stmt_1968_update_completed_
      -- 
    cca_3367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1968_call_ack_1, ack => transmitPacket_CP_3197_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Sample/rr
      -- 
    rr_3375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(61), ack => CONCAT_u65_u73_1975_inst_req_0); -- 
    transmitPacket_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(60) & transmitPacket_CP_3197_elements(63);
      gj_transmitPacket_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	66 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Update/cr
      -- 
    cr_3380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(62), ack => CONCAT_u65_u73_1975_inst_req_1); -- 
    transmitPacket_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(64) & transmitPacket_CP_3197_elements(66);
      gj_transmitPacket_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	58 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Sample/ra
      -- 
    ra_3376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1975_inst_ack_0, ack => transmitPacket_CP_3197_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/CONCAT_u65_u73_1975_Update/ca
      -- 
    ca_3381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1975_inst_ack_1, ack => transmitPacket_CP_3197_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_sample_start_
      -- 
    req_3389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(65), ack => WPIPE_nic_to_mac_transmit_pipe_1969_inst_req_0); -- 
    transmitPacket_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(64) & transmitPacket_CP_3197_elements(67);
      gj_transmitPacket_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	62 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Update/req
      -- CP-element group 66: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_sample_completed_
      -- 
    ack_3390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1969_inst_ack_0, ack => transmitPacket_CP_3197_elements(66)); -- 
    req_3394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(66), ack => WPIPE_nic_to_mac_transmit_pipe_1969_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/WPIPE_nic_to_mac_transmit_pipe_1969_update_completed_
      -- 
    ack_3395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1969_inst_ack_1, ack => transmitPacket_CP_3197_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	11 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	12 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitPacket_CP_3197_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => transmitPacket_CP_3197_elements(11), ack => transmitPacket_CP_3197_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	14 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	8 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1943/do_while_stmt_1944/do_while_stmt_1944_loop_body/$exit
      -- 
    transmitPacket_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(67) & transmitPacket_CP_3197_elements(14);
      gj_transmitPacket_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	7 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_exit/ack
      -- CP-element group 70: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_exit/$exit
      -- 
    ack_3400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1944_branch_ack_0, ack => transmitPacket_CP_3197_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	7 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_taken/ack
      -- CP-element group 71: 	 branch_block_stmt_1943/do_while_stmt_1944/loop_taken/$exit
      -- 
    ack_3404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1944_branch_ack_1, ack => transmitPacket_CP_3197_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	5 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	3 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1943/do_while_stmt_1944/$exit
      -- 
    transmitPacket_CP_3197_elements(72) <= transmitPacket_CP_3197_elements(5);
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	3 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Sample/cra
      -- CP-element group 73: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Sample/$exit
      -- 
    cra_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2011_call_ack_0, ack => transmitPacket_CP_3197_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	3 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/call_stmt_2011_Update/cca
      -- 
    cca_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2011_call_ack_1, ack => transmitPacket_CP_3197_elements(74)); -- 
    rr_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(74), ack => CONCAT_u65_u73_2020_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_sample_completed_
      -- 
    ra_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2020_inst_ack_0, ack => transmitPacket_CP_3197_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	3 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/CONCAT_u65_u73_2020_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Sample/req
      -- 
    ca_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_2020_inst_ack_1, ack => transmitPacket_CP_3197_elements(76)); -- 
    req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(76), ack => WPIPE_nic_to_mac_transmit_pipe_2014_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Update/req
      -- CP-element group 77: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Sample/$exit
      -- 
    ack_3445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2014_inst_ack_0, ack => transmitPacket_CP_3197_elements(77)); -- 
    req_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_3197_elements(77), ack => WPIPE_nic_to_mac_transmit_pipe_2014_inst_req_1); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/WPIPE_nic_to_mac_transmit_pipe_2014_Update/$exit
      -- 
    ack_3450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_2014_inst_ack_1, ack => transmitPacket_CP_3197_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	3 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Sample/ra
      -- 
    ra_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_2028_inst_ack_0, ack => transmitPacket_CP_3197_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	3 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/EQ_u8_u1_2028_Update/$exit
      -- 
    ca_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_2028_inst_ack_1, ack => transmitPacket_CP_3197_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: 	78 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029/$exit
      -- CP-element group 81: 	 $exit
      -- CP-element group 81: 	 branch_block_stmt_1943/$exit
      -- CP-element group 81: 	 branch_block_stmt_1943/branch_block_stmt_1943__exit__
      -- CP-element group 81: 	 branch_block_stmt_1943/call_stmt_2011_to_assign_stmt_2029__exit__
      -- 
    transmitPacket_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_3197_elements(80) & transmitPacket_CP_3197_elements(78);
      gj_transmitPacket_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_3197_elements(81), clk => clk, reset => reset); --
    end block;
    transmitPacket_do_while_stmt_1944_terminator_3405: loop_terminator -- 
      generic map (name => " transmitPacket_do_while_stmt_1944_terminator_3405", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitPacket_CP_3197_elements(8),loop_continue => transmitPacket_CP_3197_elements(71),loop_terminate => transmitPacket_CP_3197_elements(70),loop_back => transmitPacket_CP_3197_elements(6),loop_exit => transmitPacket_CP_3197_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_1946_phi_seq_3299_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_3197_elements(25);
      transmitPacket_CP_3197_elements(28)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_3197_elements(32);
      transmitPacket_CP_3197_elements(29)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_3197_elements(33);
      transmitPacket_CP_3197_elements(26) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_3197_elements(23);
      transmitPacket_CP_3197_elements(34)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_3197_elements(36);
      transmitPacket_CP_3197_elements(35)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_3197_elements(37);
      transmitPacket_CP_3197_elements(24) <= phi_mux_reqs(1);
      phi_stmt_1946_phi_seq_3299 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1946_phi_seq_3299") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_3197_elements(19), 
          phi_sample_ack => transmitPacket_CP_3197_elements(20), 
          phi_update_req => transmitPacket_CP_3197_elements(21), 
          phi_update_ack => transmitPacket_CP_3197_elements(22), 
          phi_mux_ack => transmitPacket_CP_3197_elements(27), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1952_phi_seq_3353_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_3197_elements(42);
      transmitPacket_CP_3197_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_3197_elements(49);
      transmitPacket_CP_3197_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_3197_elements(50);
      transmitPacket_CP_3197_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_3197_elements(44);
      transmitPacket_CP_3197_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_3197_elements(55);
      transmitPacket_CP_3197_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_3197_elements(56);
      transmitPacket_CP_3197_elements(45) <= phi_mux_reqs(1);
      phi_stmt_1952_phi_seq_3353 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1952_phi_seq_3353") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_3197_elements(13), 
          phi_sample_ack => transmitPacket_CP_3197_elements(40), 
          phi_update_req => transmitPacket_CP_3197_elements(15), 
          phi_update_ack => transmitPacket_CP_3197_elements(41), 
          phi_mux_ack => transmitPacket_CP_3197_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3241_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitPacket_CP_3197_elements(9);
        preds(1)  <= transmitPacket_CP_3197_elements(10);
        entry_tmerge_3241 : transition_merge -- 
          generic map(name => " entry_tmerge_3241")
          port map (preds => preds, symbol_out => transmitPacket_CP_3197_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1957_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u1_u65_1973_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u1_u65_2018_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u65_u73_1975_wire : std_logic_vector(72 downto 0);
    signal CONCAT_u65_u73_2020_wire : std_logic_vector(72 downto 0);
    signal R_FULL_BYTE_MASK_1926_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1963_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1974_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_2006_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u36_u36_2026_wire : std_logic_vector(35 downto 0);
    signal SUB_u8_u8_1950_wire : std_logic_vector(7 downto 0);
    signal control_data_1931 : std_logic_vector(63 downto 0);
    signal control_data_addr_1918 : std_logic_vector(35 downto 0);
    signal count_down_1946 : std_logic_vector(7 downto 0);
    signal data_1968 : std_logic_vector(63 downto 0);
    signal konst_1949_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1956_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1979_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1984_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1995_wire_constant : std_logic_vector(7 downto 0);
    signal last_tkeep_1939 : std_logic_vector(7 downto 0);
    signal last_word_2011 : std_logic_vector(63 downto 0);
    signal mem_addr_1952 : std_logic_vector(35 downto 0);
    signal ncount_down_1981 : std_logic_vector(7 downto 0);
    signal ncount_down_1981_1951_buffered : std_logic_vector(7 downto 0);
    signal nmem_addr_1986 : std_logic_vector(35 downto 0);
    signal nmem_addr_1986_1954_buffered : std_logic_vector(35 downto 0);
    signal not_last_word_1997 : std_logic_vector(0 downto 0);
    signal packet_size_1935 : std_logic_vector(7 downto 0);
    signal type_cast_1923_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1925_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1929_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1960_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1962_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1966_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1971_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2003_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2005_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2009_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2016_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2027_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_1926_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1963_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1974_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_2006_wire_constant <= "11111111";
    konst_1949_wire_constant <= "00010000";
    konst_1956_wire_constant <= "000000000000000000000000000000011000";
    konst_1979_wire_constant <= "00001000";
    konst_1984_wire_constant <= "000000000000000000000000000000001000";
    konst_1995_wire_constant <= "00001000";
    type_cast_1923_wire_constant <= "0";
    type_cast_1925_wire_constant <= "1";
    type_cast_1929_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1960_wire_constant <= "0";
    type_cast_1962_wire_constant <= "1";
    type_cast_1966_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1971_wire_constant <= "0";
    type_cast_2003_wire_constant <= "0";
    type_cast_2005_wire_constant <= "1";
    type_cast_2009_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_2016_wire_constant <= "1";
    phi_stmt_1946: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SUB_u8_u8_1950_wire & ncount_down_1981_1951_buffered;
      req <= phi_stmt_1946_req_0 & phi_stmt_1946_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1946",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1946_ack_0,
          idata => idata,
          odata => count_down_1946,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1946
    phi_stmt_1952: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmem_addr_1986_1954_buffered & ADD_u36_u36_1957_wire;
      req <= phi_stmt_1952_req_0 & phi_stmt_1952_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1952",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1952_ack_0,
          idata => idata,
          odata => mem_addr_1952,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1952
    -- flow-through slice operator slice_1934_inst
    packet_size_1935 <= control_data_1931(15 downto 8);
    -- flow-through slice operator slice_1938_inst
    last_tkeep_1939 <= control_data_1931(7 downto 0);
    ncount_down_1981_1951_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_down_1981_1951_buf_req_0;
      ncount_down_1981_1951_buf_ack_0<= wack(0);
      rreq(0) <= ncount_down_1981_1951_buf_req_1;
      ncount_down_1981_1951_buf_ack_1<= rack(0);
      ncount_down_1981_1951_buf : InterlockBuffer generic map ( -- 
        name => "ncount_down_1981_1951_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_down_1981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_down_1981_1951_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmem_addr_1986_1954_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmem_addr_1986_1954_buf_req_0;
      nmem_addr_1986_1954_buf_ack_0<= wack(0);
      rreq(0) <= nmem_addr_1986_1954_buf_req_1;
      nmem_addr_1986_1954_buf_ack_1<= rack(0);
      nmem_addr_1986_1954_buf : InterlockBuffer generic map ( -- 
        name => "nmem_addr_1986_1954_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_1986,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmem_addr_1986_1954_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1917_inst
    process(packet_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := packet_pointer_buffer(31 downto 0);
      control_data_addr_1918 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2027_inst
    process(SUB_u36_u36_2026_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u36_u36_2026_wire(7 downto 0);
      type_cast_2027_wire <= tmp_var; -- 
    end process;
    do_while_stmt_1944_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= not_last_word_1997;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1944_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1944_branch_req_0,
          ack0 => do_while_stmt_1944_branch_ack_0,
          ack1 => do_while_stmt_1944_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1957_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= control_data_addr_1918;
      ADD_u36_u36_1957_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1957_inst_req_0;
      ADD_u36_u36_1957_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1957_inst_req_1;
      ADD_u36_u36_1957_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000011000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_1985_inst
    process(mem_addr_1952) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mem_addr_1952, konst_1984_wire_constant, tmp_var);
      nmem_addr_1986 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_1973_inst
    process(type_cast_1971_wire_constant, data_1968) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1971_wire_constant, data_1968, tmp_var);
      CONCAT_u1_u65_1973_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_2018_inst
    process(type_cast_2016_wire_constant, last_word_2011) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2016_wire_constant, last_word_2011, tmp_var);
      CONCAT_u1_u65_2018_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : CONCAT_u65_u73_1975_inst 
    ApConcat_group_4: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_1973_wire;
      CONCAT_u65_u73_1975_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_1975_inst_req_0;
      CONCAT_u65_u73_1975_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_1975_inst_req_1;
      CONCAT_u65_u73_1975_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_4_gI: SplitGuardInterface generic map(name => "ApConcat_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : CONCAT_u65_u73_2020_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_2018_wire & last_tkeep_1939;
      CONCAT_u65_u73_2020_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_2020_inst_req_0;
      CONCAT_u65_u73_2020_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_2020_inst_req_1;
      CONCAT_u65_u73_2020_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : EQ_u8_u1_2028_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_1935 & type_cast_2027_wire;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_2028_inst_req_0;
      EQ_u8_u1_2028_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_2028_inst_req_1;
      EQ_u8_u1_2028_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- binary operator SUB_u36_u36_2026_inst
    process(nmem_addr_1986, control_data_addr_1918) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(nmem_addr_1986, control_data_addr_1918, tmp_var);
      SUB_u36_u36_2026_wire <= tmp_var; --
    end process;
    -- shared split operator group (8) : SUB_u8_u8_1950_inst 
    ApIntSub_group_8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_1935;
      SUB_u8_u8_1950_wire <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u8_u8_1950_inst_req_0;
      SUB_u8_u8_1950_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u8_u8_1950_inst_req_1;
      SUB_u8_u8_1950_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_8_gI: SplitGuardInterface generic map(name => "ApIntSub_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00010000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- binary operator SUB_u8_u8_1980_inst
    process(count_down_1946) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_1946, konst_1979_wire_constant, tmp_var);
      ncount_down_1981 <= tmp_var; --
    end process;
    -- binary operator UGT_u8_u1_1996_inst
    process(ncount_down_1981) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ncount_down_1981, konst_1995_wire_constant, tmp_var);
      not_last_word_1997 <= tmp_var; --
    end process;
    -- shared outport operator group (0) : WPIPE_nic_to_mac_transmit_pipe_1969_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1969_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_1969_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1969_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_1969_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_1975_wire;
      nic_to_mac_transmit_pipe_write_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(1),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(1),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 73),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_to_mac_transmit_pipe_2014_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2014_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_2014_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_2014_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_2014_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_2020_wire;
      nic_to_mac_transmit_pipe_write_1_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2011_call call_stmt_1931_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_2011_call_req_0;
      reqL_unguarded(0) <= call_stmt_1931_call_req_0;
      call_stmt_2011_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1931_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_2011_call_req_1;
      reqR_unguarded(0) <= call_stmt_1931_call_req_1;
      call_stmt_2011_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1931_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_2003_wire_constant & type_cast_2005_wire_constant & R_FULL_BYTE_MASK_2006_wire_constant & nmem_addr_1986 & type_cast_2009_wire_constant & type_cast_1923_wire_constant & type_cast_1925_wire_constant & R_FULL_BYTE_MASK_1926_wire_constant & control_data_addr_1918 & type_cast_1929_wire_constant;
      last_word_2011 <= data_out(127 downto 64);
      control_data_1931 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(1),
          ackR => accessMemory_call_acks(1),
          dataR => accessMemory_call_data(219 downto 110),
          tagR => accessMemory_call_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(1), -- cross-over
          ackL => accessMemory_return_reqs(1), -- cross-over
          dataL => accessMemory_return_data(127 downto 64),
          tagL => accessMemory_return_tag(5 downto 3),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1968_call 
    accessMemory_call_group_1: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1968_call_req_0;
      call_stmt_1968_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1968_call_req_1;
      call_stmt_1968_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1960_wire_constant & type_cast_1962_wire_constant & R_FULL_BYTE_MASK_1963_wire_constant & mem_addr_1952 & type_cast_1966_wire_constant;
      data_1968 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end transmitPacket_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity updateTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    updated_total_msgs : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity updateTotalMessages;
architecture updateTotalMessages_arch of updateTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal updated_total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal updated_total_msgs_update_enable: Boolean;
  -- output port buffer signals
  signal updateTotalMessages_CP_694_start: Boolean;
  signal updateTotalMessages_CP_694_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_749_call_ack_0 : boolean;
  signal call_stmt_749_call_req_1 : boolean;
  signal call_stmt_749_call_req_0 : boolean;
  signal call_stmt_749_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "updateTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= updated_total_msgs;
  updated_total_msgs_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  updateTotalMessages_CP_694_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "updateTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateTotalMessages_CP_694_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= updateTotalMessages_CP_694_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateTotalMessages_CP_694_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  updateTotalMessages_CP_694: Block -- control-path 
    signal updateTotalMessages_CP_694_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    updateTotalMessages_CP_694_elements(0) <= updateTotalMessages_CP_694_start;
    updateTotalMessages_CP_694_symbol <= updateTotalMessages_CP_694_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_749/call_stmt_749_sample_start_
      -- CP-element group 0: 	 call_stmt_749/call_stmt_749_update_start_
      -- CP-element group 0: 	 call_stmt_749/$entry
      -- CP-element group 0: 	 call_stmt_749/call_stmt_749_Update/ccr
      -- CP-element group 0: 	 call_stmt_749/call_stmt_749_Update/$entry
      -- CP-element group 0: 	 call_stmt_749/call_stmt_749_Sample/crr
      -- CP-element group 0: 	 call_stmt_749/call_stmt_749_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- 
    crr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateTotalMessages_CP_694_elements(0), ack => call_stmt_749_call_req_0); -- 
    ccr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateTotalMessages_CP_694_elements(0), ack => call_stmt_749_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_749/call_stmt_749_Sample/cra
      -- CP-element group 1: 	 call_stmt_749/call_stmt_749_sample_completed_
      -- CP-element group 1: 	 call_stmt_749/call_stmt_749_Sample/$exit
      -- 
    cra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_749_call_ack_0, ack => updateTotalMessages_CP_694_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_749/call_stmt_749_Update/$exit
      -- CP-element group 2: 	 call_stmt_749/call_stmt_749_update_completed_
      -- CP-element group 2: 	 call_stmt_749/$exit
      -- CP-element group 2: 	 call_stmt_749/call_stmt_749_Update/cca
      -- CP-element group 2: 	 $exit
      -- 
    cca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_749_call_ack_1, ack => updateTotalMessages_CP_694_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u32_u64_747_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_742_wire_constant : std_logic_vector(7 downto 0);
    signal rdata_749 : std_logic_vector(63 downto 0);
    signal type_cast_734_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_736_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_742_wire_constant <= "11110000";
    type_cast_734_wire_constant <= "0";
    type_cast_736_wire_constant <= "0";
    type_cast_746_wire_constant <= "00000000000000000000000000000000";
    -- binary operator CONCAT_u32_u64_747_inst
    process(updated_total_msgs_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(updated_total_msgs_buffer, type_cast_746_wire_constant, tmp_var);
      CONCAT_u32_u64_747_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_749_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_749_call_req_0;
      call_stmt_749_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_749_call_req_1;
      call_stmt_749_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_734_wire_constant & type_cast_736_wire_constant & CONCAT_u4_u8_742_wire_constant & q_base_address_buffer & CONCAT_u32_u64_747_wire;
      rdata_749 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end updateTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeControlInformationToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buffer_pointer : in  std_logic_vector(35 downto 0);
    packet_size : in  std_logic_vector(7 downto 0);
    last_keep : in  std_logic_vector(7 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeControlInformationToMem;
architecture writeControlInformationToMem_arch of writeControlInformationToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 52)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buffer_pointer_update_enable: Boolean;
  signal packet_size_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  -- output port buffer signals
  signal writeControlInformationToMem_CP_1185_start: Boolean;
  signal writeControlInformationToMem_CP_1185_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1113_call_ack_1 : boolean;
  signal call_stmt_1113_call_req_1 : boolean;
  signal call_stmt_1113_call_ack_0 : boolean;
  signal call_stmt_1113_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeControlInformationToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 52) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buffer_pointer;
  base_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(43 downto 36) <= packet_size;
  packet_size_buffer <= in_buffer_data_out(43 downto 36);
  in_buffer_data_in(51 downto 44) <= last_keep;
  last_keep_buffer <= in_buffer_data_out(51 downto 44);
  in_buffer_data_in(tag_length + 51 downto 52) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 51 downto 52);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeControlInformationToMem_CP_1185_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeControlInformationToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1185_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1185_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1185_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeControlInformationToMem_CP_1185: Block -- control-path 
    signal writeControlInformationToMem_CP_1185_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeControlInformationToMem_CP_1185_elements(0) <= writeControlInformationToMem_CP_1185_start;
    writeControlInformationToMem_CP_1185_symbol <= writeControlInformationToMem_CP_1185_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_1104_to_call_stmt_1113/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_update_start_
      -- CP-element group 0: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_sample_start_
      -- 
    crr_1198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_1185_elements(0), ack => call_stmt_1113_call_req_0); -- 
    ccr_1203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_1185_elements(0), ack => call_stmt_1113_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Sample/cra
      -- CP-element group 1: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_sample_completed_
      -- 
    cra_1199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1113_call_ack_0, ack => writeControlInformationToMem_CP_1185_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1104_to_call_stmt_1113/$exit
      -- CP-element group 2: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Update/cca
      -- CP-element group 2: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1104_to_call_stmt_1113/call_stmt_1113_update_completed_
      -- 
    cca_1204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1113_call_ack_1, ack => writeControlInformationToMem_CP_1185_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_1102_wire : std_logic_vector(15 downto 0);
    signal R_FULL_BYTE_MASK_1109_wire_constant : std_logic_vector(7 downto 0);
    signal control_data_1104 : std_logic_vector(63 downto 0);
    signal ignore_return_1113 : std_logic_vector(63 downto 0);
    signal type_cast_1106_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1108_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_1109_wire_constant <= "11111111";
    type_cast_1106_wire_constant <= "0";
    type_cast_1108_wire_constant <= "0";
    -- interlock type_cast_1103_inst
    process(CONCAT_u8_u16_1102_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := CONCAT_u8_u16_1102_wire(15 downto 0);
      control_data_1104 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_1102_inst
    process(packet_size_buffer, last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(packet_size_buffer, last_keep_buffer, tmp_var);
      CONCAT_u8_u16_1102_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1113_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1113_call_req_0;
      call_stmt_1113_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1113_call_req_1;
      call_stmt_1113_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1106_wire_constant & type_cast_1108_wire_constant & R_FULL_BYTE_MASK_1109_wire_constant & base_buffer_pointer_buffer & control_data_1104;
      ignore_return_1113 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeControlInformationToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeEthernetHeaderToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    buf_pointer : in  std_logic_vector(35 downto 0);
    buf_position : out  std_logic_vector(35 downto 0);
    nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeEthernetHeaderToMem;
architecture writeEthernetHeaderToMem_arch of writeEthernetHeaderToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal buf_position_buffer :  std_logic_vector(35 downto 0);
  signal buf_position_update_enable: Boolean;
  signal writeEthernetHeaderToMem_CP_886_start: Boolean;
  signal writeEthernetHeaderToMem_CP_886_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_966_branch_req_0 : boolean;
  signal phi_stmt_968_req_1 : boolean;
  signal phi_stmt_968_req_0 : boolean;
  signal phi_stmt_968_ack_0 : boolean;
  signal ADD_u36_u36_972_inst_req_0 : boolean;
  signal ADD_u36_u36_972_inst_ack_0 : boolean;
  signal ADD_u36_u36_972_inst_req_1 : boolean;
  signal ADD_u36_u36_972_inst_ack_1 : boolean;
  signal nbuf_position_1012_973_buf_req_0 : boolean;
  signal nbuf_position_1012_973_buf_ack_0 : boolean;
  signal nbuf_position_1012_973_buf_req_1 : boolean;
  signal nbuf_position_1012_973_buf_ack_1 : boolean;
  signal phi_stmt_974_req_1 : boolean;
  signal phi_stmt_974_req_0 : boolean;
  signal phi_stmt_974_ack_0 : boolean;
  signal nI_1007_978_buf_req_0 : boolean;
  signal nI_1007_978_buf_ack_0 : boolean;
  signal nI_1007_978_buf_req_1 : boolean;
  signal nI_1007_978_buf_ack_1 : boolean;
  signal RPIPE_nic_rx_to_header_981_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_header_981_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_981_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_header_981_inst_ack_1 : boolean;
  signal call_stmt_1002_call_req_0 : boolean;
  signal call_stmt_1002_call_ack_0 : boolean;
  signal call_stmt_1002_call_req_1 : boolean;
  signal call_stmt_1002_call_ack_1 : boolean;
  signal do_while_stmt_966_branch_ack_0 : boolean;
  signal do_while_stmt_966_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeEthernetHeaderToMem_CP_886_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(35 downto 0) <= buf_position_buffer;
  buf_position <= out_buffer_data_out(35 downto 0);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_886_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_886_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_886_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeEthernetHeaderToMem_CP_886: Block -- control-path 
    signal writeEthernetHeaderToMem_CP_886_elements: BooleanArray(66 downto 0);
    -- 
  begin -- 
    writeEthernetHeaderToMem_CP_886_elements(0) <= writeEthernetHeaderToMem_CP_886_start;
    writeEthernetHeaderToMem_CP_886_symbol <= writeEthernetHeaderToMem_CP_886_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_965/$entry
      -- CP-element group 0: 	 branch_block_stmt_965/branch_block_stmt_965__entry__
      -- CP-element group 0: 	 branch_block_stmt_965/do_while_stmt_966__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	66 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_965/$exit
      -- CP-element group 1: 	 branch_block_stmt_965/branch_block_stmt_965__exit__
      -- CP-element group 1: 	 branch_block_stmt_965/do_while_stmt_966__exit__
      -- 
    writeEthernetHeaderToMem_CP_886_elements(1) <= writeEthernetHeaderToMem_CP_886_elements(66);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_965/do_while_stmt_966/$entry
      -- CP-element group 2: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966__entry__
      -- 
    writeEthernetHeaderToMem_CP_886_elements(2) <= writeEthernetHeaderToMem_CP_886_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	66 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966__exit__
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_965/do_while_stmt_966/loop_back
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	64 
    -- CP-element group 5: 	65 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_965/do_while_stmt_966/condition_done
      -- CP-element group 5: 	 branch_block_stmt_965/do_while_stmt_966/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_965/do_while_stmt_966/loop_taken/$entry
      -- 
    writeEthernetHeaderToMem_CP_886_elements(5) <= writeEthernetHeaderToMem_CP_886_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	63 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_965/do_while_stmt_966/loop_body_done
      -- 
    writeEthernetHeaderToMem_CP_886_elements(6) <= writeEthernetHeaderToMem_CP_886_elements(63);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	21 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/back_edge_to_loop_body
      -- 
    writeEthernetHeaderToMem_CP_886_elements(7) <= writeEthernetHeaderToMem_CP_886_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/first_time_through_loop_body
      -- 
    writeEthernetHeaderToMem_CP_886_elements(8) <= writeEthernetHeaderToMem_CP_886_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	62 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_979_sample_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	62 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/condition_evaluated
      -- 
    condition_evaluated_910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(10), ack => do_while_stmt_966_branch_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(62) & writeEthernetHeaderToMem_CP_886_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	54 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_sample_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(9) & writeEthernetHeaderToMem_CP_886_elements(36) & writeEthernetHeaderToMem_CP_886_elements(15) & writeEthernetHeaderToMem_CP_886_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	38 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	18 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	63 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_979_sample_completed_
      -- 
    writeEthernetHeaderToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(38) & writeEthernetHeaderToMem_CP_886_elements(56) & writeEthernetHeaderToMem_CP_886_elements(18);
      gj_writeEthernetHeaderToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	53 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_update_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(37) & writeEthernetHeaderToMem_CP_886_elements(53) & writeEthernetHeaderToMem_CP_886_elements(16);
      gj_writeEthernetHeaderToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	20 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/aggregated_phi_update_ack
      -- 
    writeEthernetHeaderToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(39) & writeEthernetHeaderToMem_CP_886_elements(57) & writeEthernetHeaderToMem_CP_886_elements(20);
      gj_writeEthernetHeaderToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(9) & writeEthernetHeaderToMem_CP_886_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(9) & writeEthernetHeaderToMem_CP_886_elements(20);
      gj_writeEthernetHeaderToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_sample_start__ps
      -- 
    writeEthernetHeaderToMem_CP_886_elements(17) <= writeEthernetHeaderToMem_CP_886_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_update_start__ps
      -- 
    writeEthernetHeaderToMem_CP_886_elements(19) <= writeEthernetHeaderToMem_CP_886_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_886_elements(21) <= writeEthernetHeaderToMem_CP_886_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_loopback_sample_req_ps
      -- 
    phi_stmt_968_loopback_sample_req_925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_968_loopback_sample_req_925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(22), ack => phi_stmt_968_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_886_elements(23) <= writeEthernetHeaderToMem_CP_886_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_entry_sample_req_ps
      -- 
    phi_stmt_968_entry_sample_req_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_968_entry_sample_req_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(24), ack => phi_stmt_968_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_968_phi_mux_ack_ps
      -- 
    phi_stmt_968_phi_mux_ack_931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_968_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Sample/rr
      -- 
    rr_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(28), ack => ADD_u36_u36_972_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(26) & writeEthernetHeaderToMem_CP_886_elements(30);
      gj_writeEthernetHeaderToMem_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_update_start_
      -- CP-element group 29: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Update/cr
      -- 
    cr_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(29), ack => ADD_u36_u36_972_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(27) & writeEthernetHeaderToMem_CP_886_elements(31);
      gj_writeEthernetHeaderToMem_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Sample/ra
      -- 
    ra_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_972_inst_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/ADD_u36_u36_972_Update/ca
      -- 
    ca_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_972_inst_ack_1, ack => writeEthernetHeaderToMem_CP_886_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Sample/req
      -- 
    req_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(32), ack => nbuf_position_1012_973_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_update_start_
      -- CP-element group 33: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Update/req
      -- 
    req_967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(33), ack => nbuf_position_1012_973_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Sample/ack
      -- 
    ack_963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1012_973_buf_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(34)); -- 
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nbuf_position_973_Update/ack
      -- 
    ack_968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1012_973_buf_ack_1, ack => writeEthernetHeaderToMem_CP_886_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(9) & writeEthernetHeaderToMem_CP_886_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(9) & writeEthernetHeaderToMem_CP_886_elements(39);
      gj_writeEthernetHeaderToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_886_elements(40) <= writeEthernetHeaderToMem_CP_886_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_loopback_sample_req_ps
      -- 
    phi_stmt_974_loopback_sample_req_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_974_loopback_sample_req_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(41), ack => phi_stmt_974_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_886_elements(42) <= writeEthernetHeaderToMem_CP_886_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_entry_sample_req_ps
      -- 
    phi_stmt_974_entry_sample_req_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_974_entry_sample_req_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(43), ack => phi_stmt_974_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_974_phi_mux_ack_ps
      -- 
    phi_stmt_974_phi_mux_ack_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_974_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_sample_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_update_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_886_elements(47) <= writeEthernetHeaderToMem_CP_886_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/type_cast_977_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_886_elements(46), ack => writeEthernetHeaderToMem_CP_886_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Sample/req
      -- 
    req_1006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(49), ack => nI_1007_978_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_update_start_
      -- CP-element group 50: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Update/req
      -- 
    req_1011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(50), ack => nI_1007_978_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Sample/ack
      -- 
    ack_1007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_1007_978_buf_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/R_nI_978_Update/ack
      -- 
    ack_1012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_1007_978_buf_ack_1, ack => writeEthernetHeaderToMem_CP_886_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	60 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	13 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_979_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(9) & writeEthernetHeaderToMem_CP_886_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Sample/rr
      -- 
    rr_1025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(54), ack => RPIPE_nic_rx_to_header_981_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(11) & writeEthernetHeaderToMem_CP_886_elements(57);
      gj_writeEthernetHeaderToMem_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_update_start_
      -- CP-element group 55: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Update/cr
      -- 
    cr_1030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(55), ack => RPIPE_nic_rx_to_header_981_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(56) & writeEthernetHeaderToMem_CP_886_elements(13);
      gj_writeEthernetHeaderToMem_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Sample/ra
      -- 
    ra_1026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_981_inst_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	54 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/phi_stmt_979_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/RPIPE_nic_rx_to_header_981_Update/ca
      -- 
    ca_1031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_981_inst_ack_1, ack => writeEthernetHeaderToMem_CP_886_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Sample/crr
      -- 
    crr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(58), ack => call_stmt_1002_call_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(57) & writeEthernetHeaderToMem_CP_886_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_update_start_
      -- CP-element group 59: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Update/ccr
      -- 
    ccr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_886_elements(59), ack => call_stmt_1002_call_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_886_elements(61);
      gj_writeEthernetHeaderToMem_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	53 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Sample/cra
      -- 
    cra_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1002_call_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/call_stmt_1002_Update/cca
      -- 
    cca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1002_call_ack_1, ack => writeEthernetHeaderToMem_CP_886_elements(61)); -- 
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	9 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	10 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writeEthernetHeaderToMem_CP_886_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_886_elements(9), ack => writeEthernetHeaderToMem_CP_886_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	12 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	6 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_965/do_while_stmt_966/do_while_stmt_966_loop_body/$exit
      -- 
    writeEthernetHeaderToMem_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_886_elements(61) & writeEthernetHeaderToMem_CP_886_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	5 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_965/do_while_stmt_966/loop_exit/$exit
      -- CP-element group 64: 	 branch_block_stmt_965/do_while_stmt_966/loop_exit/ack
      -- 
    ack_1050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_966_branch_ack_0, ack => writeEthernetHeaderToMem_CP_886_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	5 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_965/do_while_stmt_966/loop_taken/$exit
      -- CP-element group 65: 	 branch_block_stmt_965/do_while_stmt_966/loop_taken/ack
      -- 
    ack_1054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_966_branch_ack_1, ack => writeEthernetHeaderToMem_CP_886_elements(65)); -- 
    -- CP-element group 66:  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	3 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	1 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_965/do_while_stmt_966/$exit
      -- 
    writeEthernetHeaderToMem_CP_886_elements(66) <= writeEthernetHeaderToMem_CP_886_elements(3);
    writeEthernetHeaderToMem_do_while_stmt_966_terminator_1055: loop_terminator -- 
      generic map (name => " writeEthernetHeaderToMem_do_while_stmt_966_terminator_1055", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeEthernetHeaderToMem_CP_886_elements(6),loop_continue => writeEthernetHeaderToMem_CP_886_elements(65),loop_terminate => writeEthernetHeaderToMem_CP_886_elements(64),loop_back => writeEthernetHeaderToMem_CP_886_elements(4),loop_exit => writeEthernetHeaderToMem_CP_886_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_968_phi_seq_969_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_886_elements(23);
      writeEthernetHeaderToMem_CP_886_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_886_elements(30);
      writeEthernetHeaderToMem_CP_886_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_886_elements(31);
      writeEthernetHeaderToMem_CP_886_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_886_elements(21);
      writeEthernetHeaderToMem_CP_886_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_886_elements(34);
      writeEthernetHeaderToMem_CP_886_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_886_elements(35);
      writeEthernetHeaderToMem_CP_886_elements(22) <= phi_mux_reqs(1);
      phi_stmt_968_phi_seq_969 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_968_phi_seq_969") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_886_elements(17), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_886_elements(18), 
          phi_update_req => writeEthernetHeaderToMem_CP_886_elements(19), 
          phi_update_ack => writeEthernetHeaderToMem_CP_886_elements(20), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_886_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_974_phi_seq_1013_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_886_elements(42);
      writeEthernetHeaderToMem_CP_886_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_886_elements(45);
      writeEthernetHeaderToMem_CP_886_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_886_elements(47);
      writeEthernetHeaderToMem_CP_886_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_886_elements(40);
      writeEthernetHeaderToMem_CP_886_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_886_elements(51);
      writeEthernetHeaderToMem_CP_886_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_886_elements(52);
      writeEthernetHeaderToMem_CP_886_elements(41) <= phi_mux_reqs(1);
      phi_stmt_974_phi_seq_1013 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_974_phi_seq_1013") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_886_elements(11), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_886_elements(38), 
          phi_update_req => writeEthernetHeaderToMem_CP_886_elements(13), 
          phi_update_ack => writeEthernetHeaderToMem_CP_886_elements(39), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_886_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_911_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeEthernetHeaderToMem_CP_886_elements(7);
        preds(1)  <= writeEthernetHeaderToMem_CP_886_elements(8);
        entry_tmerge_911 : transition_merge -- 
          generic map(name => " entry_tmerge_911")
          port map (preds => preds, symbol_out => writeEthernetHeaderToMem_CP_886_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_972_wire : std_logic_vector(35 downto 0);
    signal I_974 : std_logic_vector(3 downto 0);
    signal RPIPE_nic_rx_to_header_981_wire : std_logic_vector(72 downto 0);
    signal ULE_u4_u1_1016_wire : std_logic_vector(0 downto 0);
    signal ethernet_header_979 : std_logic_vector(72 downto 0);
    signal ignore_return_1002 : std_logic_vector(63 downto 0);
    signal konst_1005_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1010_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1015_wire_constant : std_logic_vector(3 downto 0);
    signal konst_971_wire_constant : std_logic_vector(35 downto 0);
    signal nI_1007 : std_logic_vector(3 downto 0);
    signal nI_1007_978_buffered : std_logic_vector(3 downto 0);
    signal nbuf_position_1012 : std_logic_vector(35 downto 0);
    signal nbuf_position_1012_973_buffered : std_logic_vector(35 downto 0);
    signal type_cast_977_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_995_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_989 : std_logic_vector(63 downto 0);
    signal wkeep_993 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1005_wire_constant <= "0001";
    konst_1010_wire_constant <= "000000000000000000000000000000001000";
    konst_1015_wire_constant <= "0001";
    konst_971_wire_constant <= "000000000000000000000000000000001000";
    type_cast_977_wire_constant <= "0000";
    type_cast_995_wire_constant <= "0";
    type_cast_997_wire_constant <= "0";
    phi_stmt_968: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_972_wire & nbuf_position_1012_973_buffered;
      req <= phi_stmt_968_req_0 & phi_stmt_968_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_968",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_968_ack_0,
          idata => idata,
          odata => buf_position_buffer,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_968
    phi_stmt_974: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_977_wire_constant & nI_1007_978_buffered;
      req <= phi_stmt_974_req_0 & phi_stmt_974_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_974",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_974_ack_0,
          idata => idata,
          odata => I_974,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_974
    -- flow-through slice operator slice_988_inst
    wdata_989 <= ethernet_header_979(71 downto 8);
    -- flow-through slice operator slice_992_inst
    wkeep_993 <= ethernet_header_979(7 downto 0);
    nI_1007_978_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_1007_978_buf_req_0;
      nI_1007_978_buf_ack_0<= wack(0);
      rreq(0) <= nI_1007_978_buf_req_1;
      nI_1007_978_buf_ack_1<= rack(0);
      nI_1007_978_buf : InterlockBuffer generic map ( -- 
        name => "nI_1007_978_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_1007,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_1007_978_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nbuf_position_1012_973_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nbuf_position_1012_973_buf_req_0;
      nbuf_position_1012_973_buf_ack_0<= wack(0);
      rreq(0) <= nbuf_position_1012_973_buf_req_1;
      nbuf_position_1012_973_buf_ack_1<= rack(0);
      nbuf_position_1012_973_buf : InterlockBuffer generic map ( -- 
        name => "nbuf_position_1012_973_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nbuf_position_1012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nbuf_position_1012_973_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_979
    process(RPIPE_nic_rx_to_header_981_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_header_981_wire(72 downto 0);
      ethernet_header_979 <= tmp_var; -- 
    end process;
    do_while_stmt_966_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULE_u4_u1_1016_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_966_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_966_branch_req_0,
          ack0 => do_while_stmt_966_branch_ack_0,
          ack1 => do_while_stmt_966_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u36_u36_1011_inst
    process(buf_position_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buf_position_buffer, konst_1010_wire_constant, tmp_var);
      nbuf_position_1012 <= tmp_var; --
    end process;
    -- shared split operator group (1) : ADD_u36_u36_972_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_972_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_972_inst_req_0;
      ADD_u36_u36_972_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_972_inst_req_1;
      ADD_u36_u36_972_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- binary operator ADD_u4_u4_1006_inst
    process(I_974) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_974, konst_1005_wire_constant, tmp_var);
      nI_1007 <= tmp_var; --
    end process;
    -- binary operator ULE_u4_u1_1016_inst
    process(nI_1007) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(nI_1007, konst_1015_wire_constant, tmp_var);
      ULE_u4_u1_1016_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_header_981_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_header_981_inst_req_0;
      RPIPE_nic_rx_to_header_981_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_header_981_inst_req_1;
      RPIPE_nic_rx_to_header_981_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_header_981_wire <= data_out(72 downto 0);
      nic_rx_to_header_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_header_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_header_pipe_read_req(0),
          oack => nic_rx_to_header_pipe_read_ack(0),
          odata => nic_rx_to_header_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1002_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1002_call_req_0;
      call_stmt_1002_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1002_call_req_1;
      call_stmt_1002_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_995_wire_constant & type_cast_997_wire_constant & wkeep_993 & buf_position_buffer & wdata_989;
      ignore_return_1002 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeEthernetHeaderToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writePayloadToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buf_pointer : in  std_logic_vector(35 downto 0);
    buf_pointer : in  std_logic_vector(35 downto 0);
    packet_size_32 : out  std_logic_vector(7 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    last_keep : out  std_logic_vector(7 downto 0);
    nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writePayloadToMem;
architecture writePayloadToMem_arch of writePayloadToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 17)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buf_pointer_update_enable: Boolean;
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal packet_size_32_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_32_update_enable: Boolean;
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  signal writePayloadToMem_CP_1056_start: Boolean;
  signal writePayloadToMem_CP_1056_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal phi_stmt_1028_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1038_inst_req_0 : boolean;
  signal ADD_u36_u36_1032_inst_req_1 : boolean;
  signal phi_stmt_1028_req_1 : boolean;
  signal do_while_stmt_1026_branch_req_0 : boolean;
  signal ADD_u36_u36_1035_inst_ack_0 : boolean;
  signal ADD_u36_u36_1035_inst_ack_1 : boolean;
  signal ADD_u36_u36_1035_inst_req_1 : boolean;
  signal ADD_u36_u36_1035_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1038_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1038_inst_ack_1 : boolean;
  signal ADD_u36_u36_1032_inst_ack_0 : boolean;
  signal ADD_u36_u36_1032_inst_ack_1 : boolean;
  signal phi_stmt_1028_req_0 : boolean;
  signal ADD_u36_u36_1032_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1038_inst_req_1 : boolean;
  signal do_while_stmt_1026_branch_ack_1 : boolean;
  signal do_while_stmt_1026_branch_ack_0 : boolean;
  signal call_stmt_1065_call_ack_1 : boolean;
  signal call_stmt_1065_call_req_1 : boolean;
  signal call_stmt_1065_call_ack_0 : boolean;
  signal call_stmt_1065_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writePayloadToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buf_pointer;
  base_buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(71 downto 36) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(71 downto 36);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writePayloadToMem_CP_1056_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writePayloadToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 17) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= packet_size_32_buffer;
  packet_size_32 <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(8 downto 8) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(8 downto 8);
  out_buffer_data_in(16 downto 9) <= last_keep_buffer;
  last_keep <= out_buffer_data_out(16 downto 9);
  out_buffer_data_in(tag_length + 16 downto 17) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 16 downto 17);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1056_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1056_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1056_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writePayloadToMem_CP_1056: Block -- control-path 
    signal writePayloadToMem_CP_1056_elements: BooleanArray(49 downto 0);
    -- 
  begin -- 
    writePayloadToMem_CP_1056_elements(0) <= writePayloadToMem_CP_1056_start;
    writePayloadToMem_CP_1056_symbol <= writePayloadToMem_CP_1056_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1025/$entry
      -- CP-element group 0: 	 branch_block_stmt_1025/do_while_stmt_1026__entry__
      -- CP-element group 0: 	 branch_block_stmt_1025/branch_block_stmt_1025__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	49 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1025/do_while_stmt_1026__exit__
      -- CP-element group 1: 	 branch_block_stmt_1025/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 assign_stmt_1078_to_assign_stmt_1093/$exit
      -- CP-element group 1: 	 assign_stmt_1078_to_assign_stmt_1093/$entry
      -- CP-element group 1: 	 branch_block_stmt_1025/branch_block_stmt_1025__exit__
      -- 
    writePayloadToMem_CP_1056_elements(1) <= writePayloadToMem_CP_1056_elements(49);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026__entry__
      -- CP-element group 2: 	 branch_block_stmt_1025/do_while_stmt_1026/$entry
      -- 
    writePayloadToMem_CP_1056_elements(2) <= writePayloadToMem_CP_1056_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	49 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026__exit__
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_back
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	47 
    -- CP-element group 5: 	48 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1025/do_while_stmt_1026/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_exit/$entry
      -- 
    writePayloadToMem_CP_1056_elements(5) <= writePayloadToMem_CP_1056_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	46 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_body_done
      -- 
    writePayloadToMem_CP_1056_elements(6) <= writePayloadToMem_CP_1056_elements(46);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/back_edge_to_loop_body
      -- 
    writePayloadToMem_CP_1056_elements(7) <= writePayloadToMem_CP_1056_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/first_time_through_loop_body
      -- 
    writePayloadToMem_CP_1056_elements(8) <= writePayloadToMem_CP_1056_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	45 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1036_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/loop_body_start
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	45 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/condition_evaluated
      -- 
    condition_evaluated_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(10), ack => do_while_stmt_1026_branch_req_0); -- 
    writePayloadToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(45) & writePayloadToMem_CP_1056_elements(14);
      gj_writePayloadToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	37 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_sample_start__ps
      -- 
    writePayloadToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(15) & writePayloadToMem_CP_1056_elements(9) & writePayloadToMem_CP_1056_elements(14);
      gj_writePayloadToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	39 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	46 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1036_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/aggregated_phi_sample_ack
      -- 
    writePayloadToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(17) & writePayloadToMem_CP_1056_elements(39);
      gj_writePayloadToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	36 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_update_start__ps
      -- 
    writePayloadToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(16) & writePayloadToMem_CP_1056_elements(36);
      gj_writePayloadToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	40 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/aggregated_phi_update_ack
      -- 
    writePayloadToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(18) & writePayloadToMem_CP_1056_elements(40);
      gj_writePayloadToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_sample_start_
      -- 
    writePayloadToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(9) & writePayloadToMem_CP_1056_elements(12);
      gj_writePayloadToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	43 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_update_start_
      -- 
    writePayloadToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(9) & writePayloadToMem_CP_1056_elements(43);
      gj_writePayloadToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_sample_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	41 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_update_completed_
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_loopback_trigger
      -- 
    writePayloadToMem_CP_1056_elements(19) <= writePayloadToMem_CP_1056_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_loopback_sample_req_ps
      -- 
    phi_stmt_1028_loopback_sample_req_1095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1028_loopback_sample_req_1095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(20), ack => phi_stmt_1028_req_1); -- 
    -- Element group writePayloadToMem_CP_1056_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_entry_trigger
      -- 
    writePayloadToMem_CP_1056_elements(21) <= writePayloadToMem_CP_1056_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_entry_sample_req
      -- 
    phi_stmt_1028_entry_sample_req_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1028_entry_sample_req_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(22), ack => phi_stmt_1028_req_0); -- 
    -- Element group writePayloadToMem_CP_1056_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1028_phi_mux_ack_ps
      -- 
    phi_stmt_1028_phi_mux_ack_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1028_ack_0, ack => writePayloadToMem_CP_1056_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_sample_start_
      -- 
    rr_1114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(26), ack => ADD_u36_u36_1032_inst_req_0); -- 
    writePayloadToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(24) & writePayloadToMem_CP_1056_elements(28);
      gj_writePayloadToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_update_start_
      -- 
    cr_1119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(27), ack => ADD_u36_u36_1032_inst_req_1); -- 
    writePayloadToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(25) & writePayloadToMem_CP_1056_elements(29);
      gj_writePayloadToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_sample_completed__ps
      -- 
    ra_1115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1032_inst_ack_0, ack => writePayloadToMem_CP_1056_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1032_update_completed__ps
      -- 
    ca_1120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1032_inst_ack_1, ack => writePayloadToMem_CP_1056_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Sample/$entry
      -- 
    rr_1132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(32), ack => ADD_u36_u36_1035_inst_req_0); -- 
    writePayloadToMem_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(30) & writePayloadToMem_CP_1056_elements(34);
      gj_writePayloadToMem_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Update/$entry
      -- 
    cr_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(33), ack => ADD_u36_u36_1035_inst_req_1); -- 
    writePayloadToMem_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(31) & writePayloadToMem_CP_1056_elements(35);
      gj_writePayloadToMem_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_sample_completed_
      -- 
    ra_1133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1035_inst_ack_0, ack => writePayloadToMem_CP_1056_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/ADD_u36_u36_1035_Update/$exit
      -- 
    ca_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1035_inst_ack_1, ack => writePayloadToMem_CP_1056_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	43 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	13 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1036_update_start_
      -- 
    writePayloadToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(9) & writePayloadToMem_CP_1056_elements(43);
      gj_writePayloadToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	40 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Sample/$entry
      -- 
    rr_1151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(37), ack => RPIPE_nic_rx_to_packet_1038_inst_req_0); -- 
    writePayloadToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(11) & writePayloadToMem_CP_1056_elements(40);
      gj_writePayloadToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: 	39 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_update_start_
      -- 
    cr_1156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(38), ack => RPIPE_nic_rx_to_packet_1038_inst_req_1); -- 
    writePayloadToMem_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(13) & writePayloadToMem_CP_1056_elements(39);
      gj_writePayloadToMem_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	12 
    -- CP-element group 39: 	38 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Sample/$exit
      -- 
    ra_1152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1038_inst_ack_0, ack => writePayloadToMem_CP_1056_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	14 
    -- CP-element group 40: 	41 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	37 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/phi_stmt_1036_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/RPIPE_nic_rx_to_packet_1038_update_completed_
      -- 
    ca_1157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1038_inst_ack_1, ack => writePayloadToMem_CP_1056_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: 	40 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Sample/crr
      -- 
    crr_1165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(41), ack => call_stmt_1065_call_req_0); -- 
    writePayloadToMem_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(18) & writePayloadToMem_CP_1056_elements(40) & writePayloadToMem_CP_1056_elements(43);
      gj_writePayloadToMem_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_update_start_
      -- CP-element group 42: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Update/ccr
      -- CP-element group 42: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Update/$entry
      -- 
    ccr_1170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1056_elements(42), ack => call_stmt_1065_call_req_1); -- 
    writePayloadToMem_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writePayloadToMem_CP_1056_elements(44);
      gj_writePayloadToMem_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	16 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Sample/cra
      -- 
    cra_1166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1065_call_ack_0, ack => writePayloadToMem_CP_1056_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Update/cca
      -- CP-element group 44: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/call_stmt_1065_Update/$exit
      -- 
    cca_1171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1065_call_ack_1, ack => writePayloadToMem_CP_1056_elements(44)); -- 
    -- CP-element group 45:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	9 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	10 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writePayloadToMem_CP_1056_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_1056_elements(9), ack => writePayloadToMem_CP_1056_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	12 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	6 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1025/do_while_stmt_1026/do_while_stmt_1026_loop_body/$exit
      -- 
    writePayloadToMem_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1056_elements(44) & writePayloadToMem_CP_1056_elements(12);
      gj_writePayloadToMem_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	5 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_exit/ack
      -- CP-element group 47: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_exit/$exit
      -- 
    ack_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1026_branch_ack_0, ack => writePayloadToMem_CP_1056_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	5 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_taken/ack
      -- CP-element group 48: 	 branch_block_stmt_1025/do_while_stmt_1026/loop_taken/$exit
      -- 
    ack_1180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1026_branch_ack_1, ack => writePayloadToMem_CP_1056_elements(48)); -- 
    -- CP-element group 49:  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	3 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	1 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1025/do_while_stmt_1026/$exit
      -- 
    writePayloadToMem_CP_1056_elements(49) <= writePayloadToMem_CP_1056_elements(3);
    writePayloadToMem_do_while_stmt_1026_terminator_1181: loop_terminator -- 
      generic map (name => " writePayloadToMem_do_while_stmt_1026_terminator_1181", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writePayloadToMem_CP_1056_elements(6),loop_continue => writePayloadToMem_CP_1056_elements(48),loop_terminate => writePayloadToMem_CP_1056_elements(47),loop_back => writePayloadToMem_CP_1056_elements(4),loop_exit => writePayloadToMem_CP_1056_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1028_phi_seq_1139_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writePayloadToMem_CP_1056_elements(21);
      writePayloadToMem_CP_1056_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writePayloadToMem_CP_1056_elements(28);
      writePayloadToMem_CP_1056_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writePayloadToMem_CP_1056_elements(29);
      writePayloadToMem_CP_1056_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writePayloadToMem_CP_1056_elements(19);
      writePayloadToMem_CP_1056_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writePayloadToMem_CP_1056_elements(34);
      writePayloadToMem_CP_1056_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writePayloadToMem_CP_1056_elements(35);
      writePayloadToMem_CP_1056_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1028_phi_seq_1139 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1028_phi_seq_1139") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writePayloadToMem_CP_1056_elements(11), 
          phi_sample_ack => writePayloadToMem_CP_1056_elements(17), 
          phi_update_req => writePayloadToMem_CP_1056_elements(13), 
          phi_update_ack => writePayloadToMem_CP_1056_elements(18), 
          phi_mux_ack => writePayloadToMem_CP_1056_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1081_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writePayloadToMem_CP_1056_elements(7);
        preds(1)  <= writePayloadToMem_CP_1056_elements(8);
        entry_tmerge_1081 : transition_merge -- 
          generic map(name => " entry_tmerge_1081")
          port map (preds => preds, symbol_out => writePayloadToMem_CP_1056_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1032_wire : std_logic_vector(35 downto 0);
    signal ADD_u36_u36_1035_wire : std_logic_vector(35 downto 0);
    signal EQ_u64_u1_1073_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1076_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1068_wire : std_logic_vector(0 downto 0);
    signal RPIPE_nic_rx_to_packet_1038_wire : std_logic_vector(72 downto 0);
    signal R_BAD_PACKET_DATA_1072_wire_constant : std_logic_vector(63 downto 0);
    signal SUB_u36_u36_1082_wire : std_logic_vector(35 downto 0);
    signal buf_position_1028 : std_logic_vector(35 downto 0);
    signal ignore_return_1065 : std_logic_vector(63 downto 0);
    signal konst_1031_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1034_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1075_wire_constant : std_logic_vector(7 downto 0);
    signal last_bit_1043 : std_logic_vector(0 downto 0);
    signal packet_size_8_1084 : std_logic_vector(7 downto 0);
    signal payload_data_1036 : std_logic_vector(72 downto 0);
    signal type_cast_1058_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1060_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_1047 : std_logic_vector(63 downto 0);
    signal wkeep_1051 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_BAD_PACKET_DATA_1072_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    konst_1031_wire_constant <= "000000000000000000000000000000001000";
    konst_1034_wire_constant <= "000000000000000000000000000000001000";
    konst_1075_wire_constant <= "00000000";
    type_cast_1058_wire_constant <= "0";
    type_cast_1060_wire_constant <= "0";
    phi_stmt_1028: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_1032_wire & ADD_u36_u36_1035_wire;
      req <= phi_stmt_1028_req_0 & phi_stmt_1028_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1028",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1028_ack_0,
          idata => idata,
          odata => buf_position_1028,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1028
    -- flow-through slice operator slice_1042_inst
    last_bit_1043 <= payload_data_1036(72 downto 72);
    -- flow-through slice operator slice_1046_inst
    wdata_1047 <= payload_data_1036(71 downto 8);
    -- flow-through slice operator slice_1050_inst
    wkeep_1051 <= payload_data_1036(7 downto 0);
    -- interlock W_last_keep_1091_inst
    process(wkeep_1051) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := wkeep_1051(7 downto 0);
      last_keep_buffer <= tmp_var; -- 
    end process;
    -- interlock W_packet_size_32_1085_inst
    process(packet_size_8_1084) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := packet_size_8_1084(7 downto 0);
      packet_size_32_buffer <= tmp_var; -- 
    end process;
    -- interlock ssrc_phi_stmt_1036
    process(RPIPE_nic_rx_to_packet_1038_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_packet_1038_wire(72 downto 0);
      payload_data_1036 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1083_inst
    process(SUB_u36_u36_1082_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u36_u36_1082_wire(7 downto 0);
      packet_size_8_1084 <= tmp_var; -- 
    end process;
    do_while_stmt_1026_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1068_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1026_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1026_branch_req_0,
          ack0 => do_while_stmt_1026_branch_ack_0,
          ack1 => do_while_stmt_1026_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1032_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_1032_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1032_inst_req_0;
      ADD_u36_u36_1032_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1032_inst_req_1;
      ADD_u36_u36_1032_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u36_u36_1035_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_position_1028;
      ADD_u36_u36_1035_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1035_inst_req_0;
      ADD_u36_u36_1035_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1035_inst_req_1;
      ADD_u36_u36_1035_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- binary operator AND_u1_u1_1077_inst
    process(EQ_u64_u1_1073_wire, EQ_u8_u1_1076_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u64_u1_1073_wire, EQ_u8_u1_1076_wire, tmp_var);
      bad_packet_identifier_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1073_inst
    process(wdata_1047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wdata_1047, R_BAD_PACKET_DATA_1072_wire_constant, tmp_var);
      EQ_u64_u1_1073_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1076_inst
    process(wkeep_1051) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wkeep_1051, konst_1075_wire_constant, tmp_var);
      EQ_u8_u1_1076_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1068_inst
    process(last_bit_1043) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_1043, tmp_var);
      NOT_u1_u1_1068_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u36_u36_1082_inst
    process(buf_position_1028, base_buf_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(buf_position_1028, base_buf_pointer_buffer, tmp_var);
      SUB_u36_u36_1082_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_packet_1038_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_packet_1038_inst_req_0;
      RPIPE_nic_rx_to_packet_1038_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_packet_1038_inst_req_1;
      RPIPE_nic_rx_to_packet_1038_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_packet_1038_wire <= data_out(72 downto 0);
      nic_rx_to_packet_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_packet_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_packet_pipe_read_req(0),
          oack => nic_rx_to_packet_pipe_read_ack(0),
          odata => nic_rx_to_packet_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1065_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1065_call_req_0;
      call_stmt_1065_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1065_call_req_1;
      call_stmt_1065_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1058_wire_constant & type_cast_1060_wire_constant & wkeep_1051 & buf_position_1028 & wdata_1047;
      ignore_return_1065 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writePayloadToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    AFB_NIC_REQUEST_pipe_write_data: in std_logic_vector(73 downto 0);
    AFB_NIC_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
    AFB_NIC_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_data: in std_logic_vector(72 downto 0);
    mac_to_nic_data_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_data: out std_logic_vector(72 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(11 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(5 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module AccessRegister
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module AccessRegister
  signal AccessRegister_rwbar :  std_logic_vector(0 downto 0);
  signal AccessRegister_bmask :  std_logic_vector(3 downto 0);
  signal AccessRegister_register_index :  std_logic_vector(5 downto 0);
  signal AccessRegister_wdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_rdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_in_args    : std_logic_vector(42 downto 0);
  signal AccessRegister_out_args   : std_logic_vector(31 downto 0);
  signal AccessRegister_tag_in    : std_logic_vector(4 downto 0) := (others => '0');
  signal AccessRegister_tag_out   : std_logic_vector(4 downto 0);
  signal AccessRegister_start_req : std_logic;
  signal AccessRegister_start_ack : std_logic;
  signal AccessRegister_fin_req   : std_logic;
  signal AccessRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module AccessRegister
  signal AccessRegister_call_reqs: std_logic_vector(5 downto 0);
  signal AccessRegister_call_acks: std_logic_vector(5 downto 0);
  signal AccessRegister_return_reqs: std_logic_vector(5 downto 0);
  signal AccessRegister_return_acks: std_logic_vector(5 downto 0);
  signal AccessRegister_call_data: std_logic_vector(257 downto 0);
  signal AccessRegister_call_tag: std_logic_vector(11 downto 0);
  signal AccessRegister_return_data: std_logic_vector(191 downto 0);
  signal AccessRegister_return_tag: std_logic_vector(11 downto 0);
  -- declarations related to module NicRegisterAccessDaemon
  component NicRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module NicRegisterAccessDaemon
  signal NicRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal NicRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal NicRegisterAccessDaemon_start_req : std_logic;
  signal NicRegisterAccessDaemon_start_ack : std_logic;
  signal NicRegisterAccessDaemon_fin_req   : std_logic;
  signal NicRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module ReceiveEngineDaemon
  component ReceiveEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_call_data : out  std_logic_vector(35 downto 0);
      loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
      loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_return_data : in   std_logic_vector(0 downto 0);
      loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
      populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ReceiveEngineDaemon
  signal ReceiveEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ReceiveEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal ReceiveEngineDaemon_start_req : std_logic;
  signal ReceiveEngineDaemon_start_ack : std_logic;
  signal ReceiveEngineDaemon_fin_req   : std_logic;
  signal ReceiveEngineDaemon_fin_ack : std_logic;
  -- declarations related to module SoftwareRegisterAccessDaemon
  component SoftwareRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
      CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
      AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
      NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module SoftwareRegisterAccessDaemon
  signal SoftwareRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal SoftwareRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal SoftwareRegisterAccessDaemon_start_req : std_logic;
  signal SoftwareRegisterAccessDaemon_start_ack : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_req   : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module UpdateRegister
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module UpdateRegister
  signal UpdateRegister_bmask :  std_logic_vector(3 downto 0);
  signal UpdateRegister_rval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_wdata :  std_logic_vector(31 downto 0);
  signal UpdateRegister_index :  std_logic_vector(5 downto 0);
  signal UpdateRegister_wval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_in_args    : std_logic_vector(73 downto 0);
  signal UpdateRegister_out_args   : std_logic_vector(31 downto 0);
  signal UpdateRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal UpdateRegister_tag_out   : std_logic_vector(2 downto 0);
  signal UpdateRegister_start_req : std_logic;
  signal UpdateRegister_start_ack : std_logic;
  signal UpdateRegister_fin_req   : std_logic;
  signal UpdateRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module UpdateRegister
  signal UpdateRegister_call_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_data: std_logic_vector(147 downto 0);
  signal UpdateRegister_call_tag: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_data: std_logic_vector(63 downto 0);
  signal UpdateRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMemory
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemory
  signal accessMemory_lock :  std_logic_vector(0 downto 0);
  signal accessMemory_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemory_bmask :  std_logic_vector(7 downto 0);
  signal accessMemory_addr :  std_logic_vector(35 downto 0);
  signal accessMemory_wdata :  std_logic_vector(63 downto 0);
  signal accessMemory_rdata :  std_logic_vector(63 downto 0);
  signal accessMemory_in_args    : std_logic_vector(109 downto 0);
  signal accessMemory_out_args   : std_logic_vector(63 downto 0);
  signal accessMemory_tag_in    : std_logic_vector(6 downto 0) := (others => '0');
  signal accessMemory_tag_out   : std_logic_vector(6 downto 0);
  signal accessMemory_start_req : std_logic;
  signal accessMemory_start_ack : std_logic;
  signal accessMemory_fin_req   : std_logic;
  signal accessMemory_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemory
  signal accessMemory_call_reqs: std_logic_vector(13 downto 0);
  signal accessMemory_call_acks: std_logic_vector(13 downto 0);
  signal accessMemory_return_reqs: std_logic_vector(13 downto 0);
  signal accessMemory_return_acks: std_logic_vector(13 downto 0);
  signal accessMemory_call_data: std_logic_vector(1539 downto 0);
  signal accessMemory_call_tag: std_logic_vector(41 downto 0);
  signal accessMemory_return_data: std_logic_vector(895 downto 0);
  signal accessMemory_return_tag: std_logic_vector(41 downto 0);
  -- declarations related to module acquireLock
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module acquireLock
  signal acquireLock_q_base_address :  std_logic_vector(35 downto 0);
  signal acquireLock_m_ok :  std_logic_vector(0 downto 0);
  signal acquireLock_in_args    : std_logic_vector(35 downto 0);
  signal acquireLock_out_args   : std_logic_vector(0 downto 0);
  signal acquireLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal acquireLock_tag_out   : std_logic_vector(2 downto 0);
  signal acquireLock_start_req : std_logic;
  signal acquireLock_start_ack : std_logic;
  signal acquireLock_fin_req   : std_logic;
  signal acquireLock_fin_ack : std_logic;
  -- caller side aggregated signals for module acquireLock
  signal acquireLock_call_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_call_acks: std_logic_vector(1 downto 0);
  signal acquireLock_return_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_return_acks: std_logic_vector(1 downto 0);
  signal acquireLock_call_data: std_logic_vector(71 downto 0);
  signal acquireLock_call_tag: std_logic_vector(1 downto 0);
  signal acquireLock_return_data: std_logic_vector(1 downto 0);
  signal acquireLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module delay_time
  -- declarations related to module getQueueElement
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueElement
  signal getQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueElement_read_index :  std_logic_vector(31 downto 0);
  signal getQueueElement_q_r_data :  std_logic_vector(31 downto 0);
  signal getQueueElement_in_args    : std_logic_vector(67 downto 0);
  signal getQueueElement_out_args   : std_logic_vector(31 downto 0);
  signal getQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal getQueueElement_start_req : std_logic;
  signal getQueueElement_start_ack : std_logic;
  signal getQueueElement_fin_req   : std_logic;
  signal getQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueElement
  signal getQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_call_data: std_logic_vector(67 downto 0);
  signal getQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal getQueueElement_return_data: std_logic_vector(31 downto 0);
  signal getQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module getQueueLength
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueLength
  signal getQueueLength_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueLength_Queue_Length :  std_logic_vector(31 downto 0);
  signal getQueueLength_in_args    : std_logic_vector(35 downto 0);
  signal getQueueLength_out_args   : std_logic_vector(31 downto 0);
  signal getQueueLength_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueueLength_tag_out   : std_logic_vector(2 downto 0);
  signal getQueueLength_start_req : std_logic;
  signal getQueueLength_start_ack : std_logic;
  signal getQueueLength_fin_req   : std_logic;
  signal getQueueLength_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueLength
  signal getQueueLength_call_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_call_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_return_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_return_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_call_data: std_logic_vector(71 downto 0);
  signal getQueueLength_call_tag: std_logic_vector(1 downto 0);
  signal getQueueLength_return_data: std_logic_vector(63 downto 0);
  signal getQueueLength_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getQueuePointers
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointers
  signal getQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_in_args    : std_logic_vector(35 downto 0);
  signal getQueuePointers_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointers_start_req : std_logic;
  signal getQueuePointers_start_ack : std_logic;
  signal getQueuePointers_fin_req   : std_logic;
  signal getQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointers
  signal getQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_data: std_logic_vector(71 downto 0);
  signal getQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTotalMessages
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTotalMessages
  signal getTotalMessages_q_base_address :  std_logic_vector(35 downto 0);
  signal getTotalMessages_total_msgs :  std_logic_vector(31 downto 0);
  signal getTotalMessages_in_args    : std_logic_vector(35 downto 0);
  signal getTotalMessages_out_args   : std_logic_vector(31 downto 0);
  signal getTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal getTotalMessages_start_req : std_logic;
  signal getTotalMessages_start_ack : std_logic;
  signal getTotalMessages_fin_req   : std_logic;
  signal getTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module getTotalMessages
  signal getTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_data: std_logic_vector(71 downto 0);
  signal getTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_data: std_logic_vector(63 downto 0);
  signal getTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTxPacketPointerFromServer
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_queue_index :  std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_pkt_pointer :  std_logic_vector(31 downto 0);
  signal getTxPacketPointerFromServer_status :  std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_in_args    : std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_out_args   : std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getTxPacketPointerFromServer_tag_out   : std_logic_vector(1 downto 0);
  signal getTxPacketPointerFromServer_start_req : std_logic;
  signal getTxPacketPointerFromServer_start_ack : std_logic;
  signal getTxPacketPointerFromServer_fin_req   : std_logic;
  signal getTxPacketPointerFromServer_fin_ack : std_logic;
  -- caller side aggregated signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_call_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_data: std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_call_tag: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_data: std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module loadBuffer
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadBuffer
  signal loadBuffer_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal loadBuffer_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal loadBuffer_in_args    : std_logic_vector(35 downto 0);
  signal loadBuffer_out_args   : std_logic_vector(0 downto 0);
  signal loadBuffer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadBuffer_tag_out   : std_logic_vector(1 downto 0);
  signal loadBuffer_start_req : std_logic;
  signal loadBuffer_start_ack : std_logic;
  signal loadBuffer_fin_req   : std_logic;
  signal loadBuffer_fin_ack : std_logic;
  -- caller side aggregated signals for module loadBuffer
  signal loadBuffer_call_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_call_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_return_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_return_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_call_data: std_logic_vector(35 downto 0);
  signal loadBuffer_call_tag: std_logic_vector(0 downto 0);
  signal loadBuffer_return_data: std_logic_vector(0 downto 0);
  signal loadBuffer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module nextLSTATE
  -- declarations related to module nicRxFromMacDaemon
  component nicRxFromMacDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
      nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(1 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(1 downto 0);
      AccessRegister_call_data : out  std_logic_vector(85 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(1 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(1 downto 0);
      AccessRegister_return_data : in   std_logic_vector(63 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicRxFromMacDaemon
  signal nicRxFromMacDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicRxFromMacDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal nicRxFromMacDaemon_start_req : std_logic;
  signal nicRxFromMacDaemon_start_ack : std_logic;
  signal nicRxFromMacDaemon_fin_req   : std_logic;
  signal nicRxFromMacDaemon_fin_ack : std_logic;
  -- declarations related to module popFromQueue
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module popFromQueue
  signal popFromQueue_lock :  std_logic_vector(0 downto 0);
  signal popFromQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal popFromQueue_q_r_data :  std_logic_vector(31 downto 0);
  signal popFromQueue_status :  std_logic_vector(0 downto 0);
  signal popFromQueue_in_args    : std_logic_vector(36 downto 0);
  signal popFromQueue_out_args   : std_logic_vector(32 downto 0);
  signal popFromQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal popFromQueue_tag_out   : std_logic_vector(2 downto 0);
  signal popFromQueue_start_req : std_logic;
  signal popFromQueue_start_ack : std_logic;
  signal popFromQueue_fin_req   : std_logic;
  signal popFromQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module popFromQueue
  signal popFromQueue_call_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_call_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_return_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_return_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_call_data: std_logic_vector(73 downto 0);
  signal popFromQueue_call_tag: std_logic_vector(1 downto 0);
  signal popFromQueue_return_data: std_logic_vector(65 downto 0);
  signal popFromQueue_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module populateRxQueue
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module populateRxQueue
  signal populateRxQueue_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal populateRxQueue_in_args    : std_logic_vector(35 downto 0);
  signal populateRxQueue_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal populateRxQueue_tag_out   : std_logic_vector(1 downto 0);
  signal populateRxQueue_start_req : std_logic;
  signal populateRxQueue_start_ack : std_logic;
  signal populateRxQueue_fin_req   : std_logic;
  signal populateRxQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module populateRxQueue
  signal populateRxQueue_call_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_data: std_logic_vector(35 downto 0);
  signal populateRxQueue_call_tag: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module pushIntoQueue
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module pushIntoQueue
  signal pushIntoQueue_lock :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal pushIntoQueue_q_w_data :  std_logic_vector(31 downto 0);
  signal pushIntoQueue_status :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_in_args    : std_logic_vector(68 downto 0);
  signal pushIntoQueue_out_args   : std_logic_vector(0 downto 0);
  signal pushIntoQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal pushIntoQueue_tag_out   : std_logic_vector(2 downto 0);
  signal pushIntoQueue_start_req : std_logic;
  signal pushIntoQueue_start_ack : std_logic;
  signal pushIntoQueue_fin_req   : std_logic;
  signal pushIntoQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module pushIntoQueue
  signal pushIntoQueue_call_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_data: std_logic_vector(206 downto 0);
  signal pushIntoQueue_call_tag: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_data: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module releaseLock
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module releaseLock
  signal releaseLock_q_base_address :  std_logic_vector(35 downto 0);
  signal releaseLock_in_args    : std_logic_vector(35 downto 0);
  signal releaseLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal releaseLock_tag_out   : std_logic_vector(2 downto 0);
  signal releaseLock_start_req : std_logic;
  signal releaseLock_start_ack : std_logic;
  signal releaseLock_fin_req   : std_logic;
  signal releaseLock_fin_ack : std_logic;
  -- caller side aggregated signals for module releaseLock
  signal releaseLock_call_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_call_acks: std_logic_vector(1 downto 0);
  signal releaseLock_return_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_return_acks: std_logic_vector(1 downto 0);
  signal releaseLock_call_data: std_logic_vector(71 downto 0);
  signal releaseLock_call_tag: std_logic_vector(1 downto 0);
  signal releaseLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setQueueElement
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueueElement
  signal setQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueueElement_write_index :  std_logic_vector(31 downto 0);
  signal setQueueElement_q_w_data :  std_logic_vector(31 downto 0);
  signal setQueueElement_in_args    : std_logic_vector(99 downto 0);
  signal setQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal setQueueElement_start_req : std_logic;
  signal setQueueElement_start_ack : std_logic;
  signal setQueueElement_fin_req   : std_logic;
  signal setQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueueElement
  signal setQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_call_data: std_logic_vector(99 downto 0);
  signal setQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal setQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueuePointers
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueuePointers
  signal setQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_in_args    : std_logic_vector(99 downto 0);
  signal setQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal setQueuePointers_start_req : std_logic;
  signal setQueuePointers_start_ack : std_logic;
  signal setQueuePointers_fin_req   : std_logic;
  signal setQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueuePointers
  signal setQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_data: std_logic_vector(199 downto 0);
  signal setQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module transmitEngineDaemon
  component transmitEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
      getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
      getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
      transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_call_data : out  std_logic_vector(31 downto 0);
      transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
      transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_return_data : in   std_logic_vector(0 downto 0);
      transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitEngineDaemon
  signal transmitEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal transmitEngineDaemon_start_req : std_logic;
  signal transmitEngineDaemon_start_ack : std_logic;
  signal transmitEngineDaemon_fin_req   : std_logic;
  signal transmitEngineDaemon_fin_ack : std_logic;
  -- declarations related to module transmitPacket
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitPacket
  signal transmitPacket_packet_pointer :  std_logic_vector(31 downto 0);
  signal transmitPacket_status :  std_logic_vector(0 downto 0);
  signal transmitPacket_in_args    : std_logic_vector(31 downto 0);
  signal transmitPacket_out_args   : std_logic_vector(0 downto 0);
  signal transmitPacket_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitPacket_tag_out   : std_logic_vector(1 downto 0);
  signal transmitPacket_start_req : std_logic;
  signal transmitPacket_start_ack : std_logic;
  signal transmitPacket_fin_req   : std_logic;
  signal transmitPacket_fin_ack : std_logic;
  -- caller side aggregated signals for module transmitPacket
  signal transmitPacket_call_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_call_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_return_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_return_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_call_data: std_logic_vector(31 downto 0);
  signal transmitPacket_call_tag: std_logic_vector(0 downto 0);
  signal transmitPacket_return_data: std_logic_vector(0 downto 0);
  signal transmitPacket_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module updateTotalMessages
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module updateTotalMessages
  signal updateTotalMessages_q_base_address :  std_logic_vector(35 downto 0);
  signal updateTotalMessages_updated_total_msgs :  std_logic_vector(31 downto 0);
  signal updateTotalMessages_in_args    : std_logic_vector(67 downto 0);
  signal updateTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal updateTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal updateTotalMessages_start_req : std_logic;
  signal updateTotalMessages_start_ack : std_logic;
  signal updateTotalMessages_fin_req   : std_logic;
  signal updateTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module updateTotalMessages
  signal updateTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal updateTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal updateTotalMessages_call_data: std_logic_vector(135 downto 0);
  signal updateTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module writeControlInformationToMem
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeControlInformationToMem
  signal writeControlInformationToMem_base_buffer_pointer :  std_logic_vector(35 downto 0);
  signal writeControlInformationToMem_packet_size :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_in_args    : std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeControlInformationToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeControlInformationToMem_start_req : std_logic;
  signal writeControlInformationToMem_start_ack : std_logic;
  signal writeControlInformationToMem_fin_req   : std_logic;
  signal writeControlInformationToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeControlInformationToMem
  signal writeControlInformationToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_data: std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeEthernetHeaderToMem
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_buf_position :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_in_args    : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_out_args   : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeEthernetHeaderToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeEthernetHeaderToMem_start_req : std_logic;
  signal writeEthernetHeaderToMem_start_ack : std_logic;
  signal writeEthernetHeaderToMem_fin_req   : std_logic;
  signal writeEthernetHeaderToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writePayloadToMem
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writePayloadToMem
  signal writePayloadToMem_base_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_packet_size_32 :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal writePayloadToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_in_args    : std_logic_vector(71 downto 0);
  signal writePayloadToMem_out_args   : std_logic_vector(16 downto 0);
  signal writePayloadToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writePayloadToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writePayloadToMem_start_req : std_logic;
  signal writePayloadToMem_start_ack : std_logic;
  signal writePayloadToMem_fin_req   : std_logic;
  signal writePayloadToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writePayloadToMem
  signal writePayloadToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_data: std_logic_vector(71 downto 0);
  signal writePayloadToMem_call_tag: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_data: std_logic_vector(16 downto 0);
  signal writePayloadToMem_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_read_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_write_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe CONTROL_REGISTER
  signal CONTROL_REGISTER_pipe_write_data: std_logic_vector(31 downto 0);
  signal CONTROL_REGISTER_pipe_write_req: std_logic_vector(0 downto 0);
  signal CONTROL_REGISTER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe CONTROL_REGISTER
  signal CONTROL_REGISTER: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe FREE_Q
  signal FREE_Q_pipe_write_data: std_logic_vector(35 downto 0);
  signal FREE_Q_pipe_write_req: std_logic_vector(0 downto 0);
  signal FREE_Q_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe FREE_Q
  signal FREE_Q: std_logic_vector(35 downto 0);
  -- aggregate signals for write to pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for read from pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS_pipe_write_data: std_logic_vector(31 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_req: std_logic_vector(0 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS: std_logic_vector(31 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_read_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_write_data: std_logic_vector(145 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module AccessRegister
  AccessRegister_rwbar <= AccessRegister_in_args(42 downto 42);
  AccessRegister_bmask <= AccessRegister_in_args(41 downto 38);
  AccessRegister_register_index <= AccessRegister_in_args(37 downto 32);
  AccessRegister_wdata <= AccessRegister_in_args(31 downto 0);
  AccessRegister_out_args <= AccessRegister_rdata ;
  -- call arbiter for module AccessRegister
  AccessRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 6,
      call_data_width => 43,
      return_data_width => 32,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => AccessRegister_call_reqs,
      call_acks => AccessRegister_call_acks,
      return_reqs => AccessRegister_return_reqs,
      return_acks => AccessRegister_return_acks,
      call_data  => AccessRegister_call_data,
      call_tag  => AccessRegister_call_tag,
      return_tag  => AccessRegister_return_tag,
      call_mtag => AccessRegister_tag_in,
      return_mtag => AccessRegister_tag_out,
      return_data =>AccessRegister_return_data,
      call_mreq => AccessRegister_start_req,
      call_mack => AccessRegister_start_ack,
      return_mreq => AccessRegister_fin_req,
      return_mack => AccessRegister_fin_ack,
      call_mdata => AccessRegister_in_args,
      return_mdata => AccessRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  AccessRegister_instance:AccessRegister-- 
    generic map(tag_length => 5)
    port map(-- 
      rwbar => AccessRegister_rwbar,
      bmask => AccessRegister_bmask,
      register_index => AccessRegister_register_index,
      wdata => AccessRegister_wdata,
      rdata => AccessRegister_rdata,
      start_req => AccessRegister_start_req,
      start_ack => AccessRegister_start_ack,
      fin_req => AccessRegister_fin_req,
      fin_ack => AccessRegister_fin_ack,
      clk => clk,
      reset => reset,
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
      tag_in => AccessRegister_tag_in,
      tag_out => AccessRegister_tag_out-- 
    ); -- 
  -- module NicRegisterAccessDaemon
  NicRegisterAccessDaemon_instance:NicRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => NicRegisterAccessDaemon_start_req,
      start_ack => NicRegisterAccessDaemon_start_ack,
      fin_req => NicRegisterAccessDaemon_fin_req,
      fin_ack => NicRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(11 downto 6),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(1 downto 1),
      UpdateRegister_call_acks => UpdateRegister_call_acks(1 downto 1),
      UpdateRegister_call_data => UpdateRegister_call_data(147 downto 74),
      UpdateRegister_call_tag => UpdateRegister_call_tag(1 downto 1),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(1 downto 1),
      UpdateRegister_return_acks => UpdateRegister_return_acks(1 downto 1),
      UpdateRegister_return_data => UpdateRegister_return_data(63 downto 32),
      UpdateRegister_return_tag => UpdateRegister_return_tag(1 downto 1),
      tag_in => NicRegisterAccessDaemon_tag_in,
      tag_out => NicRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  NicRegisterAccessDaemon_tag_in <= (others => '0');
  NicRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => NicRegisterAccessDaemon_start_req, start_ack => NicRegisterAccessDaemon_start_ack,  fin_req => NicRegisterAccessDaemon_fin_req,  fin_ack => NicRegisterAccessDaemon_fin_ack);
  -- module ReceiveEngineDaemon
  ReceiveEngineDaemon_instance:ReceiveEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ReceiveEngineDaemon_start_req,
      start_ack => ReceiveEngineDaemon_start_ack,
      fin_req => ReceiveEngineDaemon_fin_req,
      fin_ack => ReceiveEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      FREE_Q => FREE_Q,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(3 downto 3),
      AccessRegister_call_acks => AccessRegister_call_acks(3 downto 3),
      AccessRegister_call_data => AccessRegister_call_data(171 downto 129),
      AccessRegister_call_tag => AccessRegister_call_tag(7 downto 6),
      AccessRegister_return_reqs => AccessRegister_return_reqs(3 downto 3),
      AccessRegister_return_acks => AccessRegister_return_acks(3 downto 3),
      AccessRegister_return_data => AccessRegister_return_data(127 downto 96),
      AccessRegister_return_tag => AccessRegister_return_tag(7 downto 6),
      popFromQueue_call_reqs => popFromQueue_call_reqs(0 downto 0),
      popFromQueue_call_acks => popFromQueue_call_acks(0 downto 0),
      popFromQueue_call_data => popFromQueue_call_data(36 downto 0),
      popFromQueue_call_tag => popFromQueue_call_tag(0 downto 0),
      popFromQueue_return_reqs => popFromQueue_return_reqs(0 downto 0),
      popFromQueue_return_acks => popFromQueue_return_acks(0 downto 0),
      popFromQueue_return_data => popFromQueue_return_data(32 downto 0),
      popFromQueue_return_tag => popFromQueue_return_tag(0 downto 0),
      loadBuffer_call_reqs => loadBuffer_call_reqs(0 downto 0),
      loadBuffer_call_acks => loadBuffer_call_acks(0 downto 0),
      loadBuffer_call_data => loadBuffer_call_data(35 downto 0),
      loadBuffer_call_tag => loadBuffer_call_tag(0 downto 0),
      loadBuffer_return_reqs => loadBuffer_return_reqs(0 downto 0),
      loadBuffer_return_acks => loadBuffer_return_acks(0 downto 0),
      loadBuffer_return_data => loadBuffer_return_data(0 downto 0),
      loadBuffer_return_tag => loadBuffer_return_tag(0 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(1 downto 1),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(1 downto 1),
      pushIntoQueue_call_data => pushIntoQueue_call_data(137 downto 69),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(1 downto 1),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(1 downto 1),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(1 downto 1),
      pushIntoQueue_return_data => pushIntoQueue_return_data(1 downto 1),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(1 downto 1),
      populateRxQueue_call_reqs => populateRxQueue_call_reqs(0 downto 0),
      populateRxQueue_call_acks => populateRxQueue_call_acks(0 downto 0),
      populateRxQueue_call_data => populateRxQueue_call_data(35 downto 0),
      populateRxQueue_call_tag => populateRxQueue_call_tag(0 downto 0),
      populateRxQueue_return_reqs => populateRxQueue_return_reqs(0 downto 0),
      populateRxQueue_return_acks => populateRxQueue_return_acks(0 downto 0),
      populateRxQueue_return_tag => populateRxQueue_return_tag(0 downto 0),
      tag_in => ReceiveEngineDaemon_tag_in,
      tag_out => ReceiveEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  ReceiveEngineDaemon_tag_in <= (others => '0');
  ReceiveEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ReceiveEngineDaemon_start_req, start_ack => ReceiveEngineDaemon_start_ack,  fin_req => ReceiveEngineDaemon_fin_req,  fin_ack => ReceiveEngineDaemon_fin_ack);
  -- module SoftwareRegisterAccessDaemon
  SoftwareRegisterAccessDaemon_instance:SoftwareRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => SoftwareRegisterAccessDaemon_start_req,
      start_ack => SoftwareRegisterAccessDaemon_start_ack,
      fin_req => SoftwareRegisterAccessDaemon_fin_req,
      fin_ack => SoftwareRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(5 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      AFB_NIC_REQUEST_pipe_read_req => AFB_NIC_REQUEST_pipe_read_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_ack => AFB_NIC_REQUEST_pipe_read_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_data => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
      CONTROL_REGISTER_pipe_write_req => CONTROL_REGISTER_pipe_write_req(0 downto 0),
      CONTROL_REGISTER_pipe_write_ack => CONTROL_REGISTER_pipe_write_ack(0 downto 0),
      CONTROL_REGISTER_pipe_write_data => CONTROL_REGISTER_pipe_write_data(31 downto 0),
      FREE_Q_pipe_write_req => FREE_Q_pipe_write_req(0 downto 0),
      FREE_Q_pipe_write_ack => FREE_Q_pipe_write_ack(0 downto 0),
      FREE_Q_pipe_write_data => FREE_Q_pipe_write_data(35 downto 0),
      AFB_NIC_RESPONSE_pipe_write_req => AFB_NIC_RESPONSE_pipe_write_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_ack => AFB_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_data => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
      NUMBER_OF_SERVERS_pipe_write_req => NUMBER_OF_SERVERS_pipe_write_req(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_ack => NUMBER_OF_SERVERS_pipe_write_ack(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_data => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(0 downto 0),
      UpdateRegister_call_acks => UpdateRegister_call_acks(0 downto 0),
      UpdateRegister_call_data => UpdateRegister_call_data(73 downto 0),
      UpdateRegister_call_tag => UpdateRegister_call_tag(0 downto 0),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(0 downto 0),
      UpdateRegister_return_acks => UpdateRegister_return_acks(0 downto 0),
      UpdateRegister_return_data => UpdateRegister_return_data(31 downto 0),
      UpdateRegister_return_tag => UpdateRegister_return_tag(0 downto 0),
      tag_in => SoftwareRegisterAccessDaemon_tag_in,
      tag_out => SoftwareRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  SoftwareRegisterAccessDaemon_tag_in <= (others => '0');
  SoftwareRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => SoftwareRegisterAccessDaemon_start_req, start_ack => SoftwareRegisterAccessDaemon_start_ack,  fin_req => SoftwareRegisterAccessDaemon_fin_req,  fin_ack => SoftwareRegisterAccessDaemon_fin_ack);
  -- module UpdateRegister
  UpdateRegister_bmask <= UpdateRegister_in_args(73 downto 70);
  UpdateRegister_rval <= UpdateRegister_in_args(69 downto 38);
  UpdateRegister_wdata <= UpdateRegister_in_args(37 downto 6);
  UpdateRegister_index <= UpdateRegister_in_args(5 downto 0);
  UpdateRegister_out_args <= UpdateRegister_wval ;
  -- call arbiter for module UpdateRegister
  UpdateRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 74,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => UpdateRegister_call_reqs,
      call_acks => UpdateRegister_call_acks,
      return_reqs => UpdateRegister_return_reqs,
      return_acks => UpdateRegister_return_acks,
      call_data  => UpdateRegister_call_data,
      call_tag  => UpdateRegister_call_tag,
      return_tag  => UpdateRegister_return_tag,
      call_mtag => UpdateRegister_tag_in,
      return_mtag => UpdateRegister_tag_out,
      return_data =>UpdateRegister_return_data,
      call_mreq => UpdateRegister_start_req,
      call_mack => UpdateRegister_start_ack,
      return_mreq => UpdateRegister_fin_req,
      return_mack => UpdateRegister_fin_ack,
      call_mdata => UpdateRegister_in_args,
      return_mdata => UpdateRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  UpdateRegister_instance:UpdateRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      bmask => UpdateRegister_bmask,
      rval => UpdateRegister_rval,
      wdata => UpdateRegister_wdata,
      index => UpdateRegister_index,
      wval => UpdateRegister_wval,
      start_req => UpdateRegister_start_req,
      start_ack => UpdateRegister_start_ack,
      fin_req => UpdateRegister_fin_req,
      fin_ack => UpdateRegister_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(5 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => UpdateRegister_tag_in,
      tag_out => UpdateRegister_tag_out-- 
    ); -- 
  -- module accessMemory
  accessMemory_lock <= accessMemory_in_args(109 downto 109);
  accessMemory_rwbar <= accessMemory_in_args(108 downto 108);
  accessMemory_bmask <= accessMemory_in_args(107 downto 100);
  accessMemory_addr <= accessMemory_in_args(99 downto 64);
  accessMemory_wdata <= accessMemory_in_args(63 downto 0);
  accessMemory_out_args <= accessMemory_rdata ;
  -- call arbiter for module accessMemory
  accessMemory_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 14,
      call_data_width => 110,
      return_data_width => 64,
      callee_tag_length => 4,
      caller_tag_length => 3--
    )
    port map(-- 
      call_reqs => accessMemory_call_reqs,
      call_acks => accessMemory_call_acks,
      return_reqs => accessMemory_return_reqs,
      return_acks => accessMemory_return_acks,
      call_data  => accessMemory_call_data,
      call_tag  => accessMemory_call_tag,
      return_tag  => accessMemory_return_tag,
      call_mtag => accessMemory_tag_in,
      return_mtag => accessMemory_tag_out,
      return_data =>accessMemory_return_data,
      call_mreq => accessMemory_start_req,
      call_mack => accessMemory_start_ack,
      return_mreq => accessMemory_fin_req,
      return_mack => accessMemory_fin_ack,
      call_mdata => accessMemory_in_args,
      return_mdata => accessMemory_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemory_instance:accessMemory-- 
    generic map(tag_length => 7)
    port map(-- 
      lock => accessMemory_lock,
      rwbar => accessMemory_rwbar,
      bmask => accessMemory_bmask,
      addr => accessMemory_addr,
      wdata => accessMemory_wdata,
      rdata => accessMemory_rdata,
      start_req => accessMemory_start_req,
      start_ack => accessMemory_start_ack,
      fin_req => accessMemory_fin_req,
      fin_ack => accessMemory_fin_ack,
      clk => clk,
      reset => reset,
      MEMORY_TO_NIC_RESPONSE_pipe_read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessMemory_tag_in,
      tag_out => accessMemory_tag_out-- 
    ); -- 
  -- module acquireLock
  acquireLock_q_base_address <= acquireLock_in_args(35 downto 0);
  acquireLock_out_args <= acquireLock_m_ok ;
  -- call arbiter for module acquireLock
  acquireLock_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => acquireLock_call_reqs,
      call_acks => acquireLock_call_acks,
      return_reqs => acquireLock_return_reqs,
      return_acks => acquireLock_return_acks,
      call_data  => acquireLock_call_data,
      call_tag  => acquireLock_call_tag,
      return_tag  => acquireLock_return_tag,
      call_mtag => acquireLock_tag_in,
      return_mtag => acquireLock_tag_out,
      return_data =>acquireLock_return_data,
      call_mreq => acquireLock_start_req,
      call_mack => acquireLock_start_ack,
      return_mreq => acquireLock_fin_req,
      return_mack => acquireLock_fin_ack,
      call_mdata => acquireLock_in_args,
      return_mdata => acquireLock_out_args,
      clk => clk, 
      reset => reset --
    ); --
  acquireLock_instance:acquireLock-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => acquireLock_q_base_address,
      m_ok => acquireLock_m_ok,
      start_req => acquireLock_start_req,
      start_ack => acquireLock_start_ack,
      fin_req => acquireLock_fin_req,
      fin_ack => acquireLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(11 downto 11),
      accessMemory_call_acks => accessMemory_call_acks(11 downto 11),
      accessMemory_call_data => accessMemory_call_data(1319 downto 1210),
      accessMemory_call_tag => accessMemory_call_tag(35 downto 33),
      accessMemory_return_reqs => accessMemory_return_reqs(11 downto 11),
      accessMemory_return_acks => accessMemory_return_acks(11 downto 11),
      accessMemory_return_data => accessMemory_return_data(767 downto 704),
      accessMemory_return_tag => accessMemory_return_tag(35 downto 33),
      tag_in => acquireLock_tag_in,
      tag_out => acquireLock_tag_out-- 
    ); -- 
  -- module getQueueElement
  getQueueElement_q_base_address <= getQueueElement_in_args(67 downto 32);
  getQueueElement_read_index <= getQueueElement_in_args(31 downto 0);
  getQueueElement_out_args <= getQueueElement_q_r_data ;
  -- call arbiter for module getQueueElement
  getQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 68,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueElement_call_reqs,
      call_acks => getQueueElement_call_acks,
      return_reqs => getQueueElement_return_reqs,
      return_acks => getQueueElement_return_acks,
      call_data  => getQueueElement_call_data,
      call_tag  => getQueueElement_call_tag,
      return_tag  => getQueueElement_return_tag,
      call_mtag => getQueueElement_tag_in,
      return_mtag => getQueueElement_tag_out,
      return_data =>getQueueElement_return_data,
      call_mreq => getQueueElement_start_req,
      call_mack => getQueueElement_start_ack,
      return_mreq => getQueueElement_fin_req,
      return_mack => getQueueElement_fin_ack,
      call_mdata => getQueueElement_in_args,
      return_mdata => getQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueElement_instance:getQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => getQueueElement_q_base_address,
      read_index => getQueueElement_read_index,
      q_r_data => getQueueElement_q_r_data,
      start_req => getQueueElement_start_req,
      start_ack => getQueueElement_start_ack,
      fin_req => getQueueElement_fin_req,
      fin_ack => getQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(8 downto 8),
      accessMemory_call_acks => accessMemory_call_acks(8 downto 8),
      accessMemory_call_data => accessMemory_call_data(989 downto 880),
      accessMemory_call_tag => accessMemory_call_tag(26 downto 24),
      accessMemory_return_reqs => accessMemory_return_reqs(8 downto 8),
      accessMemory_return_acks => accessMemory_return_acks(8 downto 8),
      accessMemory_return_data => accessMemory_return_data(575 downto 512),
      accessMemory_return_tag => accessMemory_return_tag(26 downto 24),
      tag_in => getQueueElement_tag_in,
      tag_out => getQueueElement_tag_out-- 
    ); -- 
  -- module getQueueLength
  getQueueLength_q_base_address <= getQueueLength_in_args(35 downto 0);
  getQueueLength_out_args <= getQueueLength_Queue_Length ;
  -- call arbiter for module getQueueLength
  getQueueLength_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueLength_call_reqs,
      call_acks => getQueueLength_call_acks,
      return_reqs => getQueueLength_return_reqs,
      return_acks => getQueueLength_return_acks,
      call_data  => getQueueLength_call_data,
      call_tag  => getQueueLength_call_tag,
      return_tag  => getQueueLength_return_tag,
      call_mtag => getQueueLength_tag_in,
      return_mtag => getQueueLength_tag_out,
      return_data =>getQueueLength_return_data,
      call_mreq => getQueueLength_start_req,
      call_mack => getQueueLength_start_ack,
      return_mreq => getQueueLength_fin_req,
      return_mack => getQueueLength_fin_ack,
      call_mdata => getQueueLength_in_args,
      return_mdata => getQueueLength_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueLength_instance:getQueueLength-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueueLength_q_base_address,
      Queue_Length => getQueueLength_Queue_Length,
      start_req => getQueueLength_start_req,
      start_ack => getQueueLength_start_ack,
      fin_req => getQueueLength_fin_req,
      fin_ack => getQueueLength_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(10 downto 10),
      accessMemory_call_acks => accessMemory_call_acks(10 downto 10),
      accessMemory_call_data => accessMemory_call_data(1209 downto 1100),
      accessMemory_call_tag => accessMemory_call_tag(32 downto 30),
      accessMemory_return_reqs => accessMemory_return_reqs(10 downto 10),
      accessMemory_return_acks => accessMemory_return_acks(10 downto 10),
      accessMemory_return_data => accessMemory_return_data(703 downto 640),
      accessMemory_return_tag => accessMemory_return_tag(32 downto 30),
      tag_in => getQueueLength_tag_in,
      tag_out => getQueueLength_tag_out-- 
    ); -- 
  -- module getQueuePointers
  getQueuePointers_q_base_address <= getQueuePointers_in_args(35 downto 0);
  getQueuePointers_out_args <= getQueuePointers_wp & getQueuePointers_rp ;
  -- call arbiter for module getQueuePointers
  getQueuePointers_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointers_call_reqs,
      call_acks => getQueuePointers_call_acks,
      return_reqs => getQueuePointers_return_reqs,
      return_acks => getQueuePointers_return_acks,
      call_data  => getQueuePointers_call_data,
      call_tag  => getQueuePointers_call_tag,
      return_tag  => getQueuePointers_return_tag,
      call_mtag => getQueuePointers_tag_in,
      return_mtag => getQueuePointers_tag_out,
      return_data =>getQueuePointers_return_data,
      call_mreq => getQueuePointers_start_req,
      call_mack => getQueuePointers_start_ack,
      return_mreq => getQueuePointers_fin_req,
      return_mack => getQueuePointers_fin_ack,
      call_mdata => getQueuePointers_in_args,
      return_mdata => getQueuePointers_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointers_instance:getQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueuePointers_q_base_address,
      wp => getQueuePointers_wp,
      rp => getQueuePointers_rp,
      start_req => getQueuePointers_start_req,
      start_ack => getQueuePointers_start_ack,
      fin_req => getQueuePointers_fin_req,
      fin_ack => getQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(12 downto 12),
      accessMemory_call_acks => accessMemory_call_acks(12 downto 12),
      accessMemory_call_data => accessMemory_call_data(1429 downto 1320),
      accessMemory_call_tag => accessMemory_call_tag(38 downto 36),
      accessMemory_return_reqs => accessMemory_return_reqs(12 downto 12),
      accessMemory_return_acks => accessMemory_return_acks(12 downto 12),
      accessMemory_return_data => accessMemory_return_data(831 downto 768),
      accessMemory_return_tag => accessMemory_return_tag(38 downto 36),
      tag_in => getQueuePointers_tag_in,
      tag_out => getQueuePointers_tag_out-- 
    ); -- 
  -- module getTotalMessages
  getTotalMessages_q_base_address <= getTotalMessages_in_args(35 downto 0);
  getTotalMessages_out_args <= getTotalMessages_total_msgs ;
  -- call arbiter for module getTotalMessages
  getTotalMessages_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTotalMessages_call_reqs,
      call_acks => getTotalMessages_call_acks,
      return_reqs => getTotalMessages_return_reqs,
      return_acks => getTotalMessages_return_acks,
      call_data  => getTotalMessages_call_data,
      call_tag  => getTotalMessages_call_tag,
      return_tag  => getTotalMessages_return_tag,
      call_mtag => getTotalMessages_tag_in,
      return_mtag => getTotalMessages_tag_out,
      return_data =>getTotalMessages_return_data,
      call_mreq => getTotalMessages_start_req,
      call_mack => getTotalMessages_start_ack,
      return_mreq => getTotalMessages_fin_req,
      return_mack => getTotalMessages_fin_ack,
      call_mdata => getTotalMessages_in_args,
      return_mdata => getTotalMessages_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTotalMessages_instance:getTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getTotalMessages_q_base_address,
      total_msgs => getTotalMessages_total_msgs,
      start_req => getTotalMessages_start_req,
      start_ack => getTotalMessages_start_ack,
      fin_req => getTotalMessages_fin_req,
      fin_ack => getTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(9 downto 9),
      accessMemory_call_acks => accessMemory_call_acks(9 downto 9),
      accessMemory_call_data => accessMemory_call_data(1099 downto 990),
      accessMemory_call_tag => accessMemory_call_tag(29 downto 27),
      accessMemory_return_reqs => accessMemory_return_reqs(9 downto 9),
      accessMemory_return_acks => accessMemory_return_acks(9 downto 9),
      accessMemory_return_data => accessMemory_return_data(639 downto 576),
      accessMemory_return_tag => accessMemory_return_tag(29 downto 27),
      tag_in => getTotalMessages_tag_in,
      tag_out => getTotalMessages_tag_out-- 
    ); -- 
  -- module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_queue_index <= getTxPacketPointerFromServer_in_args(5 downto 0);
  getTxPacketPointerFromServer_out_args <= getTxPacketPointerFromServer_pkt_pointer & getTxPacketPointerFromServer_status ;
  -- call arbiter for module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 6,
      return_data_width => 33,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTxPacketPointerFromServer_call_reqs,
      call_acks => getTxPacketPointerFromServer_call_acks,
      return_reqs => getTxPacketPointerFromServer_return_reqs,
      return_acks => getTxPacketPointerFromServer_return_acks,
      call_data  => getTxPacketPointerFromServer_call_data,
      call_tag  => getTxPacketPointerFromServer_call_tag,
      return_tag  => getTxPacketPointerFromServer_return_tag,
      call_mtag => getTxPacketPointerFromServer_tag_in,
      return_mtag => getTxPacketPointerFromServer_tag_out,
      return_data =>getTxPacketPointerFromServer_return_data,
      call_mreq => getTxPacketPointerFromServer_start_req,
      call_mack => getTxPacketPointerFromServer_start_ack,
      return_mreq => getTxPacketPointerFromServer_fin_req,
      return_mack => getTxPacketPointerFromServer_fin_ack,
      call_mdata => getTxPacketPointerFromServer_in_args,
      return_mdata => getTxPacketPointerFromServer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTxPacketPointerFromServer_instance:getTxPacketPointerFromServer-- 
    generic map(tag_length => 2)
    port map(-- 
      queue_index => getTxPacketPointerFromServer_queue_index,
      pkt_pointer => getTxPacketPointerFromServer_pkt_pointer,
      status => getTxPacketPointerFromServer_status,
      start_req => getTxPacketPointerFromServer_start_req,
      start_ack => getTxPacketPointerFromServer_start_ack,
      fin_req => getTxPacketPointerFromServer_fin_req,
      fin_ack => getTxPacketPointerFromServer_fin_ack,
      clk => clk,
      reset => reset,
      AccessRegister_call_reqs => AccessRegister_call_reqs(4 downto 4),
      AccessRegister_call_acks => AccessRegister_call_acks(4 downto 4),
      AccessRegister_call_data => AccessRegister_call_data(214 downto 172),
      AccessRegister_call_tag => AccessRegister_call_tag(9 downto 8),
      AccessRegister_return_reqs => AccessRegister_return_reqs(4 downto 4),
      AccessRegister_return_acks => AccessRegister_return_acks(4 downto 4),
      AccessRegister_return_data => AccessRegister_return_data(159 downto 128),
      AccessRegister_return_tag => AccessRegister_return_tag(9 downto 8),
      popFromQueue_call_reqs => popFromQueue_call_reqs(1 downto 1),
      popFromQueue_call_acks => popFromQueue_call_acks(1 downto 1),
      popFromQueue_call_data => popFromQueue_call_data(73 downto 37),
      popFromQueue_call_tag => popFromQueue_call_tag(1 downto 1),
      popFromQueue_return_reqs => popFromQueue_return_reqs(1 downto 1),
      popFromQueue_return_acks => popFromQueue_return_acks(1 downto 1),
      popFromQueue_return_data => popFromQueue_return_data(65 downto 33),
      popFromQueue_return_tag => popFromQueue_return_tag(1 downto 1),
      tag_in => getTxPacketPointerFromServer_tag_in,
      tag_out => getTxPacketPointerFromServer_tag_out-- 
    ); -- 
  -- module loadBuffer
  loadBuffer_rx_buffer_pointer <= loadBuffer_in_args(35 downto 0);
  loadBuffer_out_args <= loadBuffer_bad_packet_identifier ;
  -- call arbiter for module loadBuffer
  loadBuffer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadBuffer_call_reqs,
      call_acks => loadBuffer_call_acks,
      return_reqs => loadBuffer_return_reqs,
      return_acks => loadBuffer_return_acks,
      call_data  => loadBuffer_call_data,
      call_tag  => loadBuffer_call_tag,
      return_tag  => loadBuffer_return_tag,
      call_mtag => loadBuffer_tag_in,
      return_mtag => loadBuffer_tag_out,
      return_data =>loadBuffer_return_data,
      call_mreq => loadBuffer_start_req,
      call_mack => loadBuffer_start_ack,
      return_mreq => loadBuffer_fin_req,
      return_mack => loadBuffer_fin_ack,
      call_mdata => loadBuffer_in_args,
      return_mdata => loadBuffer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  loadBuffer_instance:loadBuffer-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => loadBuffer_rx_buffer_pointer,
      bad_packet_identifier => loadBuffer_bad_packet_identifier,
      start_req => loadBuffer_start_req,
      start_ack => loadBuffer_start_ack,
      fin_req => loadBuffer_fin_req,
      fin_ack => loadBuffer_fin_ack,
      clk => clk,
      reset => reset,
      writeEthernetHeaderToMem_call_reqs => writeEthernetHeaderToMem_call_reqs(0 downto 0),
      writeEthernetHeaderToMem_call_acks => writeEthernetHeaderToMem_call_acks(0 downto 0),
      writeEthernetHeaderToMem_call_data => writeEthernetHeaderToMem_call_data(35 downto 0),
      writeEthernetHeaderToMem_call_tag => writeEthernetHeaderToMem_call_tag(0 downto 0),
      writeEthernetHeaderToMem_return_reqs => writeEthernetHeaderToMem_return_reqs(0 downto 0),
      writeEthernetHeaderToMem_return_acks => writeEthernetHeaderToMem_return_acks(0 downto 0),
      writeEthernetHeaderToMem_return_data => writeEthernetHeaderToMem_return_data(35 downto 0),
      writeEthernetHeaderToMem_return_tag => writeEthernetHeaderToMem_return_tag(0 downto 0),
      writePayloadToMem_call_reqs => writePayloadToMem_call_reqs(0 downto 0),
      writePayloadToMem_call_acks => writePayloadToMem_call_acks(0 downto 0),
      writePayloadToMem_call_data => writePayloadToMem_call_data(71 downto 0),
      writePayloadToMem_call_tag => writePayloadToMem_call_tag(0 downto 0),
      writePayloadToMem_return_reqs => writePayloadToMem_return_reqs(0 downto 0),
      writePayloadToMem_return_acks => writePayloadToMem_return_acks(0 downto 0),
      writePayloadToMem_return_data => writePayloadToMem_return_data(16 downto 0),
      writePayloadToMem_return_tag => writePayloadToMem_return_tag(0 downto 0),
      writeControlInformationToMem_call_reqs => writeControlInformationToMem_call_reqs(0 downto 0),
      writeControlInformationToMem_call_acks => writeControlInformationToMem_call_acks(0 downto 0),
      writeControlInformationToMem_call_data => writeControlInformationToMem_call_data(51 downto 0),
      writeControlInformationToMem_call_tag => writeControlInformationToMem_call_tag(0 downto 0),
      writeControlInformationToMem_return_reqs => writeControlInformationToMem_return_reqs(0 downto 0),
      writeControlInformationToMem_return_acks => writeControlInformationToMem_return_acks(0 downto 0),
      writeControlInformationToMem_return_tag => writeControlInformationToMem_return_tag(0 downto 0),
      tag_in => loadBuffer_tag_in,
      tag_out => loadBuffer_tag_out-- 
    ); -- 
  -- module nicRxFromMacDaemon
  nicRxFromMacDaemon_instance:nicRxFromMacDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicRxFromMacDaemon_start_req,
      start_ack => nicRxFromMacDaemon_start_ack,
      fin_req => nicRxFromMacDaemon_fin_req,
      fin_ack => nicRxFromMacDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      mac_to_nic_data_pipe_read_req => mac_to_nic_data_pipe_read_req(0 downto 0),
      mac_to_nic_data_pipe_read_ack => mac_to_nic_data_pipe_read_ack(0 downto 0),
      mac_to_nic_data_pipe_read_data => mac_to_nic_data_pipe_read_data(72 downto 0),
      nic_rx_to_packet_pipe_write_req => nic_rx_to_packet_pipe_write_req(0 downto 0),
      nic_rx_to_packet_pipe_write_ack => nic_rx_to_packet_pipe_write_ack(0 downto 0),
      nic_rx_to_packet_pipe_write_data => nic_rx_to_packet_pipe_write_data(72 downto 0),
      nic_rx_to_header_pipe_write_req => nic_rx_to_header_pipe_write_req(0 downto 0),
      nic_rx_to_header_pipe_write_ack => nic_rx_to_header_pipe_write_ack(0 downto 0),
      nic_rx_to_header_pipe_write_data => nic_rx_to_header_pipe_write_data(72 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(2 downto 1),
      AccessRegister_call_acks => AccessRegister_call_acks(2 downto 1),
      AccessRegister_call_data => AccessRegister_call_data(128 downto 43),
      AccessRegister_call_tag => AccessRegister_call_tag(5 downto 2),
      AccessRegister_return_reqs => AccessRegister_return_reqs(2 downto 1),
      AccessRegister_return_acks => AccessRegister_return_acks(2 downto 1),
      AccessRegister_return_data => AccessRegister_return_data(95 downto 32),
      AccessRegister_return_tag => AccessRegister_return_tag(5 downto 2),
      tag_in => nicRxFromMacDaemon_tag_in,
      tag_out => nicRxFromMacDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicRxFromMacDaemon_tag_in <= (others => '0');
  nicRxFromMacDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicRxFromMacDaemon_start_req, start_ack => nicRxFromMacDaemon_start_ack,  fin_req => nicRxFromMacDaemon_fin_req,  fin_ack => nicRxFromMacDaemon_fin_ack);
  -- module popFromQueue
  popFromQueue_lock <= popFromQueue_in_args(36 downto 36);
  popFromQueue_q_base_address <= popFromQueue_in_args(35 downto 0);
  popFromQueue_out_args <= popFromQueue_q_r_data & popFromQueue_status ;
  -- call arbiter for module popFromQueue
  popFromQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 37,
      return_data_width => 33,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => popFromQueue_call_reqs,
      call_acks => popFromQueue_call_acks,
      return_reqs => popFromQueue_return_reqs,
      return_acks => popFromQueue_return_acks,
      call_data  => popFromQueue_call_data,
      call_tag  => popFromQueue_call_tag,
      return_tag  => popFromQueue_return_tag,
      call_mtag => popFromQueue_tag_in,
      return_mtag => popFromQueue_tag_out,
      return_data =>popFromQueue_return_data,
      call_mreq => popFromQueue_start_req,
      call_mack => popFromQueue_start_ack,
      return_mreq => popFromQueue_fin_req,
      return_mack => popFromQueue_fin_ack,
      call_mdata => popFromQueue_in_args,
      return_mdata => popFromQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  popFromQueue_instance:popFromQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => popFromQueue_lock,
      q_base_address => popFromQueue_q_base_address,
      q_r_data => popFromQueue_q_r_data,
      status => popFromQueue_status,
      start_req => popFromQueue_start_req,
      start_ack => popFromQueue_start_ack,
      fin_req => popFromQueue_fin_req,
      fin_ack => popFromQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireLock_call_reqs => acquireLock_call_reqs(1 downto 1),
      acquireLock_call_acks => acquireLock_call_acks(1 downto 1),
      acquireLock_call_data => acquireLock_call_data(71 downto 36),
      acquireLock_call_tag => acquireLock_call_tag(1 downto 1),
      acquireLock_return_reqs => acquireLock_return_reqs(1 downto 1),
      acquireLock_return_acks => acquireLock_return_acks(1 downto 1),
      acquireLock_return_data => acquireLock_return_data(1 downto 1),
      acquireLock_return_tag => acquireLock_return_tag(1 downto 1),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(1 downto 1),
      getQueuePointers_call_acks => getQueuePointers_call_acks(1 downto 1),
      getQueuePointers_call_data => getQueuePointers_call_data(71 downto 36),
      getQueuePointers_call_tag => getQueuePointers_call_tag(1 downto 1),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(1 downto 1),
      getQueuePointers_return_acks => getQueuePointers_return_acks(1 downto 1),
      getQueuePointers_return_data => getQueuePointers_return_data(127 downto 64),
      getQueuePointers_return_tag => getQueuePointers_return_tag(1 downto 1),
      getQueueLength_call_reqs => getQueueLength_call_reqs(1 downto 1),
      getQueueLength_call_acks => getQueueLength_call_acks(1 downto 1),
      getQueueLength_call_data => getQueueLength_call_data(71 downto 36),
      getQueueLength_call_tag => getQueueLength_call_tag(1 downto 1),
      getQueueLength_return_reqs => getQueueLength_return_reqs(1 downto 1),
      getQueueLength_return_acks => getQueueLength_return_acks(1 downto 1),
      getQueueLength_return_data => getQueueLength_return_data(63 downto 32),
      getQueueLength_return_tag => getQueueLength_return_tag(1 downto 1),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(1 downto 1),
      getTotalMessages_call_acks => getTotalMessages_call_acks(1 downto 1),
      getTotalMessages_call_data => getTotalMessages_call_data(71 downto 36),
      getTotalMessages_call_tag => getTotalMessages_call_tag(1 downto 1),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(1 downto 1),
      getTotalMessages_return_acks => getTotalMessages_return_acks(1 downto 1),
      getTotalMessages_return_data => getTotalMessages_return_data(63 downto 32),
      getTotalMessages_return_tag => getTotalMessages_return_tag(1 downto 1),
      getQueueElement_call_reqs => getQueueElement_call_reqs(0 downto 0),
      getQueueElement_call_acks => getQueueElement_call_acks(0 downto 0),
      getQueueElement_call_data => getQueueElement_call_data(67 downto 0),
      getQueueElement_call_tag => getQueueElement_call_tag(0 downto 0),
      getQueueElement_return_reqs => getQueueElement_return_reqs(0 downto 0),
      getQueueElement_return_acks => getQueueElement_return_acks(0 downto 0),
      getQueueElement_return_data => getQueueElement_return_data(31 downto 0),
      getQueueElement_return_tag => getQueueElement_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(1 downto 1),
      setQueuePointers_call_acks => setQueuePointers_call_acks(1 downto 1),
      setQueuePointers_call_data => setQueuePointers_call_data(199 downto 100),
      setQueuePointers_call_tag => setQueuePointers_call_tag(1 downto 1),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(1 downto 1),
      setQueuePointers_return_acks => setQueuePointers_return_acks(1 downto 1),
      setQueuePointers_return_tag => setQueuePointers_return_tag(1 downto 1),
      updateTotalMessages_call_reqs => updateTotalMessages_call_reqs(1 downto 1),
      updateTotalMessages_call_acks => updateTotalMessages_call_acks(1 downto 1),
      updateTotalMessages_call_data => updateTotalMessages_call_data(135 downto 68),
      updateTotalMessages_call_tag => updateTotalMessages_call_tag(1 downto 1),
      updateTotalMessages_return_reqs => updateTotalMessages_return_reqs(1 downto 1),
      updateTotalMessages_return_acks => updateTotalMessages_return_acks(1 downto 1),
      updateTotalMessages_return_tag => updateTotalMessages_return_tag(1 downto 1),
      releaseLock_call_reqs => releaseLock_call_reqs(1 downto 1),
      releaseLock_call_acks => releaseLock_call_acks(1 downto 1),
      releaseLock_call_data => releaseLock_call_data(71 downto 36),
      releaseLock_call_tag => releaseLock_call_tag(1 downto 1),
      releaseLock_return_reqs => releaseLock_return_reqs(1 downto 1),
      releaseLock_return_acks => releaseLock_return_acks(1 downto 1),
      releaseLock_return_tag => releaseLock_return_tag(1 downto 1),
      tag_in => popFromQueue_tag_in,
      tag_out => popFromQueue_tag_out-- 
    ); -- 
  -- module populateRxQueue
  populateRxQueue_rx_buffer_pointer <= populateRxQueue_in_args(35 downto 0);
  -- call arbiter for module populateRxQueue
  populateRxQueue_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => populateRxQueue_call_reqs,
      call_acks => populateRxQueue_call_acks,
      return_reqs => populateRxQueue_return_reqs,
      return_acks => populateRxQueue_return_acks,
      call_data  => populateRxQueue_call_data,
      call_tag  => populateRxQueue_call_tag,
      return_tag  => populateRxQueue_return_tag,
      call_mtag => populateRxQueue_tag_in,
      return_mtag => populateRxQueue_tag_out,
      call_mreq => populateRxQueue_start_req,
      call_mack => populateRxQueue_start_ack,
      return_mreq => populateRxQueue_fin_req,
      return_mack => populateRxQueue_fin_ack,
      call_mdata => populateRxQueue_in_args,
      clk => clk, 
      reset => reset --
    ); --
  populateRxQueue_instance:populateRxQueue-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => populateRxQueue_rx_buffer_pointer,
      start_req => populateRxQueue_start_req,
      start_ack => populateRxQueue_start_ack,
      fin_req => populateRxQueue_fin_req,
      fin_ack => populateRxQueue_fin_ack,
      clk => clk,
      reset => reset,
      LAST_WRITTEN_RX_QUEUE_INDEX => LAST_WRITTEN_RX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(11 downto 6),
      AccessRegister_call_reqs => AccessRegister_call_reqs(5 downto 5),
      AccessRegister_call_acks => AccessRegister_call_acks(5 downto 5),
      AccessRegister_call_data => AccessRegister_call_data(257 downto 215),
      AccessRegister_call_tag => AccessRegister_call_tag(11 downto 10),
      AccessRegister_return_reqs => AccessRegister_return_reqs(5 downto 5),
      AccessRegister_return_acks => AccessRegister_return_acks(5 downto 5),
      AccessRegister_return_data => AccessRegister_return_data(191 downto 160),
      AccessRegister_return_tag => AccessRegister_return_tag(11 downto 10),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(2 downto 2),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(2 downto 2),
      pushIntoQueue_call_data => pushIntoQueue_call_data(206 downto 138),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(2 downto 2),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(2 downto 2),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(2 downto 2),
      pushIntoQueue_return_data => pushIntoQueue_return_data(2 downto 2),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(2 downto 2),
      tag_in => populateRxQueue_tag_in,
      tag_out => populateRxQueue_tag_out-- 
    ); -- 
  -- module pushIntoQueue
  pushIntoQueue_lock <= pushIntoQueue_in_args(68 downto 68);
  pushIntoQueue_q_base_address <= pushIntoQueue_in_args(67 downto 32);
  pushIntoQueue_q_w_data <= pushIntoQueue_in_args(31 downto 0);
  pushIntoQueue_out_args <= pushIntoQueue_status ;
  -- call arbiter for module pushIntoQueue
  pushIntoQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 69,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => pushIntoQueue_call_reqs,
      call_acks => pushIntoQueue_call_acks,
      return_reqs => pushIntoQueue_return_reqs,
      return_acks => pushIntoQueue_return_acks,
      call_data  => pushIntoQueue_call_data,
      call_tag  => pushIntoQueue_call_tag,
      return_tag  => pushIntoQueue_return_tag,
      call_mtag => pushIntoQueue_tag_in,
      return_mtag => pushIntoQueue_tag_out,
      return_data =>pushIntoQueue_return_data,
      call_mreq => pushIntoQueue_start_req,
      call_mack => pushIntoQueue_start_ack,
      return_mreq => pushIntoQueue_fin_req,
      return_mack => pushIntoQueue_fin_ack,
      call_mdata => pushIntoQueue_in_args,
      return_mdata => pushIntoQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  pushIntoQueue_instance:pushIntoQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => pushIntoQueue_lock,
      q_base_address => pushIntoQueue_q_base_address,
      q_w_data => pushIntoQueue_q_w_data,
      status => pushIntoQueue_status,
      start_req => pushIntoQueue_start_req,
      start_ack => pushIntoQueue_start_ack,
      fin_req => pushIntoQueue_fin_req,
      fin_ack => pushIntoQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireLock_call_reqs => acquireLock_call_reqs(0 downto 0),
      acquireLock_call_acks => acquireLock_call_acks(0 downto 0),
      acquireLock_call_data => acquireLock_call_data(35 downto 0),
      acquireLock_call_tag => acquireLock_call_tag(0 downto 0),
      acquireLock_return_reqs => acquireLock_return_reqs(0 downto 0),
      acquireLock_return_acks => acquireLock_return_acks(0 downto 0),
      acquireLock_return_data => acquireLock_return_data(0 downto 0),
      acquireLock_return_tag => acquireLock_return_tag(0 downto 0),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(0 downto 0),
      getQueuePointers_call_acks => getQueuePointers_call_acks(0 downto 0),
      getQueuePointers_call_data => getQueuePointers_call_data(35 downto 0),
      getQueuePointers_call_tag => getQueuePointers_call_tag(0 downto 0),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(0 downto 0),
      getQueuePointers_return_acks => getQueuePointers_return_acks(0 downto 0),
      getQueuePointers_return_data => getQueuePointers_return_data(63 downto 0),
      getQueuePointers_return_tag => getQueuePointers_return_tag(0 downto 0),
      getQueueLength_call_reqs => getQueueLength_call_reqs(0 downto 0),
      getQueueLength_call_acks => getQueueLength_call_acks(0 downto 0),
      getQueueLength_call_data => getQueueLength_call_data(35 downto 0),
      getQueueLength_call_tag => getQueueLength_call_tag(0 downto 0),
      getQueueLength_return_reqs => getQueueLength_return_reqs(0 downto 0),
      getQueueLength_return_acks => getQueueLength_return_acks(0 downto 0),
      getQueueLength_return_data => getQueueLength_return_data(31 downto 0),
      getQueueLength_return_tag => getQueueLength_return_tag(0 downto 0),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(0 downto 0),
      getTotalMessages_call_acks => getTotalMessages_call_acks(0 downto 0),
      getTotalMessages_call_data => getTotalMessages_call_data(35 downto 0),
      getTotalMessages_call_tag => getTotalMessages_call_tag(0 downto 0),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(0 downto 0),
      getTotalMessages_return_acks => getTotalMessages_return_acks(0 downto 0),
      getTotalMessages_return_data => getTotalMessages_return_data(31 downto 0),
      getTotalMessages_return_tag => getTotalMessages_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(0 downto 0),
      setQueuePointers_call_acks => setQueuePointers_call_acks(0 downto 0),
      setQueuePointers_call_data => setQueuePointers_call_data(99 downto 0),
      setQueuePointers_call_tag => setQueuePointers_call_tag(0 downto 0),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(0 downto 0),
      setQueuePointers_return_acks => setQueuePointers_return_acks(0 downto 0),
      setQueuePointers_return_tag => setQueuePointers_return_tag(0 downto 0),
      updateTotalMessages_call_reqs => updateTotalMessages_call_reqs(0 downto 0),
      updateTotalMessages_call_acks => updateTotalMessages_call_acks(0 downto 0),
      updateTotalMessages_call_data => updateTotalMessages_call_data(67 downto 0),
      updateTotalMessages_call_tag => updateTotalMessages_call_tag(0 downto 0),
      updateTotalMessages_return_reqs => updateTotalMessages_return_reqs(0 downto 0),
      updateTotalMessages_return_acks => updateTotalMessages_return_acks(0 downto 0),
      updateTotalMessages_return_tag => updateTotalMessages_return_tag(0 downto 0),
      releaseLock_call_reqs => releaseLock_call_reqs(0 downto 0),
      releaseLock_call_acks => releaseLock_call_acks(0 downto 0),
      releaseLock_call_data => releaseLock_call_data(35 downto 0),
      releaseLock_call_tag => releaseLock_call_tag(0 downto 0),
      releaseLock_return_reqs => releaseLock_return_reqs(0 downto 0),
      releaseLock_return_acks => releaseLock_return_acks(0 downto 0),
      releaseLock_return_tag => releaseLock_return_tag(0 downto 0),
      setQueueElement_call_reqs => setQueueElement_call_reqs(0 downto 0),
      setQueueElement_call_acks => setQueueElement_call_acks(0 downto 0),
      setQueueElement_call_data => setQueueElement_call_data(99 downto 0),
      setQueueElement_call_tag => setQueueElement_call_tag(0 downto 0),
      setQueueElement_return_reqs => setQueueElement_return_reqs(0 downto 0),
      setQueueElement_return_acks => setQueueElement_return_acks(0 downto 0),
      setQueueElement_return_tag => setQueueElement_return_tag(0 downto 0),
      tag_in => pushIntoQueue_tag_in,
      tag_out => pushIntoQueue_tag_out-- 
    ); -- 
  -- module releaseLock
  releaseLock_q_base_address <= releaseLock_in_args(35 downto 0);
  -- call arbiter for module releaseLock
  releaseLock_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 36,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => releaseLock_call_reqs,
      call_acks => releaseLock_call_acks,
      return_reqs => releaseLock_return_reqs,
      return_acks => releaseLock_return_acks,
      call_data  => releaseLock_call_data,
      call_tag  => releaseLock_call_tag,
      return_tag  => releaseLock_return_tag,
      call_mtag => releaseLock_tag_in,
      return_mtag => releaseLock_tag_out,
      call_mreq => releaseLock_start_req,
      call_mack => releaseLock_start_ack,
      return_mreq => releaseLock_fin_req,
      return_mack => releaseLock_fin_ack,
      call_mdata => releaseLock_in_args,
      clk => clk, 
      reset => reset --
    ); --
  releaseLock_instance:releaseLock-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => releaseLock_q_base_address,
      start_req => releaseLock_start_req,
      start_ack => releaseLock_start_ack,
      fin_req => releaseLock_fin_req,
      fin_ack => releaseLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(7 downto 7),
      accessMemory_call_acks => accessMemory_call_acks(7 downto 7),
      accessMemory_call_data => accessMemory_call_data(879 downto 770),
      accessMemory_call_tag => accessMemory_call_tag(23 downto 21),
      accessMemory_return_reqs => accessMemory_return_reqs(7 downto 7),
      accessMemory_return_acks => accessMemory_return_acks(7 downto 7),
      accessMemory_return_data => accessMemory_return_data(511 downto 448),
      accessMemory_return_tag => accessMemory_return_tag(23 downto 21),
      tag_in => releaseLock_tag_in,
      tag_out => releaseLock_tag_out-- 
    ); -- 
  -- module setQueueElement
  setQueueElement_q_base_address <= setQueueElement_in_args(99 downto 64);
  setQueueElement_write_index <= setQueueElement_in_args(63 downto 32);
  setQueueElement_q_w_data <= setQueueElement_in_args(31 downto 0);
  -- call arbiter for module setQueueElement
  setQueueElement_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 100,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueueElement_call_reqs,
      call_acks => setQueueElement_call_acks,
      return_reqs => setQueueElement_return_reqs,
      return_acks => setQueueElement_return_acks,
      call_data  => setQueueElement_call_data,
      call_tag  => setQueueElement_call_tag,
      return_tag  => setQueueElement_return_tag,
      call_mtag => setQueueElement_tag_in,
      return_mtag => setQueueElement_tag_out,
      call_mreq => setQueueElement_start_req,
      call_mack => setQueueElement_start_ack,
      return_mreq => setQueueElement_fin_req,
      return_mack => setQueueElement_fin_ack,
      call_mdata => setQueueElement_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueueElement_instance:setQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => setQueueElement_q_base_address,
      write_index => setQueueElement_write_index,
      q_w_data => setQueueElement_q_w_data,
      start_req => setQueueElement_start_req,
      start_ack => setQueueElement_start_ack,
      fin_req => setQueueElement_fin_req,
      fin_ack => setQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(2 downto 2),
      accessMemory_call_acks => accessMemory_call_acks(2 downto 2),
      accessMemory_call_data => accessMemory_call_data(329 downto 220),
      accessMemory_call_tag => accessMemory_call_tag(8 downto 6),
      accessMemory_return_reqs => accessMemory_return_reqs(2 downto 2),
      accessMemory_return_acks => accessMemory_return_acks(2 downto 2),
      accessMemory_return_data => accessMemory_return_data(191 downto 128),
      accessMemory_return_tag => accessMemory_return_tag(8 downto 6),
      tag_in => setQueueElement_tag_in,
      tag_out => setQueueElement_tag_out-- 
    ); -- 
  -- module setQueuePointers
  setQueuePointers_q_base_address <= setQueuePointers_in_args(99 downto 64);
  setQueuePointers_wp <= setQueuePointers_in_args(63 downto 32);
  setQueuePointers_rp <= setQueuePointers_in_args(31 downto 0);
  -- call arbiter for module setQueuePointers
  setQueuePointers_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 100,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueuePointers_call_reqs,
      call_acks => setQueuePointers_call_acks,
      return_reqs => setQueuePointers_return_reqs,
      return_acks => setQueuePointers_return_acks,
      call_data  => setQueuePointers_call_data,
      call_tag  => setQueuePointers_call_tag,
      return_tag  => setQueuePointers_return_tag,
      call_mtag => setQueuePointers_tag_in,
      return_mtag => setQueuePointers_tag_out,
      call_mreq => setQueuePointers_start_req,
      call_mack => setQueuePointers_start_ack,
      return_mreq => setQueuePointers_fin_req,
      return_mack => setQueuePointers_fin_ack,
      call_mdata => setQueuePointers_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueuePointers_instance:setQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => setQueuePointers_q_base_address,
      wp => setQueuePointers_wp,
      rp => setQueuePointers_rp,
      start_req => setQueuePointers_start_req,
      start_ack => setQueuePointers_start_ack,
      fin_req => setQueuePointers_fin_req,
      fin_ack => setQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(5 downto 5),
      accessMemory_call_acks => accessMemory_call_acks(5 downto 5),
      accessMemory_call_data => accessMemory_call_data(659 downto 550),
      accessMemory_call_tag => accessMemory_call_tag(17 downto 15),
      accessMemory_return_reqs => accessMemory_return_reqs(5 downto 5),
      accessMemory_return_acks => accessMemory_return_acks(5 downto 5),
      accessMemory_return_data => accessMemory_return_data(383 downto 320),
      accessMemory_return_tag => accessMemory_return_tag(17 downto 15),
      tag_in => setQueuePointers_tag_in,
      tag_out => setQueuePointers_tag_out-- 
    ); -- 
  -- module transmitEngineDaemon
  transmitEngineDaemon_instance:transmitEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => transmitEngineDaemon_start_req,
      start_ack => transmitEngineDaemon_start_ack,
      fin_req => transmitEngineDaemon_fin_req,
      fin_ack => transmitEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      FREE_Q => FREE_Q,
      LAST_READ_TX_QUEUE_INDEX => LAST_READ_TX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(0 downto 0),
      AccessRegister_call_acks => AccessRegister_call_acks(0 downto 0),
      AccessRegister_call_data => AccessRegister_call_data(42 downto 0),
      AccessRegister_call_tag => AccessRegister_call_tag(1 downto 0),
      AccessRegister_return_reqs => AccessRegister_return_reqs(0 downto 0),
      AccessRegister_return_acks => AccessRegister_return_acks(0 downto 0),
      AccessRegister_return_data => AccessRegister_return_data(31 downto 0),
      AccessRegister_return_tag => AccessRegister_return_tag(1 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(0 downto 0),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(0 downto 0),
      pushIntoQueue_call_data => pushIntoQueue_call_data(68 downto 0),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(0 downto 0),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(0 downto 0),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(0 downto 0),
      pushIntoQueue_return_data => pushIntoQueue_return_data(0 downto 0),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(0 downto 0),
      getTxPacketPointerFromServer_call_reqs => getTxPacketPointerFromServer_call_reqs(0 downto 0),
      getTxPacketPointerFromServer_call_acks => getTxPacketPointerFromServer_call_acks(0 downto 0),
      getTxPacketPointerFromServer_call_data => getTxPacketPointerFromServer_call_data(5 downto 0),
      getTxPacketPointerFromServer_call_tag => getTxPacketPointerFromServer_call_tag(0 downto 0),
      getTxPacketPointerFromServer_return_reqs => getTxPacketPointerFromServer_return_reqs(0 downto 0),
      getTxPacketPointerFromServer_return_acks => getTxPacketPointerFromServer_return_acks(0 downto 0),
      getTxPacketPointerFromServer_return_data => getTxPacketPointerFromServer_return_data(32 downto 0),
      getTxPacketPointerFromServer_return_tag => getTxPacketPointerFromServer_return_tag(0 downto 0),
      transmitPacket_call_reqs => transmitPacket_call_reqs(0 downto 0),
      transmitPacket_call_acks => transmitPacket_call_acks(0 downto 0),
      transmitPacket_call_data => transmitPacket_call_data(31 downto 0),
      transmitPacket_call_tag => transmitPacket_call_tag(0 downto 0),
      transmitPacket_return_reqs => transmitPacket_return_reqs(0 downto 0),
      transmitPacket_return_acks => transmitPacket_return_acks(0 downto 0),
      transmitPacket_return_data => transmitPacket_return_data(0 downto 0),
      transmitPacket_return_tag => transmitPacket_return_tag(0 downto 0),
      tag_in => transmitEngineDaemon_tag_in,
      tag_out => transmitEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  transmitEngineDaemon_tag_in <= (others => '0');
  transmitEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => transmitEngineDaemon_start_req, start_ack => transmitEngineDaemon_start_ack,  fin_req => transmitEngineDaemon_fin_req,  fin_ack => transmitEngineDaemon_fin_ack);
  -- module transmitPacket
  transmitPacket_packet_pointer <= transmitPacket_in_args(31 downto 0);
  transmitPacket_out_args <= transmitPacket_status ;
  -- call arbiter for module transmitPacket
  transmitPacket_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => transmitPacket_call_reqs,
      call_acks => transmitPacket_call_acks,
      return_reqs => transmitPacket_return_reqs,
      return_acks => transmitPacket_return_acks,
      call_data  => transmitPacket_call_data,
      call_tag  => transmitPacket_call_tag,
      return_tag  => transmitPacket_return_tag,
      call_mtag => transmitPacket_tag_in,
      return_mtag => transmitPacket_tag_out,
      return_data =>transmitPacket_return_data,
      call_mreq => transmitPacket_start_req,
      call_mack => transmitPacket_start_ack,
      return_mreq => transmitPacket_fin_req,
      return_mack => transmitPacket_fin_ack,
      call_mdata => transmitPacket_in_args,
      return_mdata => transmitPacket_out_args,
      clk => clk, 
      reset => reset --
    ); --
  transmitPacket_instance:transmitPacket-- 
    generic map(tag_length => 2)
    port map(-- 
      packet_pointer => transmitPacket_packet_pointer,
      status => transmitPacket_status,
      start_req => transmitPacket_start_req,
      start_ack => transmitPacket_start_ack,
      fin_req => transmitPacket_fin_req,
      fin_ack => transmitPacket_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_write_req => nic_to_mac_transmit_pipe_pipe_write_req(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_ack => nic_to_mac_transmit_pipe_pipe_write_ack(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_data => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(1 downto 0),
      accessMemory_call_acks => accessMemory_call_acks(1 downto 0),
      accessMemory_call_data => accessMemory_call_data(219 downto 0),
      accessMemory_call_tag => accessMemory_call_tag(5 downto 0),
      accessMemory_return_reqs => accessMemory_return_reqs(1 downto 0),
      accessMemory_return_acks => accessMemory_return_acks(1 downto 0),
      accessMemory_return_data => accessMemory_return_data(127 downto 0),
      accessMemory_return_tag => accessMemory_return_tag(5 downto 0),
      tag_in => transmitPacket_tag_in,
      tag_out => transmitPacket_tag_out-- 
    ); -- 
  -- module updateTotalMessages
  updateTotalMessages_q_base_address <= updateTotalMessages_in_args(67 downto 32);
  updateTotalMessages_updated_total_msgs <= updateTotalMessages_in_args(31 downto 0);
  -- call arbiter for module updateTotalMessages
  updateTotalMessages_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 68,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => updateTotalMessages_call_reqs,
      call_acks => updateTotalMessages_call_acks,
      return_reqs => updateTotalMessages_return_reqs,
      return_acks => updateTotalMessages_return_acks,
      call_data  => updateTotalMessages_call_data,
      call_tag  => updateTotalMessages_call_tag,
      return_tag  => updateTotalMessages_return_tag,
      call_mtag => updateTotalMessages_tag_in,
      return_mtag => updateTotalMessages_tag_out,
      call_mreq => updateTotalMessages_start_req,
      call_mack => updateTotalMessages_start_ack,
      return_mreq => updateTotalMessages_fin_req,
      return_mack => updateTotalMessages_fin_ack,
      call_mdata => updateTotalMessages_in_args,
      clk => clk, 
      reset => reset --
    ); --
  updateTotalMessages_instance:updateTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => updateTotalMessages_q_base_address,
      updated_total_msgs => updateTotalMessages_updated_total_msgs,
      start_req => updateTotalMessages_start_req,
      start_ack => updateTotalMessages_start_ack,
      fin_req => updateTotalMessages_fin_req,
      fin_ack => updateTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(6 downto 6),
      accessMemory_call_acks => accessMemory_call_acks(6 downto 6),
      accessMemory_call_data => accessMemory_call_data(769 downto 660),
      accessMemory_call_tag => accessMemory_call_tag(20 downto 18),
      accessMemory_return_reqs => accessMemory_return_reqs(6 downto 6),
      accessMemory_return_acks => accessMemory_return_acks(6 downto 6),
      accessMemory_return_data => accessMemory_return_data(447 downto 384),
      accessMemory_return_tag => accessMemory_return_tag(20 downto 18),
      tag_in => updateTotalMessages_tag_in,
      tag_out => updateTotalMessages_tag_out-- 
    ); -- 
  -- module writeControlInformationToMem
  writeControlInformationToMem_base_buffer_pointer <= writeControlInformationToMem_in_args(51 downto 16);
  writeControlInformationToMem_packet_size <= writeControlInformationToMem_in_args(15 downto 8);
  writeControlInformationToMem_last_keep <= writeControlInformationToMem_in_args(7 downto 0);
  -- call arbiter for module writeControlInformationToMem
  writeControlInformationToMem_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 52,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeControlInformationToMem_call_reqs,
      call_acks => writeControlInformationToMem_call_acks,
      return_reqs => writeControlInformationToMem_return_reqs,
      return_acks => writeControlInformationToMem_return_acks,
      call_data  => writeControlInformationToMem_call_data,
      call_tag  => writeControlInformationToMem_call_tag,
      return_tag  => writeControlInformationToMem_return_tag,
      call_mtag => writeControlInformationToMem_tag_in,
      return_mtag => writeControlInformationToMem_tag_out,
      call_mreq => writeControlInformationToMem_start_req,
      call_mack => writeControlInformationToMem_start_ack,
      return_mreq => writeControlInformationToMem_fin_req,
      return_mack => writeControlInformationToMem_fin_ack,
      call_mdata => writeControlInformationToMem_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeControlInformationToMem_instance:writeControlInformationToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buffer_pointer => writeControlInformationToMem_base_buffer_pointer,
      packet_size => writeControlInformationToMem_packet_size,
      last_keep => writeControlInformationToMem_last_keep,
      start_req => writeControlInformationToMem_start_req,
      start_ack => writeControlInformationToMem_start_ack,
      fin_req => writeControlInformationToMem_fin_req,
      fin_ack => writeControlInformationToMem_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(13 downto 13),
      accessMemory_call_acks => accessMemory_call_acks(13 downto 13),
      accessMemory_call_data => accessMemory_call_data(1539 downto 1430),
      accessMemory_call_tag => accessMemory_call_tag(41 downto 39),
      accessMemory_return_reqs => accessMemory_return_reqs(13 downto 13),
      accessMemory_return_acks => accessMemory_return_acks(13 downto 13),
      accessMemory_return_data => accessMemory_return_data(895 downto 832),
      accessMemory_return_tag => accessMemory_return_tag(41 downto 39),
      tag_in => writeControlInformationToMem_tag_in,
      tag_out => writeControlInformationToMem_tag_out-- 
    ); -- 
  -- module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_buf_pointer <= writeEthernetHeaderToMem_in_args(35 downto 0);
  writeEthernetHeaderToMem_out_args <= writeEthernetHeaderToMem_buf_position ;
  -- call arbiter for module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeEthernetHeaderToMem_call_reqs,
      call_acks => writeEthernetHeaderToMem_call_acks,
      return_reqs => writeEthernetHeaderToMem_return_reqs,
      return_acks => writeEthernetHeaderToMem_return_acks,
      call_data  => writeEthernetHeaderToMem_call_data,
      call_tag  => writeEthernetHeaderToMem_call_tag,
      return_tag  => writeEthernetHeaderToMem_return_tag,
      call_mtag => writeEthernetHeaderToMem_tag_in,
      return_mtag => writeEthernetHeaderToMem_tag_out,
      return_data =>writeEthernetHeaderToMem_return_data,
      call_mreq => writeEthernetHeaderToMem_start_req,
      call_mack => writeEthernetHeaderToMem_start_ack,
      return_mreq => writeEthernetHeaderToMem_fin_req,
      return_mack => writeEthernetHeaderToMem_fin_ack,
      call_mdata => writeEthernetHeaderToMem_in_args,
      return_mdata => writeEthernetHeaderToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeEthernetHeaderToMem_instance:writeEthernetHeaderToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      buf_pointer => writeEthernetHeaderToMem_buf_pointer,
      buf_position => writeEthernetHeaderToMem_buf_position,
      start_req => writeEthernetHeaderToMem_start_req,
      start_ack => writeEthernetHeaderToMem_start_ack,
      fin_req => writeEthernetHeaderToMem_fin_req,
      fin_ack => writeEthernetHeaderToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_header_pipe_read_req => nic_rx_to_header_pipe_read_req(0 downto 0),
      nic_rx_to_header_pipe_read_ack => nic_rx_to_header_pipe_read_ack(0 downto 0),
      nic_rx_to_header_pipe_read_data => nic_rx_to_header_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(4 downto 4),
      accessMemory_call_acks => accessMemory_call_acks(4 downto 4),
      accessMemory_call_data => accessMemory_call_data(549 downto 440),
      accessMemory_call_tag => accessMemory_call_tag(14 downto 12),
      accessMemory_return_reqs => accessMemory_return_reqs(4 downto 4),
      accessMemory_return_acks => accessMemory_return_acks(4 downto 4),
      accessMemory_return_data => accessMemory_return_data(319 downto 256),
      accessMemory_return_tag => accessMemory_return_tag(14 downto 12),
      tag_in => writeEthernetHeaderToMem_tag_in,
      tag_out => writeEthernetHeaderToMem_tag_out-- 
    ); -- 
  -- module writePayloadToMem
  writePayloadToMem_base_buf_pointer <= writePayloadToMem_in_args(71 downto 36);
  writePayloadToMem_buf_pointer <= writePayloadToMem_in_args(35 downto 0);
  writePayloadToMem_out_args <= writePayloadToMem_packet_size_32 & writePayloadToMem_bad_packet_identifier & writePayloadToMem_last_keep ;
  -- call arbiter for module writePayloadToMem
  writePayloadToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 17,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writePayloadToMem_call_reqs,
      call_acks => writePayloadToMem_call_acks,
      return_reqs => writePayloadToMem_return_reqs,
      return_acks => writePayloadToMem_return_acks,
      call_data  => writePayloadToMem_call_data,
      call_tag  => writePayloadToMem_call_tag,
      return_tag  => writePayloadToMem_return_tag,
      call_mtag => writePayloadToMem_tag_in,
      return_mtag => writePayloadToMem_tag_out,
      return_data =>writePayloadToMem_return_data,
      call_mreq => writePayloadToMem_start_req,
      call_mack => writePayloadToMem_start_ack,
      return_mreq => writePayloadToMem_fin_req,
      return_mack => writePayloadToMem_fin_ack,
      call_mdata => writePayloadToMem_in_args,
      return_mdata => writePayloadToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writePayloadToMem_instance:writePayloadToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buf_pointer => writePayloadToMem_base_buf_pointer,
      buf_pointer => writePayloadToMem_buf_pointer,
      packet_size_32 => writePayloadToMem_packet_size_32,
      bad_packet_identifier => writePayloadToMem_bad_packet_identifier,
      last_keep => writePayloadToMem_last_keep,
      start_req => writePayloadToMem_start_req,
      start_ack => writePayloadToMem_start_ack,
      fin_req => writePayloadToMem_fin_req,
      fin_ack => writePayloadToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_packet_pipe_read_req => nic_rx_to_packet_pipe_read_req(0 downto 0),
      nic_rx_to_packet_pipe_read_ack => nic_rx_to_packet_pipe_read_ack(0 downto 0),
      nic_rx_to_packet_pipe_read_data => nic_rx_to_packet_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(3 downto 3),
      accessMemory_call_acks => accessMemory_call_acks(3 downto 3),
      accessMemory_call_data => accessMemory_call_data(439 downto 330),
      accessMemory_call_tag => accessMemory_call_tag(11 downto 9),
      accessMemory_return_reqs => accessMemory_return_reqs(3 downto 3),
      accessMemory_return_acks => accessMemory_return_acks(3 downto 3),
      accessMemory_return_data => accessMemory_return_data(255 downto 192),
      accessMemory_return_tag => accessMemory_return_tag(11 downto 9),
      tag_in => writePayloadToMem_tag_in,
      tag_out => writePayloadToMem_tag_out-- 
    ); -- 
  AFB_NIC_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 74,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_REQUEST_pipe_read_req,
      read_ack => AFB_NIC_REQUEST_pipe_read_ack,
      read_data => AFB_NIC_REQUEST_pipe_read_data,
      write_req => AFB_NIC_REQUEST_pipe_write_req,
      write_ack => AFB_NIC_REQUEST_pipe_write_ack,
      write_data => AFB_NIC_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  AFB_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_RESPONSE_pipe_read_req,
      read_ack => AFB_NIC_RESPONSE_pipe_read_ack,
      read_data => AFB_NIC_RESPONSE_pipe_read_data,
      write_req => AFB_NIC_RESPONSE_pipe_write_req,
      write_ack => AFB_NIC_RESPONSE_pipe_write_ack,
      write_data => AFB_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  CONTROL_REGISTER_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe CONTROL_REGISTER",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => CONTROL_REGISTER,
      write_req => CONTROL_REGISTER_pipe_write_req,
      write_ack => CONTROL_REGISTER_pipe_write_ack,
      write_data => CONTROL_REGISTER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  FREE_Q_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe FREE_Q",
      volatile_flag => false,
      num_writes => 1,
      data_width => 36 --
    ) 
    port map( -- 
      read_data => FREE_Q,
      write_req => FREE_Q_pipe_write_req,
      write_ack => FREE_Q_pipe_write_ack,
      write_data => FREE_Q_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_READ_TX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_READ_TX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_READ_TX_QUEUE_INDEX,
      write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_WRITTEN_RX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_WRITTEN_RX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_WRITTEN_RX_QUEUE_INDEX,
      write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEMORY_TO_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEMORY_TO_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req,
      read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack,
      read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data,
      write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req,
      write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack,
      write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_REQUEST_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_REQUEST_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 43,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_RESPONSE_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_TO_MEMORY_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_TO_MEMORY_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req,
      read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack,
      read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data,
      write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req,
      write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack,
      write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NUMBER_OF_SERVERS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NUMBER_OF_SERVERS",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => NUMBER_OF_SERVERS,
      write_req => NUMBER_OF_SERVERS_pipe_write_req,
      write_ack => NUMBER_OF_SERVERS_pipe_write_ack,
      write_data => NUMBER_OF_SERVERS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => mac_to_nic_data_pipe_read_req,
      read_ack => mac_to_nic_data_pipe_read_ack,
      read_data => mac_to_nic_data_pipe_read_data,
      write_req => mac_to_nic_data_pipe_write_req,
      write_ack => mac_to_nic_data_pipe_write_ack,
      write_data => mac_to_nic_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_header_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_header",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_header_pipe_read_req,
      read_ack => nic_rx_to_header_pipe_read_ack,
      read_data => nic_rx_to_header_pipe_read_data,
      write_req => nic_rx_to_header_pipe_write_req,
      write_ack => nic_rx_to_header_pipe_write_ack,
      write_data => nic_rx_to_header_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_packet_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_packet",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_packet_pipe_read_req,
      read_ack => nic_rx_to_packet_pipe_read_ack,
      read_data => nic_rx_to_packet_pipe_read_data,
      write_req => nic_rx_to_packet_pipe_write_req,
      write_ack => nic_rx_to_packet_pipe_write_ack,
      write_data => nic_rx_to_packet_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_to_mac_transmit_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_to_mac_transmit_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => nic_to_mac_transmit_pipe_pipe_read_req,
      read_ack => nic_to_mac_transmit_pipe_pipe_read_ack,
      read_data => nic_to_mac_transmit_pipe_pipe_read_data,
      write_req => nic_to_mac_transmit_pipe_pipe_write_req,
      write_ack => nic_to_mac_transmit_pipe_pipe_write_ack,
      write_data => nic_to_mac_transmit_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 6,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 6,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
