

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AFl2kw3wjuupeEJWAVRMjvI4n2F9ZwKYCyTdtTbrj99jYEYTJx3fm7Ch7UNHIYnYCZk+hug4a3M6
XIrSFOf3lw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kJIX1i40eaci6RDbcVVzg1fYaa68r2QTZ19EbYvWyiO0MSVCOi3GfcyJJxOR52/mcv4FD0GrKyok
p1d2616K9ikEjuEHDsOkFkQxSSfEgbSNAEkwJoywFb1NEza/LgnXq4wCMserYGd0Ho12V4osIEdI
exWoz7u39lGc9ZiaBS4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2kMqoMFPLn7FsBBTsV6uCri7uN+peyfxKN5B0t+cAsrbL+lDiZoUrv6niJBSapyempvdNVVmTzxI
0OOKA0SUZL7oQT5S7r5QAMg9q0wHtWdtsxsKxFyZXOcUUs3IkLwLNJ9fExPXmVlCDUNWWyZ/Qtik
1q9ZynUcX4DCv1pUeRs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uW1nShxn5xYxSfsiNvMbC6cL7GFjn45B3GrJxFfTPdqHxW6l/7kPGVqMN4yc97bwWb5swAmg1/ia
P9L6G5Lmjygww+NIedzfhB4znXCEs1F+LwtP/Eo4UZuH4rQ55XUhLKrRNEqAJ5lTqYxfdIa1JIeg
6YgrU98QHKeOeZUeearBuTROZ6q9d2QFGZhc5MxjU8pwV5JQ++j3EkUIuMZJi3DVdwnYj2d1DzSG
tEt9nWmDzn5rqjvrP0c2GlNBg1tCMJxGfC7y54n+J8H6ETagMe97uL4QvKLTEhjArVfHkKedz6Hw
BLtL2VPOf8fCVrM+AsqxA6SscLteiE3Y/tcuqg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IV462y1jHGYFO6K2VU9zTKlfXJZ4kSNvewSr8uczSbz2qRhu1urkppbYmZyNPMNjUUiJfr+4xl1K
sPX+MN8CN040mI1y/WRE8sMEH4yPflkbYjeDH/AX8AZf0f51eUS3cIc3p5KYvECdG8h6xmZ6jH0F
7BqDcSAL8OaSnIetqzLPr2v1rtYXH+RRlVWmvCK2nFZ02kt8pCYkp8L5RKceyNIKFWCdOT5JdjZY
4tvHtPn6P1gVHsYV30mBGWhvJczj5zrLjwFlzuRt1FBD773q8FliSEnvM5VLjXeYVAshW6krIgcC
JRjJFfG2fLeH0eKFVJ7kqIzwNNYB0nt3Mho0og==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gxKMu2AB/FASbqvyKO7D61/XUsdMsjazR7APgUWhLu8z6ePEw4il1OmWHsQOCjylECfctRxhrNKA
ZkqobGwUpbLybNlM8OLmxSq7gFftkFYAAbUlTfr+gHIvTw0OHQ1EytNPCAXJ3C16VMRZRtIOMhuu
qWzd7JSTNzsFNMOGqUkbAJ25aM5fSFIBT9RqdtK6aDtxz+XRgnizFyeXsqGdP7bY03KX5HgTMa9w
sW64LQcPjQEuBBRxSfYreUKE1jQbO9XuIjtoOmZGDsEtv2KkhTAdFbwHWRiiIzAO+Bx945pksp3X
TfC9rKLaXHs75mi0HkNR/3vshocjTDFwp+bJaA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 122928)
`protect data_block
j9BFrh6O5oslkqRv0KMueh1qETdYle+IJ/lFALBIb5xqtxbBC83qETaMSNj9O16WumBA3TVEjBU+
isBmPrh6OyzWj/ZPk3feZNFKusRudaeRmNuJbolbPqsgTNtoll7NTONHC4MvkP8BFwu+rsHjVKhv
BMNKsot+pMrxXf5miv0m+3WZY+eHMx+1TT0C8Gm2xLB29ByNEopTWyUNNuvOzhdbuWtfxlMOLYOG
+W7XvF5C1YYs+8R4gWxnj+/vadGSIQ4H44bfezT5EZCPIQCEiJBIF+s6LSbbR2UAFyB8pPIS0FRy
8kXhYFBB+WdASEFe371iOUwJdXkNZ2hn3mznBLKJERkll+V9GNpXIr87T7kmg24CZRUb7QAB8tkc
csHoUfQk6cQYq4ge+SHDxJa6KncM8zL/GeLCyy8Ttfa+S32l2yns/dQ0miBBUROPKN0gAflQogVO
/H3chJFUHX7iXh+H/72WnhO2eh/rVOKnMEhhxspjpHJ5Z7/LbbSa2RmOoOeLln92koiF4mDtgDwA
noexEzRn75F8BSnaFRab9DTaBV6d6fuo96K8Fm0Lh50lFwTN8pQslCw6vQlbetMFRDorJst0ktRw
+59SL+r3UxRRn19M7QjBgqHMs1dqqzJJNZrViIIwlvj/64GCrS7SPuYKLkoiP3mtW1aa5AjurdJ5
t4QyPVrFEfW/UEoYlfV3fU0eo2m7/47CquHCxqUYaXS5ngoMnK427kGZ2GoPMeyOYczNRiaNQvO0
9g1g9y5bh020J0wMdOGYrc5pmhoBK1cd8xEwXy7CbgAfL/3HYsfZzKJiEuIyOz5aSwNQ+58uyYeK
Iei/dzgJzr1zpwfu5vBjyO5yl/g1c36dTW1YhP0pf+hx+iO9bQNsN6TOs5srsdphFTUYsaYxyoQc
5agt+KgM48DZJZHtWIkFd89iubc9dHET+VUx8YqCxkJR+uo+ZKgLOUXh+0Vk1NovnSLttbZUV5gS
oSstcz4KqAsaB7J6910oxRRxsUJyvgHYSOapi4mim3/WOn9Sa5354oKJgFf+Fee9zMV4Z0w7gr6v
JWFQsxONxB5ULMZ9nZoKiofn8vPX9GsbkfUQiWPJl7AcZVZhLPv/SxuP+ENoiBTHg0hF/Ul6+u1l
k2UAKkVRGOQDaUS4hM35EWiDdf2ReyWRmheR0W0avrSvna3Gec9/pVpR5hQIj+BYiPwUf36vHGW6
qg1NuXImL/c8u7qrIN0bI1FubX0uEdjLf2VCpNlpfwHmL4cAkr2kThLrOI/n6K4kWvnRmtHD+PK3
6DUwmOIV25Y/eifacfFUVgfUuEtH70DgvafxrU6iKgwrPc1TfeXXORssMCNGIo4CEOsUkgAnxCeN
W0GclBy92tiggEcIy/YZ174dxflTgXLv765mnDFsm2mk3uqr+eIg6IKYd3QoZsREVa3sJ8uRz+F+
edVaO0QVk/StoUsAJUWptQa4v20GQW3jJGrk6bv9xzU0KUnSxhXUG32ebGJazPfFpnf9eDyZzycR
N8gJ7j1mGwg+nMYWPoXnrBDb6NPfwylqwf74xI9I/3IZxLcBm9wmn9nZg34277Yw7zJyhs91X+/P
VlTHEWdLXwFnkMvLTDuN5we4ixCdHYdf95t8DKBIovz0beLtAS3feLQhYNHNmjBCSIG7m+yoFf5+
BzLU8ESluvjMmcM1mXWcS+mQ2orvHQYWAk/hKQNKbA6zSDtYl1cSBUT1TtwE5eMAS3kYe3KaZR16
ATxAG+5uBfojzRaAQpMPk5yEKqkTd0MuC8mtKCh4KTscjWvqvGbglhUUqUWkJjvRya5/6thnselg
XaqxQlvUakLSpnV6nuoQ58ElF6UOKhw0zex4xyxoxb2d+Qre+8qMLL9UgdPoxscK/m9n91IyD46U
ShuUNtr2ffslE9Vv1X1+Vbuta0Dot+ppr+LbjgpUNubNH7B3Z01Fpw6l1k1V3f8lNq+sCOy6pn7Z
b25u2k1derclRQTEKc/lv9SoEfro7EfTmeueRsDpq+kj9uXlOzwX0BvsE7eJgN/RtN0au1uNk75v
mlkh3pyZd9Eiczu4rmPDDhETUvw4/wuMhb2Eyy2It1UOlo1ODbd/FCY2Xgf7oLuBq8RyTjIElATH
Tq4WomwJYOEw/DMpq5kXCaahgbkQlsCVR4H+lP0EXsR0Fh7m3Cv20WyIS9zIw0lWmYOcdaFLHloK
SDm6wVJDc8EXTHii2GA+8flgyZu/ySPJyFJjjEfnqchnErRHj5wEbnQ/uJ7MRL5+jLRYgPCeXsOP
UTjRSJr8/TApNeK8cfg/hgMqgZkDAv2YZwGXJFjrG0Vdg8CQ+LqutK+asDKb/2UVvtW+fHXRgKdx
SDpM6IpXoBK1ihY8uQdEYmZ3QPAGOkgT+osXPcRkCaF85dsENDOc1k1kpn9SlcwsAzbi6VBBZMb3
dLU38PnQOpbXR67IhwEiVHGmeDsbWhIBoOTJr3qRjQxF1fDtWeiO+n6jdv9+l25JGKN1U64bsN1H
6E/JVzpsimWYMbbQTqRhEQ9pRQXTFVvblJkbVk3CbhUElfjAVZdGWY3GU5ULSaEm2fepIg6+fE1m
pKt6QczaEkuAJHUs5VV9niGVxkiwpbR+84ourgVYafUe5/0syvTvVN435eyMZHgTIgsC4Y75FWrd
rgdcFbAFqEPGD/B3f4YeO0xto9xzy3eejNN+KzZknjgaBLwjp770z5ANwiEThMO8xYBvDuiL94fk
x5OS341JHnIYN9LDS45oYuiLr+oVITVLjlL07A/0fo7opTMDl4cFKCLAas43gkBEWH2U1JcMEe98
CGfTdktc/9uSsZHabhgQ+fuTG4Pu8r2D9hArdL8EFRDpN0EqD3Xx1fPzeZoD7Om5VeQTcCNTIkON
/tMcepbYl7+J2rVoyhfvUkkqrzmiH0oaV4so3o8kr0umWf2RhwuWgU7BGr2JSZ0MXEvL4RdS04Bd
GoFMEpWbQu+PtQQtgUExZGTnhRQvXMB7kT6J4GqIPbbRP9XVhRjYRJMIYUkUjjPz85AItiWob1Kt
7QDAv4jirIehKqYqCBfe11hKzib6X3sfjGpkNr924qvUOjvz7hJC1aex82YvOJmlItGcz3VVwjvW
HN60rLDtpHXDhjpIYmTuz3myv+Jp75b3sRDdlX2xaRG6K/5JT/Urf3XoacSFVnH7IakUHLXkBLiR
HSwDHPOf9z+Oe1kDxi+DI4A7qECDw8qgHdhX1DL7yRsU3dfph27NcPcQOzSBJ2sNDz0gAj21LqEO
XKfTkGtE0QzRdOLR2anaX4RKqXvl/HYj9ZiBiI+8QB0XG9k2H8ff5TdTPQE/XLZOdgy5deITAw+a
QRVBekAfRSoP0NucENJn6+F3v6ok+LFwg0RNfkU4fWO5xqUMGAREQLV5Ean9IRN+E9/bC9KMEDBp
PYQjCvjm9m8e/WzJPydv3H+7gxXSzFMxqz59NwBSWw4VJ+uBxV5dqht3VS/XB7tsC2iVfEjc1TTM
sWCi+pm/ndRdIfRSSwJtmoGHAStZpRKFkOEAKdvw6GTssuQR6n2RX3oEavVNZrgYUFEzol+KJPm9
VVF0nOIiKZG/crp6b9WGOTgpAfEwR6gWhkaR3nLoS7qycez1yWLTyKeyxxuIvNQeU8UsJ555t8j4
mz8otxnXCdPDQhrX8W/SQgAMHFCe+yuo0LvWGflD7uCr5F89Dmtb2ipdMpxARzw4g1hQDZCeBgRG
UhG9alHHU1aLFHRAYb6UJxkj/YHXRMkfRC3Lu4fBjc4q73UdEEBOyc/wYXmu3S9+ELGypFVgKqn4
1IvZeywK/fDoNFl+dbtmrjy0WYqaQ9NiJ1onx0NnQK3Osv8hcexYCrRxv+q1emNU0fQHsGfDu3Ao
xwNRzCNDUijIVUe8+MAEcWsUZM9mYKH96T2nhueMiEjERjz7NvHcEQqj+N4jVnYTh9wyeJmgtKSZ
NAHTbqX8khJcmvCRupYtbQgrKRj21Goc8fo2YWO6q9oEV8Q9cZlL5XBe22+lCV5ZTWBr5hzoTtNN
A4L7FeMDqMVXXNM19r6qhh/PILvgVBcYtMhauc4T1batc5IV2sEtjUwjtgrcftxbqrTQwZZFGUJi
GHzUz+/VC7UMitnHKbLm8pya8AGtWYnhEUaEiEP3h3w+B3MoR4YaKgDrncCiLfJhnQqcNQABzcIU
mCui9gZLdx96FxebJmj26qPBjHuTyiuvnFK43+iMoLYpGCCvNNoaoSYLuMx/w6b5Ivl4xUV6MkV7
+o5o+aOUgHcvh8S5zzFwu8rDa8/qJ+MWfnkqHmGpbghK/ei75MBuncM1jdHnZGVV8CAMO8arAdC5
gB+e7/9oXK4gdjltKiT4AityBIcaW9qCQACC0c/S18yx045ylWd59WvoEBWGfKHOMdKnLRonMXEw
OvhVKWgIInIsya+NKyTzA9VTcn8lQ+BcDq6TD6zIGcQW8CLi6RMb57+XFmUSdWgQTZe5uHKC2xE7
Q2n45o2TZx0a8ylE50yFYFEWS5Sg919s0Fpxy0gCLOly8VcSvf4s4wkYiV75SwGy9gCC/5nRqYJx
QSTdygWLybGIhYpQ5icOlRrQtCDcrrSDBzf3kWFMqAJIh8grpjQdz6/GzSyzvNkfaLS0k2RmdMGN
eV57eqTzVQyGms87m1xlMdE720yko/XYHgyow+eOBiAlQYlC6pziNt79EvwPJRGfwPxrkY4oGY2q
vHNJ8pNpYokVmexVRQD//fokDvphZp1FGNULFOLU7t+cEhQEK0+OlQjI2WCQIUcilBfVWR5rNu7R
oK+L/uVHm6aLQFHxS6l2k7LyzlvK2qH3vMjrMWnWk3xbBrwC71qEDBonHIDBQi4Q1krodG9vrXU9
raN53VhgWZ/rFmOSwxsqKYIyY76U1bepnTZMunq0l/M0gcrdIYr/8YPxQObYFwOYsVCOPkS4HL8R
3Y9fBj/hpHiWuFm8204xO+DE35d9h+fgGUE5mWQKK1IDY5tAL3ob4ogcPeaswJB/FNoHiqZDRDPw
1qxu1eJax31uR9LvgI+qx6jmtqqU5v8OGS8IDyqWK9asfUC61Qa9Qpd8RJp/A0G24KhUo68fhQwJ
atiLmg3VkapaA92qHA/SjfRuKpHC1TLV2Nsp/gdIvHeofGWUUWjpjQaminl4U8AdK4fA0cisEmdf
DoTObGOrPyjsDjuAbgGiSLiKBgc+zSBo1RKG3Imq3hshUooTW0Ur3TtRjGBh94XcLMfT+IVhJ0+Z
al7vlzCXpwfP1fZVxgmp8IBrEm4ZuKbPklNA7fwM24OVVR5W/NoG/c630Ya+ecrazShtqzoT4VpZ
iG4HbIRnNFIuAi5gehA9NkJ8Y3crokYwta2WHvc+DUY9mqVUoPJ2qkb2tzdAD1MRklI8QB2jeCpX
D/pqxE7upcvReS3DfKrp3O2w0MqUvhcOwHSgYbE5tTZIuNQOhVDq/jukNI7+HjZM2dEU45CKnj1I
KqUJ6BvPqY4fkxXzSm3pRp+Z0dOeEjuI9d1O/0VXF3S8E9j0JrAVYrS5vAdYP+l89akUf1jweE4n
D4kjM2WJVIAkoM6YWMtT+oLTzFEUSW6/IWHRydeIBZmNPo2nuKfvEmQXK7eQGpIxFVKbAKLaoL+o
wTAi1GduTbxzouF1d6Mje2FSjeoVDUr24hi9kTKRGnPjypaCWv117J3JdJe3xV/fMZLx96ACARTC
k4wqjBQiPNZAaghW7kD6y4O1ojEA1YYg8W/vezZFMqlCxl32XPHoz0pPhniznglbFuTLHHwE+jy9
+kbLdCVLE3TkhCP3df82R6Uw1DsotrcZFFvucWdoM4/yF1oC/RlMBY9d7Ma5paDTP7dJH8XqXhvT
NZffEz5G9xN2ByXvJDlUFGwVYSQnzFify5JIbNOYDECHwuViXx1GlkvNFkiTrAvQtjmBoNvKElZY
BIjYk7pa8ZqgWuChHLGIyuMWf3px0YyUjX/Hn0xyhvNbqqVMBRE7SQhoXg/tERGbZedczVO0a1s+
xpK7py6CF+rId3qFxncM+bc8VZl8qUGzS9qlIRlGzEL1JIsHxgmbQdmlIvAN0vopto/0hb4adovf
HWZlxEbFM5DsNSIJCgPgZjFvciXxBVCEU78wp2APFLReA6Dz9WxpcxtX1hJfv3Neu1HYlEpZ++Vw
SjnX0EvKecc649FpO1PAC5HghkncKvllCwYNxir7KYw0l0ajZ2s5XenyE57cOgyKdJwto5lqlqOf
4OL/8+DpRg5O0pbxI8hF4UE0CRnN7cTsl99kX6OaNA5/l5F7bc0cgVMksL7Z5ilEVdcgS6AAvouf
rXhflmRjLFOQInzOEq6ZrrlCDkKOiA1kjQRTIr8Wfk/H3e4YDOJkE5TYvdByirDdiCpTiDdA0SSR
ac6DaVVovJ+W3KJOMCHxt+GPldGS24wkrbpmTlBqu9F1vfnXaJ/0PabiiCJ47NZiGha05kUcl/uO
cgMOxJjPzVwkMSP1h/3xi9pfwdlcm9kJuMvWkWI89hOa4X+NW/cbN3okCFaGdpwpBj94kpCRFw2B
0nKZwdMkqsxc6+WDurPqtdPsylLSuWg3nPW71lyxFjkvsbiMrQF6ldDMu8vt3YpY+Qx0Kgle3v8Q
6eRrYjG8yuSMdCVmuj6lpZqG7CHHg3a7O6S2a0CQWtWNVfr5jTzs+kpZVM5jjYmh3OVKAZ1cC0BN
J4HH1GNZcp+x/Wa38lY5W06otWem7s3myXuQnOoJEbNurJxi80WCytG7SS8Frv3C9Ma8U5jI0LMX
GGSmmQD+tHoJI7j3XXQVaWfn817dM1TUK32eruw8yscoMd4FALBgDKqdyWHcM+JcKqDYAXMWlhl0
YfaCHoAF8VepyTv1tYwIrq81gWgMogjcE9x1SjkJqdqjKLWNyb9ej9SFTnjbwxf/2u65H2UBEjTG
MFQTNf3RHmXxhfATYSjK1yvvldEJOLSUF+LaoCr1tVKXpyynKeDpXUS6mpqLxLClJ30kC9/y85Db
OWbbtxW159IZwoqUVCZom8nM+k9wgRoOF6BfVP+musSJbcvdTNU3g/2iXkL1/XVqiUMZlr6v3FB4
mQCZmnq3m07YjhN19/lc5Y2vggpO+Z2ZIm6zmSYIe6ucAHGB+cafpsGqFapAJKCnpidsqGHaFieZ
0HbB0hpUmxFVPfvo2xfLTbGb0ETzLEDL/2WIkpiaVB79at1000ZU3xqAWnhFKvaf5TkbtsYWhc1b
JG4bimtlM9osqd14I1HZ/zGwWJoJBTp7kwTNGbi1FK1/wFe5EL/T0KUbMyCscxbO6IhMKQL5Doiw
u5qK4jZjiMAHGa/hbWvcQq48kEgEB/AZvf6wS5jQguPe+XpxO1ou636mn28JsXLVtHGRDneKQMhb
xlqMTd6FmJtsAYOlyARWFYWb9J0GD3f1zl4f4NqtXm03vONoa6pNZvGocjaompQ3drwaxnvy4F+u
s8RTqmSFXMT2xzmNUh/aA7K2C6wHKZPPbDebeg7ffwJ5ui8Xuy/l0GMXp9OPZYU5RIK6r8scuo48
eX3ONYdEcg/ZSXwglng3qKw2HqoL1GYJmMSpK+g4YKvpdQ+j9IqSaDZqQtfrjblhhR0Wnui8jGnd
Lh6QLTN68/IuinSLrn9R9H8MVwWrU3wc4MSdCwNWNig6JI1Hnj4ger7WovfcGK9o5p+nmyNFx1A2
3xdOstMRAnQso3gxKsljM9WzaZRCXelRiwU1iIVB32bTtCv9M/qWmHqepdPiSPLu5FuCUUoV09zp
xvP9VnOvJGF1AMdSBHmQ9qGu8JRB63ro8rK8Cl6RzY1KrODO5uXmfB+xVZsIKxOrRro5D9OVRrhg
tnd8SCW7Ia5qXDR+jUnK1t2MnqlMlaZf1/1vC3qA8jDbYw32Q2NDuftSEV/lF3T4xUFbe8t+m3g5
wxMT8gib0qm/h3nhQVl1yrel4pQnM3ZvVBMvXJYLHw1N36mzotTX7pUy2xLKG75PFFWUOLA1OBw8
ZnR0zy6MH4pe9WTwTGzZDW9sJXB9GaWZL7EIVPrHhpzZ5HGhi7niO8uw/cWOY2Nk/mBLwFVDnPFU
txy/WJlLvidnmkCHvTrsYvccJBEtGiP3o32sfUJc5WgvXNn78ODq2u0Yz0ODYAFw5Qz/AEkYBRrX
WfbgFAAydWKrMoNlEW+yTH2S0q8ELxwgLTfByJr9JfHDVnVU96i8xnXRTjXGogJ9NHsggJWF/Lng
7CEC73q7YTJzkjSb9N1KFWvvba9HEaFmVLo5QubeFpnv//gr7daqkDJWQLJXp1HwAkWsljqoO7TB
2Uw6HZAq9dRemFaym8IImAUvhW6BkcXvQRHdcj3HvCms/JOtvb4faYa3nh6QD1iaLfVYTEO47B9o
nwNtSChcuPzhnbrwfnXFIiGxW/Wl6kLWZzCqN7e1ftoFuL0PfoHHMi8piXqgHtusP4ZCCMN2/A7m
1monGcm6FrZw6gZr/Hwd7qMvEq+WG1Z8TFBUKaGkt0QR18CiLxbqObhaxFMOCbxwxfROhA2jEb6I
ecH8X4xUl5+1vwpwkgDoXzdIKfhy7/IINCJvDjeK2sGFysIUUDcrYZmCpOY1gf+BXA903mDs1yvY
cBr3dtN2fDJ+QCMJfsiZ63GL5RjNkNllabBZDpOO47XRCyjnbdFSMb/E0Lax5VzjVSfOT48pLwQV
Y3nLs752z+5j8tZy8jznwl0YXqiGW71Tpn875YAlW7tHQ/jwAV0FXvjXazhmrrtqcH3NrfHRNtvn
mBkEL0dDxKdQohasqXqz6+XIUcmwxW1K3Mu/+g9aque+c5buhrQELhtnzxHdU+ZMZ8zA07nIce4j
hGFFoM0H3jd2ufQR0lZLvXj/msGbFQOZaStEOjn7846gUTusMcLHWC2SbB4V+qYOCEgmlOqbJBk4
0c/ilAnrwPlskffNJXsiwJhbjGtHoMsfG+IT6xtpFFckKZTEvV+nq1qwXUujbX0Q5DyPaOE/HTWw
RVLVMm0p31XX6CYPfkp97Qao3T2nUJOvk10HjeJXkJzqQl9uaTbuIwXqj1xVW+RynCaKOaS4ahaf
T5KXs1xmdgOh7vtmu6ge+yXAEy7Wc5JDIrJFaHgE9BqQ+48969XIH9IZcSKLHrlPnH7Jqtg9ijaV
53GY03vDdHQYngOtb9x0r/TZeW75UP1s2Ur/OlKq4qzyUfzdz04EmyI7v2DwC5hy8qj0gXK3hQJc
lqqr73SKrGTctQ+D8dZz2am5WJc7zt+yetamulist2RjqiQZmNCHFWFLrTk3CKbVINJYoNMmG4GG
9RbqpeG3JZpXIKfr8glraPV/9DDvSmNDn9NVALdYRD1kH/gJH8THGmZTRP3DuSwDhpGDTfJ2FvhK
XdK9Uc+3LtrQViUdOezaOLNNOUCbXTCltMmIuGxMc2f64fc0nNY/am3K9/xv2Vl8TWb5oIoHPIv5
lt2PAj7cS7qA1lZW6Y7+0omCtSf4SQaFswbd+pLj9Qe2K7IUf9JelwQLjY5dEDclgb2rt9Dxiszw
oGeWmf8vbFyl/8CJbNlUylkeSxnu57xawDd6KXYokiSqS7pZrOPDWrBOrs2zzYW8YL18gxsnU1Jj
o01AhOCPZfbtymMoV+ZH0/SeslPlmWgVikdJ8Wi5Ybmq+C1EAZOICa3Z4RpBkJhvwD6Syy5WMBgP
4aVFXTBbQJbXVzrA/NyZ6LHKE0VKpKi8HocdqAstxJXQUWxHCLI6F4w0QKFwXofFyk+woPQnwO4G
AFybf8RWnRZWoFAUe+3RQXORuSoldqF/sN+TBm43lTPwFZKBw2SFyKHO3nuArb+BbV0ruohAUw7i
vUI9hbnrWLOrWXHxAhT4QfpL1JKD1JrGPcFDzCN0xq6wmP7ah/37GUXFiLJdQ8I4+WCrLeBYvp4P
CqsMRnanmxpVOtA24pDHr5V1tEHJKeSPMWSN/+iJEPZxJ5F80BasimKK8ZOYxcq5EJd0HcNBrVbo
Vec/6e6SFgOPMKan9PtKMFlal2CXVT0BzAQe9G+9ACQ8308RgaUo6yb0Ij5FUxLC+ZfIeYaEwmvi
USj9JBJM2MwQyz/hd28Lf2Jon4VEbscXnFa/Q69rydEB4d+QJ7nyPmCLQ4npqC9wfXOW26mStUye
kdWsK+mo3qc7fdKDPO5mBUMCXM/Dm319b1FkB+fqscvhis4O9szlm7O05EGatsB4yqk4caMJquRf
pcLQDuTgUSFA7Eo7gbuCeZqb+DU0oQw4CrvdUTKMx8cXdnslS2u3y67zpy39+68deZngk/TWpGqs
hXem7IAF6uJCpfy1TWG87jryEmT1LivrP5WZijw1gzVGIcpEo4Ug7/MOLo0QJ6yBdcyEtR2uSl/K
CmmKNZ0SyWnnpNwVw8z1tteuiNcLtKAG3jN+zNYL8twqLu65N5Nskk6AwIHjC2t2L1OVF14BKmWC
I1fyGRfo8qIloXbs3DmlqNE8AsBna2kJSrkQF+RQOCWsMVmpllUcwJ8Y+nQLJywJZG9wjwTOGUEl
GglvoCJ4stwXc6VVLbB1LIkC0hM+zw5ZV7Zs6Ekut9Fva/6Gc1zvwkFGNKvMpSQOPVg+O+erfbz0
u991sXlImnHI6YjGvhDkoV65DgL+OEhDncRW30ONfKWDBVH4uCDsaQZ692HRnHQuG4bFBJszKI3J
5cHxJfgjQ1ftyksJkZow78Oo7BZYhhEsp3kP6puoMP+KLPjvgMbincUPruNyGVKAbuxJEmMbprnE
EEKupXZfE9fk4vq3xe4rjt6H5lyCIlc5+BAHjwrMZvAaHREIQQytXYvAOKHbqP0q+orEUqn4buJ9
Q+yPbRa4M7QyVhe55fGQkFYe0tWeG5EsMvbC07yGIpwAycLGG+XLWF/2h8qyp+3TsGs/DPj96kza
/RcXxv+7Git2kAef61kdv1eTM1WuWceVR/sCgvQN81Yr7O/PWLqx3ifYW2RHYecucINWp/V7m82H
nNxrB2a73YVnVZ5s0xLmkw9HLyxhPZNWhywh3aaSfajzjsLAEKKBp0ML6AY5itPI/gkIohKHL45J
5NFdyhA9KV1za+GVNRncTlw+rfi29PfjhoZ5KZIeuSNEEv86sj8ezM0TlkItgM2kQMIzhs+ua4hr
ReBm2tG1SEtxahrMrsWf/zvuNqVp6it0+QVx/mdS7wTZhcZ5jiXv6KNSbFVJ7xMxiYLK0j8dZkcA
VvuE8oFw+C9VjONA70vngxIjB7fH1jCXQJba4xYQpW6P9gewt7gI01c2iyYbTZOsMB4qAmzZpm/p
hHm4Oc0MW8ArK7Iv9t637J2R1YeDOqh37RlfJKgw+cvGY14wy08GY+hcgKaz8qdAksUqVYvNpXe/
wSo6uRcUrNytMK5Qoz3v6GH93ZVpfiYejWUA+NNH92AiqCMNNLitcKt5rNPzFLk0BRv7AqcU7FF0
fJ5TZxfO5g9hiHR4W9Z13KlD9k9EYqO88o3EXF9MVUjDMIAO0MdhOKMBJ7hIdpAHkGT52zUNtbrd
6KS8EoML2Uxuu1LV00ORqDpW6Uh6pCeObKd5uaWckuLlB3ouxfKQg87TuAOnPP4nursuo3HYf5R6
FAr2qYnJ9pMQ713n6cNRDEb9i2IEhj6ApkLYauMFR0dwGaEROPcZv5MMMQ2EQX9pqmiyHgYjmL7x
34yCRDXGwarvMnm7F11nzXI4YphnJdUk+NwEYMlyF/qZ82LhIIkBBZsfd9mS1IRuh+tUZhzJU68Q
RAkmTE6V4FXxuL53YKWjZxmbYNe7XI5vPDCIuOp2EYxWypjLk5Oj44YKDHbEgEMM2oZHttEDW1hR
7FqMKxKZKF6zBywn+VBB8Tkf4qTaR5EZmVscLGKAGZEKNIIB+/CNA/Fr4H9vsFgXzo7yrTipjo4X
0aL1ZOA4zHbkUhCTqeasCbzOvPpctjpXAPF7e3vO0Xb+UyTBHKFXlmA5aXc6TNJUyTHonGkVLCvV
tPax6mh5Wra2fWX0j9CVsxLwLtDE08ahFgeFaYhzaRG8fljld7OFtxjsXivK0XSUDRD8OCX6gwPM
sRu84vKFOl0fWhsVrUqNyyVlJrbHzE+BWExPjhBKKTBkqwBCMjJeDxzg8+jU+/yRIWxDPm6L4tgz
l6Gn6jPuhNYPhXmsvK+YhzcBBlzIBy4apPsZGnSIvt4wKDeXutGAgsxn5ZTICsMAMZg4VgyA+DST
Fvcgnuo7TsEWjPOeycrwWsi8jPc0iX9stZUxla6y0wFnd+4rihNrnOjS89wDl6fb0PlxcKoxWJyJ
zgZ1AUtreTFOMMCFNYlVuePsX/C6cQFFyjv7zZw/YvdH6U2fmUZTV42gWAcl6HFjJF04cQDOVBb7
GH0xuf65UBjKlBGOQDQsCFtVZbKJbomlgiy1DjWbbgP57e4rrJZ5I36y+gs7JTmerGvdv2aoWbxl
vYh4cgOCKS0pVu17o5YaiHSSioMRhh4mmh5a3t5n0pRwpittTmiFzcyTwFpt3n6BQ5TBoTkRa5y3
XSoLQpZV9FDqZ/IGDnZpNefG9nQcEuRdd6/+aE56bP02jPmLLvhchPDUPQkg5j/PudD3FTpyMM+5
QW5TTC5nGV3v+Ic2UVoQQZu86paEVHRHtiEE6w66D55cuMUe7R/URnBJrslNq9S+gONMrj1KOeVe
7GSFTKZr8so4YhKIMCXCUK1ZNy7NhsMhF/IIEFi3MYAnPHdw8t3TydAGpsAdZXa//HWl9NbP75gz
S4wxKvr+VEa0TsiRdZqclYVmFbJHVVKuMBI7D9DJXyly0vjD9Ud40QCnT8Mry8Jb7dhNWxAtNKYS
VrXGLQDJS04Jb6/Nk5wF7ygrOiGZ5+92cWgBQsLTEKaP5LnbuW5Vy/00JSJW/wAxUIn58V/61c0c
5Vvsay4VxLCsbu2dVle6mEo6OyvrS48ZhIZovLS8k7OPT/bkzycXU9anRCCTLxcZG0NmJAL4E+q4
uJYDhg2kva1ZPfJGuypmFJ+LYfzg6qIqnPHj1/mvZ5hdxUZ8DlByuydNfLGVwIK75ar3viqkFSJr
ED7Z4yFgzJlQ+kJp7Bkk/0aU0lb36RWlJkzabkori5zOcjGQLRAtS5U3z+uTfXItDXrB+B0JjL1m
4MDZHn79NAUm6Qgw90QRATNnqmbaV49RJ/E5Asdy7nWH/qAxQo2tDg/M0vvoLosJwp6VZeaXLGqC
B7QbdxwLH1yPf9+JxwDszQr4+USkn7omuFHtFGJUlXvD3Efr9/yCqJM+avgWYYz5Pg77gre5sYeZ
O7r4Lh4/KJ+qMauuPTls/eVnEOtxlXbisEDsNJcRFEnbVGb6fjmMYWqdKguB9nhxT+9pFDqeOKLI
OyJpCNqxP2BBSJYqT0KgYGKuLedLKym9a3AsmhhbzOOC97TK7hhYYOVFypcg2w0L5tmiixZzhBJt
PULAMKe+H5d3WJhbUUshmRVCWw6J4nMHSHpTiASASRqWnhoVqtrVqT1yLSz7gQ3odlIi4NM8ExdC
7ZeHFdQxFdiGJ7tr2B1uj8Muo4ZiFopE1zkksbvnCdYJ2/i9bJarRPJVpLczFpuWBZmQ98Ma0M6N
fPrvbxTo1YOKDrTCJ485BE2on3P7EsBObVZR2tVqYuFrMjBA2UvR2AVRBXErd09TCn/Elxtgw1jK
FJxGHs1ZTbnrc8YrQc8fruTJ5hYkWvsvyYHcCNfdqwaFxmIJkzJvQGeKI9yggX8v0xwop2GHu6pA
FcUlSvPQnVnBJ/OgmNduOECCVzx5lSDHEOUm2WkWSd/is8szMWw03lzjSs53lnRi2ehp9yTzy5bK
Ov2L2LrNbtQRNBKYZOs4qbL86XOsQH5y3N8bkB+oogrNu0ZJw0rbXV5121Do9O/YDD0T2Wtvv+s6
v76RR+ukRcII5fIEmpJQcPi2EaDgqpxnHCt+Ozuw6CkAputlIu6lqFvX3VsFdHhuIdbZEYLug2rH
t4e3EtbDs7phk29Ytm2pQDwEgWkkCcGpK8guLLT5mf+m+/N2HedHoy98Cy3HQTJg2BMoznzat1Mi
qkqkCsl1e5Lah4SazeOiY0hrJWp6N8TTJMEXEOnFkA2AJVAhAjOTE1ySsnwuNqZO5ivO3AQHNobh
banoagJLAJnH2YfnLDtXj2p/TMCuwbObcfSdX/287HQcMNtn+fkE/FGeBZP9bb+MkyMrRdw+x8NN
70g3iJE6AFUoKNFnQUR1DGoN5VLpCc3hwyJthHR+MWlRVaW88vv/nZK9yUs0f3EF5HfX8/l0YyZ7
QVwdOd5yvtpa+TLuUq9p6WNzxYtc5QUyviCaEUx3aCiOMemMudaBY1lM9tRFKzOkklQw8LNPM9sV
umZYF9cAxLF69Fw7SGgNix2J6qFf8KGBDMfQfSt/CPS7iQKMT7hFl9g/IVwbN0JHpiuhuv2RM/c3
JZGtXagLWro9TL3KRtuC31vHDOEiAY3xvjQrJ9nt4UxGtibNq8jQJEJoR2AC7I+j0A5nWa6dZdJy
t6rWLuvJCz8QDLkNczcSU56L+R86s59krlcEFw9lIyL9GWgDZ1p5mMpbJRXJOAwIblw5ZvrgPrkp
vA/kEywIf8FD7jk8jjlp9XYiYBvqsBWfwDro72bZCli/W1dN422amVSzekwVu1S0e1PCSseNS0Xs
GMjDzoYryucsDDhhWbdmXKZC5rAy2TD+8Ph+zHcjBSjXmXjy8R+DGMK5L34haer08eqlXFj9Y2ez
fG37TIZqj132luu7dIV0MQwNVrCEro8EpCveo5bw9G91bIb9ypvogH8R8yxB+sEkBmBWtrzzFSy0
gMQosXVeFj4G4E5ezF6CKhsotVCNuwwdIHPXnfKmtutBZeDPUY6hfU12z0ugVK4kkKo/o4lYaCvg
8P549ABxjGc4x6VS98l0X5CqMAJ53eXIxdZPNGBoxSDAP49J7zQhKkFmEylbVVjGyc2jV++eTRxX
8wW7ZL7V01YCv20U1S/jIYM90VLA5M8hlag/v2kPrJVXvJZFfufg+e/+H4IXBTvBzrsdRrlEqGWU
KvvL/Fzhe5LJkhJrMLnj4RqNaOk4R0abbXI7rEASxEacecOjT+tpbKN1mr4KAyMrwXk2M6xi5nOs
E5vsF/DJOL12rWCilC6pPNx2+Og8gFX4azg2aNPbpKhWH9RCO1vCON4J19+Lhx3yvACtw6jYpp4A
MW5W5sJ3oOW5juTK71JUF+3121p1vmfk40QCv73tLiIJ7/2SJrAgMMd7kVNxvtAd/T1xpn2vrr8V
fp/BBT40Rf6YweC84RNM4EsTnBHJfnYb/04/vSHHW5UthBW9k/4FhsP+RNh3akd6p1LErowFO8iF
SFe/pkMSMlrWCJP6a+51iVS+6ZSFcwosK93qxurgnNMhRRqUdP0GifoTTjaBM1eXBcE6//rAqc4Y
7A0B9kVp0SEz9LXxRpRUZydg2R0NOjodaOmlirHRzKl3ud1r8H/GtmYBGYBCQ7QBmHBAFYakfxjO
/6lwaoPLv69tGo4vvzFtwocRbyXsQ7OQAsPtCy6UhMPOLsLHfCw07M9gKD5KwUOVXxeMHnNb4kSY
CZ7HqP0IKYR8zInyRUKl5BWxNYz0ALL3WMqIESUbn2PjSL7HD+AKviyneXlbBiMZVLvXkXAynLlv
L+HC0X5NRpuQAjNygc+jqNHhadjbWpJdgWa6vZpkw/uQv8Xy0jSyM4IS6TuAwOINQPzWlZTMqzbN
MC9O2uCo2+v7tIWLNhvWSFNASjVaXYx5wLkOD+1nPeQD2AsH+AQ9ihcu/sq45AVeTJ56TNH6hRNw
4vEs1xuhggRgAxIxvbwWqNM/xWHXLMqKh1caiuezdtnBJDO7rwmverdhahzq1A6bXQfxc4hMpQQ0
M+STVbNeMo0m7ULpJk7mjZtGMQ2xhE4YB7ZD8qN74JVjg7FwkvLiFLWu4Hmb6Fj+vxHy3pGmbUN4
oIiUq4/aS61M3FvnQN0mAq/ZA2mRTvJiWRZKFu0Vv/I2nN/subp2xh8ZML8e5APGAZ0rNhifXrU0
3u6snuMfQQDyhoW5mxCB1WXKJLr9zm2OcMFIthB1FPJ120Cmmg/nSidR0Kgd21656QuFvdvYHa7T
soaAyuU6mBPMK7tVaRJ3jCU/jD60Hk7ryC7Fdh1pqG5blpf+SX0t6AZPAkpAh2XD277Og6rB5vyE
TSYbJ4Mz9odVlnIoqMroJrd2f05sakQnr2vVgXHP/BIr5qvgCPY6c4q0cnfqt/bPMVULKVc1+cXZ
UDTGLD+C+sxuDSgsIbGQwAixqg4BqR2eKkRr7y/0se80mAPEBoMFm7N1ATicneKm5V2RQrVGHXs5
fWMmc807THIAJsJetnxjdfru3Z33EmOgO6U3f7xnW116L44Ds6gzoQdW8AHd64aZCyalbWPdnCqi
uYssla6XfE3uqOHMq4on/hjrb2dJK1M2F1nS7lpGCXAMR8qf5Q1mrqbwIHrh1qJV9fsVY+EDtqG8
RX35Lo7CwjjWZYBIEW80RUN85ZAZTjOHyRLDS/2Q9o3A8NcuD6gcfQ+uc16VQTbQ3NQIULJl8Lfz
I5YXOhEjiyPXhLMks6RqnDEdcZKLh63J3xfQcGIZmjGMLMPWffi+hvHpKaG24OHcwO6HqRTBg2N9
MeUloJQZ1zQVBa4LTPzmqz7hp0mPWcIDC2C8gDtP63hi8+K+d30X2TRStQ0/NLdHbIeZtCB5gSfW
B+/MGsJKhTkOUgld8KmzbPWKlOLjb3mz0GKZqrqgfaq2GNaKOZH9abbH//8Fl8Nnin819zPFFRNK
Uqjvad1O0p8QRPh9Vw6PYrP8DDxchQqoj3FS6IaKScSYa7VMqlm4r3s8BrTCwTp/0B/otul6hslx
3z6mmF144PnTEwRfe1lz/jSuIlYEHh/ihQ26EIJGSYQl5j0e+/4PTNXi0kNCWMM1KeDikEBHl8C3
owHm04SlxTt5J3YDnlCr91YNSM7h/8113WEIc6OJFL293SdqOQ3WoKjkXuyk2V9hQXsmhD/7499z
QSxWCxwkWGjpbgYZB8KPP3flBLtcnq4A9/QOQZA+TWcPrVas3PalSVPt9PgsPQ/NYl8bNZwYjkyo
bdHYZRGnPHK5WncviHGAMMC5MjFbZhsqlceGMvEtIdSr2tolwsaOMLG53EX6ddi2U8KC4iTPts/w
XzWDWNLtnci2DbzbQ6STdfn0RG7HKina69TJhA77sPkYv6EfseXAcwWPzPlkbvLqvKosc2LQYNCa
isXGUHJbyg6wLIIJ+rYVrhtW+p3TToLYqj+taH50Qz4sK0+uhojFctRwD2ZQ9RGD9XqmLo1EfeFo
1qBNJJ/DBHUf1ziEXN6FBYHfBQVESjbYkRNCY5geWFlEsVqHX1DB/6tlNNaANYameRDE+xzVcvA2
91Xx8qC418Z78XsWOZ9FAz+HZa+N60QVxOYkJELYn/SiS4RvmOO7JvSWmX8rldjtUmEGx9ngOeKq
lezjaJxKVkhuY/z0Oe5KdDAGhJmON9whQ/1SMP3ZWYa4POpqQA0jI1YwQ1g2hPh/eV9jFEtLZ7pI
/JfkJBirB5UI4YdYNAozrFkjOuFbURT2nWzs9P/volqhgJlylkKEVIryq0swPlwjV+4lHf0JOn49
gJPcD63BqOeKSgSCn1sz2SgsjkeaG95DCpLSwbfyQyJeAXrU9cO8sBgX+hyFkzRMTm88GHeA9GS2
/l2xEW/47lUfAA6Qeesn9tENOmVRntegeAdIrX2qiek8uC0MXjFvE+XLEbysYQBipbCfCBUedrH0
0Qz77dIZeqk439MMV/Zpb5TLeUVWQurqHSwXRyLxp/dgkmdhF2dPHQegWzpA6e6IL8I8UfK0tCkS
MtuQuzexKmRCKKY+Y3Jwxc8T6m7JmuJFjGgFeXXc/7zzeQrt5m0RCUiWaf9MuzIG+B25THfUGIUg
WBVul9X4C+lBm4sdmY9oth9WZFcEAWZ3P1cMytuMApfQfPjyrrgVnmXJMLyYfe4M4VBn8u/Eoygs
sMXaSlR+CtEfjBoJ/A5cwBl6JtfTMgyi/N6v89InBmqRKzlDt/A8KuDzJzwhdLeEXY60GBDvpaS3
1PQxiNP56shrcRek1yjoA0aj7MI4rkHIs/epjI9Iry/XbFzP0+l8S9HqSgV6MugGRzLxkrqRliOQ
FKHjofxeDxZzysxllvkU5NgYx6Zz36PD1lDgcWLVQzoWSbIvq4dMTxUvRXu1wKadp9Noa6wmUpLz
8QnTeqhpVz866f2Ky28aBbZg8PJdPF7RXZ4QRVk6R6pU0abpVxW9Qm40uwldmjTJh0GnZxE0eJwg
xbBtWIsdgohbDB4q9peNgtbBOEEfrkU7e1g5brf29AolwMXeTXFA8SiixSHnok6Md7155LrilyEV
o+dgLIRID2TfU0QukYeN8LyeO1tT5tWwpNQXrEYFiwN6Nf2wLJiLVz+34NVFVI4iT40N4KdyJ84b
2cj2lXo0TihXPutulKaZ1pzTJMmD/s8C/dVrrRBsYN71u+pvuRhoc95ebIWB2ORfoiK/UgDqGQ07
ddOQqB5qDcUr6Xc0TG6sZgVL4ewJ2RgUzzn6L/9yHFKCQFtTSaZHiNAvOGI/i7wlOuembi0+9slB
Q4hjiYs/se2HjwxaD5mBXs0TJ+kXHzh6aXurrFu9crb66lD8l9+QuhS1nUR7Jo+AzQuTCaO/5hET
kq8MHdnyoqVKW//n3WLToZ3eSS2OVguu9peI5kzqQBdrBVFAiCAq86wUC4PFmPqOJRQiYOErYumO
f+jG3zk2uYWMesViBofxzt9SGFKo7g127DilcuCpKT1P7CGFnco3afD7gExQYb0Ml11V9n60UlTY
yFdrDh+a6lS2JfUh+EGV3V44eTvjdtkprvWmDA15ApAzwBmp48+70btLbtn2nhgCckyK3Da4milm
8yj4cZe71K7JKXcXoOCj8nOojidjS9UEk1C7kKYbbpOkTTjK5dwtFJlZD7dgwIHVJSHapqeUFVWG
eXjuDq56adm0dtYV8ZkvX6Ur4ULVwbihGFOC2VxNAHDv0fo4C9xr9MlQ/KVnANIN9NsgNfWtMR9r
tEGlq9nlsgtII3T+A1GR5nNQ9b8m5jWLCI9tPbzl1T82x5DQJ64TWWlhh4prF0kmBI1ngz5RZcD2
jd9lqDSEFvWsmcWpVRmMGdLzSJE8g/yNYr6ADFIrozPLtxH/Xp2iaihJhq09zMHC7VnPjpZfqVIQ
Q1k/5/PcCOaZowcDpliArlzuUKaln8cM+1tZ9e+EXQZAUlD7MwTLkfTIQdi1f1Ey5oNR81Qe8j5c
FXFQ0csqki209pOkJFD0gOzkxsQ/AjML2CovURkB3PApAAsOSHVJyXjfKSTl7IJrwHWNVvaokvKT
aas9uKhgVW/EOEBm9yWHrm42K8IBPkjdUVsrofpdwwzLkn0HSks6Sn883g3XbjE2YH1bFvdC0k+H
SC3CaQJ7bsXzVilVFDHFccn9FoYMFnlFhHMSw8OCUbhuJBYE7IAsJVKbPsGSHFoeFEOK5kjnUseI
jxdvKatpZ3Ln/mRCOb0xSU2PyGU1RMBfHADiUH9B7RY8txu6x+55Lznj9k7fUnIK5sI9yk2x78rD
0CBgefEvDy0LScZ8dCH0YnfG2+OaSiH3CHvcM7zfEgWCY0GqodKBOUVwwzUB9SEZix+92x4Eofyp
+iB0o8zCEit3VFPr3bLISHrbb+ZWl2WWrTmFXOIHDA4gLFa52BboWPCvU0z0ITxRzzVk1wJsEF/F
naVvt//N9PRhyghHPhK/T2mke7rRPBiVwtbJRbvQviSuYu9v1OUu5mLu80sr6eGx/xNXbDgaHhJZ
aUOFrG5t5+Bk/UJZh2hYuITM58w476pSt+7/lOq62dAcFllFq2MeUfgMo4+nt66IGS87vuqqrFqB
ZGrnNP4giDn7veecbSnEfaw/dZOLOX6AXmGYF0Wg1eAZyw9bqiGlbUIGcCZT3k8bGwT1pYR9qnG0
4GP9Mh5H5FJ6C+tQs2g0XOnYKRqrgYN5Nh4B+R6TsV6pqH5epOYLcmQPFA1+EFBTDr7sPVr4+5M5
wMsUTFiiK4mVlkVNv6saxyAmUV2i3F5zzM1e4wFS9wQMWArZs2LZ0i/GLYJ3lpsYnXqHmbdJ/F9w
oIUdcYkc2rAVA9ibS/97F0GuA8OVAYmrUxmdXCTOj7dhwDfxfMUxQodm795MFLc7NUv9Dj5HGfF2
xftn1vHiGJr52tBuCxQASOzqUWj8zwx++3hd8ZKGiTCtVBbh4YFdcUTxK5ps1kf06xlUDWNs6jMq
UlAz+h/B6kbxGaifWWW6JFQPTClf29FKoHJixtd5N1PJ2qYha2riR2YejebCi3EUHOExEf54vtup
WS/UvPGJfq2jF2uY9eQP97ZG9pY4S8hTJkQfFJ7OTeFbrK0nOywKuob0+LSOQ48zuwt9e8uJ3O83
hfeGVA3gvkVlMWjivuN312q9ihW0sCxuTU5uRgVoF5VyFffFR7lRvDLzm7wVbmfpRjN2NVg7LZ2h
iMdyzxjZX67DkkgSCuCwv/31DawmOMQQKWXS4nkL4Nww3rChbFsiRPRUVHVDfIr+R7oMgg+R137O
bKyZrR2q8PjWF6S66Gn/Sa5LAZ0mCqiskzaK7pSivPezb+03mPToTiKBHYTvb3+3OBzcbYKbRqzh
0ZOS9+WV8sOj02QK40pZda3QyWSvQWrJKycpOmkLMetBWA7iydJP/tpkZj7uBgPRPXh9kum/Gw3X
pwWfl4GUW3656sX2POGpKbgKRw7wE7+ZusgfMXOpadvSnKuaAFP2YSpbx/dcIypKTRsRBNI8fbyD
Szl57INitPyzea1Ztf78a79ELXGY1r1z25kl54jzrsXL2eS+dGV1ICtl2lB5fYIExbV/wlRqjoLY
lFwDrMUHr7yTEANhORD9d1wZ/gNPlTlp4Kqvdjl7lrWDxM6sIuhwekK4pC5kOiF6m7YkZ0zykrND
gAsZzb4cqK0tT9CuvZzjFLswzCRCFSw/ZQUCID/rCkTy1hsstMIqdjyNUXG2rvf6kcZN4UqDdF/y
UhFAPlQq5TRtTwi1lNGhZXVjIcIzG/Equ4gpeBgORz0YjiLuMIkq2baZJ115Hgy4k6ai6vSXJgoL
TkeLUO/An/PtqaMQbotS9vGpFkvaBGOY0FXqjXHbx38lQoYIhhW3Ww4xJxtSnBfje+ZxgutU90s4
wZZ/RR6tSAYr8cIhzeKwAhHFAELoXTDNCRQ2uxydUe4bg4K3VYotGVPuIXRpC6xBU4TNLhZdCIEs
DmRVmAiZpplI66HYMOt765yJ202yen8dpaZzQn3RDgCpSnazZP+hPMvRW+Wc/xhjTcgvdyf38pKi
RCcG9yL8ddqMrTYFQXBP2GUPH1YDTxn7dLyP/ttSSDfVUNB0RqeSyGiKR2IoGBhaDT3IPSjb85mp
ceBI1cwPWVsKUtE/2zqhz/PyyJXyco4b7k5Bv7LqaqK13PxJ99hJkR5oT4Q45yXSx2KlW6+pP/S/
JNPddX8+/bVhBGTnE3qBeYCvtI59rYwyTVM8rfRjxlwvwVyENWbaqoO4e23P45L+BbSbLVnF82HY
1fsc9OqO4IMWNm/Y5sNAc7XZqURIpeCM84u0Ti8HNuIWjSJjHfsLoZS/I3XfCuEJmfGcMUzTMe2w
K8p76eN8XSL4ST52ZS2DKPtqOEqlvAC/bdACOcV2djarVbEAHLVpLbCDkRBRUuj4BsfM32xBNNLt
vRlzon+QByCaBRqPEOVRGrooQ1uGyapAm4ax/FqVMnz0aWAboAo/Ho8xEVKSySmb3MjFUlMd7A3p
IcKCG8MH7MA3f6/HO8VBleGxmDmHJWxMRhqtL/jWNzCJpsH2lncJQg4+KNhAnufSGfbD3XhI0o0D
2XC9owN+O7A6eFHKv3DR+gDWOSwX4uDNf0V15XRepwcJqAYJR+9NxxRP/ZWU4bx7/B7N5hjsQ7KM
wIzLJpZrB9I1NI0iP85522F0K9xapAIyikQsCvqn52GkMrt++vgKStT0quiy0RBC29904xRAfZBL
YVcatElJa68b1J8WVROu7ebx+CnsoTUi9CkQ/pI8Qq9bX4b+YqFvJUtKInybpK0E+rTlM95TgaAp
UjHR6FzgzLSPLhDSUtkwYOFcG4mDDyMqC4XiOkLVm+MmjyXrNzEUxajzY9wGwTpB+nm81wzc9bVC
QKVRhRMibeXMfXp0J9jlSulQWfiT5nxDEc1zpYkx1v+7l/EOTbDWNcZM3WDxp06vvchLi4JqNeYu
A8GwH8SjIjGZ4Qk8XvAEtquG9M2/JssT9OvX7DylfdRgLgHjj+X3ddPWvM6jKU6APO550Qot4KZX
8/fSaXpk233jwV+QrX3zQ5oRAp8r0TWojmCZAM4/sOETVnuZbkf3OhLrD8ClyJvwZ8ORX1WkgX7M
MTTwe+83cN8mVLQctR7HtJe94Ppp+DYn8/M0wo2mrE8dGqD0PqDfiOOC/+OyWIsn3hstvxPju+oV
VPFiqp3i9Ry+fiwSHWoKpximXwh7pRpc4zB1emldRK5NUR6ssPGEvnKukExaeeuFgb/XdFQUSMx6
O/8hbUVpZEpGfVpERQp8vsktFctdcy/ObM788qHmCWPXc6QsVu8Wz7LMaYT1MxzRPDxqLe8r+8cX
szkoa8KLMt5fEVrWEsewsaKEIN4xFc0k7fqx+R7aDGVNB5OYyuDQLZZ73Bl6218MrrD9o1QYjdOG
GXlL7ZnAmm5YCOf0fKd/50yeLspoZRAUS7V2cedVW+LcZqGtwLeOwpjShWptSfrV4OSjlWyiHuOP
gaqtplF+vHuzlIwfAHDCDBLZuPNmQexqIGpjY4f0XT6MkFDh0yNQD4uEsUEKThjnccu60mzrXyzB
3zNH5GxSRvMmnZKB92gvfDeIRdpX8MA9giXsnAFYfAowZIINjuaKwMd71VHBaIzWsysF+dULNGf8
9LpWs2uXcpcBW79hCh3zRFaIcw9PNrY3Zwl8kLS65j/S8vZ+QGipND88uXqgr0F1jC0u4naZaSdn
kwk3QnWbHBevzqMWibg5iXPAgQjaShf6L5/xpbTo53ipqXKGZJCLzvfVjk1PbnV3vocimlRtSSF1
V7X+no2jo2GaaJzwdWZ7jmJvjZ6YaCKINZfv1Um7znEbIewfecP6rxzPiehUq0NaoGbmL/LR2Jpp
GLaksLZS6Qwtw1q9nTRwvPl4lfArgZZW/GwffETP2Bm1DNXKQpxXd0MOjXnbtGe3HGgMzMTNJOn6
LxBU6A3GkmckFhiEQPVI695Rl7GMCUqILao+/r/eY7TXAN2K51GhStbX/epFTnse5WfOA7mPkgQk
96fVlcU1YNoR3dSeJ1b4oQHMnTQV5T80qUeiGfjKPIIQUvp5EUDisGptMsaReKKVtbWuZMn7ea+B
yrLSRoUptcr2EbvzSrf498aY6xhAJwXX1tQK/nGSiMlIT2ZoP4GsSqd3sQbGsgByK5TP7WtHVQRv
dn9rL/nRQ7n/g2hCvoF7K7F62jq9D2DDVmR36wsWfvsOTnB04ZtZm9idW6pK9Gmi/V+hg7+k0Zkn
aSa09jCU5cR1nKJuK5SnisokBzcPyuRF+IMKfDnbS3oXbjeygBhVoLSB5kAtLFISlzKKGVaYClL+
ndT9PVgrhYqbEV4V5dx9m9T04YGY6/VnGEVG2OvQbrOPSiid/BqVvC+5z2qASEIklYwP6An2L4vC
Miygp9nBIqv9sjJLa7dbBUvmoQ5wwKyNcfnqzzHkrBOKRwQcufBUeI2yHruSbmtx1TAGLZZNoQjr
eXlJ059OfIBr5Q2VaVYE/GUNoIHVs8f7nePMdbD2G/GyMQQmt/rpTQC5Rg1DPiSJyEKiUgmNVxVl
FqROwstpFH2ZKQOgsveYXQqtx/sEo5bTZRSq9s2c/kIThm1xNhHXkQx5umQijxB416P+Vytjv2NL
XyRYYz8rJw2W104oWRKWHVXXOWUpvIroVDXEZtFU8iEX+ATJYkPu3bJWdKsHNPlYwo58S92G1Rfa
+WgovHdLYOyLOc5lYSaYj3D9LhTMJA9htLyGl/y4jTvyZoM5jG5cVLWH68gUfcpZqmx2OArfC00/
a/wouOSHgBQdNSbFOiW0QrL6GC3utsCp8LyAUjP3SlhBc0AyK2RKx/168hIpD3efZMzdf0fT39N9
6HoA+MyxDAvFnuN9ACOwGmN37xG1+nx106LnO8mc36kq024VS0VGUqoVaruD/MF7hgu9uCfgWeLk
LO0wLIUnhwDCO4uWamhgpIHZmDr4S4MWwl4R6EUUTZcWPbZYhim7B1b2AhcSyTNmWDqBvsZQ1lmD
DT+8gN/PAQL5ccVpqYvFOmRIkgavE8+jOQOn+CTn4xJuhEJyqnB9Mnw8+np4/EnDScxGcXMk6giu
cTYHFUkkpcSZaqkkkaFPOjoQ4CWUhJkKhzn6GtYPDQFZbYG473BOdOZfavGP7nvSR3bJweWe/9+G
bXITrMGmXpQOgYW3F81mhIqy8EsZg/2a88SEbUCQcSVWFZb0+VE6cchDrJr/xyyEH2KHEna5/qR1
m7/Fhd5U6BGkH+lW7FFOi+AenczaUBjtTGPSpeSBjpOSkjHIWcshCQA/UVDDdcxJfjDwX/oxEEDE
FdejHXyt3K62hhyTiDeKdk/TPOf+3ZxCjFFirJDOZvJY/1X1W9nXTCahzLDcRjhwGRuTm5wRulyi
DLU/kkFiHGl+r446hcpodFEVtg+9k70Sn4uGi1ePe3fv7kBql1JcunuTl57X2pzmZINoJQbR0HWp
fScpbUc701AZ8NN42maIZ7P7fzW+gGG34Y7+VpAVTQizgqfwOnScqb5YpWStdsyy9RdM+kuFcKq2
jkqA8x8EbgSHb+Bu//U+siRSXrjmsv3EDplTiFnU1OJHqhQzR54tqcFWdPXS6kYcZJ0wuUcQvtzq
gd1zLIZ5zFMkJKNK51Niag6FH5ItxFna4J/Ak1nzW50l1bltLyeaPHsp46/CSnyEazqb9ADZoGf2
F9QUY19LMne91rgpTUOfQwP5P9n6MQ4L8NSIw9OfJ8O+Xy1w6MtoqJv7bIMdcM5CM/+N6LsBz1dS
ukn/67tBFjEq9OkEEqJ4usGoQ37LVKIEIrU8esCAtIQYhDf/gdy7JFg76T/+JlbQSzFgMCqy0hyA
Fk7HnBBSRiA5fDCLDOnC113cAhluA2X8rj51nItb5UrBwsCxsR3Wp1VbpWjFnGpFb2PkHKFUOqV5
M6g9/e4IBDlZq2wSe3YMVneyXSyUhs+4aPq5oQ7W5kWzOA9N4r2xBnKm7lPUfzjKJw2DHHZAZKCu
vKm+UDzv0RqZc+9vqJNaXeKTYYlo01BTJEiDuEkfR9uJKc2lGpWpQD4a6dG819EyqP+PvID1civT
sPvs3iiyGItPXlf98jnahfVyUkFPOr/DBSaOfR8JDk41Gl4pGU5M7m16zWgOhud6ocj0mXCeAN4u
+jwZZeR/kKur5YuJeWI9314ntGZfkIHXpV4RJu5Qt6Ut60BbzQ0N8fz1mEdYBrt6bfFP39jc6dRx
6rborfaP7LU8xQiR5A4rmDvMCJ7yx+XzUCVBUlpIlNqvIF+i1aLyTxMPmavr6lHUYdmCNNLB4Stc
bPj1rmlTUbq6dV+mdukP7VOus2r6eOtaBM23wUpqj+hnsX6K9By/EbPbapkozkbfm6ymPS9s/dMw
Xlt1/rFM/puhpbyfeAXm4OrXP8RJgz9qzPvahOBk7A9nlz+nv3L5uGIBbyBdCLkZhLALVEPxarQ0
v0h5EkuVcYUyuQCW162c8o8R8Ugp+pMFdYJpAZaF/niPJkh0499FS62RnCf/SwnXecVZX2fYHGjv
yFVKAvb8/OooMFFqswjLFhl3FbmWpl/74l6SxaJVAd6L+V3PROwOaXVHaaEJy7LFXXMLEJBTCLmg
lqxMpdwGzRH/ylWTl6R9k3IyehCCKInSJxJuteb9bJ3ziBUYUfyyfvu1lCBPMI67DUIkcHdJlLTD
0NPdd5qYpJTTuXxGGIU+nGc2NkQmVz6JzPuSqhTGiNh+zIK1RerOfu6QonjC9TW4Z9GCqVo3yfAP
kaAhcaXWvyKqsa7e5BgZyJL+rumMlJ56m9ecoO4Ali8dgLBX1dS1kZmBDF0T2QbSbzFVmE6wwHRx
glBzt7Y7dHcQ8IevRwvkB6pB3zOsUH5nYDE3oQjl6e6pYdhiG38nDwDgUyKSrwwM75QZG/oExBxq
SGIgs6AXeETObEnnlN/3/cf1w8Npa57XhvDC7ffSPssb58DXyk+cOl9MX9n+DEe/cpW/JGRNpff/
5P0ieCDZwjufY7w+Zb4IyNjDbsZfhKPLrFWpu7IRMzwTBecEvHWyXKiTG6D0DWqR95strjdVoJgc
a10tJQeXcCBu8oWbVwKWGCHVkrmd4RblrqyoFsdhNC+EAOlp48+ZovtebI+31UQCHZkqRitWdXd0
sAQrBdqoLJ6wNvgxbOMTQyweve8tBUpifveF7LiOyTo0AXgFx0YqJcR97gg/RKSyBW5O4hLKXIr/
/KYs4gsW/9LEQxNdFGfbAOp43Rkd6gsqB/VP0Z30pC6Shpk6anLvBGsz9pVw5U0URumH4rCTF6d+
TWuCqK7PxGInL8fbvU+PC6XJ/vMnvg/5TL1RdT+HWqTfHrP/WQiKqUD3OZSZ7kNZuT4jEzEZqLjZ
qLbI8tmabbNMyaM5dYVMNr8aCrWwg2bdgYXAu87eCN1HfcgIk4b41oTdXE/HKHZMcNoXya94p0cI
Q/wH42ljIzAekxoUEYnfo9e+WAcrlFoRydpWmxwJtj6nhYX5gjX2fOPDkOnzXJf6Yv8MkB09Mdfb
wApIfvKiWgEikAD5QBqUbq7TsFkKdMjSdb1PWr5CX5UO0kp5ZLKwRizAfvXlAikmzaIWCgC9fxmA
/lWnNo4Ey1GoxzjObs5I1Z5WJAM5LXWUwjPa5dNUlGDLdUaXeKlE28K0TX/W9WGF8kr+eKRo/DTw
vOEZwF2bSU+2t8oLzrWKnVgga2O2I8sr0bN/lzepIlzgnqbL3hZJcVtw0s7Is3p4bEVwcroHFM/+
X14eAu0jLLxfOVNJTSNMs7CSJ9uue59E18FgLMMXujSaJFXvbr1cNWlc2sffsX5H4ct/Ms0Rkj4j
qv8NHCaAJSnqq5i9wS7vzUPcxB8FuRcBhucXvXcm6Djbv+gYWc3ijjB4f1Dv9GZCX6lYX8MBF/Rm
5mJ0zk6xgRArHUkrx+oGqN++RoQVLd0Rzx7ZBj7TO8j0tmtwvpUcfKSFMQi5ut6MUrsxHyqLZQxH
v0afKdCn1Jj/aPiNLCtrANqZh7iUS87Eatgdtnx3W12T0OY2+1YavtRlprZVsmQpBdfRslABZqGH
9YH3qQa4X/VFXHIXTqdQEw6INw9xOuL3hZ1huxnjojg0ljKZK7Z+4ZKTTShNrM2/cpFZtQ619CU7
o60nHrQwa/mLKHklly3bRCVRQkTCTjMEm8QbZ14f1+/6Kx82sSSiCnipuzlveuGdw+IdpLbB0yy6
2TDrk8M80Tl1B7GpQEu5+EBYAyNn/6ULNEkimj40Jy/jYvjZHQmF6U4SqBAIpj9OaidQjiz0kKDV
V63LPI2zCZJisH6EuGdd7no3rrSMV19Iaxr+uk0V15UqH7wn2PS122LJutpc0va1v0MKbDxHKMve
+rzOw5oSvdYeGWEAW5ExI4SUsGcxPOhgIj11WXemkR/Nkvs0DmvHQAgJFO114liNBp5uyIPoeoUh
3z13+PHuT7exrShGfcH9p64Y1VP7a+XP3pJRbCM/K/nkMr795DlkpQ295kKOAtzw0wKD6IhDR8Yz
T367fUe1WRfWm8Cov37gy9I1y1l9uFgdQ/SfKbHOdL6awedM7y6fqDGIYY8Un1lKrfGN5I4eXIkq
egVTS/KDyFHRh9TugRB/9cDUR2EEjnigImXCY/z8bC9fboGAKBlP5b+nArEtiUX19t5zG5UpyhUu
wIVrX23q7WVtIBisFjUb0AZjXuhIifz+xhVhgpooKGsjhZdCK0Irplo0DUjQZry/wI76VxBJo5sU
q2SdHBr7ZgUDRfT3+tRyBKxxjMX2EbNUtI7MQUOMKvDcMJQ+8eEKT1qXlucCvwsvgnQooffZS/R3
XBXUgFDTuZbuT2bxACqBku8V5qVR8itRsrjGu+WjnWWVqfgyyKgqaT2PjEAIVTaOoDi4mkw3UaZY
EaA+qfem83bKfZB606lOzcDVMRsYZnNVXHxBMwyyPNMRAtoCA7/zmD+upzdpsmhCpEmaskAZdTec
DxGBFmyZaR60SRcYcLMoWLDIcxYWyavP6FE1kyP1AvZN07l3Nilx3vDZiTo8tT5SBCYvQMA+wrLA
tvR5RAgrU1oepxpaS8Q1/HGmC4sASXXVzhvft6eXboyLeJ3+MqeAHpOLmvmGPUbHxSTC4SVdmjLD
DYrFslpNnwlKekhpFbB2LB451U+OpMtOkZx/YstEK+FXDNrr3zbEhxVvXIBEE9ewFBl+At/T4f8B
CuRt7CeIgdXfjHGbBsg0g/t9+UUsqMGHVO5Dkt9NRHt81uhLLIPFSfwcKJR8HdvwdKEDMDF4BTlj
33WwevbmKAr/1nK9f5flGwe6wni8oScZYDfuilR13wS2UNTYtobU38h2Cl32WXcyZ0kjdZfD/69X
MtkkegoP/zTQBvDQQeNb9ar9uCJONcSlBJggXcJFXOxjlA6mYeoWXacGBhDdB5fFbxneM4QZwe47
cNpiNWwolGRRwijLLrCyoNeZmNpUUihO71nLxTXjgEDRk+wPexGBKuFtKmWGNrH6lTz27UXrcdS6
bnyq4/crM3UiH0AmsRaAJS0/1Rqzsa/0ChCanA7F0c/CBeLoLz//ntQFcmj0Gd9nZCEJwQWQt11s
cVnjiypggSt7IAxkRJvglbVwX4LS4qLvXUB6QhtMYKwAW03+ohyZONVIModC6RZFRZ9IDpS3s35h
+HgzEd67qjNTiiH+KlvqURZRRfJsJtU0s57bOpamzJF+pILezDzh67wa0/ij15GHCKJdSiJnwIrW
rtMTs8E0/B7x5CjH6dqOO12CTgh/q36/OgsODkH4wXovLAXn+hBy8CM+TqZz+Mg6jkd+xWFEJqg4
xMT7U0qaDWwny9rDHkKGuY/kastbnTGWGPVo6to07DpMwq+aSNfO2rZZ2mwVNFzRYoaAAz+RCjcY
9dzlWuWCSOt1tCjuBkhQ0iZrgL0Yy5dOtbMF6OMNKykuBzBKDCeDrvT4J3b88oK7JZ92Bu9HblMl
2uuv+VHrT7zsm3yrPEbyo8M4SNg15cPLXybOd4eFKzGf27FKtUxxZbch4jjQuBokto0VxfgTjoy+
QrBog3/h1+mZ0wGUMsd9xMVTOwlg1beBxZJ+JR4Q/Ghw5xT8THbuiMFC9xJMMS3GrJtwge+67+J2
NyioD3TZd4pt33KvixATmk/4lVJOp8IdmDMiKIYK0hodZva/Hiqspi/JvKvITTxYWEPlNtLdWWKl
HaiXpNvLxar9qrlB9e8q0NvgklZ76Wr4S7zJRutgSDXMQnWIqh43M7sXdqWApsIPWf6VJGumBXDh
l7kFczGbTxcmWwVDwj9v5yzED696J+kJ7USBqQkJSAkv62vLNL8WK641kwKYpiEk4efyQIQTAqo7
owVGAW58J+w59TIbffSLWrtr9VQeQFElzIHjDXZVi1LEbkjxR7mxP+w4dMzgoxZ/xsxV26CTZ4MV
9Kfk0BVH7rhhq3+MjDj7FdFzl+R7c8PFTZP2X2gggteBy0SATL1GX/C2gbb1NwD6NdvW+BR0Bzi3
cUBy4mgBNR1AiYvVrU5CQiTRRugN7j0b6o1OOgKS+6m2xxvOh+CBTpfFxbvu1cMnGHJ0bA2XbwhL
X4GySX0yO2cqAUwJTcmGG3STNIToBjZOmISE5uPrXs52E/LOUwYxEQUmHuwHeqIzBUiualkZ4SWF
KbZAH7Bng+HDgkMjtjEjADvT+dNx+A6MQtLAR9EkviccmdpK5c8VBhYcT+FfblLTT8u1dV7QIaGs
5XE8+KsK9Q98O7oUM/khHhTvUiSx3WEuMgXslOqc7WbMAdhch+CsZDDSJbNlYQI3XoIJpr0qys0S
nSz0HLZZtvyi8Xx/rH+6g9qYT80QijzN5XQOLsFHROLZONpJlVUbLOaEY6eCPQbRwhXNclfOauob
lxmfD7/495s2ySdbCq6eRwfAslEHfcJvMzZ2KacKhtYWtXxfMQ3Pf48tLIcIIe0Vtxs7NDayY4xj
+cScqLHYFXchpYOvGoqGVnUs0zPDZ50Ys4i2mPy/UewUocwQMofbmeRiGWgeFWBdNABTPCiqcwNo
v5tZNVOdGUK1U/pUICQyKPk6vtJzoqCkUVIAvdbSFMzqN+cjLXwlDCaB/qFSOnW+1bOVqCLaOJR3
NY7javgNjB7FjJboD07+0Ww3zTaZ3udKuJE4ryW+2n4vlH3AnYmRAmrO+AGM4HyCVhnJ7AJlymee
Kou6YjpS51BCaooxHbAJQuag5vs+nt36DmJZDhOtqbgtUiEVbZg78UnzSHfMEr41zL8Ap4OwZKs8
pwvDibACMvmbGBtmZhaoW4n/gkhf6xR3/yDsPYlvysCUxTD7nZ0Kj7Dk7R3ks3pZUlBFs3CNEfiF
YgyGPKYwfIKhBsMtGL7P2+UPTHLWRFNTgQ2HDkTdUBOI+eNN1w5EdijNcYJlP8vFk3I/jD6XrJpo
gyO/piuI34Y23UclPP2HvzBXDHIBKkY3/N1aNn6uy8ak4RqP5hopHBgyhkijco4q+8u2cHV1UHjS
oStFgOglhI69MRLsnBCsRDTxuD82K2joYyKdXYg2XDhh7B2kY+el9dELmT3uyqd/qzIaJdZlSUg6
pF9pZWM+sLVTuCcIkr2mLdivOqAkukFPbuOJD38KxhWfX97rZdB/vLe4K32ebgkdOuizLnOtMK19
TQ1hkUJw3Sy61nV7TM/ef+6Mh5fHhpQG9jn8v4mxpjQm437G8NsBWlx6Yz8Fsc/8CgzelK30NKew
RjzATo3gplryU2+ANmIaelRWSxesEExW+CNA8c6mSBW2co49LeQ+KFZ+I37EKmSViZlY1412Xbpn
l6WDgtjv8abpaVl2gLHkwF+obrrTehSkkU9Cf0VoS6Cy8iWyRnUS35YXRYCDcVhaxMPufkhZeuDK
At7EwdWPJWWDTUg2oE9LKrG3MaF+98ByQgGHglMfnAliIY6riv2LJkULLY+vXbrM7pIQhxt6MTmo
PFjYU+InZNK8Rw6vBl1a0MREKCzf30Od2bAS3dpc5VrbOZAmxc8TR52vWzzSDGzLYfv8JzbIW8LC
5n42ocynb6mUj0d/3jAAa0D3vgUvvJChcWWPbMoVZRxTsmlQRd0RWpmCy4PTGg5j6zCR9HW4o9Aw
N8uG2kNeNI+Hk7C8gP68QaqgJ9TDC3+eHKy5fU2QOk+9TE79K4f5+pf9+RbkxfVmqCxBRrLDeLZn
VFIIuaKbgQqoMOwyDu8VqgDEP+sUFyWGgtg97h3Ypgz/jXLqlDnKS+fKEsd4r0bC6AzVnRqlP8Kt
kH/qbGPcql1SBQs6WUjZG9faHithJ9jc1HGfGOOOthmAsBVytGOfHU3OFZb9nIqeDJtAXCzzSov7
zSSbPrmm8oh9SG9L/3YHu9j+5y1sgD+w+u+LhT2VfGsCHCasCsJGIXJ58J8zoIyZZ0OdY2eFdcAv
vhEvRrkYYFjA8IXk5YBYfV5KJnqBNUfTlnmCZ96YV/CKyHLyoYDSN/RWvK8XFq8fVHSqKG0uSsEQ
nM3e9fvZJ1wYDlRvNgNTL69uEOsGnJAQqWirwPS8SAOrVCm7C48T3DD6uSngUUt0fuPTQOj2Egru
CsJeaeTWSjOW2i/c55axi3E58hGwSNKn59umZVZ654gq6WPN3QNY3KwOWcg7nAd0X5J1hF+D4/j5
fBLHYTTCsPc5PcmEoSM9NZl3rXAUOSMH/CNKnIPSgSENxcJhpmfKujZVHgOH8br615kV1qgWklqT
5i/QiM+vUcflADxr0QGIk/H11BBMsF6OgLU66QG2CPTZP9Vh+Xu/f/CP7Ld4fuK53BsY87gJt5wi
Hyn7yjyFsjHiQAFlb3ZMrK/xh9m54Vg2nO2bf7zBjo2tWkxml6dgvU0Ax9neCUj/0aAupzhut7mq
rW3zOfaevHFA8rjmz+UiwPCet/rVULz+ka067rZIsal6v/+D7BaP5aheXIidC096LFkR44o3nMAD
hq7hmGYYwlRyEjju78jyM+thSR+Ap3azYZvSVhrj/3ggPJCkmHzavaxpFbdqXJ1Ttf6Jb83uwHR1
yEBeMWXRHARQyEYbh2LqYhnDdYiqqLv9cFnqfJVzJ0RF9Et/p24EiSIrOgjH9biiaUHLMqpu3IFr
iEENlqo7EJ7kYpUmsghUr/f8J45GaVTRp08YekjNrw576yAYac38Oow1pUfDxB0DG+5XvM3F8efb
504hSNioOG4YXFb0eNdPFNNX1zYcBFXJvnk6dZUhUBkTn9GvJkNrhGzmfHE7IgGwj1Lr38YNHJHt
OO8IDeCO9EEr+umz9TTuPvB+MmjOJLKDTvVa/Y8QIdOkY+DFsRMvri1uuU/8zXghsK0IhfOlIyp+
A2F9mJdQXaoAy2EF+/ENYUw+BV05pvKICXbmzn2OQe/6EqsKnLyrwnHlgadtueRKmVy3sa1EJ0qy
p4vrZz0H73Pi1TryaDD2MGWZzAEI94qzCalmmqjLwxI9x7Nm/7HFLV6XJ5SW13Lmj8Ja8q6qGAD4
VIKvpL0nprgPORK454q8F5M2ze+eJKfSCcjln8P7etNzQ4lweLWA3z8B7e5Atak1H9jq1d7gkv+A
q9AoJoY0POuz0avk/uUtW7xt2Ql8PvSwy36OQOsbpe8coCzaVxswrogCKxuAWcFs0/1hMuQx0T/J
lz4PzGxKXr3t3UFo9lxnhPnG9uESMyS6ddmmK9Z/HGLqk/1oRvrXJ5JbRCTQkhEtUSQUPrf5X0Qg
PjlLx5l3pQO0YpWKSBkJ2e4dvqOKTDABce72pSb8VpC/ruwSlGZSazM++y/Ob09vbLmXktMhx8uh
gFBqWsd3o9XU1ucrm/h0FRStBfaCoEdMdUAdXy+p0ZhcAytqO99UgzMDwNbF4mVP+q/51P0Ly2mo
62kZoL3jEMhBNxzdLWbtQGxvcfuLV0vzvB2FjbBbICP22CXd6k0/jPHeXMtKhIbppeAsoNmFsrgv
QzEhXyNHcY16QA3nelfFH3DDvV8yW+GaMLSGmaIrxilUyiPAzS28X4IvLZaDlM2JuTeZSRp343u7
guyZXdiHCNaz4zswKkMM8Hk9NygVxAMuQAUuoN6S6wbTGQ6AD0k5b2EROfx/Z4fOTarMhTT5db3R
fTRF2jwinN3cZGeH/IhS+ZeK9j76gEBA2KqoUYgLriNdMQakAsNrLKtEAhc+ulBgufTLsxsS0SKq
m7szorlkdKZHIXHQAt2PLovve/4qJtA05ymMwQRJNAloNOBUi0mBuF6WEJkWaMnerX31j/XVrihx
q4P91MTPEVk4NS0TyhH5y7DOTP4iFmTQcjj0ngsLT//If01SKYESZGLYOlUmIj5eRMOf4naT4pVW
bwKEclkDpV1N2K+ksnN0cyLWZ9gIFYObTej0u9r7XfcPTbXTg/tjpmIXvtO5w1LOL7sR+zGZYDPl
lknrEOmChoky1qlU/KW88c+XX15gU9sPQpHnRXO/OZf2oDggEOf6rkjKX5UlrffYD9G+3aPHwdoa
K192ykUQyeNKqk5MHxnxAG/WqD8GS4JISSdpqRnyksJ7cXSTSdmmkAFub/b87pGe9dpQQVKZbQUS
xteYMy3XLUQYe6SD0Vp9IHUn/fv/iqoltjt9EE/W72v9zZmP7AM2rHjcItHZ12Ba/b2PTMlnFr5V
OWvDYV8HWuG455sCDLbQIaotiKURwU5avGecrwzgSicHgvZSi5sBegrbqpOrFXNhDedOSMw0EKAc
gUfKPRxeBKtr9vYud754gP/F8kp8afehbCFm5Q94IIR1YIjTrwX17ck0Pg3dKjnw6GRRqwrlLoAh
//4iHBdaYME3yTaEbNx+ua6aTlTWpXvK3cgyXt2dexq6+5TP/G2Qn04obGGp5G561yUnge8NOa4k
l7pzIcTheygNBrZ1H/kH5dzREQD8EIX8xvXmzUjL0nCg5BKqNPgnwe2GJQpx9tORxt1SAcV1V2Us
mI579xOzXRBNQqcWVLMsBRPHAJqV00W4HvICHoRYHNDUljOrig9a9PWYZ/LfLqxj5c78c8Ie7y7Z
dNYKEqNvqK8vliJBCnSu+f/ivkVU/Z9oZr/rNA13e11gaOg3pOLPrcp6JLgmC6J09/VVTqoJxCq4
7z+6iZWo+p2bFwMv7ndYZeOOlx11rRRyislOS9RYEn0PFSwKivYMak/cgqPzSEbVB7UTsYuRhGHM
PRp9WZvN+4vZRRYirtCKW0VQ2WkUJGZKkksuFfCNjjdc3x9Kbf0DXXEDAqBPUWQ9pl0EnaSmPAQ0
j8z4ayUQbXo9Jaas6+D4rUBJobx/NH5iK24k21IrhODWcyVjYdjI65lZOnAKWDisPlgtnN1N7x15
jGI5hEgg4WFCt3h1ProRHUJW+1mTGfpfA1Y4AqWoeb2E41xY4TGkFi6Eb7APps7PjcjHfjDdbXN8
9GJ5t9EQiX386SbT6gAECcpfp9jxqNKRzJByL+LF+AsyNi6IbFRq+vyjKMo6fzTclfaVDL45S2tH
ki2pZ1xfTK9c1vQtb7IM5u4P1atL97D6Oat9PlcO6msGCratuBDBe0i4cOQAxRITYMUbWpWtIhdh
wqutk5LXF43P2IAm7UIK7CELZKeYX8ehwmil8k8dslb9FeTR6oTIyZ8LsuYdI+376SkB+w+0kZrF
lb1FpaazS84od7+hzUA+sGMJhn8rJHB/IsBzV4Vav2d6WJbsW2RzfzHG/Ek1OPv5sPV8kvE9Ee5H
yRdBs3pmMnVvdchpcgZIvqBafuWyJLJLPsYHqNnK1vMCq+LLwUDfD8futrPSyUxdq0KnyyCJsBq3
W5LvQRdcnbvyOcF0rr3rYao7xv4QYfnaUlboiz1VoTKZYsk4iU0sS5U2fvtF9ZbOxr/mvxciQ0uu
kvs90/plvVYWgFFfpEVkIT7zw1D4dhvuzjRaybwnl+N2MyCd4UuNR2RpeOH3hcHFOu+jFwB52m0F
9qj/OefJg04xsHeJZkM/MfNoqtCFQv4Pg5k2y1L0vN4cldbCyeLaW62wkiFbXO3YFXplhY6e+DAS
Q63HUynuyzyD8tSYbEWLasg3W6f5AxNmp8Y/FWn8uxp6q291EHmewJ3u4uXJ542eB03pVuuSHo3A
QWRkMv41vaKacgX2hpqFmhytRv8E7a0UDKEiRVMic+LG7uMbEidveZeKggosnU+NYyK3PJpiBMSa
eaMWGNhtZs09x7QuFneWU6KoH7mnd9Rf0c9x0Gl2tRC/RfnVOZPiA7G7ijXiXYgzubJbk/XvBqlH
Ux+6hs8u0pMn+UyjJfh8Nq6GELZdQwiSKXA7EUhc4WAoB8IHiXg76gQwmpdE2nQeamLy3dE+sxE3
JQDMSlP2Vkx4z/T0AE5B/S7Z5hjSV9sJvT0I/WlEzTMC9Z3Bya4eb87tDEQLD+wgDKq/w33BUytb
3uwvy9JckY3nHS+BPSvoz8cS+OgW4rHsxBWUfJ7uwS4jbRj2C+fIBUs59XAFxTISh2gowy11rUUt
U471dWthIkqy00/m9KwqBZ04HXYD/u94mY2b5zGrIclTSsvdJfmzhR8venKU8v02sJDDtkMhEHPO
t9jrjKfyr5eAtadSdIFGFTAO2FHXlCLRVxI/06t9cKAchOWYzBp6rsAjOYyH/OvHIIVGdnMvlH7M
WbC8DJL7mhji0sCv/w0yZGTNWcePZxp7prJl7BLVyw0PfqBsnwYkIqLWuPN8y+3xaCBZBKJrjirb
62th1qpCQABDs2nHgttbbiRQlRmATyUeYyCQAmjem8FvlhgKxl3JOev0sCOcixg74HYftvaMQ6WR
UIWTCw0M6a+2icSOMtuNN8p7KEpkVn9YHcx5q+bl94DrLzSYaMayqXvPCKTEsDkopsmhzHklCA4F
zSLVU1BrE+UiUBzmnO3uuM8Z6PcgJqviGclpdm+EpKv2lAXdVybNp4M3AaJWQAOlHZjzaHNSqWAN
5dZtX/7h1HnqfBDzSD+ohHEpKIA1WWa+WBgd+zAOPzIvfx2p5324uGMZDMheYLX3VAkjOEtKoaiC
gHcabKTFvObKhd33oDBG1yeUjdQYAkZca0vTl95fX6tXqT7FTKR9nZDxVq1IPa7QGtJRYsiqi9FL
P75TQA4+6csqL4imem9BeMFgk7m7i2noVVxVITrO5VPRBbzm7TeKaEyx7fRTRYVD+16PY8K/CkJy
woHFuYqW67AB6uFHyvCScXK6ID8Gwz3+f+hJChmsp3knTRLvfzr24IeRGXyiMaYBqwoivl8UYTi/
F7euJ33UdAb7Df1JCaTf4d7v/NwKpQmzVZ6AW1lzNjZmZ9T/w7KW6wbYKdimvwvTVjAlOAaSOS/T
52v8wFA2oSG6oOhzke67hgeBh5GL7f+weSxrSgz8/dcExxfNtNZ8EbobjU242XbiZmSwKTP6q4vM
1I9b+WNcj8rJ5JqOxgrf8otoULfXy/0lael6GK7n2TAfPTdyoQxlb+59rnsVcbAQdMiN00p2R+MI
UhZM1mdWhAjbPKEawB+KG3YFd0LK8Zy2fHpmiOfygSjQBQFtdYSDe8R5Gc8doHgPvhxd8Zl1WGuU
lRMOLbCXksYSrULxzeXyauDuO7+tqQITxdtTx+bjPrV1QTKbzFzb9Ko2e7emK/FDcWszCSP/iSrn
Mc1BSRtpO4+KW3IWfC98cpeOrvcHa+NrzfmsbMMTuViVzvu0Rc+UeZjbBLqQ7G1iDXp99udcjWZE
Bk/opH1eK5gGjItwDN5fX15Xezp7eVmvEItXof+7MlkagYRitiACHpqt34ahvL/flrVWpfh7rwz4
R0YTaqcnCnHsJqLQgWXRzPpny1403hD3HqfPpL4r7qIwUp0EYM6bYGPhSNIEAstO+1DeNaRd6ggt
O+/lcFacIBaMKHaUkPwanU02CKRBsatFcPY4JwzI/n8H8Sf30vA8Ee3DCjVCsRzuekuMtR8efTJF
CWoRP4xcHwsJlORONgJJY2/w6RVtGiSyMB5Xx/gR+I4K7lP+U5NMVKJO8Y0RDZ89bKEjKEpYoKLT
ZdNIY0gQ5wmbqPGmcEH6Rd9q9HnzsjBxdKROTtgBmL/dfzUp0uO5P9dzNuoa8jXPH0isE2QXeQ+t
EVjmkDJIj0q2zSx2+7Oa2sFoy1V+FM42PtZ+kN83c41afIOLbN3QWV75oD4suJwwqJBN4hWFHilA
h74o5rPY1PETnNCEjnEVzO5TJwVAQkSDDVZkEjUjoPRfhWaJ/nWky9WbfvwQn4JXssKtwyIJIjek
KC/GKyyNTo5LWHJnWQNU8MLiJoMqjfxQA0BXh/4JmlEvLdtMYa/MCYettfuFPGzS47OwuTaQJ9Km
V0vkpLJgJRk8JAWFUQj0TLuU+Q2WySg8nAbOlES05mvCH23BGWAnWy0kl8tXW5rLnKzoVJtDR0Ww
F/rNtyXlNuB86SLAHr+Wl4a+9gAIfMLJAqYzhBrxRYoqO0WAmUTqi2t375Kh46z9Rq2nAgAG2KxK
3pzDa5Td0aCucOCPwhW87JRxBbRn0jufxUphzRn9envubiqsewgiD2I/g+lAaHEs4OTF5PHUzPoI
q4CIzK/23Yyd98wlkgwpCIEyRThIerFhM1x/cgqC629cVQ/bCdKwCXCzvP6Rpy5H0jWLYI/Ti4xu
ivxgd24R/uBQb/n7JEcD9rCgGAqu1tMBTusT87Y7nxnOhzdLu3yhGQVEJTfkGpownVCscBMRiLvf
yWkPPf7nFymi30eMw+QmXk3i5scKHmqsxo+3Cg9vSB2HcCcHu7FoTwrq7eWGjB12x718xQcciFaT
7pvIfTYiuE/DciZsg/7iBAQ8S2v1J3APcTtmm4VnSbMOUnPtRBwG+kBxgGxBGzdBh62wgCc0wcAq
7gVkgXiCQh++4hn3y2RnPeHMgyOmrifV7LIYPs+raFnJM//EmiyWzx2EMeGjVuxEiNioepdP4rhc
je/UZ2xcPuwR9IyxuNo41nxXrV+r3n2uAhX72MSQMoFXt8fLE54WT+Fzus11WybsboCc26g0AkS+
O5Oqjb8DszcYiH0UWgHDB3VzQIwPf0M9rpWb+V/7Zx66rdJcxvrvCyw+Orts+pS+fHhV6fIAJCZL
Ssx2rccDt6H3nUALUEhdI3GmkQB5KRcLufouwzguG+D4WgMryTBlLoXOTnSeNAAbdgTMkLL+/R2c
jqb7/5QKiL+plu2wn0Wnn8qIqMd/Xi8ZImclkSxEMnl1i3fiQ7I+MQF17JFnqTol7uJolz2wkcO6
1+/NEIzht7xIh3VZfSvp9MubUnpmF5fUn3/oCWVIxScRUTwzTe3laym5KURy2AzOu5oHfW9UwoI3
Rtee2qOGPOkEBY+0hZta9Bp6ARAU6vz3cEsJ8p+O00lly4B6JCxNIPL6wXOikblXl8EY/A9fo2g0
K9MgrVHaUFe+FzTEE3+vOVMeBbxYU/NS+cWhm6Gc8of6UTDbLZHd6quKcSIXKx0GGzVwEtNbq+4H
vYTJlQW/gAWw7nDSKqOEvVBJpcCs/e64ehZ9ir+kwDe8lg3knXBnWCqbNKQDJFeKa/rlz6dv7nNN
IonDg6K9RXLL+dI48QsObtqfMhBi8zcAXf3fPbps2+LGfSRUWENcr+XDQO+CSGlobpHxYVfdvIDk
BdxUz8etLlrbFlZgiJULLAc5OzSV8r0VUCQT5x7L14QtoZuCTbhmSPteSjVLItG1QMZtWt4I8F5o
lqpi/2i6ctkMmHEzTOfnYZaMxLV5v7F/FWd1q5qFqEJE9SVJbzFS7J82oPKUHbQSRznVodoY+4zL
qYF1uMxrs1bIZPrUHTP+LAhiBY2zbe7YzSDbxVS+hiIanb8Mn7kZiEsVDGKuBhG2aZPLLJfDAk3c
PSwNdxqecF2HZFGxvY45oKTX4Qzj68r13GBvAp45zfUg7Olaqux508SVzCphdejmQ6bhZWF6VATX
D4p42ifIilKG65a173gucVSp5cNLazcIsnEbgx6zsvPWngb/yfmnVJJPfkYhB+oxEHJ6vgypOrr0
hJp9lHa8gngGxpMfv9GkmYFGxn7OEhTglWjKMr0DsBF88uMALSsB7q3xl+rtSvR60mh+OLUTU50f
kk1U24D1rexaABB0gxdFTMx+qgPuF1lNBcZiagXXpfr5h7UNHj+jfoFOrBEIvZywumRTWf6udCX0
9GLEVPdmQ8rsOwsHtIh7zkPzai21t/KQBaijF9P+uTkP+l92jlvXyLY46AGPUIN8cuRtQdDIWwXb
MeNzWfKJoyftdxr9xFcsZNoW+e8+7wU09Ek3DAvgdyjRfh4Wj1SJJvO298QsSsLfD+QLI7YsY82q
n7TViadG4ejxndZ1JeUvhQP3f8S5n7ZzdvOnUwaH8U2fXVAPcsOUgzygztwO9tO72SFZcRI9qjPB
ggjG4C3JQHhe2Ptb2MDp9JbDskWqKyl6KHUK1q5Ssh/4KB4qAcCfA2vGLQGlSUx0ofp+lLy2wpFI
kVpqP5jjnyJJ2jzFtZiwruj0O+UO7+gdQOQCwXou+G469dCWY2O1EDS+CRjSgR2G5dkuWgNC5xqM
rUFHPzgoYb34M/yMHUwJMyARKI8X5pZMa0cgbg0O9UOt27YUtJGf77o58aPS9/C/yq+XESzctvje
AG407GdPok5lCW1vOVfpOA1lNFrxQelfv2eAWOrdfCkFhaKF0JxuhQWw2OFsx/3372+woKx82Y6M
4/kTN9qtZJ5jqrdrSnjs/VxnK9M9MTWXkYS9hRzWeZ5LDFI1ei+l2gKl3BnKwrLisOayd/E/DtGk
r+rn6MtKjcz2nenYwBtGpromAbFwHILA0LQw9Bhe+namToASvcYlEFI2rYlfxLOsKCYNUhdlzO+R
bmRjujshV1OT9DsdYODMjyDMtpWNj1F9e41ullrF7Sjf/AzhU845mAF4utqNVwKbQk7UkXkOoJNd
xulDL6XKfxRFdgXe+7p/dRoHrCtg1kqhUsyCNjBTv6ylkfHR1/w3dOB/5KC6QIEe2ykwe4+MxQyF
Fx6JmzoYKW2fIDPSt0DGTyiF/Z9aGWVdt6B47BUyK/7qj8faYsWjZgqL2Fq5NyDdTyFb7qA3dJSK
RF7VI7qaQZ1xnrptWD5d5rpxk+tTe7yo0AVf/wfdpHsCTRi7Cl+dxAUTyLgOuGzdv0vAczFceqAb
YRFyjwik9s2RoIwSpUs52lYS/L2j6zWrk60OlZvhioZnhhCNgC2nX4CPxR0CweUoRHSPDCNO9A2K
AYL+e/kx/Tn366IxAgVw1X3Y2FCW10tH2L/f0Hm9SuLmV8lLN8L5R7mrOAVGcyTJuZ8biAw/AL1y
KGW84kLyjI8tvVoGWPIE17FWnS6+OvxldwWsQA5QM5inR36kOCAbloNN3dPmQ6Q48dO7x8Mx18pP
O4xNSJWmEy9Bz2DTBKd6usRzQM2zgizt4tBIzToxi6q9AnqbQ5SiXKLjgViG3PbYwIfAdrxOIugT
QnGKaMTWD5Dg3rETfHLlMXsMw7myub/z18Q+sh6oShpgDjt26ORDGwOImfK3VMlDr61cirkfd93e
Ha52g5DfYoX5m2slaTVSrTVPMAf0yoeRupFe5OdZ+y1s/+54oEv+d2mvUM03JTDCldzBUfj4swk3
DiEJ9ge84fItc1WgZzRLXkYrE288ZIjwflxkYGwigYKr7wBq50I8OquXcuB8Pus+ksUOCTDAuROu
1V4j/ARnH5ERIkBas8mEIXhSWGDPpfpBa/HeRaD2wIeSTZpFjyZGYRseIQFtYlDPHans4ge7x+9E
M9FFSvNeJv+2k/rTBMIvLMHo9xsI7mDToWPpjMmSzHibEmks5noLHEPB5IN/OSRHU+acb+GnrxmI
VIDRCrrBpCAPnpJaZavQgwN7SmAKfvBBGqiM02NqnSJ8e7fHVWnqlgCp4KP4XrIGZVXhK9m7UuTw
JqTyZZBMWjKoAPnhraIj192ZAZEz6If8ntYb1I9xb9hFSie3mfu7XiC/jJml5TN35tEDNhOBoS8D
fDaylm2y9CrJFhSPlgyQFgeUQ085MysEcB+Q0oWJFPB1ZPbmNM7Nze1NrfSJ4YfGfpWnS3zI5teJ
AghOI1642HbEupJsyLwZSIgvvoda57MACgp6F0dlPFEZ2Yi4pAU1iBOM+nRffDocNK8ItgBM/Ggw
DqpgXXLVW2wPTfTHWaVbZfLGczlmOunGTwW6WWkG2OoMaskXrh+ZVN2WBQchRHwhkfJ4v04XKwmJ
D/8bSEXu2iYJfe4y0x8jB2COqIs0pjYKlPX6k34DOcE5K4C/yioA834wY3kb1TvGr9krriEvzKHx
OPTCqo7dQwphZp8M1F5rjhFa11Za4+3Mdc6DMb/RJPJUibZ3Zh00viTXj+LJWaTGYKQ9f4s3v9nG
5lRlA/imPlGE6dQ5rZp526ZI7Bhveq1XQaVjK/WKYwJnYgZ6t7LWfC9RodhV2e8/GdE2bat0gEe5
RAssAtLSH52dr0KhyfuUZZruFOQ3ly8IfuHIiB2l4f9azDIzmRRmBFrEsjhJkw/uS2ppOdNj5n+T
tmjd9/SgtOxarbZzSk0Wb+8xgbtPnxfuoO7FhHFMfmdH4imnmbA5UJ80lYl6ZFgP6KEfo3p7mkcq
2/alBvpAN41WKHQrHXo943GMyoY/3EpVo3EoDLTHKBzyZMdwCjbC1YOEwpJ2UEP40qEqdLEy5nKD
9mv8kB29ndjPanCW1sCXRy4o5guT7zb6bETQEhym3z8o3IyBazIFwAnGRZ7bbKIfzyFt48CJ7rkm
y9+yZPwaEA6GRzZQQarx3iAPeojC0CJf8vj2LdggqUKy1rgDhN6Ux714XDaEP78B9UwZyQIU3WlE
t7xxf8RF9yqEgAD4st028hAdrcCFeNNC37zqdxUHIA1FwGI+kTPfgtYwUp1/JRPIItr3L4djC8h/
wnBg+xihcHQ+3XaBIlZ/dQV8zgg4rbjYXEXGyMrALsRx+wJmzZl/x6EwBX+GY1PcbScSMH/bh4s2
0Mfku77xblc8ik6pYWhIwkp76jqE1byjPAfmDPJs+eGwNyt4CC7hU9OnD2iycDFI5okRS96VW+kK
IfsddJ86OgC87zoyVh8Rx1uETg4u0flbYa83rc5/ZTC+smAClexTuR2RnfKjQ5tVEfisLzIKXSLF
5qXzfhnJJ5AMfBzhGVU3/NqscCtSu3BhYjrMr50H5/vJnJzx0BvqEKDfjRwlmV+UnQASoXzJTzBY
Q4B+sihen29RUkGMkjQ++VaqYvxeR4gYVVW2Z0ecrpGO2JF+6tblM9HKhXNkVjDnMjxpk7BrMVRM
A8jQsh8t7DzsBIBlNrFb4rVHZ3Gekp6S2WtRKdDt17ejmEBcqilzaYPAiuv9+EvRcKz1BZkhpYlX
/VlyEKS66vvqjLACmQfbAmTWslM5UV1kXIoDtZTpCol0sPNJ2FAT3z0WJzYZLWA8AJlIPlzv8oVf
53ULn/NzNPVJKzNEeGu8cyL/xJ2TbbaXXaHZHDL1mYjMzzvLJ36+FJCZ2KuVEhJcmwc3kB+fBX+e
pdwXrS47RbyEXu+K2jQy+9VycCIo5sPyzjkR2VP95fmKjebUVKWwhvw+6IXSu9aCJ8CelZNkiXJE
f+Iddq0//DWSdXsN9GS2yCdRfL8IGXXFt6uYJrVZJLveBnwT/IOdnPVFPR+5zAtrko+NOo6kJ0/+
ZS+XB2T5Sg4wbxh/BQV5MDvH3egmlrjB74j1Pooly3CQsrtX4eCfJbExAGl/fXcCW5Mhx1kWY6NV
1yj3Bk1hrfZTUcisBjlieamjOvlX8uL+fu3hpUTnL1vevQYgc2BQwgzakn6BlvRiSY8I+/N0yf2C
ErcjTXeBdhWhveMuqRo/mZy2LK/VjUXJ5mZYJ1zOETpo6s4pGU52+IP3a09+LH/G2f3cPbqzHTbr
WQk9bZgPfpm7BYWLqC9HeZv53x/rNALj8MPCgZWc5Lsz8In5kbjGLvYHbkvUSigBn9qdOMXsIOEw
wUWjGo1+b101+8es/WdMPmPHsAfu4qFkbCGxrNHmDwBmfa9szFiKKNTvZ3B0Ap0xRRBXEfeye8cT
4+U7rxsefF5Bxpz8gA74AUs0uPym4u4YxT4sdfBdaxLbFJs8wydc7Rj/llbs5BAXsGn0Xh/gOr26
puD5DNMUs+0bug86eHEPZClwO69617tDrQF05OHpilAlGHiXh7gRxLhwBGzyWXxake1isDG/sRTD
hDaBMBGhWtHBzznM0uVJSW8BpoqoVtjANMpZJ4nuE0aOf5gCcfnzM3LlQ9Ap1USOvWW2Z3a5qhNi
jJ6k+RCz61BjUEN1CeeS/8UG7ZvUjT6Xb4G4iP4HaBF9K/hn+5tL9GEpPn7uoDWZElaawZ2gJpTd
M3UjxTYH8CxGUXpQKAagFoknIWa8Z8UJERW9/Lkp0wsOFEgYpAhazghYZszbeF//gj8WxUTer0z8
zjFcYwl6jIGw6L9JcDZkQQOlWYeVmNSk74Ht+9qSpZu1UyfMXl+RIThyIM0/LhV2AMlo/Ur0yqX8
YIjUvzP2I0FcTFuxoEsYTobGkBIxisef2MTorxaL45ISiTa8NY6HuNOEj3G9VGYdjRIt2NfiB4lC
no+aA3iYC0Mb5OnYMPvVrDJ+pKKFncp2hKnlfR8ywljKcd3QdXvVCjgkiRKow2Ngq6awAZwhb0g4
vw5EeEWCgblzHyCd09zpMvINa/x+d9BOlxetK5yLYpvotWEW8VmMqRkzg4qUguUYqpO7McFcT+Gv
UYd1r/zJuOhb1Kk3S7y/6q15pkD+eysH+Ljrs4+s7TFsjAAUVJEw/yg1jeR9p3Pmf4iwyyRmVN2h
y54p5wvG08pT3rG6ETxFoAX6VPtJU4ioGXyRoYYqp99KyZweAq5MtZjmKoBBlZoQv8hlH31+xqmI
HrUNFSp5RWA1znrP/l25tSrJQbmq7/K60ex/AgpVo1UU5q19qDSqsBBhC32pPlu6DlI2OUEYDoqW
lw3YMZZ4hl3xCrySyA+LTJ35Q9HIHQIHflXFOgbLD1ztnpeBBIxSlEBnTypvMqLvyj/j4WNhFcCo
ScikXNuL0RLyFGzsUE6mDfegvppLllSUNjoTWm/G6H7tGPWBMgD9+8Ik2pFfpZfMrn37ElWMQCiM
gbfTlab9UmRPDZrgep2jJXWb/25szQAVfZYTjDxNOhf3vSwEraw3SvotQQGLTESlqs2xRFXtufNG
uI3btsCmlI8046exPS5oJ3SOfS239X78c2yzP7JFyLzUiJCrlqGUcoGBrDw9l9C6ymn/Pf+TGuwo
r3idYbhSKvDLi61M+faBbAiosRFmFH9Jp+bcZ16LyfwcVrP6nCCpMawOK/vlGTPW1cuS44dUCXwn
i5918QgJIX7eX1YD4ZlLZ7KY502s1h7Od61U60Wt7uygRD8SYfILj923PEjx4b/16ZMnyuAD4wf+
Q1dpwxA/enGDUw3vXY5y1NzC477UydJCPOVowkkObDWCFiLvyRQTf0wgN/u8pb3xYUA4ce3x/71H
ky815oc6OGU2DN/EjCwgPdLx4wGRn7DrNtjJ/9AHbb5FUiANI4qIEmpotc0UMMfn6PF4JI6t+4o+
z5qWDh4iMpeh0IjRGDI//uqYYD9pv39G2se1iwCJr9IXXVyAnepQ1TrDCHU2QUAb90UwX9KfEKMN
bmu7TcbxrSDLI8S8DLeL51jWUQyJXK6DoBDTn7uIf/6JttHuCMJlMKdkC0ojzbAblBnSqSF1q3jz
xu44ZN8pOCxF0GRp5N56MbEfGF7HhP12kCpI66n/Bb0r1uKX7HP/4ggekLXvkLmOKGpiGZOQ7vVV
NzB0TYCzPJrd3shh+lrqY2817rrf8gMX6sRvAgYV042vuDMAe3BGyO7GiQwFrOtkuwc0jwKcruM8
wn5EjixLMkAR7Avf/EQ4Adf7P4jGfOfa580aXvQU338aQpd4/Wb1HcUBpT7TspQxJBB6L+w/NYS4
32SqUb5mwoNRIBb8vyJl7WEHfpWhwk1ZWcB7YYx9EuqyvTBHMe7H6uGq3yQtLTfRhclQInb48mFa
5gGIfyOHqkUbdyu91bzuW3xRDiQCmpSK75CgWxLcrRT8wWZp/qyzXUaN2Wt16BJw6tiFdqEbESMQ
fHW/YqV1bBW4ygnVkJS4ySvFVph5jJGfOyEQ222JPmyu1POEr/Jm4TerFgOzWoU4nMXSKAuETqG0
H2lHzaQLXKw9SWMlAEYrCDg451IWOHEd4CrQukMr2+/EilWSHeGb/fHFFS0wFVMk6xpXYYdwJv37
zSdWqBjZDRlpze1tS869sjgcQsileMQewnd+uvttKeeDAbjTBfdsPF+iVqNEuphTrpK+onhZMIbq
pnzIV+6m9idr1rpEsXoAH9VbS+cRJGj7MR7d2L3KO+b+kSiJExHbhREAkptjlWU+fEHZSk/cQEPs
DpJrQk/YTBsLLJ7G1zNu9wyEXaLrUJM06J0Cxxj4TPYxJpQZxtLiBuiVKgIhBzJbgdmXi66KUIJw
M4kcd0Cjoz4t+swO7NApJYuCklcMqdyN1+EYvuYyPmml8n64/sqwozk9d2TK1iqJud1Fzw6RmlOo
j/SsnWKSYmM1PQKvgi9hOm5vgkPorKzSJeEPnNuOezh/7WNLXdswWIK7JB4EpQnNNGcJQ+MxbYkj
LHKezPdvZkpU44NOwYtBB/sjLdcxYuOpiW9NcwqDzb+XUkCEjiTK+bI0yKtducf1ao1PlDV5f/Rp
F79u0ZjfrUGbq+yyYNNLINCvFoLt7P6DuXmfCi7DYPVHI4UhfznH+D+wgw8SmM8JjfKfn2+xZC6s
3cD7rwMx7PJmFZryU3NrUnfqYO0G6CaaEXd8gdoID6+QHEPLn4VKMUM4AkEmPXhKRNIfFaSW4kKp
CcTdib18ln4UstaLPy2nZjfsLjJ+VyKvFUVRbf0Z2CXSFdt9W6S5meWMF3aE0I9D3XSqGFgQhAIr
MZxoaFHHjaaYApC8Khp6NX82pjI/YCZZVe3aP6636NXPtMFapYb5vcsQt2/TVFwP0aub42as6EAo
Ek7krC2WaGIgzawsoYdYyn+NMyaAW+V2Qn+1e+aRBqY/itzXXMahQvFqR3LrDIQkp7q/z6FLDS83
W7Zng6hiKKjZy0CEBpH+Xtrb8DpaIhMaLDaBXim0bIOXqVbyLCbCj/F2QVYQbwKyY2Rrr4VmOgCX
zx2np4B59Bn1mjxawfoGIumcgbeGRflCIiEz5dWu/JKu8LApD1+CkF1pPeGrZuHA7oy1y9Uvz7f8
Lz0KrjSyeGIPOmngB46L4KZD1BIZndKH3asmEaT8eC2u5BkmsY0ynt3BBLvFJl79Zc0QV4ZBfc9C
TwkalUKRVyqutsI+fLlJvvazjLE/u9hvdrR3O137NwpsNBvt5MefdppFRPAh8pGHUvNIUmDViQdC
BpywJEkvV623pqiX8Fy9yPLmcUAeM2Cv6K8I5eFjssWnmysW+vLOz5opmvHnybN1/IuhwqFAV3MJ
1YqXwJIlny9jfoLw0Gjpgh3WZNMmDJqZq5lCA75bgm3zeyzASEeD+n2K6cI7h9rP2LgQ73TKouCg
ESzFrp9KjviiF9xsxzONGnauTiQvVNb3rf4JlJqftQS8ynL5JlmcCBI+cW+OiRTG0zgcYsuROAEt
wsZkKdeNMM7tkCoMkmGhewBQw/dHx3nNgI5IEiqxYh2thItJvUweWbVGJNn7ImAMsO0UNvN5KAMN
n9FC9UE7J4EeNwnbc6qoI8cz+XQVPBKnzVxsWCXuviSNd0uvOCClALGTqH7HD1YwjvPn8zJkat4e
b1lEElCnFfwEvyaL4sdIL9QubEyh1a+5kWrbp14/BJNP4o/xhlRMiY6BR7Muuvv4KNm91E2gJ2/g
xPR8+e8Rwt0BIcuAoGVKQmY30p+BL6k5JFUwhd0XQNO8d+qfpP0FKJRMmHzaXzsyHfs82vrkXoQk
GoSc2Xf3P22R1tvuXBcHg5WC1ewcAX0xwAa399/bfk+/LQ/1gT27TiByD1lsIzy9y4IlIzpbdrx8
jam+Y5faBJXBaVMHwOpBXAQvyLlRcyWBKEh7K/HxbYlbFX09CWir/OMxOG5TAydVsOoOWLtucrxA
Be3ELe3rEdtjqn098MOi/KkX3DeSjCQ8KKUyCWgesQ8cAEcoc19Q09hB64Xj8KKg/VxnwjtLVNSp
83c3WqG0BIg3YReSSEpKi3bziFRoXo49c90h7WiodYZJiavFDHMpDxjCruV5GThksCMY4zDWdWfI
qgW4Vx92Mez2GNvIvNkBYFjekzPVtTND9zrALGFN+64FCoNdja3C67cWUgFx7Dib9AvEjhwqQ3Dm
xKOr2cM1dmLIbYs3ban6SjGRJRaUkNbVaEUpOzTzFi8OpSZJ1+CTT2cikBCSjM3CxnloeidezOOg
PCYSfrSg8gunN80tB/rFoZ2Si3rOSKJQJpoIxsSz+BLJOM8yoKX8ZlOeFZwH6VGOgO217xWPuCJu
u1PgvvEAvejir0KMNmX3JEbpCX1Vyvl47UX0O9JpfTnhfS0miAZfDyhdNk9Zf6EvLjB2hZugr2oX
wgpuPap+yy8RqMXpdVwE0cVgAV1OC128638Ve1m3z93DnORxzNlR4GVYUp40N2BWU/9mjXpRJtCC
9DbtM+ihP79iG7o9NphHcsaCI5muBlePdwAHdViJAHHMMpUR05ERnFJSy7x16NCQPrE/1yq0+r8C
p9iCdwEVCNCBAmbw9vg0Nr0wTrP7fBXdMa7ROK/l7vXpNlhvKqSUZySPy3KtJL5+Ay9lP6EjyGAm
PsSKTXth4THVbnbzW4TsRhgwiVWVfGLGt3wgregKQbEXdyBKLhM8GKXnxyyqy3Z9psu9HKcRwp5U
r8nofOao19lm0T3nuWKNujjLPmQNAFD7Z8/kps2vimlQjZ8ZQXbANmjQmPVKQ8Xbr3R7TAYJf4kg
nxtt8yrvY9qIdIA7gCPz9eq9LOEqKT07Ov54qj0JoSAMghrsD413G4PNCDRUmB3AGD1TyOOShI3P
jZN0pwGimecyY5bUuIwoGCweEyn4AJi+xO16ElmXfVoYILFQvrxBUSQiput/yFKVhmjG7p6ymDZi
Uo6c7RGfQjo24ZdIe85vtdOp1oOu8isPyV1oIEQvd3pvnARecxqnymCXMJYfbLIxo8vTqB1UnIy7
XslrMCOADrfcIgCtwe2ECpU7xEuZhitvkbnxJHcSHvXLxOfYRPkzloQgTfzEfMu8cs2N4xWgU+sv
chHtUWQZlKVirz3q1B/a5h4+Z9rLWqcBntPs/Ixp+ngAbjct7yu/RfkXpnE04OxJknF+2UGhUL5A
qtxIRa5U8epll/lMc/I0fZkHUlA/+zTRL7qJECBCldqsezpVdqWwmfI2Wh94xlfHv3JeoeqIiovt
nI0awhjb4qGRW7PHS07K7yJXo6CXbAnp9c6vrKdnI8+ei7lsfhp4xpDNv81ie6UwxthyELhT+2P0
WOkwvo5hn12YGUOD1fDxZ8kpuSoT55E5kSSbadVwWYSmfkCZjg+GcGoOm7PaY/dJWHE4AFRoXcye
Z718KKVN1xgqUcsimVLbIKnbfYzpUqgnu1XdgBTlfgDWPSeZWRk2oft8pEfg/Sd7oYA2RSN8HXsD
waMTzNWZdru4oIqoKOWcJgkAecwRj0uAxsOa4kLPAY11hrVmlgL0BmDsOv7O56sQIC3vTgGc242P
Eu477CWmefIRRKVGkqum0QG1g3lOHu4XZRB8QTMRy1k+efzWq5RrGKc97M862Am0qqvq36PXxZJC
/BeeIn6NLzzrIT7nAPcykExIn2cXQcFOULi5+plaSj0ti/tg9IBWJCElaiKpL2MTV84Lc9eRldjd
b6Ewk1Q03stXW0MaMzQVK1kP+9ZaN9/FAfgriOrGLCUvK/Vb+2B0/xxXksWzIodX+NlgsxXCcjOy
zj/XtLcOFQ3a7IG8CLq5YCjIch1v2S6YBIPZc6TPl3X3rNmZUOtxkaIhigG4JR/u4SprS3zwOprt
45jhnmrR2AfbsraEWApFup1VxRygUPjI5qb4DtPIwg4QbKhNR+NofOp3OdoTu16GShXfEJaR1y1v
LVRbSNBdRkjLqlewUcfXvY9lGT4oM8ZLrdr9vWX5s9jsJOw+gdhdvX4ICRzReXkc+t0wXxVBRDXw
UbCEBpT070zPd+nMZGk15hMnlQLlN20Q0TZNesTv4bibp8xnDoWAAWib6NPKxZ+MRupvd3BbU6o7
8lzJW03dUQ8nt8R6V9cKDr095MDpm15c5/mytpBugGsZ7GhhHOtQeC10IQQKkNman6CTTs/DOKkA
yuEajqHh6np16f9ZJ7f0GKX+Qnc4LyPs/9j4cp3zqQxne0v5EFteez9/JEbaaoqxk/HVq/x1VNYm
TgDR6Lp1Vja4mQUrT43gkkpnparXTzCMwwTTb4xpVTfbHjD//EZ0W3apzA5iwGqvqQobT95YL03G
pnX7+OS/M5UXvMNOL6jJ4fZ5EjOmTuqXipUEDHP4winyF3cCgO921JR88fJvGw5RNkjemGfjEsuL
Gh7oaRPWNPyPUXcS7B5+Hm+2XCqCLIhTW2/FfpgzJJUIwLrVbr/rM283Eoi5kvZqQQjIDwFYWtBj
mBCubSRALRU/nwDi4dBRoL8UIj5oP4xKoOLdBmDJD1+6gQPtS1DrZkMKlXM2fSa+5awC/SzZSQcn
ALF01sQB6RNj8FMCmBcIDG/wkz5g4vOWq7TNUmO0oxwRPlblxj1cnb/fq9yVAkPHaRcPZum1ZU/E
tuwvnVuwdJOSTgqyvhP6IKx5wCrO/9FRaAJk+5Fprl3ZVQsuYHM1fMOTzqzXwd4As25D3prCbABI
RX1lMxiJdoB92OxxlosxXdLRTE0uw6s7M4PP7dK5E9TTtJm1n5ayfhBl0zcm2U5/ugcuWIqKv8Xa
DakCku5Lmkwg4r0ijxNGwu29ck0kVpuUbqMfu2gt491J3WKCeYzsnuaTRC10k8peHdhIlVxlfVmo
98gje/7HqkFwi1fD1eSZJF5u0XOtc36rcptZ4UUNnmcF9LVxhl8JNsVTND5qh9e809Icb6tJUnFM
sjQqX5ChLqE4R1S19/IaoK6LbU2QbBjMTX2Id3xlYm4xFHcadnqiR2yiKQceU3N/BkQ3aKCI1EgA
QmgeF/1/ZSPAga8Qt7AiSK+hCpIwcXPztZiMRCG7lq4ozkjYriQAFJzaqeW/064BS0twCq3nj7bD
cUIpvi78TiSUVKW2dPGVlqtZDd3vSU44xD8QOr00DT8y3Bn6MDy7b6deuoGZx1npYY779UoB1jV7
564oUD5yKwc/bvgTreEXFVzpXh+95nWkRvnmjKr3FW2YJAyYcXXXrJYvooUoxSdwvGy4eGFckgSp
VIRIuHxlGvqg2upXmJFcD6QxAKCoGQKkxek0DVH+FpEEqjJfl2ynt4QRAWrwUtwzBwfc2+7mOGxG
Uaqi8ktSL9ADRFecJ76380Jyp2RwDVELqwSLsQgBv0q/2CXUwYwW98pYiDFXOd+YWnF1BWzGqcF/
vN/4bPW4/UYC6Cx4JaGE0UBtgMGXoowMcIR+v4E8YKg8XS7Jo9qg6Dv/Ik/pUAgrGG7CWsT+fcWW
tzIRaVq9xae+bC4We4YU25ywGGn+ulaT5FYvRBxURD1UbUH3FNsA0E6O7eofQDoqoPEK/yTgCGQ4
iVuUqAiJEmMFmX7gsXZoAyZMccXIEDHQychIj43RoRMDohu274w5M0gSL9BLCl2ghsMxxiSUR5Wx
HKZTwNiq91zYYXt9EgRyMeYa2UhLgTYynaS79746vMGiY2GbNpjPy4QDGUlyxZPzMhPnmcF+F3sC
GiB9nb3JZnUPu6fJKYy9ZW5d4vbtjdScAtfqOpwsiecDPkI2BTTzIcHYuQxQeGm5gIZsQ18JINSk
a5uQpzTTO8zuGxGAMaSo3BdP/DpVR8FAs3PhzR0wDqGSecKSXpQf83NeggyKPzlZmIUOTavm6P0M
cvJe1uvkVhulx6p4RcGddNsXxuLEXOUewzncd5w07YZoSAj4T2JcsoeS9AheiEa8K71o2eGXKaue
7ZSh2u8liZLLLZXFMdyJwNi/vbeCvnoFY/2egVQ4FtUYw5wSX0ZIUAj+ZZsSk5VH+Ne+XtT9iWyg
+NR0C2bdMJqx1/IXc243k6os0dSklAm4R8a1r5vhPbi8k7V/TyOewtIgpORw9uuOSBXcqB5l45h5
hhkXz9qX5/epTHNpssTCob53ovcpm09nDX+mOg7IK4ciemaFoUk5Z/JjupisJ8jPcwmpfSKih763
/L7AvemdKtQ+lAzUv5HSFGPc1juadlf9vAlp17CJtM+/dpqJjCtTuFNT2M6XtGHC2HFKo3THbRYh
jZ3CV7iTi9kvxe4k6CWAm+694BQzr8YzB+6QA+QakTCZC2cemWhFMWwLd+qh0bcawidFdxaGhVTK
ukeaY43LMFdaCTrCfQhdNsaegEzl9L7gnPo4c94ps0sJsK2XdnxCGQOyik5PMzaCVLs+MhFZuy01
QolRzhcQ4g1NfI3RwdYiNgqbhoyoKqLzjGt62CIAn+VQUlb4LLCVN/9ZC/dTr9fcPNjpBszZH9pF
nQVd6nAKe6Oy8u43CUvpyMTL6RORDp9v7SwWtj+qg9nzUUA8+dRAxko1huVIL55Fxqf5cWht1DsL
MA6GcsVu7x/bbNXLss1TVSJvNtXufB9oqGWK7w3txNwF+jzkDgVoYGVsYQ0IiKA6FGzW8p6PkAfu
uWBGDoCr/UZ5oNgO8jMKpe+f1fiyqNQGziWaRSDMmvCKJvHkwbvrcC2Yq2UgLbdKvM5lSg54GxDq
HKHRdza+1FarkSnm4Dhto19dPyJf0XYYfmVs8YPC8PJGT3tlwK2egah/EHK7jK8eSe1GCNiHmbpm
i82OdlUd7hzHfbLGyqcpb/de0o/B3sICUJOR5Lm1WXS0Bql9gkLzRcX2y8OQmxApJcOASSBEC1Ze
YR1fDig/Gd9PY9j+qbELWIAShvAvYgE8eZZqzyVbimxXoteeF7Bp+Pb48OsYePy2BQ6d+K52qz4r
tdx5raUa6Um1dIB7lUVsQrU37pYiSG1753o/QYD9xMvoC1XN/A0BnBAeJZGUIP62wJkwATN4KtMR
xvIGIVJwqQBthmEludPIA82MZkrTzFhevRK60dP4iT2DrDdTxhbYtfG3qDBP7yPtWfPc5Z3DfFra
Rwc2GfqO+UTDcNouEvWVYa6IwOfz92fr6pq1Ddn5Dlr3SRLdgWVJtnsOD+By732xRzXCxlXDUexG
Yk1fNaYotfFttLUTgLSlQRGE9Nk/n17afkPCJQ6+TymGsb3tpBgqZyWR2M16YmOcmJMWKA3ImFje
SNNyOikQ8bknKQaaBBB88+RkZxURuugLZgC2MUTl7kAiJsXcfJ9UsqI3b4RYCFvkD0r6qP3WHaBx
+RjYDlwmXUp6ZevJuxdLVD+KIw1fNJtZXGu+mX3sNBOJlhctKlZuRGEiramNYpoUYIgBHuG5RZjJ
ZNIHAmb+CUw1bkWtI14UpXXozRUDBDPXly/ABPmT+db8Z8WJ/0Utj+RigmIuxnBfA8fjrwjsD5av
tUHBFrIN3XMqjw5QihLZDotgFbfNx/pBgIgR/wqAD+VWlSRlOr2wKBWOGGGJSnycgoLsqipvXKT7
dF7IOST5hyTMhBxnRm22RzdW/pLnZSbtFuDXkPyoYC6kBgQOD/82Ok8x8nW4CMQjx6ym2BmQlxok
LV5NuVqyNOyj+0BFSl7ZJB0nYdYSx5V3Yjzl9oyXQNWSS+yq8AF1KTYRHsR9qomquuyJK802RZb9
FYZxzcReHCMwTSfWowPiLj2NgCoMCf0FlzkS8OBQLcHiPw8EqHhmVc/lnCSvxfxl9nDsLDV3/MQ4
1/Ae1J3XIsAtz2UAedzyDjwIvBijcRspLXTAKUS6VG+c3Ge+CSuQM3K7p3UkbY1lT8A2zrmot2GB
nT/ce5Z0igx6wRuwf0Zl5uba+EuTR+7JYTYOmflsx04sHoVkE9P39o03K6c/l9hU9prjC3IwucZ8
M5dyp8FePVFxIaSPYHFDT+JsEMMYWt8BRescjzpQU8KehKxXF+401tmk0QnrUF8+XdF2BFRFnlo1
8+ixeGFp2T48g9c/DP9vtLjvrYR5lUpsNJh7yqXvEsXbnnD37Z4GvDLr7mkn5aWwoIUsMPlDhoUp
cy66SQK6ANrryNyRZlByVRUpibhAmwC0yb5axCkYEzKQiNTvw+T5T2kUl3Wuu6WI9uN5zWLvhv/1
0hAC3/IUqYqV7Ifr5jt1eDt+2OMCDwm5lf32bXQmmk7IoFs3FmG8vC6aX5b58/WCgbsj0/LlWD5M
CIW4f8fU7vOZnyh3t7SSO0XNChVc047B/iHHsmx0nuEjga96E4u8fue6P6GaE7vFqDIk322riwdh
40Zb/0KJmZDGzB7OfE1VBvzb10TOzlESS063IJQ9VBuO/xTqxFp2fqa9s3WuommQQuS7GfRwMyzd
JglQwpbvH0aDpQy7TSTsDd5N8yk1jnbnCuVeuCjs+fcpHWB+s6V5AT0gEWqj0/LfIxg7st1/saKl
djLztI3IxQDMdsZ9wXIVlw8rgGPEhDDCMsp2nu99ONDdjXjB4Pih7wQwO7c8Qr++aejeKd0/07W+
7IE2/nhW69jo+6l6ezAH5dBTRWOZPkX/Ldwn+htrHXSjHe4w4u58WjWbzVB16ij7GKEGnG85+heN
a50TGskEW9CUt43TbNLUIEmRfPtyZBRJOKvmKG/zzqaqKGx+Z9aIvghatkGVHrYWePi3v3AEsml2
hnOfAgQm9sfVjNre6bQ0gKDMn/4waKC5marlcRNDYJc6+x4nSU0mMz8/qwL07w48CxEIzrpAcLbs
vN9dTKpuSr9BnXZA2fWmTbFMn10+hINN1qR99H6mCQro84NRTlhRXDQ2liP8t/I8pjD7LvrUS7QJ
QihtmQvI9l2b36Qcl4SnY0WwqBxOVVkXFP6Oo74Ck5blnr5hzlA1BhD2EJyr/b82zwgkOoUnJCAJ
fZHdADDn3QFBC6ivG0aKQYcXKJ4G/UBYhk+0wMqw8k3EjSg3GBix9NbRz0SUFiDuAnxT9wrXRHjt
e2WIwrV1chHILz1g9BBkfl1vjrmS0KpV3WkQomhX3bwN5fyC6cfoVsdKGMZIdee8w6GZbHqJo6aS
jl2dhm/pf1fQSE6E+3P0SSDHY4EksdQ4KnNwNEK9SrkF8NZar2ndHkWJ6RbanXtNMXyh/chuv3LT
QqC3fj2lfx7u4jhtTAHTqHqHjBgkRR2dRGn8CJvGZCNTh74axR1D6GpCotOTtnE1HFyYFKJtpAGL
2STp1CyfYSAcZxxuYyK5ssI5KFcajQxB8hHbgVFA2Xqv2oUv3D2otMyBahKefwhvO688XQ46CXCf
3BhTUNksXm+paPGavia8PozFNlLskogkPn3Z3kSY+n/kyXpvp+FrswO2q3bMPBLIUVq11MkpQEd+
/1l1BAc/GdB+SdxJ1sjn49jg3ahHUT8mgueHDezKKaqV/9H0KK9RxmJU4liKy+gaS3Gln59py5id
XjfcxgsVCLX2ExSY4lrRyCCgphxOZsd3TJDD9Bg9lk5B/tFn1dO4RoRVhB5f/COahbmfRBWT+EhI
W1SaQiT6udUQa3V19iNnrxmKarEev+XTHWJTun4PykZlWljZquCo318p+T80QmN3X1NsRp1sNf5B
HwL9b+lanmP7uOs5GV39wm7UKm6q9APUAUJM1lEn8YBanpRdeaom5Yp5DcGjnMVeSrmadzKmFgvq
kbz5WP4DEUrbld7utBlaZBOHFr1Wq6ME+iByhNyRexKFNZLV1EfIDyuj9o8onoCQ1kWmM6IsMiA8
0xlTh9wEcxdWaLtfAxs0p+r5gRXVQp9Z6aCa/JG1BM5hA/Y5hir444Co6ZAX+niLB7gd2Sh6Fz9m
veHsshTzB/yLXDwP1kGn/HXLWOS1JarkHBmXukVBqCV9iWZ19DEGG1RuRf1u3raHIZ2V5ttLzDFC
xF2FzYv9v5+Fcv4EEkxjMXHXS6Mxlf6xbbmakZRB9Hyc7HHqnb1AEfS8H6gX0ijx1B1yZJfL5BTg
qWxRfwKYnjqLGBMDbZoOimLSXaDUyeTJS97dP/AuKzFEhJ7bSZKWA5fXRroeyDnFKHxPcPXa6Whx
bfxGpbjES9Fzuv6X7aUzW6b7l7F2ZdDgrmrfKJH+sQ7sP98inx9I45rbVljQsT84Gi/GjWxjsGj5
uZKBe4nMHFhakwajtd/ufNE3qo3ra03LaeMk8ILtlnJds6YCuZmOa2SaWpxt6sK9pzkvT/7El1Pt
0iIG1rxMTSoR4OJDEsotE3WTNqbg3YgtXnymGEo9SxFWONfqXQJIXKp/6j1zt3IFJh3lDsA5EoCe
5BOhNXYXPaRHXH+ROfdBY+5b3Uted4icGEuXctpDI8pkaSTx5ShUuO3R2DYU/HiHNK6RXaQolWhZ
iTOZIPmPPjqvEK0hUHHRQdtc5T6FdLLHuRYeHLtyRcVe3hvn2hy0AG1U68eVCOQww19JekP4aBGJ
rydtF5qsMsTg+z7F4fi6MiR/vEtB3i5UXM/wZL1RY0eCFK5+t6nd9Y87N0FBeUxrye6iLiZEEFYi
hCfh1+QeAG98V2nnrmZSN7bV91MuSEbppD0fP3gpFudKb2SweBmGOJgU39y0KUEhmQCxkGOKb7QT
niHiijXl2R6XutJegSj0/HUQs9/Q8y17aTf53WUeIgVUecJdpDc6oJK8Hw/E/G5S3oWGQR20opjW
Yvsr15cGih6uYeMHBRVPL9c23Aj1wjj6GVpjMakhXW6K+QflSzF098r4PR9WpATFWudQdsz9l5QH
Pu1LzN3dwUbvoNnIqAKuJY/LTwJ3wsWMdz/zNfr08ONTNFI76makxtu1sM9KnBpPKUqV/Ullw8/h
+v+W/oye1PUGEatH3zrwFWow5Q6NAFMi2UXXj7Q9Njs+iAzWyCrNEwtH5G9kMkEBzRmMMKril7la
ifVHIL+/IpeAgX592GnVmZZ2B9HOqH20Us/Ce6LmYELLJK8Oplwwc1Y16sj5XbdUygTKYXDlWr2G
jBd+xSHn1y6feJVjgwRfc6AnCW5Z71kB6H6/98L9r0N+4ZSt7DiWf8y7dAhibGd0x7pZkJF4T75T
3TqrBd+rLG6FSCadEUTGe/MV5ulZbwme4G5N9FXkcVh2YKaWbACyvT4fbFSfx898IbHsDEInR2CW
Fj85lGDPn2GtOIddAJhgxYONb3tCzFukB/Cv4kG8XnIW8s/qU/AOlHpih2saBjVFFP5pHtf84uzn
GYwn3j+p7mmbSyxps1nvm82vjY13WJjXcaroCvjvvo4L2CWBB6c2iFKiFSgw0iai4krmas0iaznm
ppHnTMZWHyh86UiM3ovMzwwlpaiEaX4CbCiSm+KwwrapOMKVMsXSieepWy16eAufwyagkH0nfe4X
td2EvKUR4Jd0qrCXOCQvFXnmqPjcgNbQxp8Y13rg6TiuuXVopJmq5K/aK+3xCPc7mJySIf1NX0gW
VzIjvOWkUKdLr+icZ/D6pahF04XwkHitn+ibQqy5Yq8tX2s/zq2wvBkz4yOX1GNALdRB42By8FHI
n/rDLFn6FuvtsY0P58182wgKVX0e3EWsD+zcadw5Jv44PN5Jt9mWnWm29hHBfnZYDR20PTBJBKmv
Im6sPH9IadoDqSH+Ow2Kstf+t/tLdODcD9o/+Unj3R4k2SCJgZzCurB4KPjMbFyVQnGHP+w5HN6X
pdnWAPnOKkeF9tp5K87gnx9WmYNnqwQ8u4Uo1EIkw96M1DVATXGd6ASTTJIoDVA5kuMH8ay9BCmM
MXKgw+H2v2CRGz1D+Yf33HSQg4N1oXV7f3iKn1N0MFu67QOHRCodqdlIfqOL5ioh0It6oBgpASl9
dhlRNUdzFEB92HgJ4ecZ3olXcxJGYYzslflDVHJitBZu71cfcAqNcwsJgOeNo7hqlxR/7KY5+DKZ
e/4uaja1VDeWkZNizn5XANPArflibhBth4FFvr9ZDm8GBraz9rNa1XC9vI436zyXAU2ha5rbGgxd
vLk+M0WUFooYnFVnE0EOpR+0kwTa359dKZJLFU/gc6TCPF56+CfIi1p0WMVYZZk6AjIwbKSTbqne
PdvUz5YFN9tFS76rvvR275o+0L2OxTjWNXMApUuEi4Zi2IXTbEIh3aHYDsxyJgFpRjksyDuXsUew
G81kIztGq+BNTwlHy6wzdGBzSkQYvrTkIsS37lSVyzX4Jfu4xt6X3mA0CUntB44VdaTiRSu6TM/l
WVb/xryIBb3SAF1wOZcgnCq6q//X6RbFI4veXkbpcIDoolKLS+WfHopvI8NksvmRg/FgKUEbxVOa
0nnfqRDWTYUw/6acl/TueLKwVeF72YVzwLAZIvyJz5BYqsqe31FmJADWBheCbkcMej/T0ysqRBpe
PFfa/6gFhbj7CKxn4+BTR8gIuKb1jIXLnWiqSlyqdiH3/DT8PhoLsMrfRI2HLLLt7OvFvqZr2Oeg
NW3V79pQ1+fp9wDvwCe4QJhU1WiYhJSYg3qnNOiUmni1FhhbMxxRGBjrbtWNH93AF2VpxHywrVsX
xl99TcWIqxPyfgqwC3TIm7U42vUDAxk4X+RnQzkKA3S7+zMfagGnxSRXwlevvRRwHArxmYnAKrK9
kDo8PwGrGUvA/Fvtb6k8rxws4LFvuGMeHuzqdHlELSS/ZJiZwWYBAl2O6/WInDEsEmB+G7r3kLLG
p/iVCICELeRZ/7YoPncHEI3fDHTZwb7cppdZxzXGxvxLbHQq0lExllg2GteZ6wo6vIj1MpEFQjWU
XZCnrUlNCzCRgplmtebv+viiMDzkh+pGUoyXY7+bPoSvChmLIEUKdqPZt1/GZAEruzBKlVXtvbj3
rZgtM+JeANQWjImn+WfK/NcCkMOUAkrRNy3pAGoSitLVQeV8MBRIpKCE64qsd3jznC/goT/zp72s
ZGeoJq19L7+FBo2UqMZaHtHeY8Kgkp3kUNTVtsutlJ4hJt7FPm2wK3VMoqRqANP1ulilvUYjJ70z
4UJ7qGP8w6lYtzYA/rIHYZwOu+sRkt+zJU6Pyrf0qXaDBsTPiARPLtgCj3gqCGcUJ/M/Tz4mWpWW
Fe/wmGPRspyMl7lKTy7vOG5WlpnxjHu3FyspcNfgt2AEFnjkKK90ePXsGHoxq/8QP4pf1Yk7uQEj
/kiG56jAeXydn60VsnvxSXmV2ruRAl6B51SDVhaJODyx5Bkb4h20F3hPK6PUJ4kWQhfiGrGE3Z3n
Fc1hxgLOfAHlX9+mYApE5lCWv274Db4LAJbFDaLd1vgOnx+0HYd2XUrbJs8Z//j8XI8XYQy3IQZ+
wwae5NvFywH/Xd686WVIthQihSaw5mpglXul4rR+KOUKn2sqNb5orwXOfI8o6C3FFTodCOVIZkjb
nQ0LKEnnX8iEs40lFwUobXUf1bcF6EXtMrbegPktfrD6qr1zV7Pxao8pOPZok6UIm7PYiNnybeVF
xuljGbcKyoP6njRHKxT84hoks9B4eM4IoO0kR4kfNJpqIt/2K9idTsv3NoMlqD4GbQcSmetlT+c4
X4u41ohiGWZ17s7TsLSuC1uenn8fnmZIeeAt8ftSKw6jee1jkhbTmP4toj/mr9RdErIloMmfSied
sObY80TV6PYVoV21knFXhHa5L6j2wI0UEzArYWhknPFj3SsRREDxozEwFAoMg0wkzYRUqq85o4qb
/+us1i1I+gY96vvuqz6JKR4+OdY21YbTn/naMRLGi9DcX4lEf3sn7cKMSj+CMMYAcK2HA5Feia5D
LbuoEYRWrK9vZP5zfxX0cfoMzysBLF3633nio4we8/1SAT7z2YOVSFkbwZU5cNxJcQUd8rSzTmPy
quJg3heqGksC1+2kWKwdt5O/rAyRj01eGcCo/8Da4c9dlMmnT3oaTwfQ+nhw7K58cTbVO4u/Px7B
cahVhzl0kn3JIe0iKqGrZcczMt5mEzatl6Vj6mcJ1nIuFR/Az4EOiThVHrubNN67847TsP1q8kUv
P8YB+vuPeZliWHJ62MYzjsAbmD6QJ96zeAL+NPdMainI1nyLhOpIuNqGa7gBYmi7oQ/TKCwgLI8Q
THQ3AxzEiPXPTIdHcFLgk9Skm4WPgG2nhn15XFHV7C21VmM3rj9+T/jk5F/KZOKeVnPPrJxUJIx7
mSGPR8Ow+h6URlxPbxy7gb/wK8ietPCfy408Wa+UNXv1YNWD0EohqoOV+qwDdxcieIoNOeAyy5lE
BBcuQoNpqEc2eepv/Sz4sa5a6ejWsWZF/Js8mEW+RA4/nLdVQUSJ2YfjYN/GhMMZMJLkPTmtLyoC
X3znym8kTBGnM28RybN+HhJ44EX8S19yrDCtRuzGjjAcjrX17T3tv7wgDPjGNJnkepkV7jYWIgni
/8XLiOccF3h41xFb7RglxbWJLW91afAsSpUbEe1XOsiZIsXbOPQMtaEudjdYqEq2KQ9BB53zYaXR
ahF2r80zUOtaCjK6imUFbM5UNOC7gekNcA4OlnSC38TIfzy/OWKLVMevA7RcUNh15y5XVBzvohJM
1gE3COykDntavehRtYZ20TtfaJPdAavxUBldRzb16SxK+rCG9/S+kHiO38xbQN/ZfxqomS9O/Snq
Xl7Adqo2n/HhBfm+4/o/tFdtDQ0nGsyFXB1/GEr9JLFRhsMGrTyjGhyKS2WKQwNA1T+C86Ndbl4L
Ueb+wyhMLCl2AE4KeJkejed5NZkG1O7nkB+aw4P3dwCqj4ygOpx0teOzGa+Fu87DOVSaufnF3nnG
Yn0ykIzB9ottxnWq5QCNBKC/vD4r/ARK1JKf0bK9TyUWZhg4h9fkd7KFV4bKGj/5XC7Ombc+y6BH
LSdqVLuWbDaEqiO/rzv4c4tigLswKFrz7fFuo7OKfhD8S5QiXWcAF8/D/pmVfWyZ1hygclQsQS/8
T0qHnNzvAMN24E7flS+AOSwnQEQQ1brrQ4uymbT17UuNksQE7Di1xSeT8xe3Qjh99C7sDtbFbkVQ
AGC/kO0U/DlzrzxuN9r214u1EDnUi8AVY88QrDevkLeU/86z1mY6DDYW/cIlfkRkxXaeOuDh2mvc
vzvi2B6ELelCz8GJt7isra+VBYM6EUYdaaKKG2QX+1l2U8vtVb2YcLZbh57z+Sln+kDybHUEy/v7
BqJkzwtDtq4k85TnBH/tvtvg9GwjFxhgkuhfJqbGfxdu55AgKLFpQQR53lGlmCN9/RuETYoQGRgy
dlB81GtOyiL5GA8fRztkmPqdEnxRUwIC4f6t+BPJ8cuUVcG5Lw9A3q025w3LY7xLAMXhamx1OOHD
1U6WykfwNwU72ZJ9hDmtMJYZDcx8X2FJcSKuixblNOnlvU6l0+yFj9yDacTjkhah4VIU8pJ++COF
xzn/6S5Pb6p0QlbLRw8CE+xRFAekYPnXovfUcfL/5SkPUjeiKPRyoHCidYZFPvCtCsnBLrgvR8AI
JWhb6JSL4dkHWlbCO0gFLr93YVSqFPg1sx3hcOJ7MQQnT3l9frOGGnFJD+ubMkHdWW3pnhrXbglP
67/sxY5m1r3I76DqPP7uhb9WIswF635ysbik45qrbRKftnyEn2+qdcFkNR4nkh+fA0yB2AvYChaG
wTnh5JVSTMSEBKEeLqJUCIkK52go7UJruYVz81Hnk9bLoLDtKNaoWQN6OEAV0Q45esoAyhD3iJkD
fccLPIEfD/gV8rF25ZuakmptewF3ERtbz/tM50fyih1CNmZTYnucs+ZVcPga5OzI9eaTclKi9NNF
vvwUNWfsQ/aHRkEpEtjNh2aL7D5lmgAPE+7o9e5+E2vKdylQraRT4gtgYGbJ2caNBaYg/KBkrevo
TXSIbcZzxE512OwYm9CZtlZ/D2dyGh1wor3wno1EiC1wE2NoJkcZHlCXOS+dke9fw3s//wBnrPHF
FAKaVy45SU0ZBq4fsZPJlsPBmcWappnqe936FCYPrdIvuGCFooMgMelWyqtA3F3dF3xIvOAsbWlR
WhDboYHNlhxwD5YBXFI0FxJSAL+pxP6RZTxk6izRpsAMUm8VjgUWnR3kFvKsZSPXGUVKwdBr+l9K
kG+2rHmnZrAZXTLqol6xpg1oxjgm0uf3PiHqAcOXhNjFYfsyKRGM+5Y/VMtVBkl6Wi4/Nre6WLMs
9KAc924ukWsVoUnW4rAhpo7um7d7xSxSv0UAKWOgdYRH0vYLKvsu+6bezGR/FwwZmhdgp8h36zvi
WSycE07Rk7IArBVjAqMA9CIxkiK5SVbtSzl8I9IStFp5oOY4dbd931XLF5p9J571TUW+aueX4I7a
x6aykMxTxHan+UadEgE5dZJZc0ZzP/Kwia3KmiRxmbKrSGEljMt5R9M4BUxn3S5mPKL19iUz1E9u
5Rq+lz0j0XGVTDXO7nWe9r/Mo2xONw2n1HBlCjaoqleZ32y1NPTSNWRxEWjqIGJpyJN7oMNmTTSk
3Ehwu6pixAA+4YvsslIzJqHXIRFdaD+Lerinr+VZ2XK8G9xKcVeE7xv7V495ge5mV754xxVl0WFu
2JOrTri8rcXtyA9/95f1715eEj0RQLpG32lQVgTAEwRMUoCAe7OrUmtkSNsfhCu8vS998ucEjc73
69Un9eLsviUMFrHuAMfsWY3PCvc7P6VkTwsuyS3j4noMjWtTYSY9dTrjau94vkBGLq7FoRQMPCIE
1+zDoObxUhq/GPsf9OgH8spgjriCiSPRKjTAXKF2/2R9f8Y4WS3mYVUtAMbDW3INoLgimr8C7Uvx
Q5v4qz3m3PLVv6wXe+waKHqycErBwEE7Rk3qWdqX8v720Am+JS9/UncSmDOa+o7xw37o2sYTN5nJ
/q1TYlqOBoX73yQ2nKtX7pLZjG7J1SYrHbuvP6Jxcc5Di5MWr77LVM6LQtpH9AR1D5PBO/vrSF/o
63VUFK1Bz1ZYyGz86NTcZLWAsdmxIZ30SE+TL/CCyE4IDGIYRw2ufnKoIFYP/jcRXZN+yWcEerf9
kP69sak+xFGnUY4OvOYu5MGkjVPtbVeSkXMHZPhGPRsEMn8w57i9r1Qt47xdlP0TUNrJGpnGk/W+
NYCOl9ojjW8ik73tkI0wuglbhHhbVBgSvPfgR4CE5u9jxJrzP5Wlke8/S/G9uXKEnPyV9x4P9jVm
TzGTjfeW3hPuq23Dki8tKXtCP4kPGWdWeWSOQ9moHHF4Bwp5CFpgyAf8d3KXaqUKuLRAT7E5m+pJ
VIQkxU//ore6GUS/CI1jD+jtvXXlSdhAcbDSWmFgPdozWSCZNWEpTDSAaqRqJZiQz4GckZCA7nW5
sTbXw8K/ERvBGaLEMLyWyiTJ3kjtzGGI2XAjve5Invi7UfqnC4hHIwiMR2D0Eve06U/eGue65BtZ
ddhBMe9En/w/TxM1m41ftJodCP4Whtf/BLK4LiZfOc8I465yX3fAL6VzLnJqz/vRV6xMM68B6OP6
Ov0samluEDSecayPOJN8jv91EVQmJitd1oMlt8/Pll/deNNlTYM9Ut8xFGiuX/pShjgGotuXfIWP
myWVpBzc1VlOOzFuwRy/2NeXLZJNJmAXhwE5gd6kw1v4PjCKLRUVSunQ43XLuSWc792sqvm1vKER
tvaC0PVd9QAX0GYq3bRA776plkWudL9vIisLHSwcmsjly0z2favQA6N3Hwb8ULrfea0M4YhJwyuP
deFVI/Gg/CDPPeXQa4sfxIJqbn20EKEsJTq+17YevEcqMWbhl3HRO2cr4eCtecS4UxAhpUyRHYU8
SSIry6BAZxTLN7L9WixLyphTnW6P2+y7aDKhlNhn0Ye3YBLJWjrKm7iRNyTh7FUXEnd22vb8wk2v
W2dF6ziY97MR/X+IGrYEWRClME5ZKHZaFmzdLKUP1TEZaN4XajHw9y/lXP6g9mNKntGNeY9oJ8CZ
KKVgxQ+jEPy76m/QKxVh62eBcKKHNRtC272xxfzx41UwM6zelsPLnJx+DtQknYMInLMGLHGgTEtA
tN3+Je1GWh4Cp+ByZT2X004eMF/RxfAhhCYnLM1zyptXHt7tzibgxqLDIHOtHninOk3xxdpoNonb
XcqmY5p5LRJYiEZkS5Gfm6vJMMVTmejvE7Wq1x3a+ASMp0MBsmyRrqLo+dq4zW1+jqilwoGJTmYZ
ryMPRmkV7mriGUYvr6kiJ+WOYLeo953luo198Uh6s29vjN45Xn9Qp0BOnMF3hyIF4JxwCIOEiouA
giPM0As+zrD8yBwz6mRHJdLMym2j3y3PnzZzEYz+jMwkyCqB2yI7FPhYYWp0vt7at0i6EfMYnfTT
mWVFMpxdU0180hhvJsGZUIqdyb4pldX+bh6vKq08HMKBJQLYrK6qQBLANowdg/CpCf9Lm6L/kNrI
l7YsxnSAjy7qO7Skeg1JWoHgXt57arLBAT+wwH84S/8mWeHyzmdWbuT3NJjl99d3YBgdAQ6yo+vv
m8eFfaC3fvroj9ZXu7YhRZy34B4uRAJPhPzsqFI6B1xZYzf0Zgy/pLbFb93Hami6FN4wEM94099T
HyxNQ1rwUpbUAGU8cEAJJXqe/Q/bH7dCwkEd04F1EUz6wb8Uc6jgg714N4soDEVerKuGRIe2Y17x
B/rhNmGBsSf09aeQg2NsJYiJP5n5C2e+5au2GZWSJtA3y7qpt3EeY6b6X6s+jt/S91ujNqlkpvlb
cfXBmD5t8bPT6kpMvHn8TUtPtyWGI3d7VdwGWIA2Cz/U+XPjuhik7ZjHZy0/qLMtKqkrPvqgW/Tt
0Mg2jw+27WOD+DDfhMMjh9ucX09V9Ebg8p3L/q4IDeRM+KOJP+ovue0BNzkt7O9RvmziD9mT6LD3
mdax4eesElj0jTKr0BzKNltEls04uJR1hofJDH5zrjRXixtSrqspPD8ep37astjIvsazS19Dj70I
KXf2CgdwSKpcC84yuwJmnpE4hJt3lWvZzDZwFNop5TFt5637UOWhNDKke6W/0mjTC1ZvOpldl5rG
hiCJ3uDtY36dOn1AmqNwnUGj1GPaqLUo15GXJzQLFx//c63OgFY+x8ybWkgMl+7h7nmrJYRIgcIe
+UgPnIOCxjqerp0yjtMwGHJTOypdjRcTMs6Xd7orINSxBiULUlgPgkUzL8ztZT9VNRbl9gJWFzK7
B9lY6QGPpU1jgUwXzR9twzuY90aV2St7xf0AtrM9cRFXmCqdVeTWYNt+dGDFxrLdjF1ck6bhVrny
JfKq9QAzIzsyaWKVS2mBEtfjbbGJS4s7HRtCgWXxltMZppUJ4PEbFpGim44CJNzTgJIiKOvP8lFy
2uhS3Df9EV3sSP8Wa0hhPnyMY6FUd1GdZmR/ZyiqqdGOBejpdLjGA6UTN3yS+QTfH+HuJ99XlXgT
rMTBPNqXEOxcqnSuHSktr0fZtLAHCTPv9sY4J3cl63YBFFmuz0AIfGIheE6bqmZYhXVZentmtc/j
kAoAedcOct+QDPU54RiKJHQ6PPnzFeUD/UJ6kZaeSRqrIMxAUFXIxNZmCgCt7MfgwWzOftALMrk1
S56cT4Sv1IKLy8ECKAiYWaKhUYK6wS5WYXLKfFXJvPUbwWDJo3WiVIQPDfwgoV44H/t8s9w5jG0R
7eiZoLRqyjBwUeJByWWdg8VCSkED8NuYxXTU6zq+qpquwceWEwvpZqS3ghUKGycKP62O3kObnKhA
B3LPQR6SnSG9HfVDbEkoV7ltJ5Q01pYUR+CDPzld11jB6O2fjD0AUAMURiqPNSr/Kekv0l9BqbKG
62Rkoi/YMrkpVjvX2U5nBpHxNvEFMFq4vDT+Uo2q5/bjj7U6gpKr/O9nnLOu4wE3Lefw7iNtzzP6
gMlHQp+IxFt3WmTQXkf2hfMwN/ULW4cDzqlMVPM0TYVqDPC1IamHVyJstMU2sVtDch61J2l7zUHn
rJPHmXFzsA9yAtjaNFma5sqcI1t6z0Zb+F2Gs1+uNpaVhLW2xMvDX2R3zxXOERKn4li6L+UTtsio
VSk9XOhWCI/4yrEsFWse4EOBRgJo5ehENpewNgYQbgIlayJw6TlOJaFTDlYMaePHtyVYtvbGT2dt
xKEbAbnIRJTxw/yXX0OaF/jvS5qU94Yi5irHNZ3rCpjWpY9PR0JEZ06MRzucQYxK1JRKPedL5uGS
qHTpQyBFX4/gKBygonKVQ8jeB1+atPZIWRZvfMh6QVwOWekUq+ZCYuecQ562SlNDhelEHuJgYe+M
79X7RGVhMC8VCmL66XhggvVFl5YNGTLz9+TEh/wbus9uKX7Nieiw+WKq3HZuQIC0qy1qVnIttF7K
rVXInVIY1VweD3blkfCEi/VRagg8Wohad1Sdvv+7jmfNgu7s20H/E9ehnhp0eRoTJQB7KD3+cneg
gVlEs+gjeTYITeor8r8sUEtXBVvmBeawINEfvIHgf2IH99g/X+hEFM4p3L6ldexkXVfuCg9Rk2pV
UYhJVUbqMD9WAH1oDAmZHCBP1ATaIkE5adbwEaVJ2kVelZ4f/p+EB5OkjKLRIWIepu0EonFK4um7
SnhiAGlEiQd8FblimAO12KDVHSi823t/sOafQZ0AqTx+XRcVAhHC5ZmsIH3ZmeZZ4VXY+mXBwg1X
7dRyfvxZblEHbajOGDQmsyijb63iPS2MIHE7Ey+6QqhMGjDmTxe4uMzQZEEyP3IeXVYpbXODreOK
S3zCogGQg900NZ4QXWB/OGU6L0/5bqp0iIlhi/oFS85brzqmMexihTm7/go+E6U7F7jDEHXAU1FK
ePhSQQokdhlwG/R5uhfcYz3yhB4ibw87SH7xBdXGvKG9oYgNt6iCAxD+PjC75Mt3W35J3AJFVJ60
k5r7KBYzHAf7lNeGyhKL7Ve8Tmz50C1C3SlpoW5EsiQAD8/di8VJgCCoOfFjBeGvRVk+2xybO5iv
Y1uXhy6HVbUrT2NM2iq2gRhZufVttMF08kToCKtYqx8dkSu34PwMyWxSSBTaudOqsawL2+OP2hsy
EH4XlMmgUYl24DwkGM/qD7v7L5iE3zJyaYxgm2lgGvIlw0vfFX7HVM8M7K30N4K7NCE15e5KhYEI
w26ofbrP7iZlf32UNtoDWplQCxyuZKZ0KO0JptTwtsyL4X52ed7lImQTuDjR2L1YUl8D0v1V8NTF
vb6EkA48ehONUZL2exnZXbq+dwFM/hMm05HyKPJ+p1HTlFvdfYI+7NwaCXIr3E8K5rxP2rkdw60C
gPi7rCMTuc4EZkVT6pybnfGotnyAHYCxViBqGStgYR81qW/zTqpjjqllgrJyC4M2HqJLP7vDlSkA
y4BMHdHA1n8/84MIkCpo66Xmbgoldh4Hw3W6pPmv073HzkIwtrD+lu3BhOSZgCdU1GxJY0QK4V3F
XXMhOVc4hOqscp9UaHQhkAbvN0dF8xs+8A/glmTTm2OX6t6QwpuoNrrVmP8aiU1yoWtWlNJpnihG
6K/zyEPbpdvWKtdIhRtB6aF7N7iB8mxnctfZ3YlmCvTy2hDFNN6wG4vqXa4e4wxjRxZfWZLT7YNn
CexyTGEQxMGvNfcq48QanrWKB0wPuPEYAr+O7F8vp4hxucdGyPoqWlyMsBlIoBPD804DlxXoLCgq
o+C+M1v+3PEWJ5UHONCB/kSyqcRVkCoEFoyCB7yrxo1W0oXCNsjVrHJc7WK9KnznZmjU/RRSbGz1
liCgrJp0pdlY21ePPigwk8dj4v8Xt575VKYXF5eDpabHwOQWEOUOyGI54BVGFFSYB9fIEHOuyc4+
8qIU9xSsj1HmwipB67gcvFk0J2HYhyzGh3JjAlM3vaGXLDfJ4XTszPzNkwiioSRwxMmzVrrBeKOB
WQMLXxKH5wDS3F2C6KzXy/hIEVnbTK6fn1m0ldzsLlN7JEiuBUZt5aMyHJbKdHLlOBQ/lFn72pt3
2gkzU1Rvl5Jmspg91/DYmb6xtJrco5WbdhLf/n6B3FqMedKrDHhHE0u0sSjiOBvgXWXP2LTRJbQx
/WVsB5IdFYPb6wjmz6mnAIdARxV4MTbP8I+h+CYFKqxKDPForsicbNYOng0jT4FQlM3HvLSJWz+1
xYWTLSEuSZOrTNh7ZOXw7tE2dIWl7RB3IvT5/xsZn5Y3AbDwaJK7iDQndomzPq7qrX6bYKIAaAwe
PNx5evAWH2G/U+tY/H9uECeh9E9lxsHSdXOvZ+95Fv6JKVwGagdb3qiZe+MZ/wgeAf4zrpCGF2ps
825fLUYPdeEEHadvMnGBvv/1nC6kaZLUH4rcpcLsZKPPZhwqRqCaBkquNP6ujvrPCjQKWZbr0j3E
t8Rd+hjvWKloN04ojWg9EflFS7IfoC63nBtrFzT+lbbRFxosv7wNMh2b91HVEHU934qK0uBhYsVN
8VDvYrl2uM9S2dFgNshVEyiohKKVEbtFlrcbROYkUAC9KoHtPpnlLXzwB974YJjHO1iDwI9KH9+3
PuLZsdDdjatVpGrmy0BE3lMX4X7D8udr4iYbAfrV2SF/sCAFsace9b9uYdTx++J1fQldeefRDDur
wKRXbRxw9lNm2ohRSAYROLVMDQiYxOCvn0Prv1em/IAiCU+SQcMTF2gYkpksr7I3C/095yYHkCpA
qkjyQoWtclQHQgVc3LlgeGeK2fX5FaQszcOrbf8eWvymb2KwN8Kqx2e5xH4N1neXwklOeQWw/P/2
Vm0T8IVGSPa6DY42Upyjgo2XrReKkHExLP4dMLhR3m66QK77YDE3Nqg2qEc4Agkpbsqo42SiRozP
GNf+CJGkBGogSQRgUaYcVsdPJoRTyujMGY+E5zItRFZi8Px1YJJGTys6xKVbqWovBSRN7P4tWlQ7
psRSMB1LDPHOwN0vgKekwwoT58vQWD9kD7tiNC0Ox5O6Q7AqbviukSkzZ61hPH/lqTbQvqGfSd1O
+VPRBSouLvGRYR2BDiK3dJlYwxHvZ9zS8KVRGw2K/vn0z1IbOZKVMCmcJjKOK13Anm7xgR2/QLke
tJr5csjaP1YPOD9O4lcVsnC77WOYSvg2iY+qpR1VC4qi6qJFVZBE0xujlyasERW8dpJyiV7iWb4y
8Je+4qy97mQZE9TSe9t2YLKVvTFbouRtEo9yIi7reHdUVgKv3J1zbaRPnWlGkmaUsCjHAm6eWkML
AvbHihnB4hCpY4aPxXVL7l9+375VAqyAJP3B1f9nBDD0ljBlaQnnXqDrjS1CeD9DjuuLqgZyUi7l
x4kEFBZdHIPf0E8xosazXG5umXRVIdpxzg6XYLRviSdGtZuyhrdFhH/hyoX9siNb1pB2DB7VAKoT
qgdk4849VrUYUysVDVfNfatyEwHsaDbH/XmgbMjQWfyi6xg1ymE+KUCievqtvD9p3D6lcr6+mo+/
VRehLK28R/7THJMShJ3P0VIndCn73ClR2hFHO3b5KvaMtbnowOF0RHBXkBYhAxBSOI4ygbGlt+pk
FDYNh9O+Wjpr3wc5XH6J6t7Xq+jnb6zH6A1MaruQcSHHBqwSc5gRQYN/a2Gdl4sWgpmAWJ0rpHGr
auZectMM9arDDJ3YGIEqF5sgaiFTMfNdoP+erZTRMRHeRUZm1EbDdJ4fmpKhoDlCQ5z1J0bYXE5p
QJLVumBvMtTEcanEcV1i3/hfGH4QFrYa+JL4HOWQPfdM70lAK9TqDRdIPO3PbsLLV4ivwMCoF+bh
rXtNrDASq5FJv0wMYPHG3qOrDYxAr/3bZlXQ528Chf95Y4/ng2+vuwu6tQVEoXRzYhpw9H1nNa6c
Og5f1alfn7ypU50nJG6UmcHRjsdHbVaIe30hHTeE9PRiQieQ9ery0P/4Lur9FnfXB/E6VPcH2mA+
fFR+dNi/+IJCY4pTrbyl5x7TDjLmx68ITf1hgrIZZX3P1z5rlz5xe/M36/RG4chWF7gr6vN2lpxJ
Ip8EHuChrPNWHU7vXwCufHDpkfIbLZffnh8dj2ExASYbs2zo9NYSXyV1rNa8BKnyUQuO0VZsnpKH
tB5/V6xKkwhEx6QrYtsYr/Rx341qJmvN8LhRU+wKjOmD8oPR+LiKNmP8my1Qcu3rnp2ZGr7HfWHW
ym2HunFPMh9VXKaj7+j5/hLnXy8CfDJ7L+E4r1IulZaAds1U/KSIcPRXnc13HrrbkaAH4VC+asr7
YmseY2JkMhNPW8P5i4dAflH/4eH2bhkG+8pwT/svcmX9VWE+Q36ard/dKzOhgi9jIi7ypVoVQ8v6
AXS1YsP7qKvsCKF/afF84ZJkXdM1HM5Lceghasj7JwacGeyK+UOMdJ26nsj8cLtyixCgCV2UbKWL
7wi9S13tkf1RbEWh9n0XXvLYKZHNFmsnyssy0p/9jrXhlLH4S+8om5xJDx1HANlqHCJ+XyNrsJGU
EseFdu3G3sziuyY4igC8xW2LBPL5BNrYO85xL60MQs45aPQyUFx9u4JBtwNE2/y7vNsWLBSYoj6B
+m2ueq3IKblIe8azWFXeQvDH5Xgcd5UKmaHe9IfACut2oyYUclMvuqzyjF/ckJkGtOP+rwrF00Lh
HC1B1A3uP4hm+g4og9HuiVi0yONrG3MpFQQ1ZqQRKxzEX6OCexdaP4ADJRywj8IvTaGZIELG+fHh
NwR6F4VSqwJOzLl+TrX3y23UsXYnAu0/wanQ0tKwocCixkbIQNProD/Frbhp5CXZppWJNzFj6Fz7
3yOPD2qXGmKIX9IRHCRY06Cp0i6gapFipIl9orsneVRx76CEzatV+FmTFkEMhTtJ5rCqsUWJNNNQ
4oVlIU1vDPB5YLtWiwaMK/08az7HdYZUWxbvtE68LCLYafY6iWFqi3VvvxLo+D5Oh6vMBINOkslg
Qa5VXaWKDVZMo7OTu6GaymwIiMeKEOUzt5M3hg0IYNFoozMFzPjO+SGqzLjmMewa4uUaiNAZNAw5
YKy/WvyEunCk1GZT7m1OgKyW7MgEH0E8/xshwQcj/lh//4/JcvhiaUo2ZC/Df/AaJk7P9DwQYNxv
EAiXq58loeVwlBDVt/0lj5hwb6q2byS3fZxDpwnsBcuIiQpH7IVsGQ0HeqOxYKmOkLm+gAYqC7jZ
Y7R8gFVqXfwm9Ks9RMKEIduMqfjjp4iQUeCkud2R1hDa4of3iT0C2oa2vWkURYokOJwcvIH+rQz+
kAXZ1nYqNikLTJliJGFLibaw36vZF00X01T3jsD9y90CJEdD9Zqh0Y4hFhvKz/93oTItJmSlrEiH
L1qUBR43HKHEglSYNu7VS+xySHssgIz6Ub6jbTWH5kBrnlJFt3oejNDmb1IlkrRUVqBt66aXBJ8x
sl622FVTjGgyHdzS5c95yAHRxTJn96e2JRBXOipiZfgHqIH6JtjgOMeUySqEV/iFYoQVu8YnYug9
1A1iYq930qq9nh2GBN1pq7T2n7C8SEuJfNNUi/ndIqzbDb2b6DFlfOo7qimEvQW8YhZQAa+OtEmC
TYIaiUisyk72FaLlReS6hCV50ERDf3J146GKNYa4ZdUHHKkiVHArQ+sTJNbROdCL27bXjJLppRZA
FWj3/ef9ouy+r3a53fSj1Yq3L74rG/+FQawzH5eDLZvA9vpmBDvH2D3Iw0xNuve9nm4w366uVrsN
+/61whyYEPqakoLui+1xbSCMAe5+O6vRnuPENtCiOhRrDW93/0jojYddLhmwwvUZdINqAbgRs3KS
rvs+TZFPBqChc9Kv+QZ7f3k3Zin1M7l8oRxYy1WtaBG9/q7UqRadIfhN0G/0N9pW+dt1eoyafjtM
H1p3Vfd78iV1Q0En2L2L/rqtOQH/4J4VIp3R6rWhQL69EUzOJAixGCHSA3V2s4dW03CH4RcbyJuW
P7n2nD7rhveyEWEaL/NrqbR/0b32Z7diR2Ph4GHqwGhm7rq2CWeKe0FZn4U5s4sn9T6VjNTzgWgK
+/raYrf+biPZ5TkraoaooYWZQNWMRPR27dmyBLqwOut/x39s3tkv8YFmLSKXXhsi8Q5wyDUR85q/
7URIYo3b0/Qi6SHsjVGxt/qg0P6rUnqrrn5oUP59wnpMNadC2J2kgIho9lglc8Vz1ufaH2YzhKaL
0ELindLcagiojV6/ff6D3r3r2UNjxnqkva/kOAiN2Fo2O9Wt1loMCfALC9Lv0Cg7or5sJeYQQgXg
l1q+wBeN1CgovoPAHyvh8WKH137htgr85RCyovbAIIzPxDs97QVWsVPziAkHNQl0FjcQYeq+58IW
xYlOiUj47kAlK+1IyWNKfc5XiIhVWONgo46jGNKDokFbfr6o2UrzCESJm6/jV/qkd/uvjHOdzAw3
1QX/d7Uw0IEKMmFeg76aCJd1QCqJpGFj1F1KG50WYGiQwokqW+eAfOcU9HXKgRCmkWe3+jMSxwZX
PzM/h3mMAbuNH0tP/WWn3ZYm9YCPRgq1v0vvzXY6p3SVU5UiCyWl7ljuT4if4u9UGFYXqHVHHkQ/
IVd41J5Mh96YIgEAXP7fFeJMfzCjotZY5jCxqQr0IyjcxWVl5mznSjDKxThwQ7SaMVefNtn5fpWS
ajWqZwXgJVdcAfwjPYNR7HiEImW91Q1otrBA19j2vSdLI7p5lX0L4EvUNClFOpDTHPNia/QuKMOg
lvIasb4XoT5xJ0AssJ4xL2DvjG9yv1Apl77nxDng2o/TRWaaUnX7uXOMQJuExopBtte71By25DH0
rYLGaS6hhv6ivxF8W0jzYH+NMxZg7budZta0VtiikDOoLf1xx4qUmXAyd1+ySrs1cNfiCKzqRj3M
+PB5gSfIe4YiIA3WrgkVcBg3TOfw+FhyoWIgSYX54Bl0nNF47nJIbL+ydBFAa9dlKK7Fn3Rgdfqt
1mLjiyoPz0OBKsfW0WemGjonejecGuCYkaUF8MIdkJFVFyx8z4dMRTAXpCfEhBSZ+0XUGq/P87LN
PtALTVBQpkyup1HiTOnoVQhC2HdjF6cQL5eDj2sy0ynUQGGjQEFU8FwrLPZDQNWlqDiNRB0uYm3H
9ckYsH10E8qcyWaSisVFO7RxqwfybhjcqhLoF0pk2e54izsemdhP/4UcAt6R7837t0dYO+00MvwF
iQh0VG1E4pCdm9PT3kFSjctcW2F2fLqAVjPWreWxo0A6xOgz103pQGAgo39pOa0DzcR1jjhKlPxE
5riksdhSlReP9NM1BrKSxC0cbCtFM43SkWNQGYfBNbs/SZ7RqUugsc4qrZmp9x7L4udTOq1XfpfX
rPn8MosB+dmcLvXjLmOvvyYMRqep7dIrTg6dTeaXdHu8ewFrawmE/bHXFqK57kp545mAU/xgy4Db
dMU7ajdCPDNUVhd5oJzfZXGXA32HkkMt0ypKFVA4mQ9Xvbra4WvJVvYmJNuUedU/W4Y/447gIGff
2efZGk8FeyF3DZvFHUHVSKIEX24aXupWZ0W2q/TNnLWSN+ECH7wY9GyB6ekxU3RrTgTHKy/ODtAp
bhd0ZgEnPsnaCIFB3TxF3w28rujyaWT6hAdziARmz2Fitoy1ph3rjFQVw1SoVSEcso0Bk/T31m23
jtqWRyQAfnO2t4PA4J6eTuAuJOcGky/Rpq7OiMAF0itLCPG8rLzevEKAFF8Da0w/XSVWmQyNAomj
mBnrClyNG4LilWFULbwrXjm+33qCt+rooqgGPVQ3fFcARIAukib/doLMr3MJ5o3wb/LyD3wt0R1c
YiDLqS/8xhkjPu+FT/luzWt75P0+2pheoGy10tKRbWOvsHF/5XIqC1hBR9KuDN0dhrD/VwAEdyJO
RpsqpmuO3yIPM75mKCa2R8tTdfbg6ZVa3l9WyrrGM81ABYAipbxOzTsAKON69QG0zZm474zglPiK
OWNEJKGu8Fkr/bLvOfWe+pBPxSf3q3C8SBbuCVxzz+1+H0gjj0iLx/4dyHvyRXayEsQVlW+kKGxy
0KrR+CoWvopFF/WrwotxXnQdZUtBwhoZaHvgWQqJnkYd+7dDmcdkwpEGyAPKHXpiZ78BpBY7jw71
HLHoBU3dOLdBiUG+oRWtlfhdy6XHunglHpq+zQtEHJ9Nwc0ECXthUwVE5S0MCvZlDfioDwadaaGn
2X5cldfZ5lluSSRoIvbIIhemIlX/LBrFQFCOPF4XUBG4l36nK/9vNgZfHz1x979Bk7IpUrt42Cwf
lT8W7MvdUmdVotNHIlzGWTnLul7LNZmszrhipTf3Pe4RUs6tq8dm0ttQO8IAqAs5TPH1IaKfwNxA
axTlRA0uVm3Bh3zQxg5fZVbcqkhg3TnkvMmc0puCVZVTEEzehXmK6rJYTotLlZiQliXJC5BYk6rY
GAp9h3LAuRVD3cVNC5XoX7Vy/YmFZHR6t0IjFClEsKUywn6CshkCFIEesU0faJJyyq6eHSXxTKtp
NE95nz9zbuWbzkTYcvLLJnmqVnS5HxU85Lb/3PkAhkdLD5Ng/SOxRSQIjmG5i1gWCYLMQLtgyIcU
3C9FWaGTQ2eRolzux1LdLARxyVeteVIMWQZR5zo2u7iObCgvFFjWLNU6J/VxnCjM8SzBR3atdH5/
CpXQC4HHnqG3dquK/S7YUhq1ppbyQEoCQwrzo+I8MpwLG6zDLmn7ZLUNPxnbnirPSxtFh1Z1qacL
IGwrv/DYXLTFjpaWjQXFyXJTcsTONc/MjVNxMMO9CO4NPpdTOAMXLYPBU/JLhZ+p9+tqVzmBFG/W
DLw5C4oBFVDr93lm6GgUTLQozOwn9yoxHuSX6CDl1NIlN/TD3NB6WgJdfVqzKENlI3BLT1EHlebP
h0ldeO1V5nX2jAVP79j4402jPI1AH1P+JZA8h7kBDmZi7o2ZpJ6TX+E2SZs5fJRAy/g0Iw75+c+O
pPQs059ORFxUDbOc7vrycGOzW56+HUZ4DXoJnZ04+W6MPt+oQ9GuB4fNbDB6aW/2PNp++uwwaOoz
S3Uc+/GtaMurR6I6uARhNrCTsEF/4OBwmLwfDVsQv15YusxRQzTAbJDOfdYQIvbL5FcyziH89Obx
ttXmBRtPG1JX6ODVMBfHyf7JjjdG94vi2JurA8h0JvXX9TxFTBphG2+XghcZyg0YDSrSPRGqFTGS
7l/esAMgEahaW5jAJfa9Ld9Zg2sAv7Td57pZxggKlVjeDSdmEIakFsDI0mrLh2mm4o30p5FMCLOD
JW7svYpAtHizDnML8nq5TAHj9r57V7yhPr14kqN2QNMaFN5qkx0o2e7SD7xYOepS/ExDEfozFtdd
IuUxWuLo0Cqvq2ljrZnyPIPEQYg3CJvNSsMpaIlIU/F95OHp/CENh6SwEqoJV6g9H29H0ctxptWO
0jwUHLp4IaigMQ1arGaJJmzPRAvDII5qk26m2gmbj895jbs7SXmcKcsCrs8U/UcYbrmWZjOX3FI0
aZYgvZZTxrsPgK6CHw7x11Usr620Kkq8l04LmRF7cGjVNDuPKZtZG+5egr7TC91KQFt61cv7McmD
2lgDaLpHg3VO4ilwVWgMG7Bm/BwYR6ODHJrsoB8ys/8mJOJPnje+773xb+v0LB0Tfds0zcaBdBGb
QhPnT9T49EeXwQrsgSGimBR5z1SBix58KWtPmyF91D0MXNvFOJ3yVvEzzYLyhKhESm1rQMqyGfo7
Lh5Ste4ZYUCEj+tDmJBeQpjlyg54mczj7a3S+evFYPikar9KtoILwsQhfQfCcxFsOhKyv9L9WgrV
ET8Y8UVSTiOB6/6rdykuVOR29Hnyc6qLd5kel2xOXyGMg4Hho+MTsTenbAHAKR5Q1pjIsE6SE6+z
uYC7amaTjcLbK3EnFoqqip/lAM3yf+hds082MyR1qeKTaTiIDvMjDbyr9w29PvxNxVHpx20p+9Ih
vlCNMuHogOgXYyyyBpycPqpeDx+rXIus7Jh2UkmswRtEKmUjxxKQxMuODxzruggvvvmFl/jFdckZ
S/YPEYjtES8B2NrJ3oIdHPZnK6IoT1E91jIWl4q9IfX10pZPTl11PTfEn7brlZZR4UeGOxKiHzhP
wdGBWEH93kKU047VDMpEOvUp0eDXZWndEf+Fon9vEBLTKXb2Ecf6i/JbVE9CV4oRlWlcjGq2Nc1p
qtZOsXixm5YNGWMXkv73WqY0YoN4K0dFTnlVKr0EN8JSRaxguSYb9H3ghQZnQakaTjVRruq/wCxQ
3bq5tBF+KYzVMA3Jum+A7sz5C3LcmuKKpbn9h8qwAajHdySvpr0VCpyKu9Jup8GG0mvQAiCh7SfZ
8NFdMaCXzgRcD46IycqkdHrpXKhX+52PjYUCkFPG08WVEkfSC3GqdYU36GjdetKb9m/gvT4EBGP6
hMRrwwE4+eJ8jgqCpPz5b8ThrKAB3e2m4m6uJ2vqKI9POImD22UbqA77gi6tsc5sCQ6BvM7QvdBB
vqG8v2xSOIaUrqk1Mw7wjUWaju2j5jaFxSUMQUHMKB7FBAqjZ/aeawwWWKqMq1Mxc9oFt14wRzny
tvl1WlAEJzjDxL3ixkCEhPFAufhYRt5Iels0zZmpgM5ZJkSCrkB+W5+OgsjDF8IHILx6LR5d4LGw
t81VUo/SkorJrAAcGeIMC1v/+Kr5Voufyo6worsPVAlpWVEijzdwsS7EtmLcZE7QlV71IzkgF+9p
7knF3+2uAvmSOIqbM8P2Wpt0ZSqehpjJEIAq1gkF/ZrWTD7k5r4W6KsFyuml9ixS3Xi+r/mZBYdX
D9IqoYZF7VRQchIfQTKgVWf3VPohWV4CeWNHB00n6HoMmIx5JpzigelKdjxQXjxYnPK6QTEccjiN
2/RnQAj6ElwspfKrDl33UlIVXlf7l3oNgnImuSJvU3hKB51Kx8VdupoJl8Z1tGTaedBjXfOCs1XL
LakoUW2nwj0PZqqbw6qK5kO8hYx412BezCQbdeLahyuNGrduZXtmRy0W03Wp36DBOwlSnIXFnpc+
dSZlOfe9ifV6IE2iNQhnP9UAATTtwxBrgxqC8x8aYEbPXAfW3i5NP51Jk4h0SbIeZqxnVznP7JiH
x1Eckhk9p57/4XPqLOINHrkUZqKbHRbAnXBFkc/Tk2XuM5/0ya94rzJGr/TP0ejNSJnrm5E6juV0
l79GCvFDUQM57bXqkVvjnNPARws8pl0Q9rK+gzHobgq4gJk0NYoRXh9WRUTDGaXoKuy2cHon4u6S
BZjhthycolFb/LD0GxP7qzs0VIbp0JnPWdumquIn2Rnet8zu1xVlRGd5yChWz/9DNePcT9K6GnoT
gt8xlc3geGdNXzstbfe+RC24tpXO4Hf+828agvcZzrb6jfq0CsihJebCHRlObyeG16oQe6HuB5i3
BnzW3vEa0mO+TaTUgYbkhfWF6VBYMB9qD9i7ri+RP7lJenNRV5e6oAmUoRH/elJyUP/KXDTXPtWp
eZKvBTZYdfmQ1DeTmfK0lTzX6Q66pnZ7qPr1VQQv5WiCKqqNCTwR1uerjgg35I5ahZ6AaI2gU0ZN
1/x3hSN5QjsbFqG7RWpijRWWmTbDlPvh81KkDAahocZZX3Ii2L5jPI+WVdWAwySlhs4NfwqEQ/Gp
kfbSqwbV5mPPeYbaoMfhYXUWd9aRVSSNlaY3lcpqdL4rCRrkCh/+dQeO0V2OQUqZMn0s/ZJWZsjw
cDFcaF8YKRg4R5EqPfg6UOd7f1GKvIcpl2X+Mfa+uA08RX5MToiQAbyDkW9qBJnqgdlASozZo/fm
bcUUwwuLMmM2txb7st5hmk9g/o2o37dyU7E6459mkrRAjRMn5pRI8UGrh/9LxM1NrfT2SK9vvtRw
KkaCps5Ce/NS7XU9pWhsNGxyggKg2sGr8gqhgeFJno+EmmUA4C76QgPrXLs562iEJYQB3QsJyWCY
Cyf0cOUuuk+3rUb3KUa3E4KzdujRUAu6w6s6omsUsfx05pqtrnBdGG/hRGVSeRRhh0wTqQPlHBKH
5iaEkmt4sR6JeTgBSQTpHErhVn4omaquvG5nTszVc+GibUeY5LGlT0NMKS42XzU7aIFLRI+mZBxC
TscaQWcEiunXdOUjU4e3aIpm4e/yHkBs9YovSKqXRIBp3Yp//XECM2ROGjUE/5pnDhRvvRAjjtRi
pMd428zxn+dnBVT8CqncxhzVsKNrOIV4Ur/5kg0eORdTjuCWo4HvUDIun4DNfwa1kCTw4a4fx5SQ
VxTJOXol3SUM4FJ5Wo/4u2whPnc9Kimeo2CKkGeTp6PTCRBzwz9QMozdFBi5qFmNuZqdJLg01VSi
eQ4S2G1pzlfssC4KlxFkBd10kvsFUugxaUIkKpclLvUhTefwFbhB/LhFCclf5BnwS3vhWBtlJg3m
h7F09UpIH8I7RocoBl+Q6KgaQU+Swq7JX3pargsZvu2igvL1CXEAyQIQLxfTOY3H/zOPu05yJGLx
aAqy551ERyhUQBTrLoLMKSd8UdOYqXfQsgT+ZKQRBYTDHPKzHaB1olNy1lWIeiBUTD9hZ26XUrIV
EamLBbSMrjbaO+zBZrLbu/hvTIL9OddCtTz7t1BuKUeZMH5aGpmxZhkl7WFhEKe+WJ9baAMl/Zjg
+vkWD2LmE5xu951fhGI1oI1Jj1pSAlJYpeudqt0up02xyar3EKBKRxhJyVZHRw9kPRxt9Y7MXtJo
T3/2lZ5B/unuBb4cX2jcCT1D+144Uj1JfA67T1uy7oajBRqC2p6RMVY36B9+iRRvRrxBOEQ1nLqi
OHftOno507kbqgYikT/jISvJoFbU33NAEKPKo/z12ko+H9bsWrudZApcEv5LAmSxJMqUhf2tFVce
kurRZI+r+sFbwttyP+ECtJ+6cDGdOY0ZnVeoV3Y39E5GsXXf1IjE2/D3vulkvuZ0ESRT8kUtfSVY
1EsKKwDm2tsAfB/KoXs+HpIQvV2Ziz1JWVdzCZqTn7MU/BX56QjCvX/sepOTz7iepWcXmHP+/Wm0
d1HMFsbbIME4E3Wda/k+CHo8idBMxIodmq76IO3u+LqSLUUxZs9Ta5LNAJ3tkSaV/Q4GeB0lhDvc
MKqETf/V2FlTP5oRMWjs933pD0hKfQaS3HMYgdi6FXlUw2WUM1yTNcZ5NRNwh2uDMsThGmuaHVEE
3TAyCGNHlvNaJ5JfOfkjIarYaSniC6qGWQjjz2KUw8h7lR0JFUQbEuC8AofZ+1kA+7pGp6yL2I0p
l2p3zhEE8oEdTMDxTTwrQHlxAS5X7m+nwIBi8rEkpeojKl5jh1QsR8VwanYvliTSJZMxoD1scTay
BjdLyP/eD+1Kf1AoUR7MVg9gnHUUPA0XB/nWn2Jp7bVR1xDDFQ3AnzaoDlHSEjNrP6Iyq1Ejh+cH
reJqZtBf7MP/VYnp/0dE4WABuB2Z5n3/oZkCVAkjm2rYxhhCE5asGcCYanZpExwVN3xgYkb/YQFY
5skyY0+bmg/i+Eoqjy/RbzRzcysYQ5vXoSouhDO7izwyr7pbzgsHOt0Njhh2aos8W0aJ/Vmcd26r
gHVQVA2kMQjteccw8OGMC+BgRI18nEOG75ZTjVfWWuvPX3ZYJuHaVgJXJbmknpmXzONnjIrZj44R
taSIQeJg7mij/BLINaF+jB2y5C0xB/PgtR0dvteOC1/tqGnxbZdOU3GAmlqaLRFeRHksYZYm8yCY
U+Ge2SN83lSPh12I+qi8NIoleoiChwtcpQ9R6nbSrmwHV8191t5rb3QPBH3S6rfyxWjhYD34/rc7
8JjWb7hP4/7reHiAtsWXNG/YAlmfRxbMmIz33fLUQeYtz9Kmy2Ib6U8kxzcSPonvLlpp+upPpdrQ
/o6Ope/yZRVmSyoLP5P0KcZUzWjNhmIIP102OOd+ilkidZ8xSGigM6bYynRGI6VLsrmnHG813U+L
NlX6V5dM46A/5Ib93mkVM2bu6VlnMw9X5KYSZuNTJAtjtK4wmF6o4sgFYHKqsLhiQ2m1ARslxSZV
Szu19fqnbZ9MrLB6znDDBDELvZYtH019iXLdK5jIWToyKrM+jE7g7liYPfm0IEZRv9NJ1CIj7s07
gmVmboNhlK46NXokjVCGoXzD6hTrk74jNlRSGUIYMFxf9mBurLeMeySURvVIqV0TD5gyF7lPXPVp
m1RQ9RgPe0dQq0xROcFmRkfva8Gva249QV6HmmNuzrjXGpxufYs6iAAFc/SGLqFnuL68/1aE7g2Y
V8HQAnf4sHAo6Jmm0ZqVqy2PAwQyoywJWLg7NPvbWP+2X42ZfZHsk30IjK9sSLYbC4AnCrlbKxpq
zaX4E32YzY/Np2vIk87Q6v8tm2kJL7hqqfYtoARxu8MzjcntLxbUtrRPtq73RGFbrsVYnCICTFOX
Zjlc1foIyZWFeqcCjZ31uqcmJbinEakx94ekW55TwHJcoe20CQYL4lxdjdWI3uMN/mLQPhSw7vsS
iqzZifVO94+KFzzwWv5yjjfcPvVkj4BsmHFmYMlbK65ys7gfy3qO3lp6db1kvE+MA7cBEqiorFsg
oHrUSA0QdmJQsWKaHaGYnjDhsq1eR+W4k4bkvACLJ1xzYbWb4uiiSQI76gxVsCKsOsQDEZegk9uV
Ci4ELgY+W6df+4c+llthXUkbW8tSE3S8AxOFAjWdFFdt0uTjAA41HIsK0/hOocY+QIztq9mc3DdO
XDkR7cQxrxpgQcQ0pVgNRk34AAPSgCqbWn3FWm5vR235W6kT0cGzEpPfOZ2BEAAZqqTDUtDicfcj
reDLaJglXsQy2Xra1WYyCByZFpJHMPTAAmULevKomkrBWiEoK7ciXfKnf6BYM51n76dWj5tdM7IC
RBs2TO1SWgQIBu3Jboxs/3bC5dVFtt3g8GsOxtO0kVIn/1mNfLWZU++Egcjh1f5ggb20tJJD/7HN
8pcFqrtfGoUO4jB0Zq5lUDhmrWTDdFtL/lYT86b0ngO6AFYQ+T1LTLwH2vBrt5gf2mbGqsraE6+e
Q6KD+ZOljT2q0HbNb7YmQ8egiyZtWOijoHbACHg1qUbqCBD9NhjlBegXdr3xY4IuRPiXykI2h+7U
+GHgRq3iKw3Xr/pAgAWEFbDHS8psrh+S2TVoEYZIPRNSE67PzXbZmAwDlkhU5PObFjtyA7w6UHpJ
5V6CXuEGQ0XVmwLYk2slKfng32wHMgwFwl5qt2YiYyt7DhJn3m9HSmm58ZQkm4ARkLkIpC2GrE/7
Vjl3nEgAhGXFECpGz0nP21/JNG4o6l6zUSj/d6Z44cQ/gBd5VpKNLJ5itnhcDzgKVg8KOaYv37ay
ImSGUWkjMqirUiwLMauZFYsibSDcqKMk9ndCtktEAQK7vaYDmvmDKT8vtJhvcfnvY2DqbhgxceMM
zctfrmK6PN0K+NjqIwY+VWWBXJmJjVFP/55kheS9v2GtutgRlcvvm5XtsS/ESyT/5xhHPymEwwQe
jeTYXAMkmKCp27UUsRQHY4tXqL/cFJGhgVuQjN1jStZz7uyVBnif39jkHUmj8Z0Mkpq3vfGB69R2
S2tZQeUfpqInEhEuvfdjTGgc7VFzMLE+sISjcGeiZFJE2tqsb+Oe2jYAOTXBpl2EYDLHHT5A7QL2
Cvhk6vBzZNnLsyZD3LHBwef+7ZMRvZWcrvms6tKT2WHMK3xVXhnBX0CcXKSoaVjlEEKFvo1Gxvbj
e6Pxyx8tFW8daploNRvIBXukV+b1+FViaWcU2h9U1ljJ33ConMmjAJ/vTyEgjzBytbIHCKoEGkPx
+SZZuNoZhvHGRlcjOw5qEuQZYS1MF2H4lmUoFuWjW/iXpDl6PqVmeQGJO/YiNXA12lqgXmz0a+EL
wRwLG2qAxlKarScpA1poAOZkKLIoVXRc5FvtfKtMetbx+81eKRqt2IxlxyB18LThZqwSf8ygqtxK
aB8DSxhLCU6g439OfGcIK4OKHKeow9HT12ej55BNTrIjXnnZ+HG+tg8WfeQ+ShJxFeZunR0ImoKR
ShM3J+E9KJvg5l/zgEW44J8Isg2pKmzayr1b1olulkLBswgiYTqdWxrx2mEYP81OaG48LU2Y8F+7
pXnniGJyEj3CzOjQnTrkpqi4u84EDLenwZ80v1+BT/cCmfc4g7bH2sGu2qmeslu6s2bVTJUmKbwG
1JPtYjVaxQNo2mgTTaX23YlNvyveDa4e4h9gVJGx+rQCINR1JcVO4XMYallCMxnuMr69vbAd4Epv
ZDvHIE0Ef6RQzcxIHQe4LPPuXurbGOCJODBT1Hj+dFixiKMy8lggtV7WSROQpVTlyAX9akfnjfm+
QlYTKaySorb0XAo6kIYsthl1e3lp7RBLrMvuC3NqRtHSbjN9IVcaMlMGVp6vljO54f0tZvmFYxdg
dwlu8foDwW3673T6R4Ez+T11hBuj+hy2i2kooaGFQcG8HOwOVuUngi5LR8JPkBE9ABf6K4z8cmJp
XxLevXl6JwxC+hPcB14IbUm4/pdUgaxju2eznMS5SGr/L4gV27Oqxn84Ixyin27GYa3tKuPtFjGC
ulM03/Obu/6Wd6Xzzm/6GIQkpxlSnWWUiC1sCQXbn8nZP2G13xzHuIqR/CGFnHnS/hjeRd+e5mQk
UVuZhQjCzdrZnwXetBAA5s909MZKDKqGp2Z1jBvotsVMrXiSnspWg+lVzMUdEfMQnpwJ/2eYHnYv
Kr0EK/OSjEpyJaHDEGDtT4/wt0YJKBSG9FZwARQfNgzFg7frFyLIgBQE0elOnL/TkJ3b6a5zkEmK
/Jv95udhLDJM0p+UyCNzl5vJE+j4+uv+EZ0BmhfpXXMBbLvmGidcZWTY78hdMAs7Y41Rk3RDn9Xb
QnUwXGf97zpgEp1sSeGIVP2aDBuHLb3ZWRa79Eb2Pscq/letCuX+wojHuRQTajaOU2JYEwcqZidL
GsdXPegnkCVh1Upi6rsySTASkvKggSHYm/I+A8QWOu9M0KEsqXk8eGxpBKkWCJESs4pq4prGRPEq
Ci89WUaSQ+H0shODj1wDGgn4qg9alCvPCXJoZ2V4H8mQ1X4QjCyw6h7guga9GG5pxdc/pw562dzP
vz8LJwG4hXqA6UyZMZjK4UrFDxdlZmcM2AozFHtu9G2jpHB5UqHixy3q26b4CKBhGs9OZDAaJFd9
SJMNq3pH5bkUHrbmHpOavskWwB6b5w+bbmyUFSzmsLVPiihb9Fm4ikIgyxKS2IimZvsQnClITZcR
jOuiJ79b1fOewQxiy3VrOM2Dv++9Wlj7Pn+V81nHeatB2Bezc+WV0/RNDJr2sO2Dno84/Ln8nAkT
cM34gkqGwKlngy+wAKuc0IoiDg264hkMu9fkGWEN3FO903r9cXs7bK/TNLuyA1O3tvEMcEnWSNob
oP4sf8WppN8GQqM+75qwGlsugSrw9VHbo62cSvBsVQlBBNDSwB8YcmQsqM9Bz25ZmcwuWAsDFMcC
DctTz9tzb2QH1ZcimDBg3m6nfKontzLdeGTlL1/bMVtd6rAoEJHHhDH0WsuO2AAJ/ycO2uI9JCxL
PDhiqes2o4VODNKErsELKpvEpr+TKVpD5MDZa81qRnS1pXxzX+PtcCgGgDMq7B3U6Bi6UxCY8cCX
3CBnLnmyDTyQFc2rWehUHLAPEbYihywlmXho713ZS2fzTAtj2BESsRr1Ce6AHm1Axq6dOg3t2Ixz
wxjEdB7ipfpeZMZJrN46mVGEWKKSaHQXraayvoyIwg6X5ZF00Z4jn6iIZ1o79XMQTZc/084wgDE5
HmkMTv256gjhiR6N0OIb2pKpFAVpk9+tk9eNSCIWhMl90WEVp11wmjDA5cj+g9DTSZTsZqKBLeUi
qrZWNYprXW3do9cxA/NLhUxHIjVFL8mvhRX6zHcqmhDBTOm/pfYBUeDkzaY9dhL1lZS2SD/eLrfx
SRl1GDsW5nKuUvxRCY2LVxHKJbT/5nB/NJbweftZv4ebHUe2zgijWNLWFZUf2frlMC5dV+QArxkh
sk3mcBwOobfIb8anBX6o2WdL/LWBH8P497awnoJ4Z76iuCdhtOVP4a7cpvlOmdnowplE0VzTg9ZO
bbWTYaC6BBe9iIzu5+z/6474KcztpoZ/T/h1PmA4TwDLU0AGzvgek9XPA98qdEg8PwDREA/rweAH
rwHRV4Eg3hyecZN6DZC5fp3MsRKpG9aNUU8dbomo+S+H1vHiUTpqk97h/ChniNSSJYnQkkDOOYVK
zusDTk3+m9kvJxGbY8xVob55NSVAQ1uFEbUWv1Wm61ArBQNFmXyMjOohouY3YFRtBlSiOvuE6/EX
wU3CBCKkVXxQbQtnFQYFxml0e00v94+odJ2ykuQoOfNMYqkGvoExv5MCuyYZq/UNsWPdSuvd/jTl
WqfzNSdsokJf1d2IAL3T5O9QkG5C0rVOuTBchHsDP5Sg3BxfSTXcbOjfPCDdbi3rcmicYos2nUVN
Z6GgNqH+PJ7ZvbDy4x639IAwYmQ/tlwIWJFHJ4+2933D9g76ALPmOcbt/JCBG1W4t+zVemtGc3ki
M7DLwhKM+5d3lrDi4kIFnuc2oCtXtf89E0AoaiyEJWLK7Ldh0JIXxVpTeuDIF9f9KEnQVlr4vLiM
RYbtNSPN/CjPUrc2QT1js6FTISPHz0ulH3stwuvZzfGQpxO6HSkDHkT0jl2XF30S34GAfARU5I5t
kyU+QStGfhnAo5fbi288Pyzy/S9MmXsYpi3c0nmdd1/KcDAVYwFrW6KPYUUHYOGIKC9rAF8C/ZOp
UeqxBQUagf5RRBqMGFLfhT74zXMGbkQuNoCT4s9/5Y5gjTjrBuCp5o3CV6yDbxRgjaAO83UVSy42
eeaP640pWcDGEIyCzGa5tCqlikar2YStNrzL3BNGDcBlFUa96pAOcbK8nsKvtO4PscTazslhEu5w
YFYUTaQh8OLkzcu/FSNIr2H811UHyqmEW/IOg01AR6LTo3GpA9W8FFXOMx/8WxjUkQMwnoXTZ7Uo
Jrrx8a0ifDso06cjQIrgrFhzILtUc0yyETl5/s3Okmd1jwV2vI/ZWb0Nb6p+2sPaB/Pl8eVymkm5
B5KqsvY1nhf2VB7Sq8jFlTWYCFZWjLU+DLNGpeqRTGT0DM9AoxCaG0ySBX1cKxfE8OswQlo84Vii
QeaTDCwf09oVgpvzjc5j6rUZcIS5nMjsichSjLs+gLwo6VNP1v0uJ7JPVqiK6LIYqTi/r4xj/FVn
8qZbquGnhhgnmcT26HGzIeWK2SKs0q0WTTGtlDfLgyektMFSTdBuh5XQz14jkNCzS1Iq4QYLCtqg
8XxMjkfUHB/aNslJjaWuhotA/58A2QgigXd1C0i8389LU+krcNzHTEa4wLdBVjAN1UDrWLgrmMCS
2BGHo20+QANZ1w8X929+gLcZU5Q4Rnky9EhFJBQSPNkE9Dfy4OUIKAczGLK1pO/DUTqJ3PqqUFOM
4ABVqu1M+ySpg+rXEB8K47wZjPVSpJW5QENoO0q9TXT++gMmvgZK0Bp+90EG3xHxyz8f2Pvw9d5t
7YjypfH7Mfs7EIir1nAW0ILY9Jz3JZnd1MFW0+iRoy4TCah9vzk2PRycR8QIkq+44GDeMtUMWi8W
as7SL5ItBht2IJQjbAae/GCZlE/zm884kAFC+J99JNbS8MZMFU/INHlGhfXg6R07AvRG8Tei7bRr
tpHMazISDAdDTcZI1jKin1MRr4GqVMHrShuNd4PaW9PlXeJ/IfLAYyekWyMIE+VA8AVqnxazPlJY
xA2Ti4jFs9NMnjpcT/gz+kgvc2jylCLJzsDQ/eTqQxW4Gw2+4VHsWMoqu7kHtTDnQ48a59l7JyrD
bD6X2SqtKvl3tqf5EQdGOCksrr5m8nwKF+GKvYCfEgaSameaYEaCHelcuiH74taGpidGxPA0VrNI
/62bWNCkbwVT1J+P1oZEm0Zk1COd4vqu+mrJHszO1K5g+KR96snCzEGhT0zBaQTjBBZ0wVcddKCh
93oaLrGibqnVD8MzCIe3O0RQJbDPW+T6uas2fUAbphwA/ZZ30QOVstiTwsXPz4iiozsYvo0aYWB9
ZODANns8IWToL2ldTmx0hz92f2g2n+D+vy5iJ5eaMWRLDvxFo8I3fjTutBD9vG/wiRTby78yrDIG
+ZSrNrmlJ6LMSdqg0VlIoXGZWW1vPvBeNa3rc583nZooyAQE77Ho94u5CroOhxXNxHmB4rpk9Cwy
qT6cG6ne4U3LqvdaUjTBmwRhoDfKNjPNuGDTpPomoeyE5/HVQpYC4QrBR/h66LlqwxAWcMsiitKD
S20412CdAbzFPuW9c4xKQBgJk/F+pbOZSsIW0Wk7HAyOlO36AEnq/RlDyPQ1K2pPuAmmHqFr6XNW
wgpH9FKpI5Lf1Kr8W7ZLq50mcuj1kdo+6UBfrabJ2TtHzPAhAChUEpNHSPysdRiM1Z/KaURdUlLo
SyqCfDxkkdOUWJAt7fHTuhhiUZ/cRa599LpJG+S7NuhUS8ATWSaichE8jjTa+3/Uy96hPF4ewvp3
g3dU0Cx0rFja4jtl4vbJbxItpPrU6rtiZgxCzUPIpbDwChMPf69/IwASFe75BrN3H/SGxVM7KWLD
qBzY5xFzxJqv3OWw9xJ7xyhVK8Doyw57XS4Ps2cXMvuNKtDN9ZmXJ1IyRKCllDifhHDhAji5jB65
gGnRQ54h0Cuo04Mxg1v/OGlxMnau6HLBqYSStUH2ZML1tRyJVEy+u11v84GkIgAzei8EqGWGkUcG
1Yxq56gPfPb6hQ1X/fXezjhuGT4Z6LuwGvzZt3WNRSqM4jiaygb4j/4oBfo/Y/KIq9q/7Ja6K1CE
deemqaEVGTsXJTkZA20j3wcaDQ9ImtLJ4kMkum8XCk4t6RsChkXO5pNWa+5MR6Nn+NAtKlI1oodk
ubExmoMTqK5AxywFh1IA4Ujyxnj8IyeE9/+yr5+98/yR2fTEpewTvNnt76SpodmQ/bF+CoGW9tNP
Gsr4UgzzqwIOe+d7ArHFmV4Qqwr3f1XigPStIaCE9hRYjdkp3bPoZ9sdrTioiEiFHMBv7A7qS9mF
oyo4M4FT9F7y/Cp04ENJElXXbfBzaKdc8B/zb7GT1dZ46e83weBTRW9jxmlWJqfUktoTZX0cbHJ+
vgrt5WSdN51zMac371IA2l3b01DOY7c/R8CDDSZvYmMc1gD/y6Mv4OV8gkYBRUjTFrGjTULK94CL
X0jZWaXvH/Xpk02yBdbig5oFF0dai7zx0Tg0vKpTdcVXQxj5iVxDG8Nz3+GFl70j2KYMUGBNEW5h
xOltJOaf1AdOKfSA78ZAdS8Q8N3gnvs/xSdeedNkAEPh2ZyGhjNks3jz6j9M40MzrzZYo4KtqBM6
ZJ/w3j+EDlp+3b6P5EhSSvrZa5ySi5qre5Qi4vMKf+mA0LbK/xV5OWUYZw61Is3Ng2OtZ2+8oicJ
7eatKHxOC7/4NIi0ziqSA1Q2DuhgUL2nrFb3n+Ja5VkkcmLaguwe6ibS6BJ4N9vvUGPnw6DqFLSM
JRm/vNh/T2Tn3PdL/E/raHeoEwiPb4bH9RTpqaDJ5PSdx0QdIsCanFFnmhvad7edeEbBZ8yU93zJ
C/pI+VqeHKu6TrE/M1pm8imRnNEDd1c1XNER1NR1hvepS+IkYYzsig58/ObXkAzrVo1mtle9zIEQ
KKZ1z/3aNZ+COzUqmF9imBLRWsousMhsGJ/tZk9+Xlr9ys9J6uJRf2PZE8LHLY48y+riIWnkRq1d
O3T5jpMtt2TfkJvyQcE/cI5344GfluPBmnV4MEgN9FDI9Q/S2umFykfuqpev1gqCzDzMyI1z3ZEN
fT4SKFkntR2y5Af5O9oa7Td5xwKXzK7e8T5VzLvq6JUfFTMslkog3tTbFIZqC0Jt2jyM5amBpN1Q
X6XLf/bqgP0NzIRSrb8XEbVGb95LDFS+kkStBWtEiDoC/uP5g6pa8VCKPqsCFEVs/JS0ESP9lqGy
7MM3ysFM9/eZjshuwR7F7cxNeJUakYMc2Xq8X9ZladmUD5jgUfugtsoFr/exWBO75j/c3Hg7S/e6
eGC1Xc9+07g1McIAeOeSSYxZncQ9JHqbSbXSe1xeTw/nGi/kt5T+xwjn0FEcVz6P1q7r3D1JleeR
5z4gTwrNaddZQPyacDzSF6fZQkGRS8XYsTfR3h+suDij8x3rJGIbBSzLq2LLc89jY7s/HiTaHw1E
tvyoeU3CTqP6bKV33JN7ASZmG0Ouksqnn5RUb6GG8Rj++vrewtj9sR+EZV51L+VmdlMGIXfjG0kC
M8eKHbvmvba2iv+RxBHp2arkXBzQzb0D7qP1QML80hoSUbQ+uZSNUWhRRl2OsEfMVb0l6Y4LxyNS
hvMniC9kyn4AmHHBn+Ky9Vt6105PvRwdqS6QpZGqRl8YurSr7BGrcwVhPLisnndNZqtN77sekwWn
u4nI/SFUWWjbsaN0Vjmw+VWdsAC/Ls01DInwwDFvzi50q6lPHnj1YPTMwD3tEuKc0AuGBkCnyHnl
xjP4tUVnsLjNSqKPbIEmKdDCxKDSTT1gJ2lYN5kThL8X860j2EHVOmA/jV2F3jEUuo1q80NsyTyq
7O/ykJ56j7XOi7l3Pv2UmNip6DKmberCXFUd/hZ///eBj/7uAmmK6rpZ/ZWkitzjEaOcHyD2fA8S
IrGh/EoLLV4vdxjsIrYgXn0UvUd2SwYszsLG86GPi0ef8O3c/c+oS7xdfw994xYa6oqSJxIoDhXB
V8L2hm0OQXflytGu80QP2whY56Yjt0qiQUaEU95RaVHGYlW9HFqXD/yNU3V58wXqV23T+v3oHxEd
cqRWnSWZhK8YUFZa5Lf+yljrpYYkyM/2vXdA/u7T+rd0yFobjMd7qnvVdU8VUSoNTm3rErqf2miY
aStG4FkNUINffntLaNE9onby+KnLRF+hPD96AB3ZNvcfvaQW74M19BUFN+h7kAXe7/Fi3jSw3ivd
Mgq+pmwNK5/08fZKeGEruiSkuGP8xe9i3MPZBexutqIe95l8lpoJbL9i4u6MWa3ww8o1xRSac8fM
1V5C6mTc9aaoB8iy8BYbRxqF+mLBwI3iY8iVHLEsSwDwcYVXS05PK9oyeSw+3FTyTIwnXn93oOvM
+cyZ+gbz0Dd3XEemB82XmTTir+ezXTaKCqY5WeH8VclDG+aGHb26wq1vGlX0c3M1syfehB3NOAE3
A32fcNDLx9+TyV44Duf3bh2q0uZJilJk9gykK585XQzg/6YDivYc4a0W4wknxInGWgDQ5eY//pNv
Upxo8w8AULWoTky1VyfdYgrKIQ/GJFLsEZZtSRnfRBTT4eKdWh4zxMInwKAONffehd6sIpabCibv
XpBrfhMuJDQCjmk8CUWYeUl1Kx7YbAX6oRfe/OGNhTldxOnqG3Sgzrcu/bfRBjhJZjBPZTgT/i3i
EvGDK3/mnitsxtrWherBKqOJ+ewFChPBSzlPGiv2wzgMouHEk4rMiOMWyKkHC+YB7O3gnN9uaXeR
3MSlCwIc3e/FoRoHnDHRt8vGaiyncOWhRrFXb3WmdwoCl7zhWsSjNDAw8JTYR+bfbEsGz9pxiH80
s0Mplwbwmzzj3MDxKIh2tmlM3nqwkwGlqLrn7WAxsSW0yIZtSxfGJQv2cK4FbAr4ve3dos7EUQ6W
ElwwYGZvse2p35kkU6vAQIoc5q1EcNo681x91V9y8UJwGLu8zM5Yyig/PWpGjCYtreYh7vpRA2LN
29uJCewe1P5gO7Q92wLyptSmO85pXGPh457Wd30qnFM8hxfNr5ZDVv+fOQFA56/ooxJxDh4C245U
HY9IC+l82B6AsuC4JFH/ru6NRT47RFedWHVftOW0pz6eJgoBSZBCJz+TO3jf1+9yhDMoPKYe7QR6
pVuqSpsyhk6SYMLrHqx4k6qIctSmvA2Jp/xbHQp2EAJzwyJOxdufknQHH3kpwrD8EQmnuYxCWnlU
cOn0XxwD7DbjdKCdG15fL3lzX6uAE1pl9P4lfKJYqum6JVhzxhvWAcEdphL5HyxtpCpC8igBSzYs
WaAFkI+R872jVfY2krAZdozPjiND8C+qUcM9i+NkkQ+k8ihRCw8Xo3sm3wfhgOTv40BhfeSFm+VI
L4Bpfhoo3aElfNtYfkwdtCVrl6CoX8gDUM1jJshy6gwjzorcwDPrIVNvnjSgZW/bZYazhG64WTMP
zfPSmpBNPWIWkHJA0vgRyzQzPWPvnTXfo/y7UPxmUugpFqz/7dcRP4i028TDyPrjkz1euJKscGcr
qEa2VTJTvsXSWI9kjtp55x+pWxTqkV8QEFegLMuoRKGN3lA6XSi9nrZhTbHDrF0uNFIxigXIWzVL
W5BrWkGUQtyzw2nciclNChQfgVg7lgWUoPbOoWf8ao5w3zfVQrdu+FHXJ2lBfIgj4QBt+LKGHLE2
luYew/x7RRhLut5AUy+Un1uEcs2UKiu1iclTrwLWPAKn/gA46jBGtZ8ik7r+g5F6I2khvXj24dvl
/mISnG/Hd6YqPFmlsSKHqJP6++1SJMDg3sN8ob0CCD6DFeAcTX0+4z1u/ZaX2w72Dr+80o1XxS1z
qtG4/eTJp72Nxv5qC0jFkj8o3r/viJewYGBGO+ubT5msPia2WTm66fdENqotLfZoSDdBXR+Cf4UF
4m/xFmQS6/wU6rh8Q17UY8zTXHgQP04F0QM4IfZXCzyQAtO85mjTQo499j/8VjZRBbbs6ZneEtJv
+Xj9EInHeRko62VRbO4vdq1Y7zBiMKDJtgIj1BzcV1DSlcWvBuvIUDnHKY4QQM1k8L716SOwHSxc
lMBABHRiqYb2DQb4XGmWrU3MZwlpFg0aCHkU4qPXC0y0HDILkRlTl0G5bb6jokJ42EJopSJs2Jrc
Wk+D1WfUBDktea4B6MJye1o4kNjxtDKCsw3BvqRE/PHGWQl0SwAT7qynSpGEfyYZ2oHwQIJeR142
HLNZCFFvHhsDqOWcjkZ7Z2omEvy2YOc0Q7GIHNWXMdmwPrkoo4LGCcAmCrLPyMDR4RI1dY+Kg14/
KO0H78VgTbLAPzy6oyTcPZspoZBHn3qFz3cpLrgEOM6iGxTZh7udp+EARtHkJIDtDjjvNlPdtpm7
z2DF7fod6sKJNdNjCK022jyjyjkZOwi6D7NpEaO0sNgtiE71aOZc+QY1NxGS3YVycrkgnTfewkQn
iGA8JGKGmOBmWDF6b/pubcoaVx2IwJzonyT6VY8fBcfTC2nDgycmblIxUKdM8sVvpvtKF8yagPGu
kFjxjkSoi8/pcsvXn1GiYEK8eV/C2dzWiL7SXU4JE/08m3JIG1yK7bfW2ivTCY1vHagIs7XM7MgS
ECHLA27jVkJYCXMKsy4dcM26uRMcvl4fT6Wvf0yBWH8jN+f6mpGuXvLu+FDIwtrDFHOEMh5SrF/M
2J6hfpESLw+LiN2e65FSWc+OdUgZIqGar2aCvoBl7ZytAAYi4yUZ05pIg/Q97OKzg8xSUieeg/Xl
B5zj6+ONLzUqlWydEUblN/FyBEtAZjvvT8yRoDhLeTx3dmEYXp1KcMYsfGiD1XKSWZGktIJWI/eC
KuB6G3MJ+rMEQIAKo1jGud7iua/9iJ89z4nI8McV5ertXdbAreaNAArexFMGDbKUrystYYvZG0CS
wHcCzUdCHUxz/oXPb8xExtufxexalVVVbUjD6PjvkDutwWtW4xJuK5tF8yvPKEwLiwncqqjK9xin
XIT/nYlUge3CBc+FDjRzmELxyFEZu/35kq4GtejrCuVp+ANLoWhDD6TGPwEUYqy8E0e1hbgycoKK
340OpQciX5zTdw4W84GozPle/qqRJZb6bVQbKre03PJE1coQ1zKOLqoUS86iFZyn0iOhk73Iu+5Q
7r62bri+53JtpzqjuGq+5DWCbSdG3E4ScShMTYVk895CoD2osLhsFfpcMWoWNWHUUnizhwDLLIB/
gC0e2lWKzfYg5oiK8C1EFiTheRzpeIFveDrPcP89VbjktQLDJH0sblM4iMun0NgjT0DaMhZ+FsuD
AzQ1te4omOyT0JsWwzZM0dpiFCRRieXYr7NbwlcdfcU3f0RIiEXqhF1xihe7jZWV7nJI83aJ1a+T
GkU9Rkhrr5YQwDj4Q0plMe+U7tvJqMCNJdIkomiweiJc1rd6jOToB3gsoOE56gA+N8CyX27XqQm3
21hIAuv8CARmA62DEtNZpaa9nlUw09vTY+ieMs0alB8BoNuTfOAoopKupZcPJCDVrBJuBAQhhIVg
6+4nQm2V16ooSqwTACjJswG66vP1zSzka/YIoCEkfV3vcHl3f/a/h4Cb0Wqgf9Z47XGibZTGB4Ex
+OEptQP051l6yd/EAjcM94qOIeTgXuUvn/QXRYU1jYriobRzvk6xqMl10NeKppqwekNNKmoFwuaa
OdD2wDSYNiKGrPXzZ+/g0OhlAGKMsSD+5wK1iR+JDBzCbzila4erhJE3KTbe3f3qRkBrVpFAchLQ
rxL3bGXN6NE0qGF64YWuxqLPmhStdwny9OJlmvtXBYn/3URqkzzmb455cGLL/4zcX7RbXP3I9LpG
Jdo4P3mYTwEO4kzreD73hLEhwMtfNaheDZlwhpI7w2ZTwhayfCtuxzBqU4BAKYMC39ZEZREaptPH
JSvQaQAsbId9taTzFvyAAsiqeo/bQO+xnrfpDhYuziJyLmz9voHFMEVS4G93CCnWlkVQwqNQ4ObG
MmQyS3kV2oXEaIPNiqmOYlkFRzwcyOdEqJXFIgfAVKcOxYRLvdOq6fcgfxvDrizUG85wl3t4538c
jK8q5Cs6gCBu+NcZM21p5rLFkbATibo551U5z0u8rKqLdH1bFbI2mAyl1JGmxtI86ycJeSB8zvVA
qxnlcdQsH8REPP76jELaYSbQJnH7KV4AqiSAaIKin3UTVE0kEO1oq9evp5upCVdhPCfTnO/4PDPT
8y0yWIO5Kgo3CCrNpXJj0FvOq6JExBN6L4a2VYmRBbF/KkrMezJ5H6+IqtgrNjCPVtJSz/y472cT
J86k7wEzHYl/F/o+h2XsYLe46aOCyzxWVEGqWY+O7CHFEDKK4ibs745ITRLz3tYBA19dSL0YRos3
fNY9P+DfLCR00ASwK87+4KgGuqHufdM5p4a0RPqZGlyz/9uX1LSyNOkqpyT1xB4Qd+7l48+DcGek
rkcrbUu8JSQISTJiZbSHvoNZvFRZYne312+8wT+xpPhyOwdHmcOipT1nMA2kQFDS/KY9jbYaNrH9
/dx6Pfp3SgJAh9H86lufs4lclObASxlpumC7S/3sbemk2ZbOGI7VX36b28fM86/9XUlOOU9kxEiJ
7AoAnDCm2GE6YWShWnS8Sc1T7pv7mu+3ebYCVTPGhUDbF4WpnMbcbfz9LERJIDCGrDf0wHgPhmAt
2cw9Dmzgu6HkiOhMD7s4iUogJNLRNQjBisvp1TzGLqnAKKgtC7WM34F+UTBo2XXndnzFK+tna7Xj
dX+JlTDoCT7Y8pBAdQv8TPTr7l8xPOLQ+solDogg38uWojy/LajIKPNdwxCJPqUBgjAjQTsLbPhs
CIF6IheRT80BCLEiMVA/zMWmMFiKUjJZ+G/NDJ6q3iSR+pSE13+tCZlqINYd7hEWc/4lYHA5j/hX
4J7ZDWMLp5wNJWBo3+o8IuX5Rm+/qtY1AMA4tkrjedbkQ5/kY5d5CiRL3wrBIg7OqJBqglqbmuVM
fG8ietmUB4UGdkaIiqxPGPSrHR6QlOdBqBM2K7nEOzeJ3HXMktx1+XyiORTe0QMpx4ZxrJf4zUEN
GKKkAClt7jlJmTUhS4GCQs3c5436ybo4/jZ5ruJZmdzKdu4eD9Fuy2bVikj+siaqLtzGoio54Qnw
llPXLTsdzSNHntLWkbUL/NzbcWRrr5bHtfeTwGGlSwchZZrSeLih/UvHKGMPs5fPPRht49BgnlhR
QT2OZuCSGCD2TxyqNHntbs+wmV+wTlw55n2YCR+krkjWv7Ix4LSIIkEDYv2VNUmoTMzcoqsJc/0i
6+zOJOYCAOD7ZOqeCBd58TyMWiwGujyhAlONg0eoQCN/5takuMUc2x2hcNN9IQDBgNx1+u6ewGb3
ga6beXuq6p7sFQDk6/8W7FvpCp3ADIjbPXsSEy3mRBeqavNGQMbqr9UiJyA4BrQjeD/dG2dA5wIT
c1v02XCx7WX8qQPI720Uzcas5mKtdhhFqGKl6E6koNCoFRn3zEIsUlez4zGn4Al6JbCiziO5yXKV
Dz0Ocs2X5tPL14L1Y4hjp+ltNMAQrLrPNAFj8GLlGh2gAf9Db5EXzia8b7r9Oytj+uuhtm7vYEBm
vEBNjiW7N9tkIcQWRZAjHqz4MleE08ZtQqQZz2sdpdY9DJboMr57vbwhlk3vfBGld1ID25i/6wM0
swRE/oIRA4LmhHTUkBbcFkjC3x3Mvn0IKuiG1Les99AcaQmJS9ugy/LilPl8Ybch1/NGs1ppSxNE
0h4Au4VkvB46HKH2T5kqK3PMhRppT3NLtK3ZH7cuERBKnTeKkh2j2alVnNvodKFcwF8qt1c92kvQ
pq9AErOtQdELYpy9UrHy5d87grAFNYE6i3ctL75Y2XF993yjNk7w6tR65OHsiWfwxvZJOZzwt3t2
g0xWajyBCQhR7sxwdbhDNsnzEm9PvCJZtKf0ZMhVAdsuTluoxs8CQe+n7SLz+uuIoAM//4nzQmHM
NGTCXz+nAW47IT9QB4inrKYQFGY6yXyqtb34A/A8wO1Dr7wfA/eZ7grM7oEiNaqWiDu5lhTrigNZ
Hdwh3O52nlXU3odLX5bAoFA/ETmjZDIOkOfcoO4y2hmVobo/6IP4e03N+g4em7HSrVxx8/UgNP0B
708xxH4Mr9OW/DwtLCwWX7OOhadvZmVWaECNJJ5kFw9Kzgyn2WjOrn0dYXHjhNsQj/64/26KAv6R
rGiOVKQ+lZb2MllJRbopivOZ0dAwmLsw/ado/OZALApWBbJpY+x1VCHg515d/iGltCMrc2Hax5wd
/iUh0a29JtB+YE6TgF1zqKjpTLerdfqElHDxUE7wXQbf1Pdd1ZI7mvukaDwtQX29+duNqDoWIMPo
FwqfjbFTS1DMBU89Ba3/AbILh4YzbfrH3wvfKDHvIrRf2xZE71dsns5vAr3YmTKIgj0hcpLVqM17
EvnXQl1a5Z/KtaG2UOjZNURUUonAE3zz/rfIwJ1Z3iHLgPARiu4Rhvg1NgtvlCs6lEce5HVNmTfB
fleClMPjDTKkuGUJy/JZUBcGd+ilboB5sGhYgHUl63fL7oAVwMnyi7o5rlDjXyNvxcjV3nxKiK3E
RAjJG8UIoDFxi3znJGsx1T23+/gU4/1vKF89gQ95+Qt1oB+KEv1kHMzKBy1iDUpUpzvsPj0j+ot5
E6pn+6wByK1zqtilmDOOFwWiv5wJGTOc1FQv+R1XWaJsjv71LAI/4gkk8v6Zi98CdLvmqmfC2jkN
pOZYOXKtsGQW1rDc7gp+hpVWWrO800TVM4oPuLGarC8ywmRbDDvy09qBIMCajhgW2c2LSZsc8onf
OyRDCuu6YM6JyW6zljEvL2pE+15GUy0vDbBsP6sEtiDBCcp86zc6ZjS/6RHLqd9M/NXYuKbjxMHa
dX1PJ7Dn1flfN7tvg38QFS5gFm0QL5khhceYb1gfgX03hxnNfiepp2r5OxZemLBzLM9jxr5yes/E
Ztes1t4y0ANiLP1WGWb4SPSeJf1MM6VCN3IRaohz+251K/7IaKK+CfnQw/mbJybR1zuKFxCLfkyC
ZEg7viX+LvbH9O7avr/FD3qEILe9bEZy1P6CSKuSkQhL87F1pGHUjK11zdMP2WrVP8ufybeBxQ4v
jnofdd55yWxbLlDUpADOs3Id7t+d14J9/QyjNmHDpljq8UNp/6KzvH9eRjjWw8iPvwXbrha4ytJu
NdF7Yl1stJkFMuPgqQLLicUv9Gc09AXJMdmIYLQDQO5otaQ5kYGBVLZ26oLPLtkgHPRO5SPCVpFD
5OrZVnptPMe5TEfDSwUVoiPjUMoCFh9Pd5QiZAw62Z6OQ1/kgpUWPuO1P5YqDToYEJkaFwNAirwV
l11QP6cCniCe2YeJ4sn/IgQ5G9aiz+olcmed/cIQp446ZRp0TOmdzxaYbaZTYKSYX1tiJF0kpfl2
FDNaFurVqgQ4Yql2y2lgjtS+PisdVWp960447sq4gWzFR1B7XCQNywV7yny6BVKSJ1ZVWBu5UFSa
al30mxsZ5/oUOdM1QxQMDCMGhlNs34gb8eMt8dptrNuXdEgxjc6k181x/Q5htoBnLTX30KJALHvs
anUwNYvVCGIbNJSrji3H9NNo8Ttzn1KoVs8gjf9x5dJe6gR2R5SPkro8VQ6GFukgxLjqKLSr4iwb
FSYgxC3Bn3Qby7uoHtdve42Q3XkLcG1YcoSRuSm8TRwuMpfH7M3VtdHA2OMoH6h/a7yPzTWtleNr
F435EEnBpVAgC51FLmpivhZwtXWXFIn+pUhevxhoouOvnJJrEsj0KINQ2w5Rnl3MVP1q/yUqx1FF
LsHrOU06VwFvgFtnHJwre0XnwvalEhFBsEhk8X00l6Z+2M3yHgCBlbs9hN7EEPY1sxqqYWyFCGPG
4mYTJjTMP2Fegv1ht4SSz0y1kMbRXx0KiBEVBIjvckXJT5zi6VinRarzmEHbShVkmUekuftmIGQH
y98bZjEientgFk5MZrHk8RZDJXkteM9paQm7tg2NhZPikCQSXCgiZsB9GvdBs0/txzq/PYoQQLuT
x/RDjMKbhH90FOUuSfHjRf87shtmKieoiAcXgjkg4Oan9ARLrebIkMuCLk1mQbzvGboOCefMJunm
YDBCDKUSo+/hHUGmpJRF3Ciewf2v+EpipkCaMUt7ZybfQo1/ebZ4VeqTnbtQORqAFh5THBh62HyN
FDuEhXRowjVfDJogCoSut/hi5QHFH8P8D1wKu7SGLdvbwBbY43ILO3/U25Kowe3jVeXHmVcvWN9s
+K0qTSDPOnq1igfxd85998VMxBXUF7HgL/p6XP5ok7rvzLS7ome+C/DhujD4pvELOeJKRlNxMLwQ
FlCjQRXK08A6LNHwcE205nqaShPf2XQ+ceeZzWieuKbu0xUDscs6RE6mfmoAEz2ZhuWJhK5z5QkG
tNem74P2bxW+ZvLSPfxZsuGYxFSAEf+N9UUNHlXqLgh48Nwua/wJhEsljebNmDIuMwhcAPq/3Msq
uIQmQChWYnjeqC4iApmUHTthKW4hPwlgVHNBCX+QtcVuE+19SAc+0al/dpJmNkTn0/2geSf6Z/Ln
03c3br+P0kxFgirn8DlT4/ij25CCjsxKvJxaSYM1Ezffw133qAhjjDRECOFWMedT12MpJk5MXjgO
dArYyrbIwFBk1OUAP4RfsuCzZfFbYPtOpqsn9qhIfpw3jsnPDeb0n431GyaMGF7Sw2KUEEWXplO5
pmHFkGWWdAdXeB8S4IrrY+KTVja93xXIRvET4lM8grHrwjKRX+MKueRjo3XXNvsYL5RuXNhZ+eS4
Wsb3H9Dn11jiwvPiCwNIStxMWjZbz3EDJgt0ud7fkICZ8cuq9EsmPkEeSXECSnDRrlgqpUc2jmQj
NfQz/kzCwSoNuuwkA1BorT46yMIm5jyNfwmhRJxYwBOqA26TpcuHAdPn6y0m433NgRTbB6Fnwx24
6D80/JoXrVLDwiRCwNYyISznHwKnfle5WD1xAcEti8H/qn2/cwr0l1/1fUV9KzRBVR9QutTOamcc
nKlR17ilTMeiajYY1vjlT0Mk6wNlEywSifty0ofbqHE/wHlqPkys71lLiWgRAKeiyZAccIjgvWXz
RBJiXqQLo9EqPFXGZjN/kWu4oaASP7U9DpKe2qpiUNtnIEqJKzJL1O5BuVxDvBmWUyN9/whcmJyS
jRYu7UaG7cZzsYir4YCJWlPEaHUZkryIV1owC2Nm1D4iCnQJEWNDzeezuM7lIHdvVsGwdcE7ELY4
MsWl3xvyu6zwjY2/pCglkStB5dgIkBkbf1w/S9GZ5qibhxt5gpXPupheJ/MkZgZhjEruJQ+oA9uB
DMb8nU01i5ajGWsOFFujOLdRBbqBRy1+kFFyHj003GCGqqHpfqdD/gEGNQn4B11a+UNEcrVf9sfB
PBvM0p0Odvv0z9SYXG61JbItgyRsxJGmtO4fWOSVJddVRFjH6mLlyN70+RigxOocgHCyTKX2Mdb+
wUHoX/YHqvjPO1Pi30Ct3eApHGhK614PLa5Udt14+EhbLHZA7ZPQ+VV+5I0OVz1+Qn76Bbumi3bj
kYf7LLKievkdnM5Itck3o7WJnry5MylmidH4U4NxFI4OaS+YkAga5WUircjAykXshHqg+khLlpMT
ySRhdr6Z36D5KqtrvYQjUsoVbdSovA9m4UKANqeFU3xd40egpdtSK3Zi6TMc/QB+MFs9O3337ITE
AQuHkvX31u8Kk2DlevI1ASCnEKVsvLNLYceWu5P/pQuOVT0HsD/1NO+WXCU+w8wwM6s+sy0cQI2+
XoTQvlMbThUxJNY5OesM6QzYIvGuNGefrQbhV1BCsPciny55ghbPyC+GmYOoWXs0u22S2y3hbBeE
yjt9e2Wjfr6zeK9ox1XLjK07WVqn897A384H5Mq5SkSVSP88iDpIdgQOHkyxXlX/sWa+8IASO9Ud
EJfAS2d8O9ZjW6gtqUr2qEs4GJw5Zb/NTO0TrE8VKai2TOXp+mIfofqmUCM1Fo1EuV4Ai1YGyQ9P
9y8HQa960zZ4NRtXRu3DYAx9Cq1jQEqaHyuT7atg/biUg4fDiiv9m5OaezWzJjzuFVFeFXGRBZad
LhyNuO2QdzIvOwofSIBq0UX4kAkLM3z2f7Xdj8i/viP9c0pOw9lEurbgMMURB+uW4atta3GxLFtV
52w1XJAJgMuOUSnWrmJSjjkGc6N5gyUlm8rImutfVwGWRXMT53YMvyFac3ZLZGmts9mQrDjkFlYu
N3/KkGsjdfVT3OghEDNTUyEw9ta7CFQqjl3VmoCEdmhDzrqoFtVfs4JeYpCFuioWBmToRLyIpvdY
3u62rLmVZBSCrkLnvMgpuN82uj1qFBqEF1RBhQrSh4Q317zrUoVgeFfUVeJP28P2SP7KIIaIHJH2
Pi0Tw1oiqDhUNufc54rqEJtPTOTbCUi79iE1Ll5uXBwIwayaXyiXYidhHgWxV7/VxcrI5+Tl08H1
RA+IQdJ4iwDwe4b1PUFiGqDZO0gbapEme95xHY7npU5Ta7c8gY7mh8htLDBt9bOFja/PUfvmII63
TqD2J7jSPson/MpEtmsCsBAYHYgffY3qvBRH5XmdSfH3AnY0BdAwQyX+1WS6n9om20EIxpiEdtAv
MTK5GJYTSD3JaPvIfNe3kwEUHUEAh0nHhDHe4uH13tB1XdC297rdRmpDO2sRu5xqy9AVY06bh1j+
6Dnupl3lRqW2AI8h2uxUpJ10h6d+DemaOxWuTtKOLhdVHPzqVC/OnU2c+OWruA14MYLV6ObhKuND
Piw9m9GrdnHyAFRij+xGlz0aSnU9rtZwubc3LlLYIRoQQB4uBWGmL0YiefH2VQK3Dnt13/XuPoMW
SQXMUNqk5qyUhEajNOanr5uIhgk3QO/xCoL0wUFHKWa5w9upzAzOsB904tBH6KPjzxa/whoM8AeD
PvRGYG5v6P47cwLgLm6vTF12dxx2xfQKw6kcop1K8Odb1Xh0WZhne1YJVubpUitm487/Ttl3O2EG
4tEif96DpisIJbdFmoR12acJhSBGYYJZNzm4Mb66ykz7SYvO3nP1mkPWREFA+4zer9OwBz4nDwH6
NM2JyhEnM4L4tjheVH5mh9m1pp/N8s6HvBHb2aqY5I66wD1AlBjE/ELY1bxkXDYIAHUh2HxwREJu
HJL6BQI63PCGKmY79RvuMrwBEKgKaTDe1GkymrxSGpA01zF6R9znSH5bAR3PcHBorVEyQn7waNDO
08OABej3I7SeDTC7MYEyLUU2xSQyDH3yhm72EJg83X6rVTTw8DErOfNOaD5vrClcxvQe7vLUJYEq
fnVQzRsLnSxtDKp1zeqxmDZ+GTyJ1iYzM+mBHZirM1sNSIBB9scOC9E7Av3EV9QxIgQHPKXLl+26
uwR3UFntIfwkxf8vdm+Q5wAqaZBkFY+JLlAiM12kCLY6YwFAPXfmblntRB15Ti31p5bAQPt/TETJ
ZCvnaAhcH4xWhe5MVr9afOayfPj0oeG8HGrUt3GjEQJrzWpcK4JuKV0vGYzJFZEBsiQf0H2U8VI6
rN1rdZyMWAvFZXplxEqdFAtoQUneZ2GKA+ut14KdSftqGSMGcSaIXj+0T5S0INNNMGSuBCp6BPbk
JFu28S2KQuylCMQ2+lQQL+r94B9T1lGkeRBV8IWfrcmkS2cXE74arK15Mt6lIzLw8gXERn4ksb6N
2XyFQ5VaK7F6/oBY864oZg8ha/+QuGq9c0LMyaVKO6H5AM1KR+4yYYzHv2pr4NMbxqz6O6FGnIKf
4JMPecnBpeoqOlYzKlDuJz9vB7cLqeCmbTuvgE1LdWtH7XLDm603RsAxF0ia7LtLrp/9ReAnSlAq
eKZ4DmKgA4myeXRZucZfg+IAT6Pdre0hFhy53xXF1MDvF0urY4AzmNH+HMcLnXtw7rkDlOquXJzb
YURQVuM9WxuuEVtkNsDE48I6k6LeJ9HVzhsXR8FVwgBk4Qni4Z/fPuaWB/YjsMX9JLRtEcu1F1QO
uof7sRUCBal1w5W2xf5jn/0usm2a9jh5sjSomRHUeFO+7ANF5zd7+GEo/pSo3gvNrxHYYFvgcTOo
ZocQbzTOk8fol+8KFocAwgdnbsLbMT9FTdofcFAm+pcj0DyBd7tVomxKzcyp7FvNcGTRSozCn15W
Y4QdKUYoYLM5Wv3+bETRodRWTcXVZ8hJwqBdc+tjSsfLhHFecleJi3sQ/mfzA9N+q2hS2ZiOKMBK
svKWSRj7IQL67W5vOwUzFoQ5BVThD+La7cNqAEZGPHzTNReJRs2yruWyNuL2I5oz8O9wqJx/Cv0W
gJDBAdHjkzCNZjiSWXFoxTc1fzlGIdywHu6gqOdJGP78liKMsdwJZoraZjq8ck/zZAGtDOMHfxGJ
MXSce53uPKYA+FlnbybZ2ruRvtUoqiNS6/rc527sTljRpZhXVIJPqzE0W+Qn+8IeoDqBCya2nLt8
Rs2EAHD8EMlOMO3t4aOH4JIcH0zm9DlfV+qOVdnpEh1+UrTwYLyvOqYZUv1zIzy1wRMi5I7citio
h+utj43+2RcK5GYiRdiD4jUhg4eF6wvMMdV0UqmliJL5scaumAoLWREfR4YvcP3FHckw6TKHeofF
ffNcAYyg2gy9sG+maBhz/Nd36paLGhEUKmbV0gdcfB5LSfwzkLty7O0StJAugp/XD5bPr8KgP8v3
TvWCyyLpIaB7u5Uhe7SXtiTFvMUWKAiOSFH00Q5M1sdNjGWwlfuK8txQPY8mmE6foAYOk0/SrdQa
SspUk+CXk6vGR/F2h/lImajuQ5n4EGOMc0MUh0tBPdH8RcuHhAKNReQ26rER16qwylucu0MKP0Je
5OubfEKbHmmJOXosP/nVq7md4P5WIbRTwrDl6ZvkCUb/fsmpUrX91uxZlYCSv2PqAfZadNxxT9jp
azkgiKcB0nAQvqDKO+jkyT0yovxHIZe6PRvyo6rLs3pwcBSgRWflbuUOvXOUPl3Qnir1+vPlb5VF
CcegmaJhWh8HED91zdqRVhwoAx79QzKZNfU8cnDZaWcIFq/7ZsLcJDCIJw/BEeRrUi8nFHlyDnai
QWkbgC9bBiLihVl+7NjiRJTIM8u9xnAWLkHQdOJdRDxjPAmS7Qn6oF+Ywj2a07SdPwNCjqfFxvT2
ml731lrD2V0CV4MWTl2k2/MVFAK5+B9lHB+0UjDRhjrwYf6RRKiaVpCe1WS2FevMUowjRCmvJVMF
qiejz4f9Pbq6F0Hnf3qv5aNuWyW7EyP5llVWG+lwxEXyFYAwdRwdM1ZTJ0lsB2RwclOYDt47B3nH
T5rLW+DyLtlBEGm/Src4asQ+AG+ugbyPMyA8w2Fizu+lGS3Eo6TDByCsQUpUjyCZsbq8WmrFYNf9
gpUdBwlJZc2yb2mPAzzBjBWt0PolaK+/Goi3EdDyYgzV98SsQQi5+DJJVC6N9P6fomYgr5VRmxS2
H4g31F0QFGrIFyVTt75M2jCLoCb+MWmDmXBlKgpYVZ42SKhvzSOVjOwlMpu3rNWU+GzB9HZqaERU
rs7iTDMOlmaTjlLZ2nOmZ/neMb5Ge9aV3WANQ/xHDOkIyukAqYxAr7qvhH/dGoeFXuyajbjE89G6
d5MSxBKwys/WNVMicy0b32Mq5Xm+u+c1nkmtAl/M/d+tO9uVAUGMl/draGRzktT1oL6An7GMiOJl
QwyjP4qvnjvFR15RO9ZI7tMm5U8zOJpGn6Rs2bphbI301sCQg+WbisaDvf3jhihnqU91WvuiA7SU
ianfYFCowQV12kITlfyO7ki7CJrFfJ89lBZq5y666xZGoGMaWbnVOj4PmBQ+w7VKuT/v/WSZscnG
Bv/U1noYKhih0lUx3rHJzaAzKheU+BDJEhVc7lND7US6BwyusMOv2KMEA78WOWfh3FQqvSm9jg13
k9fNrK9tXu21GYjzHmCRsM3mY7f9g6mXIxA8OaSiNXU2mujYLJms4bJ4HNuNSikVY8lMSzEZCqJ3
+ozIkbaAtyjo+Fo71QkJqxjM0xRAgEOZzPte/t7loR7MUULcyyMmpSftYSk+kLE9VXGGGOpeZZth
AZVHGArC2pL00KIJnFJAMUrt/QClRTghds56fr00nkgHZtmhBFz9Sx65w0S8GwqdmJ8i7PmcxiSj
dd4onAsa18hbZ2lq01oLyBCkJqeOULD8Q/HDZkjfQr5k8oO+VegW2EMBJL5HKAJUYNU/y4e+FVX5
cWoNx2qjHDcMt35rJA3AkbH2+9T4OVfNBB1+swvvj/DKAu/twOLrEfGPmVxzpAcO3auQtASdojNT
8pFfUi38hteyV6ELkZpHtZhtfUacX0JHzcm2GFSxUiM6VjbdHAGx+1i9wI0lIYq9aW8zqEKVdB27
5xNr20qiWxOsTEcgxsKuEykUKKs5KQ2erxdFn2u2Fqj9v0neyLiCyHCWFNSHE7It4ivkd1xXqJXe
tEyIWS8HHFPupP1LRhi2XWyCU86rquLVU0X1/OLd4sV/lgZVYAW3vNf3FX46vcYGdtlYGmChAkAS
9yEezMlgKUoHGP0TBB6/6Csi+He07JosyZoSDkiOM1maccnowEU6bhFUnouwvulWX3gEks3zS3so
G8Lp8AZufb4C2u1XCfuEWKD3HvDb+2Ao6rHy2IAKdiPYMUQcz8cLGQSpcs+9ZPw/fXFHAdWahBw+
nfL7ZdLy2KGsEjjRmta3lJ5bKvG9FGx8QXjIK3ACdpTXziOyRYvCUFr5GQvh0lu07hFduAaN157G
KxHmaDr5d54MlMI/WCpOSzuoDWesgXCWZUPxG/3x3o44bagoc6Qq+PGTfcCuqwmyuKCIBFIoz2QL
Y8LaFmK7Vn50151b7+fCGtmvX1/L64Wz2TLWnMtbZhrLdZPiUznFoA62o9zTLrVRUvFhcEDze/9M
QtiIdzb+TOndgxRcMo5WgAOySLRDxW1ZbYto6nEw3rnDaP8cDofeet4uW0ZYYFoIrY/Qb8+bhhh3
dVVxHET9myb12H8uq6Vyz7NoV0JpSxxWKiZqbD/rq7TeUefxLRuJwYUuQ0vNoubJbnvwpp3skVRv
Eg1c4dEvHCGLba9i/efMNj/aS40v4Xikx1IKcwqRLWp9kYSE78ei7LdpFdylii0/ZFlTxrK971Ps
VrxIAJOPdez6+TwIuM5gV+/BMl6dxCXclwlBlYXXp5CNWdK1CYFbHKpEbzyV5oAJ3h3hVFJPVgas
YEJ2vrn1x+hUQjsTCcelY/PyE2NRjGIhjA2hD8tc5qTML39541H06Z40BkvlzhW5Y5QC4EyFAsQk
zy1A3cwh0u2wytnUP5TQ9BOat9ZyKyn+5S0apfygE1/RQvtJx9bk+OUcfq7rV7uksOZ5Km9YD6N7
KcrEhFVA7aNzI4xyBbyLed7t5sW1C6pWxUq/2jfu9eC9+69unuvcbpZ9V+HzFf6PnVIikdKx90Y2
S6SiAlgmWv+Es4cP5swLS1JWgFsvKWNnREtL1ZyT9W67WkE8+L2hJm2K9W4XYTmQ9eFW4YYdcvk2
SyLggYkLxDYoidZ482SspCgBbJzGWdEDSOH2W4PDN0RBXfUCHbhI57fgjUrL3H0fKcwqydonuEf5
djxbk1kxs2VtbbIBTiOKjR+ai9nLGPWX5FQaDnruHWMG4eIUarKfnBbWsVfXxg8RA6d83uOIThlQ
dHylFbn+KmUyBEiR8ciUnXHX6dFMZtjbwAwx65+nbc+rTiQeAxLypy5a8dy6SEumHnEis+DRkWLL
dkCUsFZW57cQxO2DMoqjnjVsC89WP+9qYI4oeRoyyCBiZdmp8e+xQotc6f77Rf8qoJ8O3r7t6Neu
0SSbRMTbij1UU21rJlVnbS/FOrmoj1kQGRseWfjerwNZgb7OFCoiGZKpzWlR0qgce1BnGTbpawuU
e6MQf2yXohURdGTOf7sg+FSshQHf2v02drTOHHvX/3cPs/Drwp3vXkzVKDbNCLw/eCoBX/D+GRRA
TC2jEFVPIDR6q5GEfLHNljhuMxWBVRn4d5YHgiMZVU9H9LPqzaNXKSY8GULBkiSKFSLGAcugep14
B5zSrHTl1Md2pMHpEqb1TzOg3yQP7uNpSebK2rIsyuc3AGvzYRDJPv1RF1Ey43jMpCqLCWr+eAoC
mc41diotxtzn6weeufFSdzt8tbJRw5k0GrX2w13TzRPxeKuBGaaFRNGVLiVoaJOLfuGW3iHdJDqC
kF/sPZDjj45UVQfOxFniSK8KTlWjXbZ7cV2gR61CF0vK5xWsLbM2ip/KUmYkp3A62274ntexigS0
t2Eho992n94knP4iR+Y0h5exsniyk4gXFRsuoywGh5VH0hc3B4aY04JRlpdc8bD9ysW5vvl3N9JA
m5DMqCzPAQm3v62egN/Mcj4C8y/QP7UUVnEC5vQ4K5bQZrqIZrApcv20W4ISv09dkCLXyFfB52Qi
Del2cuN3w+GjrSS9gP2BnH5/nV5g2AeZpK1Wa/Fvw7MIP1EBdB9vgqezGcM11I0oNoBxq7DgqotQ
qXl3F1T+0oLMiAGfC1hrwSQ9vImrLsM16DBVnSfAuk3aVUP0CfYqtP1bnTI3M1BbPRzrP9KutfrZ
7os23JudayXyP7kfDqdlErybydLgYPvPqnZ5e8w11z2S/LoQIOuAF8F4j4vyfx+mMqC2zz3c6mR1
QQKI4+lOkqJvEaYFDSaXjDuzwBXHYKrXjJSNwnqW7RluyNC6cYrvD963iUeWRJ/Ev94a8zU+8bda
QOBd4WoYUWnfD05Xc3Q8uR8aQDSA2wzPN5QtsfV15n1/D1BnhO1k+UzhdFup+s8W2czg6sSczP1s
uZFLVhYfBETqyZmQ1cJG3xUXXv81KkQ7U66aNuhC4NXvsLA8rSZ1g+p+SugekR6+dFdmPkCyKxR5
jQQLZrJ/IegpOd41kRuwU/tSorp1xTajZLfpjLVMRylX8ReP3q4RSyXHzhQj6ZESw0dIcpNe9PEF
J6WQAE3vuavjkQtapQArYNlOZw42lriDTgwb5sS5fpAQ0aPj57Boc9Su8ROIP8aDJ95PRChXaBJT
0Tai4qNjUZ2cxgtbbk/LDsl0wG0izZtWJIN3YMXUeq2V0r/rWXGBifNdI3VpFc14rNy2e1RbG97U
ftNXnBBTlpFJrjhw23B6hDQnulyl9k0BBriqrUyGY2p3DchJSSFWEaXbX0kiNGHz/EEN9uiJK5Gb
NJiV6BvCawAus2zIo01lGfp+3dnf/Z6xfO4SF1ROsF1sBSVaU6lWV999dkOOecUQIzz3TUrf6fP0
+RQxBLaZQn3b62GYPc9YrW8d5r0O9Yl6/oAYe8voCymUkfSji44kpWu0jWo2t/mpKs2eMNsp0GVm
KR5bE01BkuJ9XJw1GAoKmt0ZBOzGuiHUfsfX27uM3cNLjrvc8jqEj/hbMB/6JLQwt30amUbhcoQr
d6nCR60qnIVLYDw5DpjTSk2Nu46Qm9BnymUS1LHAxImK++udelLM3WFnchehsCPzScHXXKkkH952
R+SM3rN5kRYD3SD9R3VKLw31LTrL/0rG0Hyw4zGovikaS30LWPW+XzRd35ksu5HL+LydkbmLJ0g4
JeGPcqIUP4DGwjAy30XkdPpvfL2rN111+4Y6/EMt8O7Ul0OiystWRS721n//EaQjaMOgnnq6A4EW
7tCwR7H+6gdwMNeQ1xqclkey77Mzdd4RaVWGDiOvBGCxA2vyJ0uKa/gVqUIngXbhwg+juPG72iMC
E5A83nNzBjSObHyhnRif2/6cHrjvyOtQ3VW98ok9cF0AwPLm21eautlG6HHu+ZluIvAdTsYiDCsT
ecNDnArNLIOcpiwyL1wN1bQ3uY20NULMfNpfMRac3nNXBNXVH9bhieGRirkwtRCu4DI/B7FAE+7w
hseOnRgosEH5pxf7JQLDOKXXboluvp9INCOPWN5mECPj3/qtTWvbC5XLAyKZzPUARiuhbrDCoXK9
phaKmoE9GeDl5JG0fUgIdF3/i4mOLzQw6AFvDG4RxctbBon0ZxYWu6eVuMnt8lGsL+A6z/0RKMt/
WCuChyrVnl15QHZhUA/IME2y5V5leEKhBZtM3hkkVUoNCM6ePvM064/QZ0CunNev1AYNuh5I8rXm
VTOHBd4fPPBmiegApSPOF9mdYyczoxkZznBb88Rb3/7X+0HosBA42hEuhSSThD1Son5TJPLszaYj
2Ns8LGTo0GSJTNIwsZxSiy2WAYoOcOaSl0oBw0jUNMJNobSlYP5kCFqCA2sJa760ge0OeatDvERe
juJ2f2tTPFVKYoLaAIDsN+bMrGbFXNKnK/ZQsI9Um5DNJru7KmynvN39M/LsltzoAUnZbFqSPnWf
eJ5PimZkmC0mAAS4Vi/KCVKHHaneEm2CwsdhFMbtwaIK2Cf+ibpLVIxypFdfG7TSAloGobEQYpfH
ZvLswosO/bOxUoLTasgqK7URdfYHl4giW52qxxpyJ+Pt2BX1UwDMviMWpcf3blu1JZZjdX3In6sy
b3wnZkaZV79oiJod2LsSFSqO7PyBwplYwAzpBgXfUsG4C8YCxAYPhruR1uK2ZtT4EJEsBL5pra3V
8nznbss0EzvrVsnRA0STxtCruruNZwVKwfMeQSeeTiRaF400TLObW9kPhSgp+ohb6t3W8oXPjeHa
sqxkvRklsSHFXsYPQPAXkUewl4/hvIRGf0GzsXg9/aSyoxy0Qt2PDI6WLBAgzRvQtVVwgNef13ms
nLjakILKOafhTCXgzAqHlIbSw+xIElRbXQ87e8sR17z5agGH1gchkQ+05Z9dWAMY/5jAXPI/GCJM
B+RGGOXn24KEKLINVYZDYCdbOhpzL4/+9wZJ6/4ae8yDtqBe4xfEsjB1Z8ktMjQEiKocWRca2BDV
3jt/5hkZMie+Aguj/tyBM9LAhTekVst5JKOZICly7cy2wkysMh7IF1GNHK7qB6z6MmsZkDN+XlIc
L43iZ8qP2WqREmiwg6kV42DORUzacChmy61w5a3ZEpRkvdOsbSJdNV8tUDYGBOuv1+bnzv+niixs
E5kn83zPokBcfJ2ERC1u74kRYcU1bLmlA8FWWDAS3EJij8Kj1k9pvV+H1WV2Urxfxadzl3pG593Y
T/GVzzbTsOCbkotwf5tDQebIjaJwz9qC0p50EFWBtpPjTrXEfyEvlPYidj2mEHa5yMZPCRzSmv9k
ryEraemAQ9tnh+PQezXktCFbKYMjNOIOLh+P6jkZGzGs+uS8JjDv9UDFLakHaXhwen8WXE4TGT7s
HnVMPsGfkwBgZVCXW2My+eEMAq6lklbVVuLTHQwLCVj3z7n10XxQBJwG/Aaz8Kw16LX9FbpKnt0Q
Bv4sV//CK8Io44FOsg4HeZxvZwy/B/yuQBeC+qkrOG8QatxNxqR5XZCn9IqdV+BFl+dnj26REX4/
k2V5qH9nCAcZrxCEDvbjXU493HxPvRAX7GTscCWgNcMLDqoYQDzFVBt8sSJa08t+5g4h81ezVsIq
V+uu7gVHgt4OEpgG6n16IIRuDAZ16os4+zrxnA7RxzW5sXME+iQbIZPzD5jxHdHhHbGRSI13d5d+
FixDSyJkVwOvBmH8mwZHtrZ2kVqzzylD7sXOtmP+zwMFGBxPtRWzEeRpmDMVaGi2GFdI0EM4U2iD
l9G/bWXsmRHxMwyyOLZ95tZePB1rmbcAdJ1nEELRGQXFDsevxMxzQ+zNkK+moOckpuUIBoRGIFf8
we2NDIrkYu27nlOiV5VevZHxXg/9jvGFtaqueafIGRz+ezisfqC2wd7vVn7HKkqaPi23QbDHrhcv
u0OaTwYP6fl6AONYMevANKnsFFVWzHGG2juteKkzXMy4bmn08og93GEHJiZtNoUdwzNJ0wFq3EkR
OK9ducjDKiTAv55pglJqntfwxMJGulV+gq/FGvOcr2TlhvSN2myDqJZrJIRfkseIp45qZU4vzlvW
u1umDnn4CEN7YFjheRnfcsIUdkpAsyhUcZ1AuWVjEVxeExW8BiH8vkXLTYoTvyVF8ZG7fzPlswTl
EVPJDEZiW+8bBYQmUZn84Ktey5imnCb7Mf6ccTCJyx+C052ITELcw9yR9VdHuJxqbExdW8V6So72
xl75lhyCsvrBwr3RAGjy6nh/oBopPRjTZ9Osbk7Qq21hEVsp7s2Os9tI2KfS78IeqFfVoCmBU9LF
syqbyZFGKJcKoQG37++6S1E8cc3R7vKYmgNVaXsdPPW8Gc+6Qqbt5H+S6mJ/qKVyM623QKuye8Rs
L+g/Nz1t6U7nh63ozSxDx4KIrA5BmK+SMGGuFIG3irwwJjMR2mcCYzHbvmbcnzU7GShjscYWNKs8
1pu9XVh7g+Vp4zuH8jAzv+U/IWveEP1YlgPxWmloiOXOd0/S2bZNl/UIaQym+A1p0Es7OMmBooNA
97VF1ypDcFyMrrlzCmIHszBcPbsbxl7i6Sz3iPbhOfbSBbRECf1ltmsNhdG1p4rpA2Y1L2Dbdqbv
+5fgWBcuwzs2kji+UKxAQXs8oqD8E5GL2tIXADJE0kns22F0piAkB4xqv+CNAjE73Y7T6kH6xgju
3oaZVizogD/hORkG/iI7AvLnzfx1rAG66aSaYh/Vr0PUYK+JCz8Y1CDyJHXwFny+KMryISuWEpUZ
23Vrh5fvRDXjpwkPnSwD7wMd1oiU4YW0k3T/Ly50czT/N+XOfah3XQyKoFUHj1tMzHRcXi+ExW1j
uayg2drgWhOGujgSPWa3kE2omwfAFYB5MOxenPYaB1gR6kLJSzXua89XqJ/nfOhOdNgvrz2ideWI
4Ba9a7yZJZNoYSB7r0XNQUeBfVTKstNv3hD93kikEWA03JSBCXTDqaMc6NbxkTaATIGTvCUP0rfh
zqwM745U0+s9/1L2ssh+p4Kq1NefDYMiSFeKrokE1zn6TbwlspVNRNO1SMAU9vG4klLix1sdqT4Y
Rl7d49RNjsnzZ9QuQvmd0eZbDq4G1UU1rTiabMUWAWyZc3RVakHQoMgnfpA8yKC44vH/slBTDn6y
M6Q7iTYE5PKPlrvUuEusiw425pyVb7tdBKe+44/jdNX//t994qhf5Iy1c/SS5Mg9DMHXhlDmboI6
KGo3JFSpPGuap3LjlYNiH3fnrUJKbCmyAnaCaNx2xsAIYbcdI+plpWsJ7qUCRXe/MxEziUd+IbQc
Esb+mWHN0BdYsh5nNAHy4n+P7wEci5ydjqifEV1W+G21sZoknDyXfcT2UZew/NdRQKqO2dbwLSZs
9hEpPOsjVHOupFUwG8Q5u5jUNRHivGQbbDxnjr2/VsRWhnTZdkgUh7oC32og9lt8QxCkDRM7M/SW
DZUXJtUdCfmcBfsFTcg12Dq4IpFsL4pm1+Uct+H9jecDZ2retjW3vD29Js9j6LRWYSQCtCCh9gbZ
MWjRGRQ9FxyvC00HPwsKflUn+ZOFNXRHE/crBRS1aO7mc2HLca52ygMbxgLc1mzAtlW7UvJp2z+i
3r+6/4vp1vuBCdx0/t5d8ONZAVBI1tfl2ZtjoTZ3oASurXoc7EdvyBKjKFgIPXLjaEK7qKsMi6c+
Gus8bmfQt5eXvuUUTSapKyfr/lD7JpR502YSyBWr/p3VCul1PgLGcYklyRpV++DFdwvxDpWBn0iR
8xTY/XqK8heRCPAtcgu5JDRNFvgG+a3S/h7H2qsWutUGyb1pE53RRU6B9u1th7IfA0ogpqDLY9iw
YKvsB0u6PgWOulz5lP49XJiu+ZS+Ep72kdi93XDvjmtPVKWhzCmrOC0Mn5Yof2Bch9VYqeCJ/fJy
6AYwqvf84BXXka3VBIT6ptedu7LPwc3jjTL3s8SXKtBKTEQRjpwuvHKDFPtFzAv9ykU8oZQomtTu
XWn8yZZX7b9cYc3nJDvCsMUTk/txXe9gC2wvdCkfTreDZevfcHWOnp71Y8hoJIOO2TFkNeRxWmN1
xhfqF8F6xxvj62IzgWTV//57rMTJj8vSoMoUF0TYSLKKjp/FMIj7aIUjquQfk628ZRuAG4yFZLH0
Ai25ZedSgtj8Pm+rXy2h8yX5KGR/L0INXYoc1J9BKU3dO9mH5P2jS/aPrwoM/7QwfFtaCBmJBiK1
8IjrUyikFgtpCJeGgNVgyq7RqjYs0ho1QV5BOBuXhptqghmQGE4hvGwvU0OjvISdlTXm1VAyrfvb
N0mgPhKgwFDmm7JJwwwy7zzcQ2QphGM5brRpJaslEIFO8wUAy2pdBNlf6JqLlO6bcjYx/yBF0aFq
7NwM54PTYon3ZqIFV+75r2yEmPsUG4wWyBdiuRPZWjMP6m1AZJApVYvWSpTxPQTfwDMK+ZKc87fo
SU/Q0OA0YJLpqVSAxT7gTaZD8hbaili7ZIhbkFERsmjj0Bh5cmrzyKeeoi1Om7RH0nNK7AOvW7Mu
AumN9o4ErElgy0nbkMgmNrQPRhT4uzp8UFmiaXBU/pLUxc5n6eGok5kI1s6Tb2nX52gWQA1MM6wx
T/1RSzkTAl1KbIZO/DuwQKhRZpfpaYCyMSa9i66hZ0ItM9SMRh+RSpatX+pFUcPFvaq7fQfeAAy7
ziS1jBgjmil8qjArBFWx9JSVewJQD3xF7Mo/c99QxwJaTzRH69FXyUdxmVZ1euh/IIc7wc0R1JvM
Wy98MDiLXzdx9L9oDLtXSf7+lxUu2jjSgpttkv0o2R9ngtC/QgjSxd7BQYDHHKIRSk8LtZ3+US+f
UAfydlk3aOIBBasquWo/G5FD6ke7x/YZIUG5PrfmVB75ht4S4teygjugvg1kzgdVL0NER5OWrizn
JqdNaQPxl2eu0FZUn+qApYiGjNetI8mxyRLuJ20Xizib7+IUxX6Ar4YfEYma8lSwLEHUCJOLEH7X
0/1Y3sr5KZ+78LjlgEiXCFarOHIRymXSNtw5xvfU6CeWmWy/Xd0223TelKdn063InUyM/u9utr2a
swRpUhBUrqp8/nxwpkiaGfvu5QGoGggD0QC+dSTpSowR7Hsgb9pVtZV040d14tVOsLD9mqP0vQ9/
lE1yFeZhgb1XbqEJdB8f5sC5S6yBMXNv4CqxpKhyixBixcXokvXB80eolz9mgCbHF5CDiv4yjIV7
jh9fYY3wMav4Xs8Vji5q2ayE5HF2hdOfNnrzXu1GqxTCRaLLu+w0PQzfdiKjx77hCnKS4lE1hVho
iNco4Mmrr18JyFx8b1EiCJE3udCsFXSYKJIiLwMIPBw75tD6AESUQIKgoaRgSseh/onOm+HRXXee
Nnq5noK0WEwkZxOcrFxEjEv+idCxLtZoCIa/m49hHjYct7JQLXLeC+Pzp1f8JFVe4T62cZtvuDTW
8yRuDzojWLAT4ZSdpdlF7oCEI9nwYbdA5rj1Yym0AjzUv1AXLEHOh5EnDOMny88PUxiEomvFJnaf
dUK1CfSxNzyLTytyAoZOXgMAvsSjscot8FM0i9DOKNE4Pdd7TaGjvgQlkHmLV1OS0Pfa41wXiiri
Yo9m6Im8J1qFNsemPJx93c/5uXRxNY/0MJOQShxZH6lFK9a0pHcWRrnMlercUyVgv7T2ucyInerG
jgWVoQuKiiVZxY9aoVf3bSelCjY3LRolhJ0fc60BV5t/HLmiSaMDtaEsUPvR06J2i2wSQUCuUjoK
QlErCmJAeSLPWULCXlS4rCJddl13ad8FL8YFSxSY1eTqhXgd6b80hk9MoKUrmknu63zi45eympSB
Atqj5Dt6KTrsS7XqOf8ZQwWkbDLi5BMI4a55XIC+kwUOQaiajOsgSFeNVSdJKGOU29B/TyAI/LLm
WiiabkIvycngh2fIexeUY6T/v0ZlyIB55nape1VPnrrYsL7VWGAOSRZtj5x+AeDMCNX+dNrWFsd9
ZPbl5NbkbAiHWJ/wc4jFpRUoBWuYBO/A9PLnCH01rtbj4w7/a5iv2vtk85ijBeaUDt0d6d7cuEKt
fchwMOhs2uF3pEUFsu/CCoUNZQAyIouqlOPgYu6RR65R1dVl4o60ycibGlAzQ1gGNkkJi5/cNOYJ
HIc5Fv4sn4T1CYyj8pjOnsT9zrhjuw/fN0CTh7UUAa8Xbe97BHKT9Map4eNeFvl0w2NsLOI6XjDE
SU/LIB85BmbJToXnFf66mdLQ+q6UZihEed476vii97Syk4h4prutucPYpYk6CENRgWdiTszIXj0S
4vpULNqhAAvqCA2zdpzZ4cx6cL2Vdo95Owpolplp9XcrNTpdIRRJrWVD9fWRKViFoqE/4tK/WTr+
gRWHufqJcYM6HfierGRWY2o4bwvaveEyxPhXuM8x5U2aTghWHZp2jnEaVPxtsNIuEvoq4+g2RzQO
nVfScP919/7VLIosKZYI9D8ol5BGyAuCL46h4cOIdQ6kQB8IssHlpdn5mKe/Su8Ay2Sg/cd6kHIN
L7Q489zKLLCSvTpSgKoLnk8GmwJ6yDdY1DYlMMWdlrd4jifjSaEf+j56UBi1xi4tFBToQWooaumh
7ReDVVgppyHofVxNYR+WPE0img2OHfCI2ohZNN4HqxnCq2Inv4GloKLNtgjAv0/ttVaNq7/peHkL
BHEjS3TscA6sPc/WSeiRgSu5ZJEP9KOptaBNudWxPKhY9QGeB8MrmMZA8G1LUV3TOjcY/iZQEqdZ
YRM9bSHa/iE49KCe/lcS2FW2jOHcKRqhjQ5KlAotUnCoKgo/gu0m5bZS+lbE6rPS2oXi+PhJBU1+
D9wO9VkA2x+zCkUoHlHIz6B7o7w2HY0gqFXK+y06re009Ghj5vMFTbWqdPW+jOtPJpHY5Nk7CeU8
2hpgN8y1rqtnXgDeUJVXTpfGVgoCWb67hxCTqLnUGqorzFuVOwjbChg54V30bidszccJVz5NfGXU
bic6XNQirLAjwGWI5wtQZZZcttU1uPyI/+vXaTGsVbTucra701vH+UCYmzzSEGpcrfEauR+FwESk
1kmGJflUbkxmB4Ac9r8nYWCHQdmBuKU56DsjBa0mjDAjN163YywI3OWk+qFbpevLVwCNDXxU6t7Q
Zbu/WLrdUSUt0KA3gnfRbJCSzD7xqcx6FmI08/vYrvBCmrHOgGJ6gskPxs5iSavBc31qV4ZvxRdp
eN100/lUts8WgM/pBfWOXc/izATrED5zSGriGLEF9YY3+Hrj03Ug0RrS0UUoSIS+TQ5bPb7UW+P8
RwWumBvWCwsvx0HjxBoZs4sEE2dpPTzCm3/+Kc6sPK5Z7KHovvDE+KZ8kRZ24CwbroTxrGsWQntf
qvfIpyc1AmIfGPuBlwJ5F0NqpO3x6ClCx9FnfdFR74Qfzj423m9kJZuBeOjFnOJRzqiO+PKE0tP8
eyQjVaG9NZNelu1tnLbJv34B2ZJD+LrRcAePvFKveHwmwCgZr54aBIFHVGH/P1jO6SQmd/MGMb7b
m53UG4cRxktBFMG29De1Y1TgcBsHTKEZG+CKoHNnkoIgND6MCWvK4uQUcwXAxrLpWZTK7gxDksX+
09TjA0CFKy4riP6OfE1MWwqghz1OlL+QYYvtwS/fokx5aG1PALSMN+deNg5dlSk5m3MW/kr40MPW
45lcGKMLHw2J/6SumYZkJCmbHXcXEhII6osS8sCJzE/UL7kPQa6fSgIx0nh8WdQKp/XhXy4Tlf9b
2TcpA9NQ3FUB1SJZoL2WAiH6DB8NDsRkNsrGUHbH3sq26gvOvj8FPKN8rSiABAWY2L3H6XJCfOva
ctnMIkrqmz1zn31eKGSxubTHuOx4GKVvXmULJ4Y0kZr7rPTXyr2nxde4x0Bo5ZU84zXqPtxzx6U2
VtyQY0FV/wHbq8rJjgmigb0bKP+Hj7yFcBr9nM/FNjGBXn/bmWEDMzjIds+yxdnLOD9/yq3eIeTF
teJPHo6qUPNqWbA9nO2rStBxjFZod1mce8tRV4ekSKs3yTzdf2auU3drarV/VDipaKzyso8l1EPE
KJ5wxPlwDqF/tVAwUe/9IqZ/zaxnDMyHrlK7yLuFh1aUOYPky8nmIBY5ZQFmO8awIlBYddmVgapk
x/XKil2mnjTrO0aME3aROiNPvsOrw9wpjcxYmfbajiQ9gT2jcUQVZ+J19On5zTh8XrP0C5cxhhIl
dTWub9MvblKAeAwI9XkOtkPa3H6MQtEV84DWLaa77d94UYVC5RFBeBZ5XIKXUfearszwVlfkU+Ch
G1/Dmo394gOK+kYXhqotuQrjqocHsCSOP1sRY4PkvVeyC1ykSsT66MGU1vQPf0cnkHyuY9KjwqxB
xu46Oe5k/m99e3II/kwQ+R57WsS0lpbYOTztJTn5CEXME762QCmh7H8LQaW9euMaX6DW27uNKEjh
isL3VVcpwyZlZlUN2+kcWBcXPh+9YwVLRJ6llJzd3GK2vxKe/7b34LP0j4ZQ+ZBMpXHiLhOFhjTh
whf3AXaC5yw8y+IVnAhIrEhPWDP8cBfDSI1Nj9s1RwIKt85FXeMNAZBoHvEyC1sKhGQz8EaZ4kv6
RyIyOTGWZ7rXfJvCwqKmF0srR6WEC3fYlJccz3zwOaWAT43z2vAXzGuMGwEnFQ4032b+tCyQ30WA
ngZPHrsIe7IYg4uG8mJcOkkM4BjcAZOj1N2TDCUE1E+DCvG4MpgEIW7IjbyW+5xsxRfp1+hzQgCz
pOunAyYkOZeep9N2H8HDUkuCrpqhXNl3gyw43Xo3/y9Xk5RaDa9+CJexaDUm6y8qIX+4w3eYrcdV
/jrRaaw0qhhuGrFP+VH5TXv2mPBtADFydIogoI28v0+iXmXhbatHKeUSTtNTM1N8uBLgyKRd/6aa
hRnjiRTiTiN2XKX5DWMbAPfYQ6mn93xZg6WFGDZliqcKFdjrNoRUHNt5I8XhssiScevB46tr/bKV
YOU/yznAlsX/GwYKDZ52cGmC/DdA779wewQDEECWnZZMmw8CB5nBxeWr4n+vKW0iVUe3KAD5qm8t
rXwrBF7e4p9CDeUCDfzQuy21LLjzf1S7UrXTHkmNZ5YIgxhOBmaAx0ueJHaKUiiSaAfroJdxX58g
Uy7AT6FumjjX19ufQWUTW6usB/0xNm2PFX6UVmf/ibv+5e9Zms4AzhMZdqoVvxHSzz2UoGsUqUlV
a5TWRK8B66F5BpFKmWENhEto2iRyLzhx9zkJ/os0U0HGTfiFzDs+u2vsYlVjL3pACEyCpt/xiLy2
M1aDYz+NH5KdqTzezHCEaP0SyG2wzqMU1BVykXF55wjbosXOG0dk69i9nLUqNF9u8WlYZl6EU8jE
5D9BIvP8CTqB6u4Cndl+iik5Ku+uwElXzWGUkc2676KHcENyjy7IpG9Kufe2OXLlLYH9yqQ4rz8X
3L96Tugh/OIHib28ddNt7DA3v5otpSnFpqnoUkAxhsLmkfEH1iVSIj90kaIOxA4FJUPcNvabcYqM
y2hf8tauVxnIXuT5XJZWvyxa031PfOekeXMprXehBQ7rMICyWa6x1aYkr0Ey20h2kDL8hj3Q9Clb
nQLsECBfaH2YsAJZ2o32nn0TQhh1W/+cNWtPY/cZflXvLyrlihW2NISLWZcJCTOyGNjay43j9n4x
E+APGauX9ujMBKZdXrAE18axfaq13gYoQc+oOC2x0veuSFit2fwAjpc0HlGks3lZ0BkxAxAyVJvD
rIz4VrLqtL2f5G3VQL+6fKav3P54k/vcqExQhjYaC6Zq1HkXj9B8KN4HeDKOuci+7v7qEx+4R7ed
ChRhf8T6RMvD8LD2K6Sf+t9mnA+KZLS5BWPXxneEIcN6B7eTmz/gUeaiPvSwlsLta+Be3Msr86SE
giUtyEoEQUCA4aTUL5E45ARmxJ6UpscT/6hyfIdkgIFAZYDQpIMs8YitMcHTm4s3f8H4pHVaZ9eW
uOPyXzweti6h7s8900PnZhgLhuYvxfqKr4eHiV8XbCj5Y9AJg0LamLypRMJTj1sUdJU6sLXM54Gd
kE2fH3vUvyF+KTQ7vOak8LEmanvB5Z99AGHyjgBXqJHBZ6nBfK9KhE9ULFk1TzUyCt5uBdI2+Ri+
644mmAIoWD/d0UazS9uI2jWuWU+Z7jLiDUly9k7+LTjnYf3Rcdr2wqkHXpsLk3j2YEgfO1QKbo2g
L2JVY0wK4vhn7yPmvq8TECk9zNVYSVQg2yNctqCVU8RRJnubHSBKAyDxZ+Pjyrd6/aWrRrlVtR13
fiqcM1VMqzz+9pc+hAtx+1/qeuWi3zkpLgEnKT3l7u0TUOSCNM92KMcLCNYVEx1cV+nJ4h9YFEWO
CCY2tnOVy+ostCkkEPzv8+GMKZJXwD/TGdQxl8nh6UF9IfbhTcoUwyWwEF8+t5un8Oh6LmwtirSe
VCwmvhF0QwOyEUDOYJqG7DyrzJPy33rNLZ0TH3f/lFgp5bIJSbhWOQt5JUPdzGJ6gNN/uzIVvPX2
vh5ulBpbK1FQb40jNs4WhpVnN98geiXC56XkoaJ+0b14xG3UGIQxZ6fP5g0VY4sCs0sgkxlHGz/7
LTizYQHC54KFMUuVwoi7jLGFwjvDWKIZjBHngetZAyZ8emw1mlYHm3uEa//bb3nOiMQUZ0CtAmg2
boh5LhHQcWnNv03RIOFMEy8waU3quN/LNZ0xFcN8Dr65Kwh4PF5gBMPvpcbLGtaj3QUjlQfeBSOD
JZJiV3pFHVJolt8QMe3Dr7+A9UU+cyty0awdfzkn+L9YgWsn6reKOyjQ2i0S+KjZ01B8EvEWjQxi
90rAI9EpCmy02ll6F2Ky6TQIL+L9yZJF+IDE595nA1zi2DPmOPG0LvEqF4I1YNmbyqZeP1A1hUdq
mC+LJzKApKWU4zJOuxfpVzYNrN0I28QPrm7PWLWNrqjIRSOTUbWFwldGeqtwFEkJYJXokjA1nDtF
8M5YvLa/nvWQzP+AQhgHvicrKmBjQhFUr7iEOMaBEcltQUBOpGxuvLG5RqiNKUSbVOzo/PsKeY1x
+nuxp8/1HVndvF77dqXKgq6GxuVla0Qj819R63xLVKJ6qFTKNdorjRshQeAan/7roHSuPcPIpu+r
O0aczm7667u/uop+jbveHl5EQq6tb02Dv1YVCrnJ8ykaLP/Pjg5ioHnUbfsCXcSIpuN79QzrD60C
30QMNs6vCJVhXmQNopMsCUJX5c9VhmKmEo1EqGmTOzCBqb/x4+u1eaqy3OfnRg2SI9xrO9xFLsEC
PjCpxZZH2Y9Wc4Hrfwu76GMwUnsZN6aECBBzB3N3p/FPn89PzjZcr62dDFk1RVBSyo8TaRT/QbnN
+hWszTsm98hpcP7J/V6BCpqTIW+0nOpsmMIChI1WP0MQOf7E/PTX45Ei+BTe29Gex+UT+FKN471W
OAged+LVU54gSBuSK2e+MzpFLP6voT8KH+6G7fXA9CWk1gWFuBa2LaNRpA75HxpjrWERMff9LR1E
oBRq78Kt+Lq78LdBh8wuEvFAkgTB/Bd42OI3sGCyXwlxLYoFFRdNbvfJbmaJ8Z9Q08JEnQ+nVU4n
azmDvTUW76ggJ7elDEdMGUx19ED0TsrynwsAjR4T6LCwACD8/Jai/DzQAMyDkuOA4Qo+Id0nKIsQ
kbyvJ93wWAEh1bT+5eY8ndETCCc6cxFIPjT2i19/5dx1CycSX0mUPENI0dICoJ4fW6dP4yXJe6uu
zKBgcgeC1GgbFFjzfbD7RYiip6R4Xgkv/sU71d3P+Cy3UFf/N2Wy2zbyIE7JxvvZkI2Jp9ClvVef
FL1TzspdeZV/8jl5QsOGf9KhxxfSl8eIYXsvn/8cslbuSen096jwP6I1OoQhXOvuBMrP+wNSJL8S
CjgcAMLfCV1Xq2KUv32B4goYllh9A6ws+OMG59I7Md7Xv+z3SUrgOWw7wQvbxu+fmmfcaovscD59
RCOdc7gLEs+otcOEvROI5I7a9GhdRPqfcgn5a8s2kmxakrnHm4dvNkUHh64gNEUfa8CQR1VeVby+
M7Xpo2q0rF8OOTfBU4/ZyZGw3h124iNYTqrn5kDSjBGAXVQiPSUhm2A9/M4YsQGKau4Ue5gAfP7H
w1zyQMEua+FKpOFmH3V27BCvHlqcPWih7Lu49Reiy3xze8BUeoS4o4TC9INM3CNGYKPDFzEcP1yz
x4xdDgcqThDvtLpa1ab1+kH+5q3tG46Xbaa/YVSfzNsLe7f5xkLRl2gjyxybb5nznx0/XCJO0kXX
3g41BpN57gRjHFzuVB1jdZQWVu9cH2Vj3Fhscxej2u+/yGBbER6iNuLj6iktl1iZo2a4WnjQtdKZ
IFoM7QesxTyoEJ9F1TtCUS/svJVAefoN761BeE87gwn6ST4yT5pP4SfICg8VhgkchktU6RtbdGj+
X+ej+NfRR+NL1bEuqirrA/TfJJMHDBv85L9SQZOCLS67F4z7RH5oJw9ppk9Oe0xfePsk87n8c9jw
dOJ6jsTrkw5lT/ZvRIO77m/AaTu6rf/yjOZP9tTJpE/dGYUp0Ez5iMrL48A1BJfUQTttbMnJ0JOO
O4tl7V/Zdyu4gfRHDtS4AlowZosQYvAKj4D4oGJozPMZvqknQMcvyA0b9UCHuwCt5a6JGcqMfiYZ
xRIJpiGpDfWvWmuv2YMNRigRQ4LSCr52+CiwlZ1WQUUwfbcJtWrvFNmrQRZuyUZyi4dx9pifWOZd
MnC6NdVoiX6J0g6ivOIzJdnx/NNGa8ykHvwah7qobYMYi0wz3bJy6VVlCvhuvi9++7WN6rv+oV+Q
BFFDxO4ehJ6hcPwZ/omOp1fxS601pPcR8pBS/QhjQEX2OEkQuzquWzEOLqDJxsE4tkPOrjbQHBxK
3KOASgrWkiCc95YEHXc+2HloInxfpNvdDQHVTtHLDKYmlp+c5lNbJmSk689fJiIOeqsDcaXkL+in
aWGo5TadJUM2XrCGNVMpQSXhWhqzZ35UJUS3m2UdJllWh26FjOD+Mw8K696GNKTjwfwivMIVAmrr
c5bIWfZvJfpZF3/a1EfAp9pPYlKnHO6d0uQx7t17l/nIjxyx6NPCx6iU2eAljGFHM+dxNz4YC4hZ
ABIHoCUDhb5J4ArLjLs8WxkxG8+Vxc58s/rdIJbJ1g3K0r/yc9F4clq9Z7Ajr0bjoJJEOlF8DAXz
zytEDm/D45iEC3haKh8DN5vwmEXDXuMkuMxj7eDc96rV623YapSp7IFt8LWpgbs7jObtf2K3nXVe
w25n0uGGmWbx7ost6n8cXRNREHi4sig8MkWckkem7RaTNXTxi30RZzkqVQrYH5Qgroq5uph11hzR
JjhlJbWPJ4z5xUTJnyZ2xJjLisAEp1fTcqb7JRAnuzo/OGD+Hya3jyjoSIHiIWgCO+ZqvQ+wicMn
AUwhF6UWHkhXbKAKdGZv28yxeQTiIJUrm1PXNJmqrpNLBj1+LmgbmyBz8/Pt2cRoiSDfPlb3QIgF
vQNZ1K3zkCUnBTnL1IbZk+FrkVC0mETqquqVbV9RFJFZKuiWxjEvw7BGaJaZZNI/HSnTDvCJQewM
VIPZm/HAhxTWQbG7uYZ4DyWyiwOw7MY7QPv/eihi/35jwi5HlkChyYyMXsrYhxHbW0ZgIR2rYHvi
GHkPdbu4H/KAhjYbh7kHmbkqtDg7kjSUYsL4Aiw+skBTh/JtFK2nsA5/mg0fzbl7a0u8IcplRVYz
xcfFVPwuLfXEUvCg7+5+89FzV4Ps/QpLJ6rhflrhFk9gxNpjc0KFGBHizVKWdko7To1MceVOsFRf
D1MJEy6NJh0JYmgo54MC/ErQPm36Zcl38z6saHKayOGpbiCaLvNIDkTy2b4oDHO+hJniHd2P35ua
SE0r5AzJRbCQU0Uijr2XFvav3JRR607bb+N3Tz27ctI1kuu1jh5C4CtMZf1nno5CuylFNd8TNQXQ
icr0sHDy90W9cXIpTei5OOo1BUqVGDoU/hXM/dKTFvtbsI9JW16t3+BQbhMMX+HOgEKCEVK5iYhI
LgAyeU7iylruK9/9d9d/9ybRSKDOICVfAWJvGgNecyQ+TMWRnEhj9ti2O1A2FJkXRN0YCRI2evl0
eEBg1swFnheWkOYn8H028BtDS72FaywSkF+ih+jcHc89tNMKxxxFfEHgXAuVo9umNQOu2atl+ScO
PnY+jFZX0U5no7S3qbEsUucicSNu8UjqBNQLjYusg4GqfgIjstYrngjO7Bgrk8jKn+KWtluDCa0q
IBFeV8LX15QSTIQAX2W9ySwWCCY2xyC6n07rengO1X+lbsVRJq8rN3qmm86KRJhGZv6JfJToH9BX
ugv/alNfUh+2uz+W1ZmNFM5URtJXp2s54fVjgwAbW8mD/9vWXrSQNVzKBplllQNFzTMZraRKT8WJ
521Fhg7BGdBOrsMGqz87gC/MVS6beR7RQpZ9m2N5AlD2QA6KzmKz3E6lxqvQbiMg2OWYMeMEJjbU
4mFw4VrQ5r/2zlfWqFnW7ZvkGyVUQ1OLIDhHWec1QDRqzpDmt6GH57a9KGa37Iow20g3ma/bFQRr
5vkq/XBF/ML/AeGkdX/YqDmdcPneuc8IjymQzdl5WhTb9YgUdJnyPJVM1ZnFBTsMjtC34hqpZnMZ
25vb/LAVs13SSXryWcGwIoFDhAbj0zSlGfeDkpGNpjCgu7Wwf/rEoyWnp1FoEo0tyJKFZLbBD82C
U6z4uac0VYOmfEdMyvgtH0qBshV24aqwCy+9/1WTTq0aYJCsl/b37W1I47qRDpWs2jQyreRIu1Pg
o/bqOUXujX89a4tzawVhlAR1uGGtoOlEVmfPj8TAqkGPOX0mUwqLE8/G9UR8cccoGCp8F0VfelwT
s4rMqVnxnP8lAUSQFf6nJPEXSlIyI42tFw+h+mBYbD+nOPvqHiaI48Wxacr9yhVMFh5mMtCWZA1+
hzIk2JRCdSrlExan5ylDP8o8Vu+09OfnU66eDi5dnRd5hflxkSOp2+zbqxUziVspqOFXvWqi/92s
4OzKz3MqYHzj4c6l4yyJt1M++ghL9SAW1lQ+7jkCrJM37aHatwcxn60RvB2eQOuRtXYh3PEQYRhs
MFhcWy1rvZuac8WTvdvcsAk709/8bluWLoaYA8l6Ojx4SMju6TzPL7LWi6pF4RvhVwZvEDo5P296
2oNAubEkDaQxgUK2EXz5BMVngpI3sJO5gDvbpqYRvHgMrl+WligOudFp0Bgc1V3/owaBfiGmzQ8y
qXPh8d2QqfnM36LfCEpy3lBs+LFZNRTI8j1fXwLMOU4h2RPn+00SMY1jrSWAjAXAh3crTimSQixW
/wRgg3yZ1KLbQCQIWNCXH/EUjS3PNBoLpbyS3fwnXSPvNPC5jMy0T9OvQXIsAjZ28usQKe+V9ZAh
7X5uKW0Qb+ETgoRIVhACE81VhRc0tGtix5cLVLSNK1ffWo+pbdTOIu1QN+EMnfrKQ6fLFBEEOpuQ
TWVh7x4AHJA2qWxdR5EwaLfnAoFtntxPLrmumZrOY4je7OGK5f/uZPKBqD2rNC7hlMF+Fa5D/fzR
yphCy1P0RNSpUuyD/Cz2X0CHzQTRFH20QuzLcIN69+eOHT+jQxTxsVjpm9C0IYS0BzmVbywphFJL
luhz0sGilf/vvS+FDkVW06yR5JAqaU09k4GYOQeI7G9anRYWrHNzM/sUC1pyy7pQ566BuwTcnceZ
TIRUr3UWmdpPw/nOCuERS4BvIpCkZ8JUnuzay4PfPmfeCmCOV1eDc5Nq4nZhQFrAmpeOzgYl50po
4m1K5kWtq2giZlOcj2VD9hfMCpWdzTGxrHj9oUxYmvmT1GI1D7e5sdELZd0aqqRr9E0SKQn3JmCB
5Useiox82uVn7b+C5TI0fY1FtsZh/0+jBbh8Du9trs5vPagni7QXq7erANI+vzzB/vKeIMQcZ61/
G6jHmjNp28u6Jo1tY7zI1VzJDPhZVvBekxDZq0aiyL1hJN8QoOGZ1GSSPP+n65c0SjeEWT7QMvL4
tDoFITb31PhsvPEmR9xLhfpqqt4TN9eLEIKrxAnOZWPBGkEYKnq/Fuz0iLN5le0mQm7aJR/MiPyV
dcKWufM4mMymIh64QGAVmqaTyMDJlxDc4P3ZQAdfkFoVnDDApGHa0onxa+h5U3X9v8vcvLG/SY7y
23jf0FaItI+FEQm5dVL53EGlcfAiiOa5w+s1z8+Ka6Z6oaW9hCibF5h3SU4g/wo5NQn7lS9sPo6L
whfjbdjqqgUKlT3Ae3fq06cJ3xZgi1mpy9uJOQ6r/ByzwOvvkECEIWobObuGWo7cg5BCCBZTXlFF
ZkQhC/1T5AqiG3EnKEs9cH/E0ZazUHxwgHu2GbOruc0IqrD+YnUIP/+MIUQi3fEMGR3orZnnJr67
kvmcF5vR5A5dH9MIKfAqfrLtCShsco2HbFNiaFG5grYyj78tHV9QmRBI9oM2oGlRYilgdFaTnuCV
fjrFLRoiyKjlKrKaBak3325aYA6EBtyBIvj6uoEkXFaRvf9iid4Ze0GBRlt2IURu2i+4t4+3xWj3
Z68kdhvRNqNaQcfPPy5BuzCVWFvwgGOmQsnpDzu+UNnVKWu7jKD5iQfXFd1fpO5YeXX+K/qhGRDe
ZJhzxjPJnDRs3z0qDe+5xlQmSGk5b5CbgnYD7MYWK7XJMJWhB2J8b1onx1xu0sNtvr73/bfGUDoR
I4j08zU+7QvkAiRvaeeFC1mf8QJJWMO9TPdDgUa6jD2jp54nFauDsN6sAW7ObH2yt3Xsl4Ul63OY
QDQ41E89eVaOMcYQ8c3P/K5w+q/hnq5r0v030F/7g65qsGka4et/lBTi6z+zRBygRW4lkGn2BByA
D2EbJPLrIcXJ1So9p/A699E2awZqN4NDYCAEzzuIXeGuXjJYfEXrK9WMjTfaQzTTdLS8R9TnMx/N
cKtn/t0uxNFHMrMKHWfN7LHXkV4cHY0T4T6luYwuEQkIEVnd8ssWP+KLbNgttQTayh6SkJfUjGYg
VIN2VaMtTdHcAgFsEoSdfw5usXJlh8lYGw27/3XHX+xVlfRNBFqfPqBt+863KJBREDCOpKhkfFUJ
pBSaRfoXeE8vVHtErD+gYLJMvTSDytGTwjIHEUGdqSodcXTdetkP/1riLPFQhoX8E5CgfozHeApY
Sf6S6GeZwy2MgQi+r2C1Dgw9ai9EGmlNuO8BkLDYKLq4y1bwL5ELr5071nvCf1o+bEwoqNdZa8fH
m62O3Y291AkZEc0keSlD3Lt1gKpDdxN03Hp6Xn3QEMxjpXse5KSqcV8wtP7DNS+m12nh8YmnsV2T
yNILLWs7w1L1jGd5LUvQRFWUNps5C9FoikbBhYwhlNJ8ZCztxZlNctkay1i8XWOD9O/3QRO7Gnt3
R8vWOpXjWVpMldqcIYc/NRmy3nJ5x/r+ueTUFnw9zr4PmrbHZgivPk4AqGrLPdrurzX+w8Na5y8h
JNgY4igXZnoD0L89YWzH/LjwBRAFZL7aR6yRDLAu1MuINbYiiQEWM88wz6800DExyaOfBXApW/ap
372OyflnIZKUW+MxApjhW/Yv5+8APMd/bFHcI242Ce+wiwDTJaz8P33rSOmlRnA/eBdGGPgiylNQ
SAQyc9A2jdcEpUJWcAec8uGvV+vwwM0XaIQ4TMfqJ7GZMukY7YlKQtbwYb3nxxhYuI4CJeRGMhnm
ZW9u+KYxHDwLfmva5yCltygrMO5l7tLWgjelHbPQWaotw7CgM7KTBrJ6t+uvgAaJLQfrUAAX6F16
3kzR/4OaH+vIzCz/UD/lXkmytA3aWI8yNKWU3TYYqKzu5Wx7GCbNb9qgRmlqcnXLjbB1s/CO9X7D
6MLO7fg/HQRUV5aPKVPMF3AHx7vIOzxC9m5sf6VttPORp9QWo8eTXGwUz7jaN9QcQdLZL02ZS/Zh
I3FvJJKhQsQNI4tHJcZah7rwDrJPNQEfV5gy6P/ABCKzevcV+TVPJafrCQ/h1IAORtuaJRKITInk
t2JIg/fGMNPvnutlv/STBjqlIDchsKO9bWFW4buQHGEcj0dXMfCBUAXFHJgeZZwwc11BahAVWoC4
eIudxTgCy3Rk0p7Z4VD+Nx/qX07rMA4TXs06ge8mqBpr2huaLStFjpyG6J9NjOWWqnkaIlQPMFsZ
NBfvA5uQ5/NI3a60rBg1xF95B80pn/HcUuhwVk/z2zdsm0WK9dqWkcZcVETU1ZIk7W+gUAFkPfOA
faQxV3J+mzngPGrJCUha41N/PR56b1Q/ob6MhVUpjcDt2063lyBikilr84VDJuCmOe/ZuixQzUMK
UuHQDzeO9I2rUidN0v7IX08/5Gmna9ulM2LIvHHsZaEt4XD3F0v3kGvs6fW3IEncevZvtqL6rnj+
blXnQ4E1ZAUb9OuZtEJ37dlsSJsTv++/fVsh3asiiK75h4tKkhA+N7BmCsEaaQJ/RCjSVt66HVfD
muXu2/1G71TLK7QNBTXbm+3hpJyjc8NVRkJL+YgRXYfMN1rF2Hhj3tIbAdEUH+/Y8beUmzVCxe4h
g5h7BzGkIwoa6TgcUlYNSaamIKqvuRYNjnO5rHgiKfmcE8mrs2SC/pAGKR/BJh38Tw1WQZUaur4R
irLe6E/S4PtJpB21C8fddTK0pH643MmbHzN5hFF5PtaZhUvmSZ15JlVykl5ZZQGOtr9GeIExUHcW
0se4YTc3i4qOMbDPPRds27ZBlIHRHUSnyy/W45f2D12EA4HgjgKdSWzzeDzN4sMKQeglljRT5n25
Wzy1NDi8Bor2Ow/j6zcyLfFWgVPeJhv2fVyXOK0EnW2PxiS9MVHi0NGlBDj5FPzLp/Z93XInm/s+
4qVhWhg+9LBocOEzk0/QY7q42HyWkkFT5RHTiH2GA2bn8DQR0RC2Uwjy8C61Xb3qg5gkZ868x+8u
tjLVTc3Lj5RWjrlF8wAiteJt1tEjX40H8qdyTx4OOMQCkMHqH83jTuITzBRFbh7N87BDVaAKhMAr
Xg0Dk2qaUYYO6R0qM+d1ZMYExnumZ/qtA07uB3V0/Wo8zdo1E8YpKahNLxRyn8ik1Vra7KGHUX5r
obb5WiT/rMQd/8SQLGyhfVwTY6J/YZ22N/UVkf2gjV/w4L4cJff9nT3HlLfswtA2532m6jbzIXow
Lfdl//yUHdvmTmtK1FLKZw+/YUbQOcii0ba7hY5B9recZDkx1BC1BpYVtGWqW5RY2IVad0ZVzLm1
mF0WALwLcEtZnfVwq9tNFCJacKwQD5/76JBLSoni5bCB4xiHILpmXBX9kZ2VPEbU2mEDJINHcsGR
0YybkY6ifBQ8QlfdgePi8OT1GhnCMzAkrwIDq1pg+vngHG/Rv9DOwrhlUkVpfPmuHbz4++zhVkUt
kh7tE5UURTrDjPgvimHE/gbFzg1sOuog040UNxEew4mV8jEgoYaZEgAhVfk8v5HyS/Vm/AC9+3vK
/5I7YLkv3U3/vOb+KNso/P3gkPnUiry13TMipTI5I9y9jh8bpNj5/PSHK3YySYTO1IDjg7pm0ajB
cblwaLs+bkz7cE/aPQ78VqBFkfM6fiqhD1bSFNqqEBk6DQXgXGitJOLezQWh23iK8lg8gKrPZf73
3pWI7FIsU7/CrqymFTPSxX0YPjyGMlD0nfkmO7ioBK0CLZDBmPBfuQJgkuET1ldMdTLV2GXcBj3A
zak32lfKpiXIx9KCBz4WBGR8vtkVYuOIe2Yn4Rbh14B0IAlDTS4MjQac4f2TslCqt6w+8bvuKFMO
O/RJKMLeS9LyJOp/O2SnlKwKIIwPf/xSToaPODB39jA/nLiWma1Kip/bgrFEzVMmDpRHsgbQB02J
4FnVr4GAmaeu1ZcTHnwqzYkhcdyJhzf87WkbLsTBMPcNbPYUNou+nwxHiBfmmVQtkjKqdiuQ2GSA
3wleU33Vga+sEyvcu2RAbNVNjQMp9nnssfVbNRqhgzizhXPU5utaKM0WyWAR9yaZ5yDrY41w54ij
Ru7jRZgn7qkSfkeqcrtI/YSciTXuNbWNQJzJSFmsQ4NNafJYGnhVLZ9mhf7EcOArVPTyUahPqsa5
u/YRwV5K4cVtvslfET0Ir+XR7NMMy5oM0WVPOj2f1swjg0MA7jQMs62rEmiUQYeXcDh1qIK9sPTb
JLKqUxs5pRPD3dYWyVSs/Ila2gRSj6MeuiBEaq1pcNc9VVqMchD0tmo3Cl8ow6aTAYEWO3xKccsF
P6aWP4RadGJfyugqFPbpCTib6aMAqF1SqHThxY03Y9XW4enb89U+bPhkujjLDogcJGcccRyjtWY8
1v5uble/NwyK/7Hmy4/bf+gClhpC8m0MI6BhNWIK87FAufRi3w3iHMUnAW2e8MgvNZ3LRPJkvvW/
yAZPZ4YyWBer784B/7Rta7Km8vKJ/wuKv7vCJgOuh6JsXdhyFkNcsGNRE4CIcZPE8rScTnOBOSgz
GrdDYSIloP5hYzN0ZVcyVVAACbaEnq7ifqS0u2y6TwfHn1nrxp0YjLm7fdF/5TGY/KICXO3RVuJM
RMLVTZYm8Y8xoFyM4uKKesdCqe2FcbiXWj0JfmUXFLrehorT08nImwqU30VC3HEj59wfUOpdAous
qJhpABWQyjJnExo+GPIDP8UqU9ns/gQmq75FrxPSlrvr9D54fFraE+Lu9yJecmo7KSt5xS63pzOq
3ovECdvvXiQLClOMNeqP8vwBSCMkOiI9pJR/H3gcK0XRugd53YCipOXsM4FCT0mzT+YWWUqj/0vV
veYpi/sU3vKeOK0nIhx0thXe7EckapeN6i2wig0JLV1JTL2Q25WB/VlTDiPn+ZKEXP1pwaqHy9NS
s6fag3az8b1HdRQGL3NOhQ5WOGIBARw62lDNdcKBmYVCYfi5JB6WZ3G5Bq+q56vcBbNX19Hm4E5B
gKySUl3jgNGF7rYue/YTtG/0K2ShZUYo8mUDtL7+N1GPz9Ab0Q+D5i/YuYEHlw+9g/tbglKYjCQl
owWVsO0VsLmoi2jSgqKjAed9C74Re4DwehaZXgS9KastZd0jBDQxa++aMZmoXeqo/FFm4viIscW9
BzEDDG0qntGkgAR/eEj/M8Lnkt0CF/SpIN5QYx/G1tvHDfmA0A+QgExueT02IjhHcY05ASNZX3Wy
41Xqz6h721ZJA65F9Rjz5XxG04E6/zPpCU5dMFau6EgTUUDO9VPG1KRPMoH+OitMbTvhIKBubDub
+8UvZe/4lXra6hL64f4s4Lrhq19uLQgRvq9X/cluVELjBtUJd0KYA3rGAP4EJ8Yr3b9tVbKzA33B
7SyAjKssAoiLREEAAIhQS3uE0sVwzO4PxjqwxGVRxNa+GRuRkCBe9OF82BzEpp80P5oTZ2tD1h8B
xl+9rDFrpZO0NvnJTeF2TdaOThBYjbkBVkZPxL00pjqZshmQoS/7T2yah5Hu40MY8jajW1NqMmEQ
7zeoWFbFNeUy8p1Nc/P2D1akmVZJ+GDefOVMfb6dXex4Lyr7Gjrt8WQhlvd0Z5eUeWRO5JG2fPi5
ce5OOnclus0qSvy1330d+02X4PhP8Q+E6Q9/Hr4aTWeSzvV1fJrdiCk6xeFYKazrt00iWxJSC6+o
1kcsES2SqofjHX1+MG+T5F50qw7H77vVjPlKuNV80lP0CBREpfXuYklE44JcTnUSc3BA7ky6PQ/5
RjPxAWq8BUvfdJaWk7JDpb1/KQPqrx61MZ/zex/OhgUpnAr7+KofA3C/lmgfZ2L/JljjdKid/n57
eO1NSPPeSL8XVSCFkKK/mzXvSfVmW20UJ88rMXZaGZlk6PAp3A7QB5J7mAjP7hqQhyvoLVt4vVyA
m0/OwFwOqOO5G9dIgNnwVoHa6741i2FJoOapqXXEiZg36MzTh+LkWexd85fO6T4xpZWMFP5YVAKd
1NBezsd4v4yjrjisdyoi4z7js7Q3HM+3Q59En7Bwsw9PqUKCgr4+5cVevOKdh6bQ6P2IfdzbywM+
LjmeLkB/WA+UbxH+06JsdKttjilYH/gocyG7lIToiedMDaU4KPfHiqICeCZO1syq+7ExV2uFyPUd
Mf5eZT9AbuoFWkCuPxxD2yOG1PfCzExR+AKSno+mNaFUCVh8GrjWxLI8mj3Ij2l5DTpdxums3+lT
XAjSW+EBDcYr3eunbK6WgNxxkeJ4yziScLzQQlHBnfckRhUqWmBBk6ExogtIpNMTKtS7xyqyQu59
WTfEqrZMrU+CPoA2CSHSDfyrD12eOXq21xE1eX4/CdBTCS4vmxeqeOm2C8yB/i4lcrkW/CT/Aawf
8oEaKAHXJ+In/AFdIiC1jWLih+LfuaPzcJR2oSoQY/qcq7q+vrj9SpqTr0+Ga3q065koEcVPP5q4
r1nxvK1w6ozvQiydvQZZQdY5XJihaxRMjDabsUft6bh88RdJAX24SiO4JoNtITYM8bB6Plg7sK72
a/Z+WP1bSi8zmUeAE/uv45cGRRJvwlPgtcwiyRl82NQHf/DXwE/jtqW645ppSEyICT37rGSl1GwU
ao/Yw0Nebuwh7EDcEXB+3o86XynRwfKdIxgyH+S2z44wzAB5KjBXKBLxUbEqSXjdyBtBpW1JUsb0
/MDrb0yLvvvu1zJ4G0cJlZDhQZSApVe0ruvNF0cbKMBeYnpphSnunNlSfDRBXyhma1JzJniOHW2E
BxB1SCeavdXWHudw5GhI830DXGr8PIEVYDxQ5qKi4xZmjkTtD/jZ91jc7CGh7yDBUtkFjguiUifF
ZMf3VO/pyA7ZU7eNFr4XZ31Uep12JiuOvaDU1csTQWZ/06QOh/m2R+9RLlISelI7INq/gIxxtFor
yNbczW8gXD+LiGT9yFsYPOf6Devqi4uGLy6VCVYJAiz2Mbi5NcdnxNX0FUheypD13ocap1q3ZHnh
K+dEgiDe/ENvKRsgbIqRII/aNUsG4z5+uq45v9mN92j12swoCKBzW5OW+EZQDsuj1UNBdI8mpmeo
WzSRm7lwDYe1/jUr5YJCRDHbJuKHlOy6RgVvDxMMaCI1oDYZ9g8aXIcklZuJFF8ym3aaolAwnDoU
IrjexRome27y6jdifoT7a7KvGinzwdY+b0WKIRnw5lDPydxmufgkMD8ItWSJ6EUBDl+yFWdgPuZ6
OEwTUnbpdR+yMlo17ZexBKDa8XYO5maKDS/HjgCE+8uZzB8s856V+9ic2VkxBBQMXPhc3Z7TQY/j
7aTMgef8bx/YqDQObBn+bT0mC/h0yF6OUQNqnnGIdXyQIcglrEPwkgBmiiOZmQdF5cFJ8ZJB5DQM
lVmhl0E82qcQGUbXmMxA6ENG3uCxmfcIWpK6Fg5xPa33BmNHAY2ZWauyJhV0AXdsc+c3skq46sc0
A7aPStZl5M0/FO/rPEGtaf86914+r1Tofyo3oaV71TV2sBul56ZQsXB/wbeed2C8D/rUs5k5sjX6
WcftINyXph/w4NKFAMxy6/MzqtHqf91pao6ROZjwR9PvclqNPqzpS71Tjq+wSxl/ou5nwDpLkmOP
kyUwyjP0uRVKMwq2iZp6oiVCpUCEedWNMWxLdbBjycGgZP0GYPIhvND9FuPr8ENuUwiGF4/ljwED
TMz8qVKwsNMRIJ8R+VuXxVebMiQd79hLiiWjts04qGUYdrh8OWVvJ4gFos54Kw/gPvaXuL0DYMUg
krQxDFEZ8pq7yuIDbCH2yVUzRed1ttKNo8dzuGEPQ3hbKGkDmuZY7ZsfAmB8/lE71QDq1sNjyw0/
L/CJ/0MJkPItDIlDOTqnevw50XGL5rOFUfIfImas9wP274adU2C9Ko+W/r6OEKcXSgvpoGTHcKK6
aqGdqzPnfaWuHi4PK3QL8ppGxCCjEHRhmTp8aPR2PwqkfRAta7MbmcZMRmP4az+V7EPXuEOkq7jw
IhE6kPYEfcNwK1u8MnCBIEMOuKEbYmAbUDH/vHaMTd13q9FkEujcxW5AjYD59mTpFhdDlkHsilGR
Oew8RLgOCtUra8pqAQ9WWS4rS6WVozsrItwg8TbUrEBmScXw7hgFgJs+XDDcte0cj3gkcgEFvygW
gxhP6kD99qNt3X7hbXXS97qXpWcDicymsN8FrOIDVx1U4cuJxisIhN4TayiN6iexsdtJMYD+KNBn
e3p84QE2DiTxsYjlUPbs1kdC6xCN7v6y14GEh/yUDpcmJe1dAMXFCvu7ceBRyXSb1amUqZskZhZS
5qSfpuZ1LU87wbdv3x/CW2bb8Mmh+20G719rYr59rkrtopHbzuniD7w2iTaW2vhpYmdBq0q7dJ3k
t0kp1W2g6KE6/7ehOWgNmrOOOuS9O+z6DWeB55ulOd+2HKCUfUE5FKG1S5wsJ4WJzpJrNdz5XW20
gwr6oxPynH+gcd/VsDUxQml/ku+HzuMnyQrQ14S+1U9Mrli6jdPCSrVvp2kXi+mRfFWdcbGdT8rf
+DXrnwllzBJlTKI7FOQSmetSxggXEcrpF7n5Ab0/ogcYVZtfIAy8IOvoSkIoLCmGbb1tw08gtZs1
bpQpPw4Tr9ZBhYZWQ2WUl0j6hFWpt4HC33irJjFpx/0YZOVv83rcu+SAd3B9TKdpKPhDk//JjivO
fPYYuXsZLkFNAopCBpJZMKR6C9LxuBdmL4TglrX5WruN+mSrF9DGb6G1MShq/bmgkZDv3/YSbfv9
1OPo092vtmZ3BibCLNTcBhFMeJ/gIH6HmOE0AtLktipQzK1hKCz96RmbklmLKQHeQBYOHusZbQdp
ruOf96mFVW5U1yfrM3fGSDybWUkwPDgKxo4sO0UutthaT3diD5uDXr33E2+kOLER0iTy8gvDdGHQ
FisqappJJ/OnaOfiQzvl3bsIvCO449YSDAhr2isszVnYYcBzBMx/b8I4bRO6H9wAPxl2mJhmcWe1
nBNlxmOEfd6ci5kXF9EKy+daX3+L2nEAVLT9B1ropOX2vqoMZgEuBEjvDvCCU9xnuEhvtT5D3xj+
ld97sZMvqC4IGkQhEMj8R3vxryKaREb2mUKhFwGC0tEzHoh3m7BCI3Ky+ya25j1FCdplbeUtSuYJ
DLa0Hf35Zh1gmfrY3fcS8F8xfk0DsOkgXPV5OX84d4NKZ8KiH8qHBVC0IA2EXdxiNnqQ4hkd/p8K
nQZrAltcAii1b3QCO++uOKfQmd7TkPZXHJGHwnoNydRtR2O0XXhm88MB1Uu+u0B/BLWEriXRlyEY
6etrrZVItObwTfUPoVK0R8oejMVAq9W1cW/r0a/IE50szCm79/Pb5fRQOlj/2FlL9MpYtZrjELpy
PHMYoEibtQ3lczyCMRuTju2kDbiHaFwZMmWuUBSURhVYvPyV2X4BQsGKdbiJpLJ+Wf95Q9lVeaYS
oZRFn+RH6hgvLZHaTvT3kHEbgmdjOWCa/qPEJ/S2oTuwIOxGIwJlPTxsEnZC14ssIAMtpLBVGyiX
MR4fj5ToAhQv3b7WLCMI9wEcmTzhLmAJ/0elSHVANvYQSJX/vmmV79hcBD13oRby0TQtGPgT4Q4M
KGsIvtRwKZW/17Sqj37mZpWWGI6NlRisJw6+o0SFoZFx+GGGQYnRdZgmmMV5sSF48UqtCLOGG7KO
UN9yfP+7wWFDdvXBcaeWg4thSSl+BURO8vSBk/53TvqJqg3zOPDxsZ3RSBM40hLSzCE2bsGYUOh1
Jdj1iK+ylcFoZV4rZsydHIr3rKCWlLXTU9YLXxbg5ddUvvb2sIjQpXvJ8aPHQlK9wCxwtHE9VIk9
1FYUQE0ah+JUfObtMQj6PenbQY+ipahhAxN3I5WrdnZTRxF+Gn8xEKjdxSVPOt++i/BliHJ++6Vz
gK/gGLBCtRv6dWjSXCHalpCMBjtEEIl3NqErEPMMK1oS6cj5vzVy7EtIMLm5RwtV0B7pTW64nxY3
Wc94pXgNPF06QTKhYHaavA4l5B1jcI9HZ7NI+ZndkYtH/tW2URLhV5OfvJps1mTuIqesGDZz6ynR
XxkE/w81kkzA452k0biWX9iTcB2G+hMlOX8pfGtbpmnZMKaCaSAZqLFzAPHu7naJWp7OG1erGxSv
fOmVw1TV9yfhZpp1ZPRQV2Jn5coCSib2ENVpMdrz+ZYueM1wM81jcN8AixAqBs9UDEXo5a4dHAXs
XWhwoqgxGAY22FnN9QQp6sRX3nT1ANv/lUelpPNRyN5yKZROCr1jgThS4sCdn88VaIZgeHrycUpf
FY2oAZ42HQKxkv+plBQYUeUztf/+y7bwegTYbAwzPPOXZorCo+DTFWvrMf1jRSi1+OsuIVeFBA6D
Cqs32Knlkg8ZD3qMvYX8LS1J4fgxijOCvild83mC5uIAAWPnUQe2MmiGgVdVYt/zxBK36CY8pd+f
5hMGhnv4uUaxlxL6l9o4sQA5689waBO7rCpoAdFQtJZprktVKy8tbb3PW1lk6p78pMLZ9JBs5wAD
Lgr4jB/YEnWghnhJNt48nDjde4d0Xx9sOtQP0DAb1hLJyLFJ1BOmqL59W6kOT4CKBTFefeDBBAK4
DDnQ0Fmss83aoAWmj9aSS4pN1BIOw3R2YavQoq6hzK1LDvNTEu7x/3dHXhYNXE+XBpNaVa6Ic40p
GzUseAWRb4FoNwMqh/L7v20acpi1/Hn50IujUW6LPdfFuNhHlcQee5LNVFBPFgDpKSNB4tsMK7cf
9H2Iezy8CKmBjbRDSRXWZJq4qpyI8jb0VGsk3dP52RGKsLalgaEa6y4U6iSRsiD1zIc94IoQd51x
y9nuoy304WIbf6evXSvE9hOm1WJE44zNYjGxABcSKfmEGQXIbd/rF6G/Wab0H9286jzi68TftFMN
t+puoS9Y/kt4VN2stsFBWcC2Ko7mgkJbB9dLlh2BXJspjClurzV0vNVv+5cDGwHl1lh+NK6uhqvv
9VPyUTiSXZm5e+oYTMKCXmHxi5k5RUjj/0ULx5fUJrHjVf06W3S60Ja9bTHAqWxO5dSkJIYNDyzI
vB+QHUgviixJe4qcg0xRQnJM5sTw4kEuOPYB7AtnpcePjGd7FuSbPrSN2yr/KgHlYXv/C5vU+jIj
qT6J0KKscLmh88pDssou4Ha+FN5CuNGTzx6Ew6hWr8buDT7MrGS4eH7cdX3H4yKNW8sQM6uhwuZy
VDXjrWufTLuMU7qZ4qmFEVCCF15nZjZhTrgZlf69Nmc81HYQp33OJToeu36YnnGqO6uxxV3gPOfz
BZR3epru1+i60+DoLOqa/+UcOGnoHYNrXhHUI6yKUbnG5VBANsDzdv8OpUnVCMuf+rTbbwXdzNas
SYhcdB0Volla/k/m+G0yviD4IFD+sukevUkrNdH2AewJwDEe/Q0SfxR/dmL8//mteTzZIKEs0VKd
Y/uUZTTYiBtlsTFnUFK+rAQs28873aqFc5JqI/axQdO3tuFV+jEksRz/PUJxPyUbNiBUSWcTLWQa
ahvk1/AdFHawemPWdYp2G88G/7fMRJwRpoS9+jzSRsI2O6AGKZjKQeYMeYHbkY4g/0T+TMJzK+1D
5n1eKqPoqrLPZSy36NUBjnfdbX85pvviX3XWnPLjiI6NJAGccUfht1FIxtP0IO/MK1xiSD1HPRaG
yvRDxb5FU36mvq/ka8DGTod1K5W+H2mEl085yQNTOpwr5f5s67jcJ1OPHU6jID/maKjjCZHZV27I
ONWyZRb6C2w9twfhAFTuQNYKf28OcAMRzfWmqnEfrZlcbmsEn2qvGF3dK7hvqulKLG0etgtS1Hce
N/65jqLLFKjKxeUsOcSCk/c8xuh6ojazECIGJ4XltZ0+dWSnUWtkgeoYolElsPAoYNTwiapK5IRk
v6Lf0dLqaRmaAOvWtAgbkvtKbxCUWqHrOHmVmgelTfLBplb/Mvx0tJJ5e9q6eE/pkKy7dIDkQ7Kk
//g9KstM1gxn8uHITMWwiA89csrBNWiGHS8MCsUB1yxjqjcPENOYO3h5N76jZyKmoZuJ81iRO1vo
1Fu0NpRohg3os39j0bkVAZtFYSIevq5w2kQmJnKlyFcQC5y9aMSTOPFhk20YYKWr5hsx+2R6ucV9
Eez03TyLj9dv256Xdqz3FqcuF2u0Wr75/05TyX7hu7lsrl/EoBPXlT4V0/ofChqNwgt35F9SIXFZ
EeKIWHeJZOj1p5RiIbaDRlGa3NZnDEJnoYC7ftAZ5/7VONktnGvbPCth69VPguc9wt3RTWmpQ0/Z
opvMhME+715kRPM2ySNEbB02WRNraXAeVJuPTZO269P965mMa2rKPLA77oi/beiNh8PXk66TLzEy
Q2nIbrnKo27GbPb5YTThNUlycB+esrXVH/XP6PIgUNt+wwYJk7/VnXhRs6N/8CEGDJZz8nci5Iyx
JyemlA0y5zmjy/41n6RgqUOA+LP5Dk/4RztGsvhOEOpB5Zilo3TLpEuEuUz80xzA/Nq/uveyTqG3
hmqKFTLwnSkWEEezeJHbfOWytfZ9er2O9QAR5E6h/IhYfXglTbVqI5xcyp44DUXaFWUTtMEzOC8U
OditnhlxfktgoXLzw53cnPrOAmnv/3ev1Aa9LgwKyRjdTnzMalmBOenc7/1on2uKy639bNgDj/P2
NWyrl1hWOddT/utE2+nMShJ9RAMqgoCvtWYXgcUjbSf0PYhmCIXiG8zRy6bWz1SHKgPICTziHXj+
azYquhcKnF3XxcL9GdLrHv1HQtlJfPZOp2P1KvKbyPIRlta/cUQH5hgIjlCIP2J+DQ275KvskEZx
QLdu5WCWakD+6gKYwz6P2+sXCdDS0Qwu98KjnTE6OZ+mho//oJ+vlp8xnFTidDIq9Oy9JESjQLg8
nyzQCMcLSkbt6pC8YuV5WvTf+S8P3wXCLz5+jmw6QAohMebKt5VMc3tNGT0bLC9SPXWLAwH6CV7j
/PTtC63Ry9u8UgXLdjmMN8UDOLrZTaHXY33hFTiDqH7zjN+plTef0QcF44y4qcXk4ycA8xeh/yOK
2Wpga8GjXNjwry9p2fOA0VOqNDvOkAmu/Ah9qWMv9A3IYCUB/0zHWVU0/HRcdeBntfZeu7GBiPcw
wwcBC4Z7x+5hUyBndxUsBIRzRujv843ztwnk0yYQUlkErXTjS0MoN16dE9yjCsHb41Vlq76CID0C
KlrgNjcWRaWyupD5P4sFmsjcMWD2yMcJKz1bHk7ES5aUnqjrnuYEOOKSmsEqQBJC695Zn2Y7xM7J
u59C07xegYf3rdq1exv4Q1uh7js4M9jak7jjpIoeEC/EkhNaXzjy8fCjf0WBYjQkaaw7AqWpeNrM
54FeVVZM9bSSLSrLRDCo3qn0mnad5KnmzYFda+4rE+8XwcJqewZTu+OGkf1ZwhWORVFrvY61QwED
EcrZdy82NJOoJMn2Soc2MOOiGlxH6JPI9O3EZQAA2MS6HOfeP9xuGwRdRSMxmk1Eb8LbpiehQ7RB
FPL/Hrtcwdgn/1LtAfGM1am/uAz/NzCK4tJD4AoNJuFPwf02xUSzoYxhD0FFz1Aezdb6bSm6Gnqb
CVn82WucZ0d2gqnxwenvJ722g1LQIJ5rMG3+xw9IuHj7aXS/b6OZoUQst5rmIbNZJHeywLHY9x+d
9SP6DNjJMlgSqxNoRAEGJ5jK5F8BZPFhgYvc1Sib0qtb+Nxy/vdoLvHq0OzagwnhQlVxHTVxwaug
fUbK/59rJYrX/i7uQ9uOzLZ/iGVz5ES/na5ryiEv9iluAzjexYXwhNiR4zyriL99O50q0f5Xch1O
Xq3XrXGTglugCzyJnCaP35ABqt8rXHM19As4eANv0vGq/bsZCO1rv2LY4LmuM0+K3UdnNRTzhVu4
aYvhkqV6JCUfvSEdFgB5kI68hs8zfqkrAu4Ej19uq6ySKpKDbLifecg89Os8rKoL+hEJ/ncVDQY3
3eVqhvErNB7P7FIVToeaWtakSBAJMQL9WyDCp2xaMs1jUqtPSoRk5WhHE9xcP/IXimniNapw3LhD
W+9kfuTXsj3J/iGUD0SrYw7jXlFcsOOhz7icbSCzv3zqOcHj7b4Nf6kdvO9tHUkx1DgU/hmR+GC5
iG1vJZRfN7ViBh7J/trTVDZOi9nf7FiO7Bnl4dA6pwZ0ge7nWgXAq2w1PH6wbyyp9EzHY0yleJBV
2xWCqCo20XzIlVlHNujctgQ6c65Q44CTXfVJRTm8CH8L/owDjDC85h5nlvbCufz2szrMeeoY8CXC
vNB11u6V8qu2ioDZCHFGZGHQkLq6YrhVCMKNLkwZz4xqVgroFpJyTKzF/09D2Br2gphQi8thz/Rr
DSUKyhLUmgVsu2hyGf0+wqAFsApoBlO99wRksJ9/9Nx5pTNl2iSkm/v/1hfeVyrfH4OKZkkMrB5C
Sf+j+0kOT8gX3ewq3Fx1B0c49K/7C/gBIYVKCmXxErG4f4kUITpQt97StRQXwZ8Yn7gM9J8NG/Sx
Prgl3j4pLathqpPVeuPBhyDPA7SzVy/Y53DcWpzbajhF5+OPiCd2rwlO3hVVTxzMggRl3mGV5eWU
+5xxi5OMPOg38lss7effpabHH+Ra1hv5trXS3UkdwlKdoYTkXIcs01zhbTkGFo0DYTAXrh+aGNrC
4U5Fe2jfMeIF8vqs8+jU8u2RR1GS47weYcvuJUpyA9mrVdGc+bCfajwqN5kqtRguql7TniO6O6/Y
stMH8zoti9yZKCZ5TBP76c8UUI/PS4sPFk4w5s+4vSY9YZQy9xvfMeAjviOh4suMrB8l9m/I/N3f
6SQUf5s3GoczUnV0+kDRZy4DGEdf+vLd51r6t6afunbBiUQ/M9jqoMTbPx1rzIfCKUNhE8CmRbZq
eTLM8B9m6RdJ+HTQSlsaeLVLOtL/CugK1acEv/sNdehQcX16YTUmycYTgGLbdwRC60MooouqeXDZ
UU1BQeCokdYOl0ld5zccMCgf1w41s42d0XUmk+YipqppG1dA9cyHcP4pSzp6dDLFrLos3VRyXSM9
oh0n86/5sMDuDSRTaChzQO2SbGviSHLYRAuoS0JlHAvUP3JZByUCDhJD82Z+m2RYWIoQe+jBu5te
X1VtVqCCrn3kf4aiOm5lJK3Jtzr5mBgTgIJ1CxHtPJ4ZJqBnSJHPLNHrtRiSVtEdZ3/eK1WemMJq
AHx3dL15DBm10PEal6N3l4Crd8JLBgO5cp8tG7PaTn7Xmy3KFzWbY/axxJZnHmFD+M9UBW2aJ5mj
XfNrFpp20j1geNgx4cjnt/o8yNexZwf4XFdCqCCmcxWEO0P0ODh5nEtJxbrTmJ699dHvIl9+TELt
AR3h5hhe4TFr1LpRsuw6e7AtvpJhKSK0LkEv3riB51O/tEHBsY0qqoWQKhgbodzGD4jDI2NU0yRy
eGlV1EcrLBdjTTe4nYJwJDkCXi7YzuoN1/GppHhU7Lf4pXQWBVhWUdSs9ft6DOw3UpnnZX8pdEvr
VH5zEUKBV0ZZLC+v9VgzrPD6An/vyTB9lwivUxBBO9PwVh4hcOTNvH/+Sy69Ggc6Casp3NWrE7aO
6b06qSzadH62ZtI+eKTlzxFJKjHwDimvfALSAycB3BNrN7Ybaio3gPxN83A3VCmUHna9FiG8wVKB
0sOPMMygq3TNi3DuxmAyd5CcRxG+VlCq8VMz2lExlaX8l0Y4FzCE/KThX7HqWdrwV33j+xbA4u/j
BPv9CbKmnI3bI1SXMwgnFidiTDMLGhxjl9/m9aWXFYFtDvDe2Zym4iLNvNmdlH+p/+tzwDS8Oy+4
BSVcSBrEPxm/SYsqXmnFTp+YfEeJ3/0mzlsemjc2yWDKmpQNyJ7PNFMsF8ydNlLUrA1nygc/v7sH
2psFh2zdW5rYRDW82oZj0urn9Ip9JdYu1Z6yQFovkAetMV7w+0cLyisIjN057pT+axeZysGezYOP
GpzEqtPpZQbMQkYqxFZKK1FLW6r7mKZdBxV9Ie8o8Y2Kcozj3qwFvV3FI8n73gCmJm4S3Tcw9ZZe
QxCwotfS+TeVkRo98nelSwDK6X1rbio5apE+CuipJFX8V/4rimgPhxZ2V/jq0004voPF330kCvGb
DFA3L0LbRvEiz+xv30bWURGLev8oB3RgPedTEFcMfqRS+XW3ii8C+44IQKthv7dE8Fa7+c9w3ngy
qZUYG9rxg7l1K8EcpzhJVg6W5ZxMu2jryLlsRIKtXEaA6UxdAQh661CGzGmXNs+K4FdyantVi2n0
ZSrWXCEPWhylTcs1oU4S0PgD+x3jV8D/Yg7nW6Fuvaq977H6wuAmZ1ypTCYj1/CH0wAfC+cZKxtZ
ax08KiUbMalEyqXtTgdpzN+H3z1X/fLOeab7twbMmkAhTftl2hhhYM57sdRCx9Sd9pEP4Q/lhZ9z
OeT2YSczKwlImsF10PvPawFsYN/2zcD4eC84pvM1228rq61OYN/PJRqrLuDaNgsCkNbygsW8goSk
zVP4o4W3MsbiFBrq+voJqXSGbKFuDQeST9eoMoCku4ZGvAlhSCJcHw2U87fot96tphbwxinNx085
PREF1nmB7xxKEVgA9DFkn2GFlWrgQxZKfA4OaQeaeyTPRqtPf0LtLzPzGVq9OpkIqh/AYT4EV6JM
d/pxP7ltuWN3SUtfzvauyEQhvZO84JTnl3QCSmnsLjcuLkejfPu72+AO9737Yw0WZKxH3NoVYCwK
3F8ki2bn3WYouhRPM9gSQmGeYY4aKwb/8tXwSquEfiRB8dcnLFZ58y1x07P3wLjdDlg7cbnKgwJa
n2OEZo0nSk05v00Xhhj/QNs2+RxiC8JgYCtO2bymDrS29kROcHmI5/NAUpOiL+l1lwjXzCZxvVk3
OQ1E9prrLjb3AnYqrrJ7SEd2bEWMAKxGhAtE+n4mlC+9jtTvtaYd8i6ooQcppe4gJmnAvzZ1SCth
l/GsJ/5B+QXC1F3XXFw4qf1cwMPFg69c9xKzjlqx7MK+o19W3E0a/r2Q6qw89YUaweY7V/dzfw7T
/uAGPk+Faltw85NfnpyhsHkKu4EwgGjxiNHZBOYc6Vi9Li1nB8TNBYvj3zerfYwU30QCr1XmWd/g
H1YBK0o738uQprTfkQ0UlD0bfqIskh/nF3hoywIyjvrBz4+FNlw9WaxXt/yTvPqZ02t+G5U8KrGB
LiL8EDo9ELoe9RJlrQYxWm42Q86vA6VynRELjoTESjuStmK2cXxGCRG6XCpB5tGEWCnvyVkUJ9iD
MOGbNpIJ2V/s0aty+jTOZk5VABairT8oLBf4Qv0BV0opKJ8zKNkhdjNQ7pWjViTDtVM1KI82P99J
110R0+/789j4ggz8B5y9V8KDN7kfQKl6PqMD6oVArXNJhXBGW5ny680UP8xjcGPeUtPlvTn2p0eE
c4iPH9/V5yMdfKGvWnwR5/6xKjhbMBLBGM+zBvmvkO8vVIEXuK7OlMob1yO5JHXDXHB25lKCx44K
h+olgW7cozJyXZ4WkBfNag1RxMN2xJGKU8WVziI2PozjCwPiNO7YGfp25HLAEXyaDey/rQDlcc5e
ICGdaI1BykYe8HsFhYXU3hh+sMPTry28gBogDRF8gR9lKajjddWbHJqjNwSrjPYWPzNx3+HiEJei
WFZ4td7H1zKcOroTVbxTKXOKmGN0DjMXKFLQKV2yuXy2Umbtd0dXxSns7yL9O7UvUYhtVvQwTfTE
PMGugk2M6Hhs8qyymW9V5Zl9+NFt/aHyX6LJZNghhUsy8av+XP5RRdqtkxVufqlyqa2LP4wT7CAq
FxSSedybI/n0Sq/kxS3CRzsWBAoEVB7tddM7VfYcg0wPEu6cLOApDn2rZp7UANHl5XlGVCdoactO
IKy5HjgUoDc9mwmgFDN8BdsI9CIoERi6VO7GSpcbQduSdyLOD/6heH24IyURz68PoGKno6VA7Nxr
En8mT0sQ9QIQvqcXg7nnmoIlKMMdYz1GU3BKHwHFsknafK4H0KyLzBGzcDp9fsCz3gn5d3sgudsC
9njlJxe3e4+NNwy59p8ceCwXzJL2p8aDGcg2/UtynHQSRW6FHup0JeBOdJhhaJiQbjB5IaCC65i1
KhPoIZALgXkh49P+nFlWFbeGFZ5RfSnHkLSU1I7JWpsgbT1iiczYlOpWMxQUESOU63hsE+aLIINo
I7CMByfwzMDYVIM30Y0hN/3XRc5NuSJZOKlrACxDNR+ft/GlnDgJwd1A8LbN1bA61giwLkcT6zx2
Eg4LAbvREIrVIOf1kVMf50hPDYt4AdQ5+q8tXwYCif3epX3PTntoefE/t+bzVHWmxJiT9RMk/+bt
v43vY61k8yynw0/C0XYUrabO1o8/Xea/fLoTzHE60+6YICqHyhSaXQqrdE9zW9iK5Htqm2Y3qRBh
VJM0xlhSXCIraPRb+Rr9sGP9saezjctthrR6LVPQCJCVA66Q76LB1zV1BsyO/q0PeNCIdMNfHpdt
w5FAzyk/8xYvT/iYyLZabpa5oMoKfdnPBR6qoob/YZXEHk/IsvQy1MKtA1N188F9dyYuBELXPAem
P0cnc0oVUmwWGSXa42xEcSsuz8GSDiHmdzle6ji4IbJLlhG8pmFJKNIW6UbrJQDXf5DkwR6qNDQ3
a68bKM5k+5IyRA7m/o+5Uk2jA7co4wQchpCQWbtv4br8Y3U1pI3ssB13ibJ9z/BjSXi9E2Jz0D1j
YvywtWj/iz1EhbW6W6qhFsnJQ4WcuNC+44sAPhANQG1oUh1UC1s6n0ypyBKsoTGUPYj4jzlpeWLy
bzoDN8M8n8/VJb+CPCqECDsEY/qtii2MJIxYjYdtyKvX5NhVpizRnfNSsDnfriMsu8hckkHDLBWd
cVvwSUQj1v9b2RwIzKiDzKgRz6CFT0dvbMS8cBMfdtwgxy+4ORdrn4ElPWH7gnnUKqCl6gejF5I1
q/4ad89s8R4UaIJ/BK0Bo3TpjjYrGO8A3+HnJ+UBWzFhDqovOQUFgz9PvNj3Be6f0rjkSDSxyktn
Nr/nnKvAa4iKMIqYIM4aRIhUPyx1ChkWdTaGFttGwHiphoxOKbcqRmtjMqdbHvXJr24pzaUuQPdn
P2nI7UGl82E8gDOGXfNbL7Sf5JmglFF9k5pvCGvcTwRt1hG9DekNx6LVwXGc05lba8VNfgPT85Xn
a9hi5cCAQeX8+8ew8WgrchW6VVYCTqiraSSE3xTa0gYNzNllj+znV8O2jQlMHemUJ/WzEgpCx9c6
TJw9m06gMcKzsZppIxDpyF1/8sPnxHLCA4SGXTxdAC02eLmVH3E1a3aJf/RSqNUeVQxSp4mTusg8
tgFvLrYfQ15ZvXim7uk1K4hB98l17ovjRaWcqVR2MFfjuHjiT4+cLK0dB6YbWBXRNZuChAPoZ+QH
5ZfjTsjtqbF4Nd4aPDrm1Gp08PczGh8rejxgeVffwWiw/+BRw42h+bw7y0bfEPX5/6pua2z7qqgu
r2SDFici0M79UhbwvUcvdMXZSpHSRTuBGHaJQxutpNCfrFJ+suCt1vQFeHcM8hSHVIzqXT4vOmeM
fu8MGvDX6w0mtyh91UlKhNMkFaNlUOQwwAFkK8JgOJxmNlby0WOC/wqIVCy2XurN18bPRRKnY6PT
4WFzmjJBwxG5Aw+71ZGa65OJlzvFwqDuTSz7Jdquyzi0vyKQaJyXa7NeGISQdd45zj3vrcpbzSL1
YlZzhd7JxJBxxskMmeNa/qq/oNkGsRuNn/OmfAnLIAtbLMZ9la9Q0HNSPIS/krx7lwwtnToazBlX
pVTpZ2UslI0P/plOZG8vAhw1A6xGGXJwQFG+Uf2hGoftnhSdqmtEIRm3kvIpIjDy5JyRYGKlCBCX
1mRp6z6QRuuDxhoCllHd5dK7iE9XIgspzo0QS61NZz7i7KSVSyBKnTtqU3XlmA3yC3PHFXUH8bCL
uF5daSEjsD46WoJZlD5VsgOkAwrVA+O2JAUEhY1NuvswEh7MfkFOJ2nbzZb5pNpVm9EIEvfBh0J0
khp22QFpLPNRmFWlQrEFbJRAqufJxLL6pQDbdDGpW/i/HkL9fsCTJpOTFCGizxR799JYVZSjsMCO
TO340pJ/X2IbqsRdWWIv9Br7AyifBurRdRK9m1zPZ0LHS+GtxgAkw8RSYYyZi6ELtaqjrDFiA2eB
zXcm0jiddufLWQlv1n/z7h1UiQ6baFiwbjofqFd0Oy16jiXKyxFgIJuizoKVT1/0uRr3fKMOUbZ0
kvoc6bBDQ+5TWytxMW4C2pKDmvdy61fsc/gI4L1RDc32mq+rAih7p7vyZGx2lrhpEqGjyvO0HkD6
3cw+vizJwAh8xHw+mYWv4c8elxYWwWYjiC6gMWMB2NbdYgIdTUJmXmnKefby4SGR4CV8YOhnvgJF
RghoLP29nYgCfoQBpZHvti5M0URFkPEH1xL1/HmM0FSzv1upe9L5QhNr6/Rnhw6K2LzclNXYb61v
RqYXvr072hupV3pDcGnB/1Pvm4qGrkjHrYZXYddw+NSQwQQbPGlB3VZGk5JY2ZuUx+AEFrxnOvL7
T/lutM4f7DSKdkEAFsXBt9pZ33/Q629vPzW9SDK/0DM6HbFh/K1E4Pffi3gvkENuoUmYJLQHHEHr
E6o2n0Q+ZO8LVdirUYSKIGUg4e/tobPV61sP+xGrgICYaMfnfQzVPlCuBmM3CPe1a13E/0UtB/9Y
3hRdiolper9lgMcXN+laSzYROHEcKXUtvxlkiuS+rnbeyXn3J/Tj5XWE0hJY5lFPOXiqQuxsTHS7
pU6V++9b7lDOxMEMEkJcto2k5W18AsXh7sXqtzZy+44B46Tx0L3lMTa55snxFntafnqge+1mKnEH
eso+xHc5n00aEwl/FVLA2jmXw1IlO8iUw8/tej+WiA8PlBT8L+m7OUvLyZV9HsyyTLJpoztQ5m8f
L685dexUO1PoOoPmNXAa5oDVndE+P1QayIIMI6U3oeksLBuOTbFrOgEeRZvmtN7yrKGhVnZF+tVD
fXuKewMQbl+Nw4pJKTCpLys40sogfIaPn3rPuIMg4Bzb9EAQ4QuJeDAuWAHwOBxT+ozdOiibry0S
5ZH4z5QbixpZkouZC4hW9HMI6qDulvU70+O0c5rjlkJSkRucAF5GvihzkSvw/MmKkYEPLIwwuGmX
qVmEhYbiXK+TxecN9gfrS9Bj3tZpYZ8GQbRk+r3K+F+RvmjavATlmEIp2fXt5Zz8w3lzuYZ4Ts6j
X1EwokLxGz2GiGJeQs7WcuTo3qsAi9bSO3RYecV/CYHtI7aGlLXH//Q5ltU5RksGWyhfbC7DFnCA
IJ+BB296G5x9kXNqzFRuxfeAl4jvs5cFkrP2kWE8CpOzxNcJJCsQoFvc1M8pXcjSSBEOVzTSmcCN
Ii7yQl1S2nGOvuoReovFCVxVhmwtDUNoO6VtHKoWU07d1sSdtP7XRZmTKQsOJFNWU39k1yf3nIfP
1l7rtBalqi9BswXRIwC+fJtWFfNIu1Z73qRhSD30pGb7vKqoqUhFDoar3G+KqYGWnAVxVQYVOOnw
SHpDDjG2CAdem8R3ssATc8/Hap5iL0r0iFVJyN8Z50gUuiFzNmgNryiUY3YX7q6rD1y/wwAErxs7
2iHvRLrCGNIP9Li7HHaruNmQyCCWd7XoLSmu0TWS2/JL3ddZx7vm+pBDozPGjNfrycm8dnfbBTpa
qKLzv5kRwqTimEoDTUvNBIEGJKN5GhsPYiKeoq2t8xAzjkUDJk9zf3ojPki1bjrUJ3WrFcXfiBaS
aCeDPJDdSTmOKrdOdbg1sZUUPMBclHJtu9SmDyECJt0BWvLhR2gGwuWm3nOdBWktmGJNrMa69XzB
BlUA0m0nHg+PN/35RrGMNz1av8cAelQwjklPzVGn7MWj2Byz3liDceoaMYjkIUiakaJteatf4Pwy
GlCY6QuZhcEImZRqXAs3XDYV2ZcOF1flWFEj8CzMlB7lmabqJHiuIEwJwpUM0E37EE/07nZ0gXuM
N8iDBQufbfxVhMnPWL8LJkDEbCP3WRGVOBbS1c7nvP7AR/h+GZkhHqW1NMEPAGex6EUwYXu2NW7T
n8EvTFprz9VrczMTu+1wXnFZccQmwe3nYuZhkVvOc/1wptILqBn7bAla3FwP1NCtXic+QHBbjuUs
tEpOyFkdvXh+FwFFTNPO+n8aT2KrV0ji0vRi0sRZe5VXVUbTRyXG225Uq0rOXw8U1iC7A2A9ySpi
25rNGgzfsCtxO8vtPirxAwRdCV97ioi8IU3LcyA4iAheCeLYMArWEywlU1ryijPhUliTJHdT1RSA
D/zxRk0qgayvQdkwZs2qMT8DtPDc3i3MP/M30zaFabCszVZSvJu2l/M1Z8LgUs6V6NNTtpywZXvL
hNXrCWjKE6JbA+1uLtB3x0g7LK+UdDMz2q0CQkw4Gzc8kHmED5GBbi2tXLIiFQfmhB9QFodFm3ZI
Pagw+rY4OWyvgGonVcnJ56DuLZKrGQRn6MqFjI3DxJP+qEsMFN6ibnH/qA6p4GgyKROO4bs85yuf
Va8oZm9cKXiEHKgfkXZ2w0XNOWJlYBA/mhRA87gOd/NXOqNi3eVDtbILO3d04i6GyHoQh26Em7V7
sSbQsOnR73dJz/YP/QS/mC6szgyhFDFBZYeq/L9QWLfRauJHwgsGt4glrHSwzaZZmRaiQ9RueyUm
RIpaD5rlG7ZJXGaw+YoE/rk6CH/auuTAzfhYNhyM+G8F7SNgpw19/3THIEwTzTyW1Gg869B9lIgi
9cOdetHkZ6qN/DF62qTOl8Fmg5Tug5AB2gueGEZYlhZK9kgK9mpL02nd4HQQQKFjozmpuD9cCDOf
oooTci98q5Pn4j7h6h49jx8CZ5kTKZW/2ZxTpuvXeUGMmcgCf8SBZe4xnaYF6eNBgK5r2Y6APcPi
PKQyzhzgwqm81BEBxXmkwqNNwOACosC4ru2KnwxR7P0tchK3xz36vXdh3mBcGrBE2c+29zp00q9n
dSQ8TYrzDoPosdFzABz08xD4OBGgK6wIrZNHFHCjj4VMaCKgMAUoztObobSvXSUcbEH520FsHRdV
sy4xzWYfEleHzsNl7dgZoJiWN97rCmwjhPJTz6Nl3F1/tP+R0FtqlDFv/3hV0FCiTx+eP0BZTQF4
wM5/hgJNH6S+zqUrlefXH3erecrS5PQbZHFwm/oYvA1UGZM9ubTK3YH/9zdVEeIs8abbKwt5TeIa
K+zJ7jPaw4XxXjh2n0BU67It9v0qaaARIruh1p6dKJETbvqJwXp6cBexcjUTJr4d4ilJJY4puKN8
uV8m0prgnWEnRq2LybRpuv/QEZNtXcgwiSNX1m3YeVDOA33iH7YKvmpppw2+lt+81J8ZGKSTxVs0
FSw2vzrXn62pPsT5QP/aVuZWpKhtB6SU2/+kuddCz+hcVTUlOxY55O5fQMvEkYa5XgA6L7gqUlL9
9CLlmTKLQRnZ5CKumCBwMVBc6DnWh1muSrZlmOfJnTxo7GMiklRJ17U44zQTFWXHacROWafUMavs
Rn7+KR/sh0FZxB8ozZr8ZynLPgIAB8lFoGxFzur77ld+m5+4MX7MQyHAauQUmDNETcLrGtH+9O4e
dsx2Pxe0vLY2m9GSZnC62Ghjw/eKiAti37BkgoJ+B3zrEdkEyabYARQb8Az118vYCdmE7g0bco+2
XmFv5Nd2/IOWnA5NT+tVdWXkEphgDR8XibdnUwps9JeJXS/PqBh8iOPN4AKJpkeUDPxYnUoC5sTB
bQHGZStjDWXUZlUI1j5g6Hf0GAb06vhluJxBVeh6HRQz1G54+51kLehzb27fhEwpup1ESS+09k8r
032nkBVTGYXsen/fvD23RL7GQ+Zl8E0y+oyMKbgih5/c86QptXbilpZHBTgpkkvmNQrc308WDUUH
3yFZuD1ig8Jh7ondLPHqkTJ3HLJ2eg5e25cLL50VqXfv4FRHltPdJdEgmoIOtECLjKi2vKAu0KwY
Sb0Ossufcc9ofiReM9FjbBKeJe5WiQ0QNFie+bdWjWTGBzvjK8kcls13DAixZa05u8c/xEcBrlzV
2VfOKeH6AMHyPG8Yop9YdHLz8x94FGXyezdjjdMrnv/VjcPNq+g6pvfggvehv9dfbTn0s9yamVvn
M8y9YKL72iThlq3dEMO5egst552hk0VUknktPna7OOIFskwTD/AxfbTXutvQUP78LBlIP8plHGLR
3EdKW1uppHyiZIjeyvRxI+N/Aurgq8AmWQ1tgYs/f5rE3igd//5pubQSFLhVthxv6Zjf3IVTS1mc
4pm4NPfus3bzEMqbogzxVM9mK6ev6nfNj6pLST3aLV8tvANr2muocZS3+4fHme1mX7hMTRoZt9Dt
TftYFwQEK949/TbWpLxnM/Emr1nW0hOG8RWgtMMs2/CznotYpU5ZpFUu1+YxvAarye4uzJ5DYdU7
gvjEHo42xHNQddSym/UNe7zmJ7ybrILjRnFGCkWvBOXKSmQC7KQJEhPEY2tDGRgy7jzcAwGmwKxE
weKpAVPw4bbCr5vocAWTmQoE4XZw2ca/XiO0lrqU5Tt+6dKn0n8O+xsk+Lk4jlM98KW9ajag3lqB
qXnPoJ2hrieKa2hSiK1dWOB3NyUdwZjR63kHahVNG8WCOunEUPE73JtjPloQesgMTzUaPGK6Bd52
G4dnUMTkJdGcJY7AXCSrTo2CkI3y0bvf9uUatZ8diutf/pb8ZK0rI8/b8z0c17geo8qpIFNtowN+
DTOhybc+v9PKhaRUjp8pbXcZdICPQWzDHHz2AaNJ8guPm0PuE89luHE2CuALrpS975drZbrSWKcZ
CaVSc4hCpDC7c4jUHt00uEpyIqNXcuGhKpc355qIRrI/aYYYdDS5aY8KrVkVnwIwSftDpg/06jP8
ax4SvegY1S19B+H9klZn17FxIxDzJLL+H4WoEGqP85+h61dbzOZ0VmBfIkwEM3rH43brC3jkAgu9
N4OJtIUPGXQFgXLmuiSyX0Jtmsmqpx2zmPdWDA0vsi+P2BhmMWWxfg/bC/PGF75yt5AKzZnYMBC8
GERa4v+w0xP9rFkDwx2dl1/l0LNQ3idoafXxVcm/APfuhXQKxnZ2yMBLu5qLf1XVbby/rnZ8CJ7y
8uXcd9XFXVxj3sztEK90rWmfCWDPcPENVbD/uNgk+zUtgUrWyHniRjRsHXk6NnIMrtxF5uq6pm7f
gmaV9XPR6rn6B96KXEVrk4NFxtcoUVFq2iKrJhmXUbyTu6zTQ2gphuvE/O2RBk9tFA+CjIgzZunu
1k/6duJhn9GlCLARLHASofDX36Hg0FNJ4vsp3XQcl8h7eFmatEnDxbttopJRKVwbG3U+cenp/2Oy
98crRHI5PNOkWzAAfCD+0NdgTyM2Zw4KQ+oSBTv19m0oZC+r0knveWg6bGZwyyxTqKeGRNsU96uy
Pdhh3mbTfqR1RhCj54fwoTNqRCOs2okHI29Xn6O2WUQydQjF4AGOHRnKRFT/kdzwYZSDw93PWV/p
4f0UE4ZeLnIyDr/As8N/C1UxeTyXvjdLTPcb3W0Pxc3s1YBD8iZliQH/K6O+/HSj/nSN400EijiB
L4uijaXj6bymFvnP+3Obluc2HkILthqG6IvWYUzdU4ak5yKEG9OdSIfdv1bQ57Gp1wgKEclVawiS
x7gp3xNo4vWs9nmRLV1D1abUuBx/VQckYQ6rXT1OG+RWbAp13CFrGvtTnmQA6+quNye32WkUGglO
dIcKGojo75v54ssrliSen+DccCEtW+QZOBph4Kis/5n0vSmX8KNHoL+Z+kpESwVlnWIzcFAs6C5h
58e/YV31SUXP5PNoyqUNoeHbN9wrgEbUC2bLawlObh1FhS/QjWhDbkPfY322C9CVuNhIliJ1oNFa
fxlBmceU0RjVnb+Yv0l4BH4I1ol7UFuKcyiJMnrs3UuT58m44YAKZsTeAy7EVH++eEg67ilT64Au
i809qg6xUeQN/co8IQVmrdYv/8wa6K09i1ZoaTVPy7uBqmNH9r/vMivmnu51TBmdYXHxKZMgtqx4
UtE9Tf0LqE6/Jmgy78o7jWEuxwo92L7batTdTZ6bzIQee6BVngJCSMRr9KtqrFiURtS2VViUT3ax
RD6l8quiAw8XKw0ZsRq3CqgSYjJKGGLoYjYn7m9IQttlF+2m8l1smi9uHgfXJZFG6JA/BIKop82a
Z67amKtAaT0Xp2lyrgLFEf+1lJ7ETS/lyQ8vf3rcBWyYqrViRRpv8DK74OPeHBws8pq910xFzkd1
Gr1MmlxpzG4HFdKYMXz8i/5VlVsltem7bTyYXuHD5lP3j2Tu1v347vT4EyhJAkepq3MJutFwjAt7
TELkQj3nipKrgjSKN7qTCb+UPxIWLm6cY5o8vZ9s8kwCUgk18PbSE2RVqUBVksVNmfDejCdbYUSi
rGEkNuJ43v77+3L67Pdw4aGjQf91AFqC7BTE9IysQaJPNWTblOt4f0OZOR+oeFdsaqNqOra/OZNV
VgjOpod8xOrNXHJHyN7ShAE/aWaqpx4V4azCP/iHjirF8KLCQueQ9PWnT/Na2Cu7qXiP7bwdjfdF
w3qZ8kX/wnlwRyxPwiq/G8SLFxhY4NAl8Qy51bS6rsYGiUf7E5mmopxow4voP2WQZk0Peoc9vqY7
T2MTF+hnssQiKg4nJcCsizBgHHm6hMvsN76yKOtgnww2p7zGKK0uB2HhlOlL1MpPb0QKCjtWyPlW
pZbP3dkqEXpyrOgnzmmIg4OxPdk/UcbcBmXyfDMQSuyhGeI2DXh8ur4Mo6AiIyn9Xov1v9cJ0Vij
24g9J1eJFq/+7ubIjU+sKNmANrjcOQdNi+8qEwJ5cdbpaMYeMageobdIzaRzMr7KiO51E50MVTCQ
6XQPZOGxHdT3zLjkJ+htLlg+sdHwqYlxQfcF7RAk/tcsA5AOivAZtI1kDttl359lEK2oiSJsWwUy
H8J910iJTeB83ntkajj6hy6bvoUmy94qm5Vq6PKDHgVcj7jR9aF6axOc7UTy1ej1BFhs9Im0mdKX
4d7Rns66R6G/URBVwxDpjAiOepdqyWI2Z89KaQgFPy+2k/D1Mv6gIHJPRdUHKxfIOFsTp7Gf//TM
mYDV5t22RBDdDLc+xdnnE2JPvywFXOxqkUQXJ/DjVEk5FyR6iwL1lNhZzITQmR3ntSnjubHn88QZ
r5aM8xEsg36uZYk/k1GWl8QUkxcFzhB0JAFmAG3WA262oBrTnCdvSLZ4RzGJD8HQmkvZxAzNJANI
56CvJRY8lCvb/isAcwvLNXNM85qq8F3T27vbnn1VRhhZz7p0YRarmDM2Rwqef3OKUr+iJsMQgyk4
QyRkgpw9K6QGyJDjeeje+PSYUj7eZP3gPnEifmRU9Ac6Fvpjx5fUSUrnzjLbLJgGH+ixOPoNPGJr
sWvQzM5np7vFEwKLsVTXKFLELvCFgjy2mQfhZkHsCrZtgAm6zlL/QRXqM+fbTGPcR8tD2x33+qb1
bzh6y1vZKEU3tQH6JXqaqG31llQAjgupqX/wBlw3GMWnkru1HOHA7gRnle10M2x9sWRMFzlNf5Jd
x3jiywUxluOdFCdywu0pdmN4h3cOpIHuJrXEgVwQbBZyFh6RmkOYZ+b7auElmasA8P74OyWAB2em
IIjxOD4VMgGJ4gZVIz3zOJwQkRKZNR45KXwZUWdqSrEoHdLJnv5zTIBhlIVxbUnQ1nOhICKppbpj
N/pbQLvQujEYOj1q6Quf00HRQMoKAoUsP7wcvCZ4Xt90OUhwZT5y6WY1OtibH7vv6dSQ515DFK9C
6ggqLhsD9XUYxf4sm6OC7q82BLRe17gGFLKAOaeq9LbzeUNSIhQaAIX43NIPQbXbROYQHxJlrQFh
mihCBg7aGkw2ABn2D5a3i818jvISQW1EJwRdKgg3n4/t2VY6nRpeeXJj9Kg3t673zxDRQHfwVuxz
zRB5LMaplljRnIrmC/+0SLyI+sLH0yuiMwrZIKw+hXRiLN7aUbi+XMiX9J6ZojOZNHQFiPh110DH
l/C7Z7NMYq8mGeEFnSQjw9sHWkmptERVyZqyMAR+D/VKMDFM03xt3okD3mCA9i96opA1XaIgd0ob
WW/HYiqz5gGfzKWPQxu/R0RBBeizHckAhNBErlbAg+7wIs+S3/iSiM6DHJfNG8yxIhOSGuq0CYne
sxfQIIKfg1WsDtM6BTDSRrAdgStBM6o5TVqYrdmBO6zNOhehJJio9EV6MeUM18BVCVqyyc27CGTY
J/Zzx8wAXNQqQamuU8iIaneNPE1fDILYzP5M/ydj4LUMYXk1o2AYJihK6NAzGVmHZnqJ0h9aOyAJ
r479qibclgfP5iwCff1RM++aSLtTXnZ82hfEpENUIv56WtndPmOXAaAKl6bc0qcgW4DFllo1+yMz
E05VFXekV2e8izX7JCIHkhfu/felHETaRfVykDB4gODOYuC4NtzBwvLrKzzpd8399lItFHMsMYt0
e/KT/5NXHdybFkg5P3BMqUiBV1BCygsy3w1joxX621oVHAUjeRAR4aE55zTdRJ39Quf7YsHX5f8x
14ojBJZ5FB4m6XIXJUKoojCCufryrbhWC/pFGE5Y1+Lf9PZD+UJWVpUxy58s+YkZxZ+a6bBt6cK2
rXdFlbzQaJF8oVl6yJnhIjGU/5Nm8fZQCqV53jW3i0KgSamklCSIHPHHtlvV0HMkiZNnTWcEBU5X
UTEFvn6h9MYzdGhXaM4aIy870VrnCr7+Ud19jKOZWLzhEgkhA0WyrtBlK5w87XRkGvnPrplM+xuV
sZgR71Ic6XxK039c5aX6zleJxxPWnqSd9EofzCTtTD3a8214MGy76x0CbjP8zwp0dD7crQdlbAE8
TNztifWIG1r7XkKK+KsU40u7HI6QG+IdUms3p1NErdMnxn8jho9OccjJIXRjvmEJFN0noX/pWN40
/pZod7gW28dmAcP70WzERUVXNNRdwHtBzCKq5FhQLUa+sda4FywUmH+a2VefmK3AMx91WLcmaMg1
GDvoYt2czD3yPcnYYD4Vchd675QCz5jVzjBSPQPSDVQjiyhESGBxxG7jTk9iIkhLvEvOvwB01zwG
MlF7Myhn0CMT0LG8R1qZ5emkF34HX7fC1cu3eFHTut8hgJcG4hl8wr2klk8OOer5xq8Ugq1u9f5B
RKUlEYGr+Rhjo3yFOiYpawP2mUOicFfOjUtxE+w4QykIxqhCL3PrY67CQydoPYhW7Q3QYUjkhmsN
myruA+UTVGcGJbwKaVRQ8yFaFStgKpnVEGqqWg4OccVDoT0dObRcktfSCMw/+PGC3Mc1bFf5DFuK
AEqolGHayD01jEJ2O57rev1eyYXjyc4RPbKjEvqLxsq36P2TFpBXSIX+3H60JUDrF3Y/FHevTrvq
BjBzTMWvIvLxy7QToE6xviCKKhptwf8ynx4I20PFasOi5MSUyv0x66yXvUjMoIdGdb6hfF7LfkLZ
zgGXgJVEuxu0mpFneCxxKd79g97ODHlm1lzqurg4kBmKmq0Jsgt0k/+fylixg4lUF/Ec+vmaolti
0gj5Coi09atY9ZStXUAUkHqPbfTT3FBedUN/lLIWj+VH/D6ipXtZTejXFBVEnVj/2Q+DhLsk5Qiq
7TvgXBUjlni4C1SrdnRwUnoudkD+Im3qYYMFZY0le+5ip42Bh/eCnGu5E3x5kv0XMmtIv0j7qvQN
9kuTq2mxfr0Up2BMI2qHKkP5I0j05KxZw3u1oeVVjIeoDhHZu5RgavhyecneS+f8kYr1taKkZV72
yBZJ/JIgCdaMvwyijIJZKVgNuB1hJ4mDd5DM+JTkoB4BEUg7Y2oyWPPf8UMnbolq1/+++KAtd9AC
5dw0JL8UlJijwspbpeS1zTYc94yZKf3pUfeCM0GfVKzwkc2TlD0LYcbSEt/UPrJpWzbOU/dQKf/f
6/00AFDtRt4HpQ19pT4EuqVpL1lybieD6Nbn6lf0UY9NM6riarH/hqvjDw+OubAofSjscva6r5Zk
9LUts+fofZvd8UeveJltxWyP7v7YHzemM61zEfk+lhmuGduaZFR2SZYsq4XJTAnnd4fPaEOnwy4b
cGHFJ39STxuV+rkSyCtEhl66cQdUeGbSd/ks71sY9O7QH0aUW/J7ZRbcjd3Y+/yoQnnPQJqxcOPG
MbP5uuPzbAmnXZmqlQQa5GtsTMs/K4zjYme7xk10TjG/QxIUfNpnAcfUMNDVl4ytzHNOHpZpDQOT
hVCwzlLEe6ey98NPHbQx/xDcOcmWpJW/tOnlU6hQXDHSrPPf/sZMJcTc/afppPKFjEDv0yPLGEQX
q0GgyKULDPCbsbJCUbD3HH5MCUsbTCVGVEt0s4LBqiCAjkQAIuACmgM1Ph1aEJ+hd4dfaGk/gvxT
5XMiQH9P599WlC5xzsV26cXkFfeBT5VA0kqe8DdD+elupKf0+J2Tx9DKY81bAYwCHZXCkywik1rN
VBGtdEPqTXjFksp3CIphCndQLQYTGq5VPi8Fbf4sii0yl8zFj1J50Zg4giXrKW9/S5ODfryNEFdt
XEFGbpwyaFrGvqqYpivQOfhTq5xdL1XbzY36/myfCMdH5gKI8ozYiIGz6Q2udsYmnb2Hj3kS+3HR
z0V0h+3Tha5PAa9mzo/pipaXAsxioGefidkY2itZ6CeWOW7q18wyKrPBUMccb1T8vc2bfk61raaj
3rFWpwGp3O7/YmaCVAmYqypOioePFv+fsKegrt02sfLPFLucxE22G5meKDvcUtJAtyIlvV/zZEg/
irXEy1NWOgRRqhhNvOiO4ibJGCp5EQvgOaEsPvcmXiarSQ4hjvCd6Vf3oCmFSPut2PDih7V1/zld
+/AsywGXhh8v3X5axKCGq2st8caEuzfEHYT0AKD7sJcPiSRakbLCHT3iyFp1XeSnrgBqQmOpZ13G
Bdr/8FFuI0iyzLUphfGjBHl/TPFLX4NHJOMvcnKFP7qwVQlWKzDPerJ4gxP92bkz5nfKMPDoWIfc
GrxyJGJidMdi23xf9mggAZ3F1HOZtoBEqBXDXCfYiNFQfToSPch/v9MqIlS0YuRsWXUYy5o/iCrB
TCbQSIwQGqp2v5JYoeEfP6n3/6XPi7ngqgHJdfaan0PEzsVe826/Z1Q3YTzBfIqk6EU30u6mEhDJ
2L13cZ0EwRmGNhmG0bun1CmlcyYYIp8+Vg5LJYGR9VuJxxUKptbH7kg+91ewzXrxierP1NTMXIyy
wO+bblooUuhS02UiY3s9srw4F8A6XjMKXDZKOED6u29369VM8VF1tYPPBGfv/Ayz69BrsguO+2Vv
ZncAherIQHKXOXzs2caHIy47TNWHBwJ8Gm8b6b5VKHFB3+dLahudjdtqFvbPvID/t1cNB0nF/qY6
aLnwQ1FYhFm5KUaRg8FiIex9I+KZEBaUgnggfye7XRbgHvIo3YhSaUfcv3DIkQOZCrKr0Lfr4pHl
GhDnCpiDtbZLjpURHUCcZCa17svQB3i9nk2sW3/FF0XFjiXwOmkw+RXzUtZ95FJSkvykFnoOoeWY
56tzqdjOrGfOCMny/cH/IvZ0Oy6EeH5+vu18ideSC4wcCl//qERc3LYwG6YK+M3jiLqcQ9jzsQlI
XvVWbweEpVA1PJtgoRXFN1q65ChAv/YB6RP0z1VpYn3/t1Q+u+kcfdhWftUbw2dA+Z3LWCrF6UH/
qREhildxcks6ZnRCm0RHsR3sNWXZwd2O5mm1t+aY2PALH4uRvjjZu7X6+NucxVA6fAiTqEvgekgU
63GZOjzowfs33V3sCnsK14+0HUSfQPkiRYJi8XbWdvrIVeK7KaF5mI2bAJb7paw575cSWXo1fTXz
Dav7WzlBgqBd8wDwy1jcwNydoGt81olMKIa+7NWhFmJXqLI/sxrDAC6427TjBfEPtlCe08sX0FNJ
JrHcL5Xx91LL2Ul5Vw6KmEnrszKdLnW0epOgK6W4HyqUbMpFIykt1zMcKbZ2rVMjuEagD8Dt8iH9
C9GM7nD9xs5hzo2lUzPWuA6pKt2HTpogwLX0tJAx9geDn/ZcpQRmypCEJTZeW7xN9bvLLCaH0DcH
48m2YwwNWIPekcgXf1apQpzxAOxVhTvBHkGLKTYZUHvfHu5XAwlqo4bUQCK6Cj2Qpd/+9Daa0QQy
CSJ4E1HAzLkeaX5r4umfMbSRlSYvVVsDYoFguuvDbpKewxueLjrMGYmBvPfOwOhcgoo3tFNBrty1
b+G/gwZF7wXfpMfCtQ9fKhf1aGt7MOOUHMu4vZ9LA0jOM8mO4SkeO7q7KpxTxEvnq1nKg3s7OYVM
aLcAPHJGzCXh2j4bGXyoDBllAnDBcAI1jH7gGeRiaSoM0G1q2bNXhD06equxrAKDTiUPdHcWQLkf
Nxbz4UyK+qlDI3ko0+swtblXYROzH5BXBTUPKuUHjKmARsGUa03C6FRmXKVEsI0uNZwx4/vsCJU/
qotVYBBH23N9UtxWE8JPIMc+9ddWEAXW5m8Cwnyv6sbTsqAUEV+6yvfjXfqgRmu73lZOFMEknA3/
Yr2pNx+s7drshJoywGIMQBOECZrCNdfQD3CdwRQ055jcLxsYuHVV9Dxk6Ebi09NRUs/ka+GhFwJ/
H2DehfMms41ZEtwiliHYp5ujMdC8TeAy2SYQY6PUVt7LE8K+VOvDOzQbBBysskcZHU53Dn7sM3Cb
v0BoQSudwWVc67aztgR+BzL6c0xLczBYMpk/hsIPVYV9dTyERK9YTyDPCVehct6xBE8XfrQPa/6x
+4hryhJfAV1zt+gwpyG6ta0rNKdjimz/N91g5kGdyiWr41tXmWlbBSPglwkKBATIVYkjpuRyM/J4
DhucL0S+G21smhXAy0DWfynnHTjH4nNwf/kdVPnuoiS/y2iD5b1skDd4AT7Ii6FvwyDtMBgTd8fo
iX9lVa0ch1HKfLB97DysYoUrij7UFw7f2bo93pWqL8u4X/FxKIKq7iP05nJMqsVO8tUdGmngVscz
lnu3t+rkLaue/yy5O/wJjEa9Awqwcn4ICnF3pPyJOZb27QVbu5ONp4+6T3H1EyHvnmRu9ujpIR2b
tXU4GTwGXij4jgCK8SjWErucPLq3SZ9AeMqC9y/d02KpB4SNbciP3I9HgSR5B3w3kri2m9y4a3cU
ilW2G9jPtUje6P+0+rEvH0EY3KO7dNvrgs6vc4oyTMiQPPX0CET0T1LXYfpmR12xxGgOIIt9C2Ax
jMg344dyrPLvAnxq6u2Fn0Xi/ZsZbtZzckmLHgOf2+Vucj1bbi01MluRZF97R37gaFfctLPdSbEZ
La53QV/bWTQ59P0X+z2aap8T679R5Jg2SSKEAaj6KTewj7nubkylVxiW3iGz2Letz9JxiFs/tPVr
/KULWKJU4xSllz2gjzPGTeIwwF2dFgwKAn4Uxby0IKWanMRDpOStU77LNtfCC313DMdRb9x3W88d
Alk4Fzpk0Qwqg3IzTrVLM4MGzFPVbVBSsofp6HQA3EjGp1pMZZLd2JNiBDJmM/MOYzD5/mB8jwWt
qf1Keum7+aiwULCzs2epmcsOefTiisRmcLeIUO1FSBLjmcZp4uviGbtOmc8rLLy6kpz66hwwuW34
WSp9TYbICElKBIkiKrroU3EbFp4uwBL8zTeOMa3JPsYfOfgFJBPoW3NHBUFvxZNg6cyBiHEoYO8a
Em66fs27cVm25jIGRhRcEkF8sJHtSGeOQB3GN6Inc9pMayDrMVKrE1Fv2Tyip4hKum120zD2DYJE
D1R8SDPzGyLTFq6OAR/hBh1fG9qH5aRATW4nHFfVMt1bvhQGo9L+btFGKM44F2GZCIQ93SYZdB5C
zED7H5AG8T90NbZEGm8KH303xy74k5dtVcRI80D5iwEiY5MeEB5eeq6xyvxF/gYVOegvZpKzftUQ
I/5ifgL1Q+HQmGlOocoB7SWf3t95EDwFnrVAdGu/1QvfwqyuBsJdrAZ667Jo7OQTebQaQr6R/kGG
ewQNB05xrU+86iNbqL/UvWMkJwWRI1tgUrxQTZfS+j3q3DFbtt4nPvyq6e4svL0jOry9PjvCfjJN
+w8dk+cgmTUiePKF2yi6xU6xfVxTbxC6D0p2GTvt0/mcfbCxCu0CfGyn+hmYCvScwUDmRiPpfqh7
Kjmhrx/+CZogFUHoAz8Bfl5OFMAaZNpkc4XOIWIKezAMFsv5xGyb+dS6wyHEO0oOW64MbxZtXNGf
N/s+jJZa6Jma8UPLMPmU6Q2nJZx1wMhCMmnfC6/f5TTllKGVLhmZtUP6mSm2xv+cLH4kbmfadfj5
KvGTD9IBkmu6KrhEN3VbvrO4Cv/eriRexmGEsG9xxKbwZz1F7TQ9jQ0K4eYEIiH5j4N2MQ3iduNT
zbljYhMeDse+NXRbtsG6XB3FaBKvnwTW/ypoC465CRZUI4+CPUl2ovJSBCEvYzaC/iYxS/FgHnN3
8OHUSWeaMV9cHtJAw14MGDP6rkyDUz5pbS5MLYDTOC0QKRHdRko2oIXc9NrIsD401r0wTDwCFp+w
AxQibKlWoClRnVERxEZK0AStrZ7sG7egJQjfTsOPKvFCIef3T7/8xxxTzBGeQR1OzxJAMPaF/T8p
Lyr/QF0TC8P5NTWWMHOX10ORhI54N/Er8fNi7Cm+lZ418+pFrxB/o8VdxtrXxsu3RidmF8JxmcIM
tXeX2TtVBoOSBRzJh1uDpDOfuRCHfNkrEJnRQzeZCUPRehuAguTL3YV0lzgE9sFDxDgW6kxPQdrL
GlrlD/VKWuoK212gDCWgnDLJkFexK0ed2KJAobDee/VrizY/YYfn3fIGh/TsGrz0etQjgZi01LaH
7eceEC71YQgRvZOALtinOcpTzZapXaOb+C5dsZfmuFoOdg9v1GQLMArDKFJcfd3RNR4xTfp2aPAs
PcorTtyJOLCoQF7KbN2kfaZrEJLWO1YXfHnlHf7JmYOt9h7Ri8grBDz4en7j0cYo7nrQa+okkf1D
nVgf9mBqF84vR0cnpf1jVizS4rzoYMxMbKJ75OEJlfJ/2PcQDp5fc+Q6VtSpmBfCqIa+a7i3nFkn
mt4KDS1AX7uChFDKCjgU0oxHvJoJdna+1tadPh99iY/9latDAke3ZDnaOKYuu5LiHs0hdzIejHuD
wnwDQjWQKrkS9EsdZcFFkUChBn9megE7KeuEtMOnx+YpvMvKZ21CBhL17YjkmhFp9ZZnqci2MkKC
QfxpiJi3bGl5oieGZHLizErxgK2d3xbnwZxDVLbVQU6TsAUAIbhl4tIQbSi4KnV+QOAUxDbrtWnC
2Mf+FOWY9XoDhdoUb/qSioO1nREvL9uh/yGsWkhY9dURPAQCF8EmcACVfAxd2Dn+RaCYmBcZlCj9
MqiMkW+JfVkcJ2x97lvKynzJG2sJiIGUSawJ+nVJDJChVLeCNXq5qlHSJEI9VCPPbQoHA+b3YRqU
Q9xG6Itbkn+G0QFPRJxfV8ktWW7HCBA2H+i5iBcIVv4PVXdSfihP88T8A6b55FbLw5tyNtHsgpaa
ldqluTqh9U2z3zpCTbmONiQoc9F/ubgk85DehNlIGhZWa8rNY4cdREBLeDL/+bYIbiEKmWaGNUX/
5MI0izByqmf4mXB/Kyg44RC4tZej5VCprI2luueGVlLdDAOJ7SQ4mOyhJgl3o31Vaj85dF0Ovful
zJdPjwXodop5vzQkUJ6IzYz1IkZ+MjbT2CH0TjclwrxfNqxKBHK3HGtIp6caVO7ZWwYeKlw2Q2DI
dYYXg/AFnq2DsBP8Q7PooULw/5SEv8/pv0wcVaQ0sgc/j2f9WSc7IzmctNYVsdW/GZ6Z4CWTQVa6
w99rBhbRfPmdx8BXl/QdyjBpUwSZO1TisdPgYkzVez5HiVigv+bTpNrTJFuhIbIirWrFQ3GrU2nN
d+PA7w2S+ixUHGtwpbXqFnjVe+qYPzOeyq1ckKTfjK5jSPnY35oWOjrmLJalopeVfVBA0URE14pC
QxsJ8qvMxNyZQGjjrV5fd98XYywWmvVzxM2bKaB971TB2fOCGe5jDkapAl5oJZ0o5LaL7P0+J/5r
nyuPBfBg3aFR8FINL953olvViInGXhN0lxc0VHsV8WbMf2u7Rk7oaMHbYzNB/s+QCOrIsfAmKV6Y
d3qIefHQKCdqbLm02XUosW/Ocghg3x8a7m47nQ8ZC1etHtpjvR2SZe9fZcTyTsTw5YdX6K4BpQHA
wHbzvHkKyCFh2kCdqrMIFSFwEcUz7SYimfUoESxja+WT1dve6GQ92i/MnywQu9vUwvmdIWOe4PcC
EBcPQ1iajgaf030vc6W/HUzTZ/h7DSzS7Vggs8b5FtOv7iyMcys88S+T+Rqt3o+drZ2VPPe0bo5n
Evf6w4ec7hVldRDI4Io92YcRw1fHzQ2RNJRjKZ+Q9DDFB7myuNf4D36nCUHW5EK1u8Ljn0rN55td
XMjukbKpqE7UUZuKcPKCG7+HU2F1bky+S4uZUlKfISWuY/WRJVRbynEEG8SiARd3lAg2GrZZLcQ7
U+okgwcMwspMrf+hNVj+RE5ZrNy2GTe5GjEAH9V5yvCrFVb74r0gsvSozmSQRsRwhIxl7RhXdayq
BD3f2wS/d99WokJmEo0ritw08GKMeHl/esUglNHItDKcRUOhKO/TW3Bh3YXb0WNAtWT5jcHnXiyq
gTfoH2OTLVd/WlEq8EmDVaNSzy1pSn6jvUVScKvtoRCV3WtBSrs29BMR10Id+zE6AdYMv3/b3ZRX
RSSsaMpsBTCACf+JEjKYpEP4q7FyTu7mqOTo+sYaXujJjj6p/0KHPS2b55jEho96wvJIlu5DPHn/
OInCm0u9R11WGvjTQw0lF6sqkDAFyCVkTKzAuD50Gc05hBH6YDUHMuw/NoBicEh3KAMA2bbhiC0D
CJ/UtZfmlOJlkzYXAr0RDZ1/5aKfOUUlRNO6uCakTqGuPSHM4307OM2UCP90XFaTyBQk9sWjM6au
W8GtKJsVqE8+iK/N78obmr7g8O9y5iTR19BfxZ9YWEGA+w7lQAhDRHgIg1HfLTSefLiG9xZoovXP
3WV+kFd5/9WKKd9WJwd3nvkRYXFora11S3XsPt8S7CM6E2vyhqlo7C7XWCbSh1tiejNJrmymiXIU
k1BukMPmD4iObe7CKe1hv5Rr2FI+E1ZTmSn4m14KauGUJfDrglZdQZo0plXfCBsAKLHF5SN55VsS
pPttQoHcxtR8PTmvnvqwvM/mBf/5gSVYfuhUPhvJvPMNgbxOeJi4KE4fW47Xju5CDLofCE8xfGpC
GdrfdCDJ+LI3FmJ+d5s142c3JwkTLRU1TFTZ4qzLGM9WrXYC4ab8ZJKfpr+Urz1R9eUJqCtEpHwI
XlQ88g2e8KhdD0beD2BJsjaRePiM9k3pySRFQQkzTwsbA6N9rUbfozIjo+jNwBBDgTM4QK37yljs
T+PCNW8bbwxGDmSd+MuxTCpjl63iACbkaiGJ9/voYg4heqI8qxL7LxCqxaPXmWg29mApS3V11gDu
1q+Ax6M7Hiyl1qKcRHkLvz/VIz6/VMKx1cYkhqhAc0nDFZ3SC17U+KTbXb2aZ+4Kc8QURdp/AuJi
dhg9l0iH5C27jTAHgIuCHmHaBiBjkTkz94yEOiYi2QzgK04cQLLH/FDWbLtCV3656oVHu6pFO9UA
s3GGrF5qLGR+LqrScTDvVkKFywV2jYpm1wQmjiPY8MUZ92lI61KbXEody1YcDzhWpBITCNkDFwEo
YrUPPXHbRyzODQHe4BxEcd/+ntxNifkF/grKWqT0DfsSU2EPeusBZw/RgarhcmGcnLS/0r+PZcC6
w05kvhl3DmNjcSXNuDevo2db4LBX/3TxSfqIj5aeAO5AbVFMYiD9ozhVi02rtuac2Fy+e4nAYDMU
i5wtDLQZF/dyFOhQsxw8MmicmczgyYsel4LtJuU9fXUhkuDAYhqiZctrZ33+bxyM1HWlfQSYpXx5
k4osHkoEYLOQTtJV1lUIT9JYMjHtGImDo/XLZpfZwZwRZlWIxy8PuUI820UuB0SmoAvsKUMWCzYt
CFw1B5TYVfrURCh0Sm4H9hSX1mHcQ7S9G3rzh9GLNCfZ2Ke5UEFb15cQcVPMMj780pwFK+iwUJKV
uyre/tS0b0cfJAKZqhNcXGjki0hxI+fOTFPNfU5v5RORGCmaUP0UmYr8l9SfE9N+yBEmOW79POBH
EM0sxD0OshQ4Py14uLwBMdNJPfJ/JaxHdJsGh0zdXMHoOn4TYNFlBp+bq1GR/WW3SaG/U7XBQZiW
Ci7gxyH+BLPhdYQ/ooAvOeuAEnxpIgv9Y1/MZRQV7gORUFTGQ6rmT/Rt4VDMgNRF90+CT8IOJ5LE
yWsshKekZwDVu4LcuKO5coudQ++qBI1xF7QKqkmUakL/aOkLkgjikZ24UgbFRVr3YjUBpWBJnM41
gSVrsjHI/edON4mySNodfrSCF30CKc+edHtr7qSY4Ts+EjpK0WfpSlIuXWcEcRj1P8uVPZdrxMMQ
3zqx/9TyZIJl1cT6AwlaPsQjPGbtQQ3dF+t38Dgpn09hgIIv0Bu/s/G93Y9BVKG7SHtCc8Vp+MUp
2fkhD2DHAoZcTgBTLzweD8czwex+ufe/xnvesaxkukPQOA/pofx2j2+Q/koNSUAjoL2ROvtNGIqc
ven36/R3l7nBY7ACHp4TJA5YDzyyWW9wcV0pPWTeXAAxbTLqhKk8kojQnGzs8YX9MhaU2oguapjC
+rFXK4ib0ynRA+ukonubX6oDV3PSfd6N7jPymyHvYuRgy0JylvAlZ8Z+Ga4a8fKpzmIs/G9o5JMa
dkjSn/e2RxfZQm+LBxTDjPn1Rw/pyHZh6nyeLzQcP23aXh4wRWAJV5h0+dGIpU9gskCF3/Wcf62l
csb4giAZdJBli3StSudcI8rbsXreYwdQiXQlHEvdM/PpVWdEtlJxsPVUdzVF2upv6zPb/r4IaTbN
D7LMfNuNwPcrUwNaAW5R8dE35FzNITVRDhPA6SrDQBaNPUbMbdEFUAn4ao6XKZCerfj+Yqr2zdr/
Lzbp4MKwGhUF+yA3mcws9i/3/F2lB8OXjlgZaozzl7Wz+/svkXb5K5spNBkaFeIq7xRw4a/2L4cB
zXrsoyN5c4QMV3EZeiabzC85uF5zI8FHZ6uucwV+WFkGlMSSSIjSIyZ2udThGEW0JgvAMsDgxET5
6j0ID5do8GUq9xbsPBRG+5I5eWrwIwbRRfsi8wzgmP5Ko1hwH+h1eSk32ZVJKC9mFBPopSAku+Pi
ISt8HKaJEebQ1F6cZ2Qg4ZQ0PAc5dJbSmwx/k9mLYinQ3dcvAG04ijUaKKArisbVxcuz0WZs8s3O
SJrSSKLZeVggLygWpZE37MbapeffioUk1p+g/kSzEBfVWnZHh4j/WX0cMCbyO3ytRgwPg8Rp4CSp
vkL5ovGmrniIfyCbtNL+3kf9LiNNd3DTfQe1b7rfJqLDL077X/Tu5ZVRcMYx6drwjommcaeEYQrg
f6OLfGsfmhRNtY9pF29TduWlVtWaxQnYLB3MszW9d4s/rni99fTxeXNTDWcusmrZa0D2RRr7Wc49
D7uzojHxaMlIBaT3pGXc3a2nSy+oaPIfNp9YwYou3NqDCFTT6cp29P2eJttnRyfkKOge7gMauYNq
RIl2xn/SHS8KWuiHMa7CZhZq4O+e/iznUhBgmbMBEP5w2hxfIvjhbpCUpcIIasFQQ0E5bFVzEWwJ
gT4lDHZ2oLwaDVmW3XUcH2SiApFUTgUiD43qg6GzPdIHXt8FgJmgGoQMeYFC4Pvhg4YmfDH+ndGE
MWUjENdr9OCPLZcTaqURetC1ZbK8gFPySxYA6rStmfMbfj1erBZn94x4nL5Tnqx5JdzoYdWabXKP
T5V3rpVdtmGr0AAd4o6dpidrXhZgwdGpSK5xV42UaSfO1kyRQ5bUAUn+3pYMcKHfAoOpaTwrbky4
fjXd9srAHbpshUTESXJF4Pz0z8MFsWWx5aAttmuNgDpuqKNhmyvEkRLiy2cMSk0i0iagQADZD/Ld
KOjeQK53S/nEn6AKylsFDrLIA5l70UO+t1WJDZHSt50Yh66bRYdRMJWQHrGLMCURTxR1Gxqs6QS6
EpqXmSuZQ/j2oK+5TuBoj4PxAUtMTX2XMjbT6YbSi0ZVXxJjXrunJK+o/QZVIsVDuf+zN45eMaON
dc2eYH7MtnnVNdlbu7e1g5P/n5U1kEAtZTvB/EMX8AqbU2Zhx5AZaGg6Kase9h8/Vjms/qWy2NOE
RDcKnxK1cNLnB4bDl4iE/RH99XeI5ugab5qoOuEFGgyHXmjlbC6JCtKvJWSJN9T9cv/Ep/WFY9V/
3t07TVhGWgklmE2MyftDZSEw/SSB/VwmtFuAvQEM0litX7ZRiHcB40iP+DNsiIvYfxK3bTZvOO5S
FxCnDOW/dzEx40G9MIYSUyx4YPFWTRWFiqyJ9vZ3X9+eAYBMwLR+oSsM4jj/iWWOk+6JnzVkGK9Z
KiHhcmz5j1HjepLYse1sOvlBlMeJaQq/lKqgFPVp7GehX74wfPea46n6+xZfz8DxqCnTDfJ2FOh4
874RsQz3Qoa07SFtSITq5mwQXT7nVuMGhhjzAmGKZ9dzW42xIvNpGbRyzZTM2E7OKH0/NZSp932k
5RIGDVMoiiXmjobUd5bX5VybUS5jaGzAGduOIvmngTxyvc7VqAjhOmffgyxN+VoSTNMqwFEeDd4g
4RmVL3K/mxOYv7kN46f2yCAre9FePGmYCr+YjzSdJmHaR7+lrWr8xliGebwhkFoKZyvpT/imNhY6
Wotd+PS7lUJb3Wfu/IFszc+8RnTz7/I5xddGgTrw4D4Xoymz/1xy4CKb5pFyMlV9I74coNmqM4mk
sros8gD03NC+Lg4waIQXiZNcp+FM99e//MNA3W07S9nZMwtPIr4OCj95qgH2cJpID0e931F3kqoa
cSeipYoRCSt/d3owLSJL8ybcje08tZbBCS+2wIOBgX44nMo85/wzFJB5Qk+vhv4PITEg/M8AqKDO
S31oOGTVLoAPIHm7CbGp7LoK02BLw40+MGyMQqI346eX1G0Zae/QUQhtBkZvTGfJxz/QJoNBGmbH
AlDgHMRx764K8juKhUA8s1JEDxgo8ocjhDYMk6r1UIExtzt5PrAAvNrKN2PHGobzB6mHK60uiXN1
QBxF+Zu5qc5xOk7RIy6pa2fc8lmpKgnFlV/IwdPjWk6V7HRbbCAW8u2U516TW1DZT36FOTY/Eh+i
UFG3cX2+hP+abdagNpy8DcmHd67juaUawCtX0FTPQ7oP3bbr0tAh/4885pqypnBem/jmRlgqy/es
wTSefOGhbKACQz+K11vNIRQxi9oLypfB0y1Z2kppALJsIF8U+7yHgV+D1MTkJvansWIhbAjOzK8j
HcCl2nTHfpFMxEsMA/drbRsrIRH39DF3aiefnqbj1Dog+2/m2qCleo1NR0Krtq1mYRKVI2zAlO4C
b9725o3vLsLsAZYN4VZ/zR7oJ7JldeAlmQoq8idQq+xVTCe04+HM6Ifz2p0LMwCDBnX6bf8Pk2yU
6HRaTCj3jvRw/INIawpDwOmDLjqyte3IQgc5NAER/TUnZ8m3Tl91QEBrM1sH+dt/K8+ecPfKNT7J
dC0COB8vwm8DA/H7tPVjzmv2EOrRbqsMkjZncERW22gsDV19WPbn6xyc2GsCElVmSjD6NcR1p7J2
aPhsQ3WQsgyJzCT6KFs6M9fGU9LdRLJRSInND6Ct/qPRiTBltmuSICVbmhZIAcyx8+DkGTxBLKfn
cpAlQjH4cfVJ6l2vXayw9qd56m8w7n3VGegTCvP9ugBSxjn8Nu/ox9tW6ZkJl/DQ4f2zM5lRhKUj
fTDaoGovu2fSZXn5kYFQbOnQLk3mWzSR3i2GSaXpwJHxoCTghIgSmoFHoAz3Ik8fmP84ZRGmBCUW
MQPv4uQR9g14XloPxW6Ggy0XO7SEOHT3W7FdIvKttnLZrFQ5uZo9gfuXOr5PCj5x8rw1LqOvqafl
T1FeTOu/6ZgFAgdDMk5yi+nDsIjle5+EIuUQfFtk4ZVFA8W19G/tNjHQCCYwxm3ZayIlsvK+bFGN
XyP0007byjMysAM8FsJrhfjPenxRvcVRXqEAXIcy2ABH5RnVtd68zvWXOLhbbhcsjDRjvq5ekZ6C
WCcpeXO77eBmuehKznxSo0mOyh1yatW1Oy7dte9olS7Dz/wOObpFdfGbuVf79vFXNXUTuwXHcwfN
1EHPvPUaZAcQGbCtY0deR+8/gtNgl9+oibxjUuQmFdLcReDUfreVtUR3OGtFQr06onTD8smG4AJP
O6wNYxwUdFTcorzSX+Y729wAEindTPZWAP9SFeGGXlJDev+i2bDGTs8pxnEzj4MypO27N+ty1kZW
0NM5a/+ZKLYCHgiElVQ7eB+Cqjjm3W9Bg7TxX2+yaB4tnKcdYqiXHxxquIN09xYvPwYmc1DGYmH1
3F7dVJrXdwZWrTXH7T+BaMqhXNJQaSvAVrVioX+ld/I9woUat4YOL8IZlKBEl2DqjF9Vr3KiNfyh
o49Et33HigyevJTXRd3gcQ06UXdBj0E6Vhe3eHBZNwj5ClWzjmFU/qY1Dfx0zvxNwJylcXFzi/Uw
rkeHMLAYa1VKkBCYyaMqJqL2If3O8ypSz1ksARexj7wHIAFx12iFLIqLugQNgpUKZIMNpRbkENvQ
f8T0GD2ZA8Sv7+Sn2abhZlGAEnWF7CqmzaKCubcgd59h4AmWHi/zBaNNbx55CFd6CB1qewT2SQkH
oDNoq3zpJpftWlAXw65VoQygTD9vThaQ9ss3x5RXj3hzyfo/auEJlVbUFuTkGgJiCaBchqBjqbuK
Am8I36BglyPw7dpuN6WjOC8QZ0ehtedFZc2tpVoj6VQs0eSHrv4mA41j0uGKf23KnTQ8eWwJ6RvR
opUJIXIq/w4vlGCE/il0bavdof22iGprHXw0ubcsfga3emQ1jA19etjPjtH7blrXJPt3DsgRT+Bv
jv3fKIjlfJYpjJu3YJZWImQlW2oNL76x/Xbd2TDKnaKL5nORn7/GaewJcWjyg+jPbrp908psI5WN
VEEV6U0I8g636NbxazblbLnceKHOZ+HRyHfI2/aLqMUD1GV2
`protect end_protected

