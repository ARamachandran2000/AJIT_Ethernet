

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AbrLtZEWaMZ9QRIEqn+KbGJaY9tnAHwhbFbsPC7WH49ehpa1EbqXv+qkeNRGupFwZ63XKanLVUyO
My0fDcdlyQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jBjvZpZ5ZMxrEO8+CEfz6CEl8aMhkYM5vXXCdl+QFohneB/4ao6UdzksCSxNPxkQX54YmGSOciXP
wgiPEkvihckzTQ7V+IwmdcU3758CZsJi1jYV4WKld6YxfbWBrziJy4pEooel9pwm0aG1jMx1yNUM
erFXjNZfwKELIgXdp9g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bNlKYiiGIQP+R/ChMF9YxWObkJMdPWBzZKUDypAuNCvFSKj2ODeFkzLXYHokfw+rz7RZe5YojYmq
4UkICxShbV1k/N1YYli9QKFi7npsW0xHaRa8L0tSoNNqAKETg1msjVmjBV5kKgQ78l19v/4te7qL
zUqdthBriU3NcZYre5k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0gJe90X6qrVRqoGU7iK/i5s05zq/0GlJ22Kt2H/04aXbES5oZ4I0aGRfiLSYUCL8istn1JleJ/n3
1/LRSIHwjesRoSy/6j9iedPDLLSSnKq+N+ZcvCJl8gg/L6B9ChU+h5YNE7HqJVfqJzqKWKPqsHB4
WVtjQ/Uh+QwxJp4Q/GXnPw1qlnDs2s6lJ8EK8000R7Any16QZ06T5S1IW5s5v9bKhWJj2Oj7lmWo
6QSr9mTUFxCIV/m+pXzsIOsSgFWqsBmD8jksQw5AorgxI1HaqEa3+sl/imtv2p//6lwEVtz8coiR
PUlfIUpZ3ecBYh1Zuc/GrakwiRgEs/Yjfe+jCA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ux0aTH3zrSOSGrjxNBhNJ8nXWhxNzkLj/DcKiIgChJ1nxm8i4YMzp0L+VdbHtn6L3ZPNF7NTEh1P
v7Gcx16JuF2FM4sw/t6m+FCjX3oHl0zUFDs/HfDB1IEXz+2hsgoR9SYF+bXbSth9Ql5SVw6WlbpS
yFwlhS2eW7RGdfH7yFg8yRwWXcYySMv+L+udV6VzSwe0SODgbmC4o26VRMdm0RBQjLnYxl3eT+4N
Qf9DbWnbFLLU2LtQWORMV3hNidJEmt4J99c08slF3izsh110Cv87/wiU6Xuvi2AB6jI3wVkno8/h
1xSxQBnRHm/fJHMh/8PrydoVk8qMhMXs9UM3dA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A3eq7CQ1ZEC2Oz4Co0wE9eavdVVL5N2w7vnxu/t08WjNVvgkDcorbVB3GWcUKigHFQo0FHxElw0D
PA15/K+npi+dagAdVUmv5cfV+KYrdhCLG+Kvl0Tcm6fhXM4RH49frRlov9a41BctZWlMEXzlO2Ei
69nxF8+cDN/RPLjSUoKp8oVTX2g6+udi83fdCBYaBZQYCaaDSNeGqephcoL2zlXyK7vU9KpsDUWJ
oZshHV12Yw5hL+4YuSmKv1aODQadN1UJ8qyFc0vRYTAqwP+hcDUwxiR48olGBo7U7czJnFk4AkkD
qULDB9rPKRIK3YJacz6Pp3GAHUDGm2JO78Eg8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
M27Xi4lqkzSMc7BZm34BkV60nL3CCXteVHLJ6dj3pqCHdoOnG8Ws0V+HkZpUxWY37pFLlSh28c3q
f8ww1qMG0QWq7Gu3bpcHEU3nbHqgjJGKREKiOt/7RrDuKebCY0nMkK8HorpWsiAWHhXN4dqLwTCQ
7fdi+H2j91MtL/xjCaU4Z1ZoAExLdSZlRIRZWUcYyyS5bcpBZzQlbl9tggWgK84lMphDQwmzruS+
uL0RddjWQxNMcBbP2XGQRBWWxk0X52WyG4RHdRA4xw7NNoWdkeRh6chZXSc9+TyWpGCumtJpHVby
VFUsH2Dj1jzCn/mlcjvW6nUVymn1vYQtvmA7Pn6A+nZRn7eTstCb1mX0Hlh3X2Kg3MM0VJL4C1NB
fhbEj7E6eFEm6YJdSdDuxojl8Z7aPR+uWaNI8YQrwhZcNlo9PnK0153StiflBR5O2mQmBJwvhYyF
2RrQIupgofOu921h1qksVpc8Jfo7aeN7kTAP3h3jNsnS+++cE9h/Fo+B52koET/dzkHzoruxnJqW
eriCzhI2ePK0avXIX4SM+A1pW12GTpIyRjxjkrn2w3eX6z/WUWSitdzThBpsTpv8H2X7y5wqPdxb
/ExOOmTcGdsJ3paCTHe/9pnFCY2GUjnzid+YGpALA0iIJca/GU4NsaTWBVtCRvg1GyY2K8AQGO4L
G9m70rYnRwvHDhcTU18G6VEKe1GwIJKGdmmMMHmg5uRGy+kAm7zUHnx0e+hjtpSLpcaMoPaRRdWM
OSzcUPVhR8iaTvTyHbiug+P0hoKN0UtIM33WlAjBG2ZJ3QpA8zBcRwLsPRcwvD6YZj882+hryrW2
GmBJqivIQeKCKe/wUD9PSYL5lxmAIHPr/rQIFQ/uCKfHicyFeVgV9bU6WR9y0cOBxAJVqEkGH7Fv
awj33KhwurW4kwwtxOK8fPXuk6FYxblIRlwCw5Zl8JBYdI9tj4w7VRCIeWHhxDUU5QlFcI1XM5JZ
ccqqRtbpWhtv6STcO4Z67fOQFk4cJcG4s+/BBg6vp+2ZcrPW/fOzpEmmHE+AmIyWw4VV5MdRBLmi
xrIVyNLgG0rOROQnOxWrW9X5/1n0tTaZYrn9m9XfY3ngkfUrM+oD2Wi9YaQMda1SUbjkkV/mgxGT
wd3GnEueMsNu4uDgqKrwXEJFzgjUyaAn1X6BXWHSc6KzC+Rjca+7wsYRYWy7OqhhF/GYj70LwibL
yjvOjfMGLIRGb1eBCWLaEpzFN6iTDwqKJ6+eKIitETX0W9V8B+lCPQk7GZPKo6/K4Ia//h5yjWDb
VlFXUKptYrKQrDmB3o+tqF5NGz844uxm60zWavpvM7N6baPQW2PjjJ6k2MzZr8Af03/dCwksouTz
afU7e7rR2jBmd6IvSmEvPCRPbrEXJqSRyjDbb/ONiWwXMV2NZ6pkcqU2n0QJntxExyOINBpMzWEx
aOMQEkgIom0d5RVJCMC1p3adX0xw3yUCLMPVvH/tEWcgITRiDihy7+YemdZ9+tgYx2Sjgc0wf53T
SWWYRq44kTVxsEZ2cjnsCTl/Z6RIw9p3antQw13tQeZyv+Y9kizevAa7idNWXpufVPq+BXP55PnO
hbFZP+T6WjjygyxvB1M9hDuRq+8vlxgxXCOjBc/4Qhl7XTXWwat7D8DCCGcfCDHkwJTDeWutVnaE
bVoRi20TB1p9cz8XjNZumXenVWu3wCQszeZZ8GhqwCkDGaOzUjmHpVkfWkHqU4gBkD+V4qH3e91k
Z+nE1zP9w+aMQdLqqyoR3O7zdENn7vtms5ECgBFp7OnXsOJg4lf59fUaQbrRcBIv7vDiP0RZ9TET
vFMDE6ur0DsrVmZv8UySIdDyEMOiU9AdB8rs03oQac9eY3onqtt0K7yb3EMXexNmsWao29AQsdWq
Z7VNVXCEhMFiDbSGeZ2jDvOtCHqp97FiFHqN0d7bicxnj6I+n8dWRNSxKf/sBY4OJPy/Rj7YbMNS
UybGvjj3TvM/7OwwQUDw/z7zOyVV5CLhjNcJgNJ/n6tDxOHwpzKVT7uUpuV8kt28FzYtXaLIDD2j
WK6O2pNQpgEDF+OK26IYLpMmn2lxZUA2uXvtYx99ZdzMibCZxUQ+FgndcPTbi0+ppGApZB6kxxZW
RWfxMneBjpH/2xHKxUd1a4zA7YUu5OSL6638ME+r3I12SQyI1Rycg3VDH7dCdhJ6iDs9fhJuKinx
Iy+zUW7WxSU+/xyWwW/w+KvoWtK7c5SrTwUJbRcSwXgcCZIbRaRRSflFgqeT7IKQiHYx66ZU15cz
Uwhwj533AkLGLgBpsnA4q2btCtcXb4biy/48yDE3x3QDGqiP9ZBhr8WyDhBSVsAzfjXuOb/eAnzW
RpsOveCLFikGyBoIdfSClSZaEBG37v0zdnNY6iacon5cPN+rqPBriScqfFExysT1XTfjJSqQ+dtN
iiprCSeeuVROYGwSBPAn0745MdwC/HBJXChkPUfHK176oWWpRx1jy1rymE0JIIGN8CGWctnMvGoh
3EDTQqQ5YVBpwUq81RNIrldqH43/PXJYo5W/BG9mUe70aVafcP4Run5wv5qVJRpNukD1wDd3FVIW
+m45r1d4d3+v0qGNO/BF9OByg3IsDgXhosP6HKd22K5jg9UDwn44YBgH6npXsbEfxfhtX11NhWBS
xA5WbcR0MRHL+973kdJYol+wqZYs5iwbWtXyWndP2G3v2GXdi+14/hNNJqkU9SIKFe1IzH20HA36
agvhWayIBAFY0NudD/2Nf3kLbxf+5k50jyWuaxzttx1pVc5Jt1rV9IClYDW12Irl/TK9OcOzC81y
HK7c0TMCmRUYvAIZuoiF1ohQNDsA6TR1OahYj4IILUklU4A8zOJ4+7frvsU+SbeQv9oagn50BxfX
2p6L+PCUoi80doUOG1HQl8sGH6oxA0emODZrvMys0hYagtyxQKsqPzFSPMMR8v2OKK30euzuIPey
LBzssItywkisTbnZ/3DWe+jd6TpQ3+KCQta3wVEiutuv0LoG2mlMNKHiPRNpayzIibiR+69ReBzO
cNGtykf5Dofc1tvTjSKi7YW7DofmRpzuRDBCM9ccoVOeD5nJjhSGo9zixXmGXObI7eTMbzDSNSew
fY+kdFo80BEkmn6O7KuUVIBYLw7lD/PGB7gY608I8i68JDY3Rr69y60AvwUTIn8ltTwLffFQPHTJ
2l0bkSe24SJCXGeYimKR0mh2xrbKfp4g7drdiejCIYyQ3A+2/UiBtjMfpTvgOVI2rbyc0On/08DL
U7zhD31mZXlCb5AlhGpIPLQsIXNUTXQpSCvs9XHkjZ3VIGdlM7P5Bt/Ck/ITjGcpDi6Nt9PnuSeu
FiMIDM9NTL1gUFMX8cUwauuzrwTE1sJMNM7ukVbN1PRhE3BRVoGawIdV3CgDbCmhDDPp8l2kBGoV
lJCp2xHxybvoVSxyroJ77kYAYwb8y2CLr5OaKABOCIprbO1Iw4EP8FD4Oy7FhaPnLOn2SBWUiiKU
Qtkt7WxkRyW3HgHctapFqDmW2Eb+0i1ajmcbFP9sUyPGV6oaj3kght5mp+QHLjDCx9V363sDUoWO
1kYr99yAlncezkIVb85E8R14i9baSVEmFkIY+MX6weaL5wwVE5rk71cnYGRPG6Cvdc5YhK6X7f0F
S/rPpJblzARswjmF6UrtbRKZafLyA7U7FtmFFzaBDBJiYzpDiOGerI5jr/8DPaxln/s7/crQYeJy
u9+dsJbXYX+9DYpTwBEKF2IV83NoE3RdsGsgmMzg81N9W9O6pXoGWe08L5QCqvse9+nqHGG5cTbU
t72Afby4TRUxTtqS9SbGdGGG7I1Nii34lJtdrZq1QUsNZyoTwDWuxz1QN+l4nzgcA/RPJr+oi3uP
PSdkuCl7vsvL0ZGPpR6aaN9SBC9aOHFqtZb8GuwHc4R5oV7DyERF2Qk+5gYbGLrlyc+fViht81bh
vvlhMrmgnxIn8Y3U+OnxaxtDfOLPkNEqlPhfDt3E8CkQX7WVHWI3Tr/8vWERU9OXHD9o4Bl4GfR/
hryukz2TzausqVrDyS/3bLlhsODbjDyioxONkgD1iG3qaOIy1QTIONpM+QXqjambqMzCxeKInbhj
SKI0WaNlZDqXq4QnwxVvB7sOQ1gNqng0ZBxO46qG2pXX5H+oNWu49XMnq9XrCiPzCmhpGOcjrdj2
WZOhVEv0JGwu0SY+ecxkWcFWv6b5zDXcTsE6vOmwyCZ+bSxA20URYdTbvSgu9alb2tMn+2kpJouu
Ur1zoN0m4+NfKIeoAog7YZXgQyMD1gxJePjkyOtwEMWJjVFFfS6I7MGS2UO//xjFcX/oJDnNY/+o
LXUeI/vvcefBPcuw7dbPh3URr14f7PWQxKWDFlu6Pbjh2x6l1TljUfX4+j0elx/Orb6xrilTImZs
vsCC1FvOjjgm3KvZK8Il2qSePCegBdzDNRZdW061L5LSVlmCu7Ee289PLn00WcwsmYbiTlA/h1pb
lSkbq4QFiS69m2RN4ggQaUd8xRZ1KwJn3P84Cwsh/dLXGM9ExBvQls0M1RHqmibW9DQ20lHyCVKM
kqik6qvPOQTLjPTRdt5h+O+nbC9TOsPW6rSC2XkYXTrk/CgTZrf0gtjaxfNKaeHWsAJT/c36EO6J
C3VYEtyIKBnUXSxGFLYJ61FfxjoPxiHSBRCa+MZca1EpCqgaoiIsaw6xTfG8xDmKnSUVqo8+fZo8
oLe9E2X5dHY962aB2+q31rPWf9ZTi+cc8JSN25mqHwDvJPiG7shgTuo5oxgIFeOX/ZeAI3ad9EIN
LzET9xIxDmP6iscE564RZ3UFmF3WvzBGxurlfBuM5CRdvhJPTNJx89OvqIeT+8svfLUUW1TbE+av
9p2Bk62/t5yaSsDDfk3NlMr7pfaIXwSa5QGJYDNT/AogpO3fZlSd2zT31/quKAgJh2GOseRupd2W
DVtSobB48Ww1s7hF7AZUFoaatn6+gK7Mkd8/PJx7pWYcbKV2Y39xyRSzmE3WGcy7WKDt9hj8qK8p
7pxkIoiqASgPyEFUh9mtuAZLnmu9HBh4QvgURuUQh3E8+cdvNxt1uh0U7l5GxWtyVGzjtONyw8hF
4bvG8irzTrz2BLTEJfnXe4hTkoKBgK1wVUET0fVRZzLTvxwQagvHyjFuEyNvvlKXZPSeSO9NNRVC
SiOixd7a4gP/LyaVGgD7n4FZSYTy7+MMuBLVhJyDNPTY0DDa4ee9/2gZHWbSrP0v3FCY65wy6BLE
B/bgY7nT9dEGEU0+7vcrwb/675NqHDUzZ+H8CBPAaABSZcqCMrbBkcrE9l4V34TkrKpBT3TisJzE
9qjM4Q8TX45a7DRyj+mTxbjZkjjl++ReX7Wpj5L+UzDwzDViSsC+wZrtbHSAqRZbDfqNl+9UqGFv
QFgsEHcwFDflpdW3+OK1WwDTuuQzw9K2SOtBkazL2APwubnQZ89DJYrkZtkz1Qp0B0KVcyrY7lZz
C1IdA1YyuINsT6iG5F/CkNyiZynRmzd1QBG0p2xcTK96QO5vM6vb4VoEEMJd/2GPrJwYe/hEnK9b
1LSAEnS0lDc7hjodnwCmOFSSw/Tt01JoA8vYxIbTgO8LaTg770vArTIe5slZWBScA+S5d5z9emR2
5IlPxBkxTlcQu8J6Kg2Glj76/81GHKYqUuxizbqpbG5ViANDMD2zYRe7d5zFsCZ1wzcQ43Z6Sw/5
p7pXzgb1UmRCZhfM9ReuH49SwW8+JTT2lJ122vnJ89GNMSu5E6yAA2Rv0TtBCeIDkVemgZPOqqk/
8JA/hVl+GR9HGSLv3x78MkUld7dI9GuxHDInq/4zDGCQXgHj5FEfTzOqLIY6KwyXsFw6FHnWXDB9
YPfkb+RnOwrtqa/gGQaJzPplIxacziRHhVKoNy86BYev+uGUsiDmnvp0bS7E/B8bjD87SnXTz/EG
08mH0pcfrGilNELrWP4Nvrnj44twW5pQ+GGLhH4XFhQU558MTp5m9Y/lgtNfbBWGiYO9xBj/yt0A
jHgArk3rz/2WR8vp+nMPri5HxT9wSA2OmNRYDU40UKdj2PNl0U4tKANKcIKzin/pEPQn0CjadLA2
UvpM98CtRWkpVXIeSBzyoPefFMDXorkoVHeOlpkLbep9Up7YP9pimmMUCD4HG1k1yPdQpTmtPXwj
cSLbQFIU7B2r3G2TFd3SzL6JZ4v1KZ8O/yta3JFZ+6fvBFSXwJWcO0os3Sk0Zicg9rFsFrrW0+dF
kDIeq0Fmo2mPAvs3rHgoNrczFj3UCpLc9bzgsOutVAAyK1Z3zCIaksUAqcmxvIor9lNodTEUEY6H
dI4opAorb3hlwQMNF+UeKYfJ4Pzr6w20JMDrYkqcvNeyoIIcwswwoHsYmGhA/eunrRQvEv3fuw2v
ik4c1wDDYrojj7hTpMpJV5UgH8WVQXXVx6E7tAFmfSrJ7S4ZNDvf8tF3muCl1KQsgjKBEJthoHDJ
2oc1UWiD7O1Nbi0SUiCMlVYoqb5P3cDxm2ngL/PS3/T7RpTE/UO5oDbmIS0u989/YgX+iVn4n6xT
hmIdElFa2dCDn9RGHAL19504gWzZ1nGy7cR4w4DQrK890d+KL9aVE6DXjkrkR1BuhVzhBoemVkHs
RfBuGGO8n/EK5Zv3FQjOjSPI4RR1QZ+JJ2KjwYWyqcu3aXS8IquCkCxB1KktfFbDXnOYb4YeCJzm
yoORySmNsU+VCM7d0rJJN6FBl4CgfrLtNaesJanUcebiUXWn4JejBIvvN8kxNhOO3fjKKJSJT4IU
GP6FENOLA11yxWEhzJ/nbyj8GqfLvWuHHvLPYg0I1+8RHVqZAmb/y2SLUPoatR+lgSNbNeh5a628
wNGJU9ooYbCDQ/VkbGvbGJlylNdQUk8dcmu9WFhDL+zn8axrTTCHV19RTq/KcbPFebzOaJbJ+atk
bnYWx46ScEcbnwqn5FUE3gBTfEKQKLPf/9HgY9HC5vcjJhNNi5YhqB5Ux/hijAaJk3WauMx/fbvJ
7pi9M5gKh90yU+hsl1KzWX5hYcEyOjPxcpsqnjJMRMBxZ5w7Zlyj/xolUz6nlOJhGRr+vhM/JYB7
uMok04+JpIWQlvJJzfhYfvBSdWv3SttYzgymOQE+RTxFh2/H+v2tUpnw2oeIf7dYpDgvjjAF4Eua
8vflSKQDxaJMTQpGfRd/e+JdKx4EWSz0637Z+cvfgyvF1hrg6pfqitrLNAvaJ722S3SbdKvlU7DV
lcNBgQLkvfVYkEGjKLY/+QWtELslxkgqOa7DWsCdhkOQdT+/AMiz4uQwP4lyYjzdVSQOBvJBy2bR
BGJygS8qrVXHZXQ7NRCvN8IVN3GincP5aaMtkIb/nnCtYN3QwaDvwALp3ER8+U7Pghp/zX/doCu+
1Sdtv8Cc78IzLF1uhziXfmTElx4+gW4OdBEPnYFmBhXsSWal6lPoMkue3b7QI2nu3VI6ocVSe80X
il5Y/uTQZ7s+/l9sBuuxlP+f4NWYmeS5IPj8E5odv0XTp3Ublj+GGGMHsqhgHWWexxD4bM0+uK8N
ip1XfGGFQtoYtz+yxs981UwcWUeNH4ptE/nQADKWjHs/JhVJ9Xx7DmGuz61uyhr6eUYEXL1ZMDa2
Ej2s+vYt+0vOepGrP89KtPBtqBRbcrbWeHE/S5ZX58TV4wmF8O8lb+UW46+7bRN7UwHtUGihkrDa
OZecW3zIfIiGPmwnSKTTAMlX9OdkBZRWBbBtKfFHSDmggXSeuIUgJTNXBwX866EvDBTdQNBqWkjV
bdTG2el5rx8op1UlU9v8GWqVJG1tHjrQPrDunS0Ccbw3IUznXSl5RqNSGhjcTS4z4+LYZYO3qdZ9
+VyJVGAWTOOhkCFeMbHJkMuhWLtpM7mp2urCDRgQ76MFO5nEbnAfyHgQ/G1Rl/s1SoE8gSho6H8G
SP/NVfci8E+jX/mnsl6sbN4JmuYg4hEMNBgrio2kawCe8oeQCtC+fdfvqjdMg2/RCdu7Iv0xYtrr
4bcTX7QK8DqzM9seH4N+bOTH0ZzR63vca9e+Y/uB/zDnEqUGa/B0KqTT+xcY8Xf4OfhqBw+Er+zO
Mwdw/j8ac83qNwhm4HbLLYWFXbgmGHZHk5u1xQjnM2LuVv6mA6MXmPlbY8oT0S81xuixLySiHpuT
kc0VOfJiv0ip7GQ/cY0pofn42IAYK5s7mnFmwz9lLFM7pbI18+vlcv+ZcaG2PKaJo642TVw+GNua
0h1M3ritBnlLj4DZIDpw30ZCWAvTt4SxCIuMqCzt7XfBmYP/ZbZEUW+b8gnoUKGfdKs83dFBT2+8
IqAIY9JNQx+1NW2j7PtWjOwnCadzWg52fSG+kb7MOMaGw6Pz/6dCLO8r6un6Q75b1rb8EHE+k3vc
niAqeqCkfVFp0TwZSuM+XpUOzEFSwsTDmYHth4P1eZyjMtcvxUBudpmQIF4SOVXufTqjnZPpRfVX
wlPkt8lUIxSUvS1gShhMDadkjNcvRWHZqMNFgcdODVqJ2Wo+zEB5KNvMyVZqyyqLvz575dRkiS6d
Ih/3HgJIvI3jgqQ8+cGfofPkQIa9OodNqIuhznlFidBRaBJspDbnGa+UEdTBJYbn1E4Cy7vnaL6U
zjigzWFAYNcm0AEWlvFRXu5EJ99cnX06cRbLWAtC0s+4EFUThqQpsm+sKuN5lc8omaCrAa8wNxr4
jR8X51IiMV0tLcK12pppsojY/KcjayiPxXh6o7br5OHEqPeZiqeXxNAvQUQ0+65L4weg7BUlcpUv
lfo6hsc/mNgmEZ0vZwGfr/5QZKpP0PYojXqfFDRk3DTQ7sBPZfGKEcdNBHV0qp94M14PR2/pKBdl
s3IVquWX5qjNOeiKJd7Wrf635cUY9p3qrRjrx+yhg9zdx1W9YrKnz5OHBRhmYg8xZtxbhtac8dAP
M/QFYipY5BiZNtPLapiHhd7TmqFYFj9Z0y+q6psarQnOhYg0ObqO4hLRDGRIuP2lqw3VmtJJq3Ry
FYn5+xi+FIlkIAhep1sqbvmWQV0HP6pvB+8tXv7YpHxGE5D7byUl4qCrNWfezkmBXOrRgWh1gO3z
aEuCRgXzXlTasgXA6LmXK1+/DEcWEUowBxW+DgAzPDXgrRhgWeJYZ79b77znezJ68q8mW2QR/ZRQ
grzJx+90/VK7svecQXYzoLGql15VjzrQrkeZGGF+eWnIFxg3mwgAv2ZfxT3bZgA1uoqQ+zsYFG74
UIl2BhkD1alC7rRXohNmmOavZfXfi4izPkySvAyWxUh18/PA2Jcj2C0tDSsMNcw68TBPUC28pvMh
e7Zm/w7thNQNSymXYdzJPq4pg7G9TdGCMuzEmMAfH/UHl1qbm717QnFeU3S9L/+ZiwW/vG2l608q
dgDW01PiLCRqfG1mwzVkuTMraKys2rKQ2zcLbEGApXgsBwdfUNHkRCweKVJMu02WuftglYrxqqQL
s38fnWUCLVzBQqLYo9OdmhdFHEAfUWy2k3tCm/SXyWNVIxR+uELgO2uEOwcJKcV+kWFb8LCD59Jj
1/2jH1vb2qcP102bhd12ZvHfERbRDqN2/4PfN7lMrCSzgBS2VqbHKnnYg0tQfwuQPSoK1RBGyqt+
QhTsyazQP/2LKKHg407JntXP65i/WBP7VtIpZp1R+oedCq0rJWg+R84z1Dzm6fWw8SkPRsiB4Rev
wmtxnO76aTJcDxP/SMLe+7FxbEBjL7oTXtzPBR4Od5Y7vo9cQ6tYj+374Q8+XdrrBrvIkFHfmIF1
V53DprMnuelvQkebc+t21VxgCXkF1mZHpZQLllTqKBA7OM/+PCmGyJeFZq9uuRBzg6VTAOg66KYs
hradi9Fg0xZDeY3j63n3Ouyw4CUV1HZwHhSSgLG2bCrZuy5cghqDRiGelTWY1bBonofs+oWX3ZWt
3UDzKeZsEQmhzfEGHWT+MvqwtXGjT6dZVmr2nTzt1Jclk9FafdIuuzwfUcf1jKtHzQ6siNO6tfeD
i6reB5dcM4kN1ahWZvX7d4rjfq249gE+6xuR6v2978YkLSjuZu5qJm67wWOqk0ae3zuT9HDmT7Kn
o79YQu41fMfIqVtw/XZH1M+5YczDHCHCIp8hwFPQzCZzLuHhkQjVtP0mGBA+VMe0TKCG7ow0YGwh
6254/eV8RtuGbvzJ4dZ+ySgbRv5DooqUYIEHGHgv9EjJHDYfy40QJekQPcxNCmIGZfzDmiAO1xvI
Let5CAcC8U4lj/RXLLYfSiR+AVfzM4Vbuz4owlwqGCHHpfYChAHJ5Ya0MQbjGGzLDsxhiihEDj2q
g1b7CFvCqTpEN+6vE0ILIzEvc0w4wQ4X4XS4Cz4fJPU5geHXEUqV0rNUhhw7Izzi6b4JIdy4TVFW
AI4fTDguFOgZLw3nwAQqYb/gX/hXbzTqw8Ss3RTX0hJBCgotEWZNRH7VGMhJFQngDN338sSA2Mm8
sPQr8+g5cwARNAw7LlGADQkYj5jlIqLpNgNk1Q8is7qGoAb1fFShfimUfjNOuBx+lnDRqInbd9B4
+lREurKBihqElN/xmw+dtFqKLgWtJPh8EcBQqRXCdiKOnvrX3DQxgXQ39T9QG2npK2yhFBU5aCYA
aF+UFCK2olhFnm6eSw00vpZDBE6SlJKt8/Df5uknU4p4jqQrK0n01H7cJb3+6/bgwI0GFWrrnRGn
XbHwBoXHF9k8truuMLk4m46Jzv6ylek/UVC5FGP0CvmbCHtr/SLcp0LX3/KUuNxA4EJLvhLy8til
SxXrnMVcBFhm+X7DmTdsmBg0pdE4fwwxoePVtuZdMzpCqtv1j2ci88I44jd8u7j6scirgYl5AFeZ
nd1amJ4/gHdW9dEXiqrNjO+xpeCmTMXaEHLa8gl12UjzNyun09ZtZWW1B3A1ZPUPm8TjAEezDkiA
v5ZsOt3PRfOPMUvha94dQKhzLQmlIhozYS0qSBbMq17/FwJoyWVuY0OW/0UQPMhqmCxWL+6AeJkv
Py4dM1eNZBUpNem5EK8RKFVgbz0fmm/G3OaK/Gk8wYNjbdIR2qToHQvoRZUisKpKZpaJuv8QrlZE
2RI0HKz6q2rN3J31dWB74vGBVD11rhAejcSH7rOfq1kd9pwroTIs1cJFv/CnUiDJAbHD7U0wh6sE
QMpO89yxpk0Q59eqRILQ8nq7yC+NzsKAWuykm0q+eparJD+0jFL/LhxJL4+aMDPLwvhtGVspkokx
gtGbxsXHEeEyGUGo0POoDimqoOXGcBK2KqOYjPu8VjTGH74xqLwj9mNpP7n+782nnkFQoVb89qf9
10IO5egLT8q3jVZzALFYqfI0vB8dIzr0LnWucLHepZaQneXK8jffFTnHVFNA0HJiE/yFfJbUkawR
TQq09lGF7mq2FdeTPoA0jJgko3vjlY7KorQifFxryP4yDonVRVKNKH6pf5CI3z5S95aQ2K979qyJ
TDGL4Hq8y4qRXkUhdRBeDsUeBPKEOxMfBKxFgHjRjQKMRw8sr6i9zM//4+9ogsQ5WOjmuCTN0umm
ozvOT0HWxAfY4ehRBbNgO1S+HcqotRuUs7m5eY1nRQ/CLtnJQbbj6wGrx/SSEEurdYnWWqxHCd+x
E5SA93lg5Rfm8MKmz5h8u5+xtUsH6hoBa82l23hekQPtTtU9fitoOMoDt6+NQsdLxt4ASvOGUZMV
XoscCReXzO4DdiRbEp9x0lxFAFcbJxQEsKrYT2GzAAQBJnIOrCQqU15paemx6etdhyEbuuP9RkKI
RXtbTStTkC+lbO9MIIdz25tAYh6wwFjZoSu4PnS8zl+pr0A077d0JFuyYAZRF/eEWDagC0G0RSpV
Altl8w7M2bertItJjhUXKQRA7+3s2W5V9nSr+FXRiZEGyAmPVm+CXCJSJMjcN7TO4cYscQnR4mWf
Suc/HVnsnZAZOV1H8+8Oq2VaKvFdd7VFandAXD/o/P/c6xDVAzfSJL7vnbLyRsUEPBiWMhrVRDMZ
PY6dak9doTXaA5/4TS8wDEahubwbczC0M3bFNYxLed31S55TMEBjc4Vvuqv18frdUcRB8ge0H0Iz
ftBIHuATm6w6k/2clNrXTlTNg/4hHWbvSh6GuqKReuPd78JYjFfHxNdVtlClkiKbK6bwhKDDg+kx
/K4EF6mIvTdvotrpd8GF85wbOeE4b/h6V7s6cc9uzwjI+UX0mhtcNELiECpppO77eOqoaqznTMXz
tDXPylzNcu/1Vuygsv2IXeYcyvvJP/hS3ob62yTrpksGNKGcLeErK7eXZrrirC3h9R4/W7EciKAR
wiPXGA1K00/Tyd5xi1Yuri4l1NjTRnCr3RL++Oyb/FTYr2uMGhKO52j2/znQHP8PGN0zQ2O8piJr
PPfkdopND/KMfvJejFOdJw6pzexecoKRrdeiUpC3rXm8leTlpRUj+mGd6N4Q60yQcBlYw1P22wx4
6XeAdkZ1SqFaBaMiqtX5o0O35ZGHzU1INXUM9ihHNFywte4nGCLSDtv3znkuIp3uDNrs+OZ2VCxg
gui9lDZx0XW+/mXY1hYg1HyzEdyRpZ68Wy2Hi1VeEr0pF44ZZT7LgsaUa11dFsHG7OGg0Ej+0sLt
KJiA4vGNu017j7Thf/SDGcUBu/NryyxyRBuWNdy9+/6uuFaZUpyJS7B2Z/USJN7wyI2wgQtVtTZA
yZztslklJJNNjisrVbduby5h07tyEKXndz49iBLdpow2UYs1yqDbFGz2l9V1kXEwIt2zVGdGN/yS
Zyl+MFDikOYHQ1V1qkcv+NbBsD+Y5Ut7yx2KwE0aY91l1PLBOD8r44xMRKs3fXyFr7dftgs5mhMj
/zE4fQppmP4GjVHaceknovQABqsZx9ddlZstMrIt7MZpn1EjEht98YPUTgj3o8IdSLAWT8NILaXz
RPuB10wRJthi/FcPvHBnj+xXuFMbEXSXIbcRw3jNwDKPIFuly/3nkvpEbSScJ/OGlL0TkxPbFOEA
w09cRzvIeJD9RSX9I9T/A83KUj+iUGsD7jGPYRFvUPQ9+DRMzLJFVmJ6dBgL1yta7+mG5sIkcQJ8
xT7XqkiM122gHeoJCSnWHX1FeNFoQAQEMwKWQkixgizEeFyG90+lgBhs40HvWB+w/6L2TcnaTTBE
6bSWoIWCYhjEPCyXV3zXMXXurTkeHhqwYaWf5vnL1p/iL6SzD6Sgl1T6I04a52S801ObfaJPEmGY
+yfXtR+G+oZ0ETM+33wZ9oRHyrawqgOYRbFa6R2+pUg8t6V+HpcLHc5V8epUHA20iOP5H9gA2L1I
W8rdiLI1vJWIndXvXXgmDRkn+FD3+ItPe1Cr6LP5/nnr+NFI0kbD4Jg0d+CnioCSPvEIeoYYUQGc
imJ0xUNSyBLE5G2GAOm5nt50g7KvRBr9ZCs0KHHyup4rmrgaoDqYLXXCfSOlevP9riP91jxAor6Q
PT7zq1GQKveITekNrjkBU8IOp0+CEjWGnT4pjzWqIRa0u7Q1gl63VIkRYBG9QpNluz8Yhio7ufm1
CUazbUI2iJW3chHrFhjezfkXqNzp7YFI55kbBan3jh938mPVm549vad7uNme3a+phxS0+wEEMvYH
BOKmN0qeml9Eo3JLlqM/XRin7PPHreYA+Lp/gM79dGMJsPkogdUNJiElQ8+6aVl6Ne0rKAutESVi
Eu2kvljT1X36QKw1bWgtSbTP/VDzOc38rwJF+mGPrZrqudcgXqJAPBd7YTlYt95CzukE5kpT9DuL
SYrzTB9ICNbvgvWL4RCNhoePrm6Smfn9P2Dh7aMCh1KCkhNRoz4ocOcQX1hPYpkyW6VhJi4IxAe8
7qqNNFhJ/1A7+COCepnxL3PEfOkMWLnEfzzdXWjcENixgmTUajftrLrrr5rXtzzmIdU9G2IovJdD
EsT6K4U4vQiFG3VslwnFqMmufviUG6qX8K0/WpjC0zouUzP2a1Kf5Agmp+RrBbRNeeYB07qhxV65
i9XeGL0rRG9ktdOWZCQ4EOzst5/jBNPyT/QMe4nWzR87fwbEOawq1uSdRbaxxxeYadJ4WG44skWE
dQu4SUJGJpjVaE1hL8gbByN3tSRT57PEeSfL9izY7mgwSsz0i68ue2DRd2meeYRHEID6tz0LmFos
ggiNGHgEEXp71Rm36KBrf/ffrZ0eNOw+xIaMAHR49kUDmtKF/sZTvg3eSwM1W5NZK30rGgSSCSGt
GfkGBTnVUUa3jkY+GxX09DtXJfDfBLl0iMbwKwjh8Y6mZGlBx4VeJaPYJZOnA1UcuEkdExDo2L15
l2j5yFehYArF6JR8pse7Kry6F2swvWpK7uk5uuDA5MURL8m7tUJ51NppesrSuzG1hvZzy21TnTuk
NmgU99or617hS+fGivPBeoNDEimb88iUcfC9D65megdh8ZuhCJW2mNAx3AtnrFn9xp/Aa5S79JGK
WRSYxOic6KE1x00OzStwG68WCE2Rp8ONPOsOrudZxcALorYaZ9Rxc5DtUvtvT0KZhxCvpsUhvsJJ
SRmxao7sK3j9wxu95sfGLtegT2cjBPUNhcSqW/5hh64A8cr3FsjhdfBSqKaBHcPURbOhZz+Y2/cB
qn8jCNnNac0ExyBRrN6C97YQoVxGbEjFAJH4P9c/AS/kSEVnuj5yJarB6pb0OyQa2vWgJbvPjDjF
LFsqecLIBTRRfbNWZ/usUA7gZfKOK0N7YHtkgjCVpuGDI4rASTW+LKmdQIQtfgu8xMajVNsSKsoE
T5ICQi7N3PO7DA+M1xkBFkoW+de8NARxpVD32TqKNhZ/SY2qtowNgmuYHt4IOM6Wx7UuFbs1oRGS
iYVJxSXgotkf/AOt0n7sRl3NUCSrmrfMrvnFmttrCtOaeXUiZh7mUEA1fqlOh/Ntc7ZJBfR7NgNA
nmDdpL597tn7gc5FRsXOgZDw9/hPrCUJXpuSnGvTMwFCvnHvCsPUHtfut5deKTW0ICqQADtLble0
Y+hN7+XD3f4hLMPRxCk9vD5Enc1KiLV/An5/YlpoUu1ToiJRucnIevClH+HtFbvo9V+cKGFfMUXZ
YcgBPdqPzTMQFzcVZFJ5Q5FwOxKurSbANEiLK7VNIKtFspxTMWocJ3m5sIq2Ep1v3Rfbhtsea46q
NS/XJZEwawZzFyDLVsA6HNeajrG0tZ23bjTdIa1VaAYDGKBzTNY+HSQq08grf+hXMV0exr1pXv8B
v+iPQDfMTfEWRcTBpDcsDH9nhQTQbB3Txmt1j/dYIxhsmxslVGtz3oR9ySfXnFEmcsPXF1BEdgFb
8PFAXsz+/6bYoIdOx2qAhXA1TuJd787y4b0LCWQsQFYsODsPA1TDvHNtqxwHU5VM6xD74KmPA2Do
UskeXmfqnN/Pc70in2l+HAeF1X+KbK0tCPMpiFmIfQQd2G+CLXx2TWgcTkhfYPuiQOvhskRIA6Yj
u13UOuzTgECmeC2Xcid2adzor8RNaa/9fyfANAiY2Rk2SyZy5xgfP4CkI5B5xPafU7LQKCOMRCM/
vFSWiGF8lAEFIZU5P0Jvx8tbb1HMOGQYNjYclqoVVc4LSH8WDV3fQZeapV8Yr1D12sd5L3Uy2cuh
WHxPBo0YC+KD8Ej9UX9H0/OvwTHxBhRvr1k+Bk/zHn1FBPvUlcHqpDwfZdq9cznSViOlKEs/6pO2
2FKp7gANPozAe76jdOQ5y8R98Xqb3lMRWU9OP2EPEPVkOjZ3hx9BkenDws1KMCJFKzYZdW1+XQYT
A8oSp99cR/2o7ihZ7OjL4akcRsgX5yJnzEPVdPbRQZ1wYKFh3OWljkb5VvgyomhmN+L6880vagoJ
auQ4RbHQwH3pHFCK84h8Exs2CJh6IbyEKKAbDPpC2dBUYuttQMg2ttF+uTccM1BV1QuigikkRHRt
WuG4RQVHIVEgO3vQgmK8lr5ZrYf6bR5XBeACFWA3ugZsQLT7cc5U3qGE27AgJ/rxzDbU9GMTzI5E
Az4r1W3nkhOgn0G0WiDc5OXvcyX+OJOXcN+mDzaEA2Vh4WOGFRacj76uiEYPlKrLh9Y94BpOudtD
biyrJNGzip2dW9Bs56FT0HdiP5MdGdBLYTgUY8ja6fHvkOYcsWDSpW0XuHJfpoikelz25nmjY59X
DQtKQiGdU4xIrk32CqOcniHf1ICmHHpLKmrhXWYbtCbBEQLOd0VuqwwfHNWA9ps57ez2QCHXGAlC
j/Lnk9q+Zsl+exnMRcqfiXteqXn2G6GXIOLuZEhqjBNzk3ylLgUldPScmRE6QTsnC4WLumd1Zm0Q
GnDuGHvy2u8OOlxH0hLMsEjLiY4pwyEW2xum4BbN+VkIS5+n/P3LALBHVunB4fdPMBOPBqAaB/eq
Ze0CwPatIq4GAJRDHqvtmJo5Yjm3rsUrw3RY8yOajKcz8OfxXHvAB4Nc6E8ttxAIHq9FI50sDjFI
hkNZfzydPWPTS3NiKFR47O/bt4ivE5boP+nl0OU3gt3+97ZL5H5xLbgojDwdayIrUvqeEkJDZ4vG
Gfs/QffaWR9tyMzqBqXMDOCNcK8NO6NcozNUi7M5Geiju+NuYiS6B3q7S5LQEjaFWWbRkcI3FrDo
BTs2T8R0X4Kl8FgpwfCGXvw7UEEorZAzGvmBjk4wRm0FWhcKtZ/eB7iEFaXNw9PL+9ebc6BjHHm8
fAlxsjk5dQojh6YSH1xoBEkFAYRpeya0wiOI7yigyGT6TV+ZFvljwtRj3zJR3BMSpNXdenNG2gF/
ZEHhx7HyKA0ypNxHoUGOhmmTupdALFy5uQqlb9bET0xz7M00lK5otfgiXzWtz3m7i+QScKh5HPjO
8boO3dTzdGcKrYA5GuFeX7iuD7QBJ2IweldHjvdxVtejzqZiRDgBgcjVCTbYCo3A7xMasMNONTum
Iqo/AgkX6LzQtFP74xKoSSDlPlFNHxsQgh9goi/3ATi+fvlzfGpXdxq62FiwJ7H7SKMH3h0t3v+2
mBm2pXukI/k2AAJbVIbYvTq+wzKtOeCcrLoQX7kslRUD74rjvvy6+YHZ4h9DtG/Bji1O2w7H1iXr
juM/0BNsuz2I+azaBcz9RXWi8AdxZkITq5YFmbLAukgaKqWc5/+mM3/jhc/yNShm1bFu+ydgyJKq
7LZExwG43BzzZxd/OataFt/pkHx6yPykN9YPc8enRciSvb2LHX+9UZD32P0/CNZpybA6U019fG45
mpKELG9OznZXGkH452mGSRDWPOhoojXwGw5d+wzXsyLwSbZrY3iP+3WWu+WfXZvfXOd1YYDqDMB6
k+zC0kdKTDsaWZtzM6rXxCKp31yRQ5TYjkHLrsJ0KS1ZlXqBVHISEzElccYjnKjht4Ft7j2Oh5mt
i//ArbdU80VCF/HNCf/fkUKotW6rqzFnOdqnJppNPHY72QFeYjEod7XDgO2JvdnwxbKmIdeh03hn
Lot9dDOTsip2uWptcZDwhsBKA42XLBEOeDkB8kyim9RTpC9DJfhlgJr5JfYDPf1TaSLqr6k5Gqnu
XtlLWx8LfOE/ozefZ8qDVnDyWqwDt+qzPxnAraKr1rQTLOomiQr0kGeNhwGsH4WLYdKalZaV91Hc
FGT1TYbFDixsFJ6+DquLEot14Qt0+R2FzewoQl62CPPAvNq523jv0OBJxhs3UqsMrrScu3GU3yJE
MXO+xQn2z+pcRzB/ck+i0E6gSd60OgfdIc+IYnORy0E6HrhoQi2PoGZ7ctN6z7oJ1S1+29hQeMaN
pXuQVpgQwSK7TO9RGImonyVwm+fJ6V+dv99swkKmSJ6mGpSEt57s8NFXsWW3sVPOQam7LPsfoAeU
8UUNjae77GZG4BixR4Dlg5Lg8lKWwovWXcp5ixwdx7nPz8rtDzCw6c8cH4WTPjlYavnJ0iK6pDj1
XC097IP9f+YFZLHAHRULp/6NUAaEduJawEaLK4fah5A02D8poFAC9/MD06F+4j7fYn8DmYM6BYcJ
IfyLhtOmwWwAWfCjxbyibBTaj6EE088CWpogjzHSoU0LoDheaGxWfCxa59glxTHgBD5ewGZ/6pNK
oB1gEBr1LZaKcxn/m6Urz6shlshaB0xj7/Fr8vR7ywd2BDB0wg7d0lOPviBFglUcXMohzjlkRq4f
xNhrvH78LvC6HjkBmJg5TGjwGMhtIsP0uP74S2vDqqAZwKAazsls/3ZG3D01ueObFQIMDuF/y9bg
qPbnIabZ0u1IIDQ9IkvsqTu//W3VHHcCzBrGI+DXZYSdh3LdvhQX+YQmm319fIEVk8oVVwTlutpv
wyL2uEvkxv4EH1AC29pClbf3UY3MIB4HLerJDj8yKsNHgeK00j9rfv0KCcdkQjAtSV7+JIpjBYJA
I25Gl4F0YJQJa+W2Kzh3N5e4sO7M+SLIXedQ8okKAz/aHPZ8ts/V0XszUWPxT7qAYX8byCPq1Ku9
3vfi2x4XCxV9ke38B3WkUYoQvAIK/c3NbVYyERYmQkRktSJqPdVq95cDyrsej7hV/VBuD0zQhfe4
AgMFqMqWnTrLJ3RKrmf9Frgx6yb5cn7XSU6eh3N3qPVTTSFxYgqZ2mNSz5PYKqr48kU4DKvOAfxZ
EuFdmHtNa/So6eRAa/QeN/6PbPpHcr8n0O8iH3IgaHJhk1JPyAP+l2Y7cgjUysuLwHwyyRpdJpCa
dEGrFKBmzYDJtvqJ7KWKea5D8xiqtfyCpLBfeWzUfPuVLS8koj54dRUvbsWjuK5kCsIYDbHtjbA3
HXJq4B/MUtz4BItTD7C/O0PFFILRM4j9WR58pEGOKYkZ48aBf6Ym8SfurSq1DMDwacW4+m8sHK1G
JStNX9WDoflNc1agLqVJDodElJxzTODseW+cO3TPDjPZNeQpOkYHD/dzni/vIk7wkPbfkR3cf49W
DbZz3/WaAxFKKBEEBocnMqYJPd35VaNxQbcrHQqbmZ048kRVNPcj13t5zvPW5v+tfaMYu7htEPhm
kXXE1cyGLQN7Sh5C6iMLB6TMiQW4ozQBJbT19hXvnEwtM7UBqhGwHVo4GOJX6uH55iCVM4Mp4K4r
1ptTb9oWmDyqZfrpuEGlxaHL1h0m8MovLCocIgmyLDZYeSlcbju6oKp9fj/vQnYoI6EWlKI7Ksbv
QbmNXOC2/vcn4TlsPRBw3BMTOqo7xtHKDCuRhfOTVHd7lP7Cf8ZcjLggyXevr4p5IHVVBqtnvPub
UKMqCf7yCBZXL5qUCVsCP/b0jqafIOb7Ur2rtg3ZzLTwyHnyMJprqxMoCVaniF0Kj9jPS/4smNEI
Nq6rHFcxNpkB1w5XECZgOGa/nZMfkHGUP7dRHPUt0Z1Bmkm4YfQpSxGWOm25fktrDkIH8vj4XSQp
1bS7zuZJL1p5RLQkEgedRyckSp1PrkS695p9CiqXQ8hUV1ug8NiJ5tijFg+T81Ccp9sIZ7kr8Qec
+z/PB0OdFUDy2KULrOBJG9LuV2kAu4UIj97bKOOXH0DeGPa5pcDHB//oLOYQsY+v4kmISk5ufQz+
ss+tzbMorXxJ7WXGxA14SChLVu1pHnV9qxbj2VY95DPhk6DiUy7EgSZD0EdWHisUjDC5+cHKWaL8
eAvkjdnoMpocPh5XrzEjJAmFTCVMYbAjPUcm4u2EOSO6xEZ8NY3UjTmDmF/ZQY2UCB9ju5UcYbn9
QsWSCSD3qdGp1RCaJ0y27dpuamBYzdCnPyO6+r1L4NSaeJgd//v/EUuEjlnhfrjdpAyGOJz9SvtM
YFufYoie93ChKpg6a0bmujqg43aDYu2hebwmcqgFqvTcFF1oux5IkCief06HX+DtV8jqc8/qihcj
m1Q6azetfxNKn444NUufAa//E9x083JfR1yafH+i5nZiadZNM9JP2sEaLIJ7ZrUynkIKQEnrDSXP
PSMhVoeN8qk4S1Fr7DLjaggT6YDS6BPZCy/DVipbQmg0LogqWA5FLtAjI9PBWDBXW7lIvNmSLEom
UmWWVOmBNCBpJarNHXLnMm6cUFY5em2uay8Kx9M9WM1qk5xzE/EXlIfK16f5OULgCqqHEAqmV/Pz
VD8n2J/KZMxyjSrLwS3Y4OhfSj/mjRZWcEK1GLhwTKOIeGttwnO4bQM1CB2E7mcQDKgvkWAub63y
hZOYhfTBdXQ8AfpTgIT4ep6+YOiw/BV9YASxF53vdj13Nc1NqBvoWl78dx0q424MXb8rJM/XDPje
OJitmy2WjJ/Gomfw8ARqUF/wfvbkWMYzw8+PyfdVi3+ZgEio/hfZSK8uGlpoQlZ6CWdyP+mmREB3
5j+tYCPGoxxIi/Vz/CFPme1uShWJ+JQGD+w7jPwgsUxKpiALqIvD0Ti9qlLWYa7VCd0d+bAha6pC
ZlW4FMT6CgO/RjCBdxHuyQVNZcNJ8HO6F2y7b99NyXhSn2Py31zjxGsqyrDEJbzep3YgftdkF5yY
Oy1qHPLr47ZtwTwtQgsz5keU29wSIpnRXnKl9MbYfAw43lW2oxlKqliQKReRieAAKGU7eqTsq2ld
xd2masgZxWVB9a8Kpj8DdrM8L9SJzVO/jgY5pCRSbVzLt8GbqdibfCAUwndxZKOdpvPFqYkz8zfX
mO1H5fWk1YNe0EH3zKz7uucstXEu4Ai7daU0Bx/gM2PPVlSDbJDW7d2t/KA1/VdTYP11x4FqeKl7
aqnkpytU9939JL89cMKYvohb+56jyZwJ2s6QmW+9tYD4dC8sWk6UnVTmTopDB/Isp3nNb+0xKg65
lDtUbwizunFM8A2+hMd1XunTU2g4B/C2ZXtO4l2XVv+YE6ikHOf+q5OD9snK3hVvGTX/B871QcVD
eTfvqogacIGh2HhTTzZ3hK2/UxQl4RRX3gDnYBZRVM8HR6HTwq+pnSeYTEyGUSmqRoMDyftI68PH
uBKj2XT1tRnZE4HfF23gC+o7j03zHXUirIT4y+avhIPZgsnKaO96QshG+DbG4YdTAdvJpMVx/0dJ
TyMnFTL6eWd37UAKcrLKVWLT2vxSbo2CDahQ3Kiy7+SKxM200cSvas4U28UTZaUr25I0eTP2Hlh2
MVbtDSd5iDHCMQXf00FZrCMgY6JS0ZJtUzs2iiybeRFBrhsGuUBB9gDw4rbG6iJxhtw0hNlYERd4
/AqCgpfYdfxfKUHiFo+pEMCh1KPkxrJY3joKtGYMBKSRs1krHwWAC96l2sRxY6Qh7R7O0xEXFshD
Am3DpnP1A4LONe6ysiwv6wI4lZajGGkZS0xzKBzPgoYrxJerpjEBc1Ar1erI7rHSOoBJOZ8hVQ7R
6kTi1utz/Ecyh5myvTSpsrJBKriXOq+MVDmx5C/F6kqV8n3EAFOGIYY4h8tElr4xAHq3/T/zzgQx
Ci8ZTvkw4woyeO/9+sQrDn0pXZQaZyh1ww4KB6eVHsNnh87wSR73y4RFMS7To3HFymoyi+uWV2gG
xauUTxQBO425kFZgy/AVOfGqTvfjLn+Ry1MfKZio+2AoGLgF3aDSeeQlLx26tCTVl2SEPrGS1pt/
zM9z2OpbapC05fly1dh0oVrBxDMAW66gL7ACtlorSzPFUUumdCBKhDqFX1dA8ffDumzNU85ar3oR
n9NsxCMIkg9CpBAeNSzZ6lWD0lXLEhORo/4oiGxPSvf/NUHzOG01H0CI6cTK9BMOX+tvxbIouMIG
A1YqGG7be0JfUCGHq/r6rtg2t0eFB4bzwIk+efxARwkX5Hqa4FcztDW7P5Um04ouPeLn6YaVqS4M
xU7zmI+tR+qhUTAzojSOSZy/fIZCd9zd+0s/0WpuTrU5TvDx4NihxHbSG1hdHj9rZMX3JKXc6PYg
cHtkvjtsaG5RCAGg9OfLL+qtR5VG41WSgkqWYSuSZeMbXlrsAz3UKboM4OCEXUPymct7ZDpcNQB1
FJztOHrr6vHfyA2Q/DRxByNT89ihS/TanfOynWzx1HCL9tkFiWhMPrlTVgkbRd/yeZ93BsHjT27I
Yl12rgGVMJG5YHe9PCtTqYqgCYsZwCYjeTDD0ITfdZvxX4dTrZZvzO8Wv7Px5ZSfnqBTiXtiODsJ
1KBj83Sji59/Mgukbanx+QwFHSi5EJEhLmq5hDDGWol/UgHUnM4bqEeFimiLqbzPFvlXkj1P3udc
rXE9Giw+KHbV0oQ4kLxHnL5htqF4Wa2aRVjMhs541D87ADpGnG1t1R+gRnRMzuzyQAmtGee25sJW
240qieKDCL5w0YuUwsrIGV0+8RMIKSjet0G7rCtk8YkXms44NqWrOUABeWenk01ZkcUMbOAEpQOp
bfLnAdmO6biKSluZuYxM1rhumFHxLduZHwQtOsrpb98z7FJZsuGTXeoY3Cy4f5YvJRcbem2pRoq7
ZYC+aVqbyWveXwzXpYd4tRYI+Nt1SXU6FQwCB81Zz35SDtvDWctLlNcYVHMAcw9wo8c63YtZHJOb
15OJGXc/k6CbgaMSnNvrhbl2bcAK2zL6odvWIxfazT9RcRETCLw7JTnk3oR1eQ+Jve+drF8G49nb
r+YPXRjX3sYneD7GG4IrtO33fOwbetzWAOjBGMvVh0Z+Zhx/P2qp55OGSwzOnE5ZXG2ChZDqk7vq
AtqrinfAXQsbmDdSKwI+T5Be++VSiQXW0BPFspe3D8w7EN19yGKnbTSXedNWke8gU19cSO4DgSRR
UOKJ/Eoj7RlKUCW/pOX9J14VAOi8kBgV32/Ns048c+LZTlfP61wQwuB9tA/1elKLwGMPFp38tjcg
K5BPMfDncI6rC25Wbef0JLHHbpc8XiwWstYjL6H/EaZlniirfyDN5+bGX6peA/fQBdOXQfPjwcsh
wb5hOtTPItAgbLSrsNONN309tgLxcg8m6UMeWHG8f/VCPIADp7ndtnI4HBKUUCPZe/whJvCuaPTO
vczejJr7Z8K1b/DF9rSKrsKU8k8FlYbtIgYOs6j3+DGLNqviXUNyuHHP3vj6J8FN8Zv5F57n3sin
rcLPi7PnoQ7PMYD82Qczrs49LMNMQowGWiJ5AK8ggcvhJplJavVcZEn/uE24djscV2tlMxRFK7tH
1TdHThUETp9M+zYxKHTIy8IlRMORaCnPMKvcX8t07kJ/lCE0pFt4y1JGpYLuhDvnZ7PdUsuGtd/A
2uR4qHisjrxjO4YHCh6utMjASLhtHR1nFgXRAamD1akAgLuLsTij0bqjPfJtZjehWdf+Mhd4mxWA
+kwjMNkWIHJ/IFQGfLkX7exST0NNk2LTp4pMBz24EsZOVe0iXjYt8EDh5SuZTmnyCoJbEPIDaxwc
HHl46cF8yoM5eEZE4T42AD4twVNlTlFY5jL4/7qOZhQvjZEPfqx8JVwDfTserlNf7fgciddov5vT
4btgI1KxeWHAgI9Yi6M1XeLC8oCyKD3j8KwcbWobw/rzPuIG9zIXk6phe9mL/AZvkk3HpqcNB29x
wM8kGIJ2avbDMyR2ak2DZPYA2N6I1tCM7AUIKwtA4pAFN0euuRbtZs+zPBhSsncXYR1XMBhOCT+T
wWpKVV+HhUx1SkvXoIfizaF3iZWPE+S1f0HXN8ZlInmxzACEuY7gcfP+mxK6S61N8s7DlpZ+Wi76
dItkQjH2pLxOLMEynQwJ7RreF97W4jZ/gldhxr4sKXO24ueH93otyd0/oiQV9F3wNsY1cwJ9b3xj
Mx8adwxxw0eWFoaCjSu4TGHD6QlM9wijJN+Ssn048b4fGCykm2DfTLB9zzw3oXTp/cut48yeoQqQ
OBZa6+fD9pR9qoZbkpMjhOO0xlSUA6KO4zPc3GHp288oboNwgbqjjyUrUQjVuPbt4nbF2HLGNhQq
qM0fIqTrg7KI0SXE6zpRvxoeo4GT8HYxUIUaVDDPDY6ruUOap2ZXiVK1zo5cnlaEkqPEySgKk+ew
0/P2zMjp+6dE5wOOEdYQ1KfBULkKTXmwHKcvjNP3AlC2DE+/NZ1KXEY+clN8wYpQsCmQEAiTNsQ/
Nzs68rAsCVKE2S3tvQe53h8sSsopX/i7Y4BgxjhHU98K+zfh8A4+2I1QPiI+XdxROx7P49h+bNdj
bpgSX2nQx7PtxHV1cx4TqPyrq9Vk+h1bBf/7d3h1tsB1M2bDSZe8FILF5d106DU+ASC0wDj2EgFl
++dNhgV+RJEWP9wlhtxV/xtbBVua+K+ODAM55AszLBXvSRL6SbI6aLlhYEmfA62nMEBfo5ZqufJP
QuGiSRnZ8X14UVsCoVnV2415l/kWndLivF//TKKJOfTTXjP8kIkIlF9wLISG/6m/PObCxNafKvjU
WE/rrwZVkYkqIkTjk7/TMtrlwUvY1DGL7iwM+UJbBSyMq38/sK0oli2CaaRJpB+qiNF72JCtZylf
bjR0F7xcgFSfCuoa4jiIO2g24W05MRcc0YfVAYz5SzUAih+tdzmp3cTiDfvXeXR1BDcEbRkQohuq
7ra0oGpSJHfJ0nZuKaSL2xD0fnN5WfRqoWKss+6swZ/06QzNc/8b+EI1pVLUct4EsJQ3n9YIkLtS
4Nt5SKhK4q6pWFFfDYHaRyw8sn+SjsMZmcw3Dt4WgwmCIE+P8kkgRyeSg0V2RNwE8D6BZA3/EVs6
cyv8M9QdY0p8pqqaZrN6xXM2OG1m5uj94suvWx4xh3205n0Xnoo05lskQb11glARdMoUC28Fi5N3
OXAEcTp1CYexDmr5FxzQebdpum5/6dFDOnmjQuz+Mz+1II+18YjVzKkqZY5MPKfzLrCv3UJCH3jX
XtYT6FS+yQxwzyHzgv07JPZh+6EKZnugJqr7KybeWcW8Uztl17GRBOyY9i3gycPxL8b+8a/QgFgN
tU1ZgXCbFH9RcRHXcRI07vWOtQmgmVC1Di9pIhTtVB8dX2C0U2RIcgtywbH7FjDnoSCf10ASE2TU
2iXCcPSZuc0vf5FaGU0ie053rr+vXUboDbas+mhQC/EVz913BAl140RM8JEhB1kn6yppmkUzRA3x
vpmYnI+b1K7FbFXObNn/BvB4fTrc+BjZwaARLMV0ulMS1NgLrB8DqQyd/gUis+L/thUVMmJS8LMo
9eg1vud0H+G2y08kxJOuw47/JN0uUO+ZA0izOzidx3Y4TC8I0eU/kl8uIStstGufx3y3HfgLbCdB
laeEp4WkIAs4OMVQsMUawkjIfJGhDrtO+j/byTr4Jq47ma+B0sfbgKD90YkQLj2o/G356DWSQCI/
/91ViehjjOTWQJvYq005q1BNYkQOEZBrMGnmd9w6lFtvbQqVpnwzlHQUhGKvnXb9kGiZI0ZPwnwC
Gmlnwjvio4oU0JrlJMQckI/H9zNoUVEUUAx5LMAO6nPhQLDr5yWXhfIV6P9vPFx2tOtxvkMidv+J
UfPG6wYUJmddlnXUA45RHsMaHIhuqD96Qep3x2ovUTwjRHlz90+O5ICGT25RtVlRT5k3wFEEuAlT
Yw18+TC/BJpNliehM1evIJiA+dpJ1K6ZWMYubRB2kj5Gq6TY9V6GXffVBJz8dNvjvjoLob7VwdXw
sfBm6GDe5lpaZg1olP0iH4dJZzot4xSUXCRNTclDh3B+cj7Vcv3RLDXtI34+KYApzzCQ0JcE/205
WUZ4WS5bo/C/xvpr+v+yu2DcNgt6ZiYjga/R2FDYh8uje/PkWOYHOHmXgtqroqPoI/YlKPteQEqQ
53ID4rcYdBYvdpzEXJqWTs1MTS50X7EeC59F82C9SYJASE0rDHTe/F3Q9umg20Kn4dPyr847IrPJ
alCpQv2JV7aD2FKhUqEIHASChWgghTCZyagb+WOIUmGIkhYmwysLKUHKxI8gGaKgqijiu6wGKlXQ
MfBUXhOcwmrHvINzr6yKfxI/BZBkOBVk3TAyr9dD/L4RtaQr4pFKIZkte1Y8Oshrw1JtHNp0rb02
0+8AQqEOsphqBloVTYVtOUICeZrCj0rLIqGjcgQ8RVB06WuLejJ2l18AsXxHQ/WOT/jSTpAptRV/
PizGF7GlCI1pEk2CKJZ0lPpOqykXP3q0m5I2hYKuknWr7728Oc9OXoU9dnFvikZaNRiFeInaYxNS
SwTG07+N2ilUQXnpm9CcuSrtLCexpTNHrRvoId0cSaC2e5+bzTNy/50Zj+8reD47qUHL9fxOwrgJ
5RxVOUswalJcAmNBdRy+IEwXneCuiGSqL49Bil3k9B8fROtTsVeL8jbuDNbClgSI0K3UwqGSb0yi
rUa1/jBo3hlJCx01xiLwkPAvREbHn0uUxY01zvyQnFFUKQNv1adnsYvw/UzB8hmn8nTWi1q8A1mn
jW2bmpp5toT4tURFhgGqaB7MHcAZdsFGvU41AjQu6Np/+o+Q06Men+cJUeAx2RcN4edTxoZrqdV4
Pw7slM5I3bcA5CvNoPsxVgF2wqaRluUVCjLMBkXom3kUnQKVeBsJvi+BGA+l2kBtVW+y+9h1ZfJn
ONVamvo0LYaeVUbAfQXVU8IJ4Pb+nNcHukNXQrvDQw/+i7rm/TrPcSLOP3mPKxYft03IJOBzu8U6
IjUpfS70cBO33qXJ6hsiAUxAj2NMi+EFLqTPEA0dc07KjCBXsZYRPunsDWkq/EOFhxEFVDvhRZBg
yo2keJoeumoAV4iJg2gGnbVzj7iC4YVysw+TJpp37YSK6YaSjoLUOFCLfNefIVjG7ZnxYHGMY6xM
LsEAQLQk8QOQCkZrVcz09b54xu/jmNUODWZFXtbhWIWe5pbtf2/6Sap56TKpWpF1crDhYgKplxml
xt6M1koJ+sykY1fpttc4BBZylkIbAFe5D6POU0Cjm4G6P1CzQLjHMiVMC9kpFUvwqeSYxJzIWdGK
DER6FBjbENzYo1to30eXAFIP0bXsqoSUeEUR/HbG//M6YT6KPJOo0vdfW5q7hELZtEUWveWWgZze
oZRMpAC00GXkz0Jm0Nugp5VBU+JQEQbGz3X0AzSsCdt4IbrDDy8Ahga6rYvArR5fHmKunbXO2NVi
FswvRHv3PP+SNH5f+9RzOXx7QxUb3ODs3cVk0WyEbh4CHu0BLSpMEy6+kNTenCkgCyZ4mRHYLVQs
DS8ulgBMpdB+X6pkNVc5oJ4WtUBChK16VdojCp6xCO/xzPTht+7Oaf6fa4blpZsO8NkvC+q0eb6f
AJ3qwwKTm3yOOgbRPg/uYWIOuh3PvrtSzwiNcTtvOos3cGCvFC5xqubmGXpvrRL8fFNOndEUiGbC
SD5NUTfn8jBMDDiaPM9ONfp/dk8KlzuKal3m2p74oed/qCoVs9AO7sfkcTXlpNQTyqi0Snz19SNV
Axoss1OaeAtF/I+k5NM51pA0etYz9ELEcEOsWSEblglg+SsS9RyrxL3em34N8B14T7XMjeQYUy64
nJQEMu0WsCyzuH/o6gpKCXCJxd9kSt3AwWW+OV+TS1kXsDzE8qaG8U9khzYoHMcXnXgvZFTtSwIo
Zgg/yZ3AV17RXQvzCk3RhekgQReDnUKg3gxNIOLJnQZ1qECvRMBjEp0iZKDW2tzsJgXvrs/XSbI+
4Ij/dpgE0JsVDKo934ApGgKlJJU7Dof+urErvr6QaKWSwuwF6eP13GCjJuVSnsuWTVF6euk3hPSy
bFpIPX8fY+hFeVND/IWp60PKDXXdk2VUm8V3GQAZKCAxJo4QX+DLqZ4XzuF8YNnF4LeeX2S/yLaP
xZQe7LW6dHwKSCxSGg37i08/1XJpl8OBeLo5dDjhMLHZhnwcQhEp0lbXVdQ1EwjpMoCK1Fc8nIaf
HH0bwXZ0EEPAFaa9fSdy9VczUao9Z5ctMTwtB4l8lZBf/tPuWoJqsbLp7SRkjx9p0T2yH2/wNN5P
hbmf40Leab0uZ5dGmrAuM3eCDTI1LHGx8vOo8X5Ff1If9mzQq1ZF6b2x+vxEhkYFUzVwV2LctWa7
3lxIMoUbp5e3cSeJ7Ssq7UjrD2Toq0nod3pdc4wnjYqKkEFCkrrhGwfWkFMcuh6mFSXastIQbuYX
ePFmnkDT8ZoM646VWQ5L7K45DmfxuQWmLeCN3QPVJxXtvyknxvsdE+9FU3B0M1BA/kJW/82/oVi3
88xRIS9PxrQ8SIf/49iTRny2bQ4U68KBa2aQUQhDQi8DqG7bp84XxkHpyY3T0Y9v6jtYvb2ITXHi
P1I0Suc4B6zGuoNwvBQbmj+qHkfFlfHZJqcRTllxsuNG/cZlSS6z19Ja5kMSaz5myK5fHEjk43vm
eXggFv1ViLccOJW1Su39aohFioagok9vhxBCT9m/FnBX/bDu2TV0/4kcM9qNVeGW6CKZcIBuOx+u
q5K47GeFABZUIjhsj3b/pehP2ODInd+FNK2YhcX4d8x8s4xR0x+9rrbHL8jbJyAQXZx9LMj+oEON
EEYHFUg0ooBLRwYAokr52imoGGiSi6R0KpM8WZSevIqkgbmG1qftykXQ1ZFSm91ErRZMbxmt6nTW
PUdgwci9MiAChOgs84S1D/IlR4fVGVdzNuiY5u3f8PlsHiqWQU+DfxY69l/uhqOJzh3X6SjYFwcE
9c8q0w7dy7za3uaLdPs/Eoo6Dcx1szoXA1ted0oDD4UOdNNjG015y3MvqMgB4hULJ+yc2QJECqKR
m28t+OcBKdDiKFMuEmUOFvUFdVGS4J7dInOKb5KzrUAdpJO+cPYzLrgpTz667zh3x7qADVfPZLii
BZSDRmrhRDKWjCPEAKqnjM0FkpFwyzT0osCTlG5XsMDLr++tIqOGQynHL1WJJvaMNjHRyWMRw35P
CTkK3O/+fGFVBZ3+enO62Qn/E1vU4OKS6LuQUKk5Hd6q4F8GBhHtfETiSAQ3wCXohaOvelnXifQF
/cxiy3qFV5SQhp99hSvpJ2LBrkiQAETDQa01XNK9Mw7+Zy7jrLhkr/dmEQpFETDSZuro1cMYe2s8
6uYDmNF3Tvtf177ojPPfqXc0BdUClr67qc6CoJcK6a7P8FmLsWQ4PUoIClTT9ClDHscQjHA8mxoi
HRV9z0tunrlV/HI9zvNddRoIg/Fg7YaorbEfxQvS8wi+KM9KFKAUjrlrGBSV3p1HLqMYbQVXdkS9
MD9gknyk9sTsU13KUOtl5xAgXYTdlgXzQnoYp1bvhQOGqoG9jfy22SWZPB4CF1ZyM8WUPMxwNwLo
Pu9yOgdGs1aOdRBYBTI+CbM9vcktM46oQ3EqhUzvlaXiNQCbo8W1z/iEOFFcGPfN6AbGJH3TCnec
e+NVLTe++5M6xPN5YNI5aS3W9ba87UzJ9GVAuCbQDCw7pnSFiKScydKkJ/tHHZzd8KZi/4JGAsO2
8SMDmwkBzIh4JorlRVoT+6yRyyfiD5OYj+ucvcxaQ/v6iPy8IC9An+d7LPwUvoJcnUSYPs9J3FmY
uZffZlrUUK6cqWOZquMKK8gpgt8YaV5qKSpiN3K7Yb0Dc7zp/ONr7RXZ8RA5e7p+Ls+z/KbZnNr/
t1r43DtpKK67uYlJPeMdqDvQhKTetQQfY+cz6Qd8HW7ZNlmSIzmuxTIs64uqYteCsyzJjdr+A/RL
gwzVeT2t6WHFINlPTtOs4wevyNYGQlB0l908l/POBccXG0AENLglSQc0gY+IBnb8P5pSE5Y3GwGE
41kevXxK2nl1/muZLDgwvsOSOxU8YKuQ0vT4uqdKvEpiQWLCPdyOjm5C62z4FqEDBw0bMNhyAulX
GhyoVq2tYeWdQDe34HuNCs0CgJ3f9IKzKm0VkSsZqzNq+LbrLQFGFSjGkFxAHTPUlKbwka4Nq0Je
NOFx9GM2QHuOyLfAUCuzypIj6D6uWreYq6l0w5ek+lyxNTNQR2DmfKD5FMiwu6RFVdVYUftcH4IX
Wp7uvB6ZDJ2RjJGJsfpCxvk2B4723uW500uaa2JppA5Gz8/cUw7Edrfh3hZ5DRkVzbM8mXwRyepS
Hxt+Q7OE3QErbW8GeH21yiMWkNWp7kNKolFp662ytIqfXcaVI0gN6Ax0jQV6IzALPxY2WzoolKE4
2YLbABSPrPLn/mWxf/2TZV4nqrhgBbl8Ldwyy5uGctfwDM9N6pltpMrLGC379rlh0zJev18rX651
R3MqA33y5CAb/6L+z7mJ20N+Wy59REn4V8mJBvzy7YO1PO/OpG+bpCr5+XPY3wEnwC4z4NmkROCr
auwZQksliUDybILQZpQONCS4q7LEs5894z2S+MpQK47zAQ6jl9tmbrJbm1454x0pk/p4JkyJCCxz
ZTFMWg3mqDzmzAhryJQVZz8G3iodTtm9yx01oGSnRPuMQmv9Fc19PqdRG8B+xlUARRVBgPXsBoKv
vHw4hJNhXo9rNfs1cWYa8XjXHGQabjIsnuR/OMEeoIDKuQ9Y07FFS4j1THbQ7C9O7Sy8hWICaMrg
6BmVlDPnjDF3n3AOiSMTC0lrHw16PmtuItuxR0dRv35MS7qX0oQVF1FcozVzvp2HbDn5klJpXZRS
3h+FGAtKhzZ0U5xMgDf1uX/sY77gHwnLVeRjsHYKAbr0w/INxLoVtLTFtcjO0b6n1njm3pB9ra4g
1PwYyRnn798H3EuGw8CqNQDHk8SJw7iNqlX9KvFyXjclhElDomrq16jUPS1lqQDyfl3lyusVV58W
esPWpvot1fZsTcq1ZVG/xdE4JwtEY23vxvzpGDCJfHMRB0Y7XrGBSYpzvnBJ/pUtB4JQBg9j+gEX
hnA1k5xGjhy+3wSt5SarZisHyZBiKlubr0+ErjHgIUDhxKW3LqJ7OZdYNdNgehGYTw1agmlliaTa
P75hDZO6acHzhGfs2e604F4py01wo3AxyKjeRCAWIgPuRHMJrjYBu2qoyj8vydcUzYv1BRgJ/6B5
HicdRdpZiPmjG4g7oxUV9ApcRoz9llsjJiybDCDwzJVNgUYl9P2BVGc48Q8pYkeohrfJXLTejiE8
7GeNvWXzAnHzvADH72L+wzkeRHcwCLPfiwdadB0XHy2qo6NNeiWxFn9SZk9Ald5gBN1PW91bvS+k
E/qLjAxzq70mzX2QdMODj8OGgJ95IpdQyIIchmGXoWjoKL1Rer+udTUh/IQdRuhRf9SK3HllPa+E
mO3jvERynZRyI771R6IYXO4k5FeNKWkcuf4e/81nwwUCm4bpV6E6TWr8qNU/FKfbyhguPs9tVaXV
6U60toJyByX/XbZf7sajIw8aGgTEC6EnvRD6f0kvFJ5FW2lQEWJPJFdUrxrJGUIWNuAvN9Gcl5UC
o5BiEn7xaX10rnFq3P3xa5/AuVAabXSSldaBwETbBuYJDlobCFaFyT2gheKCUbEi1clC5QM9YRNF
P+uhVzC+k7eZvr868GGRQfa8lR9YOqu0YuZMy8709drrGvwXetmfcAIpraHqsqcb53xFQOged1m4
VadL2Jn4kBUKcjLHXpscuoh6F1hSNNHgFLpZ3vkNtkMYGsEvBAgulV7fRkf6XyxZ+lYlY/NvEjZP
7JzRcjvT0ZBp+kVmV+YmFyXOtHg/gNqUmrRdfT+3oKEs3E8dZXDTvKeTJasYizYA6CFUhXTYouzR
m+1StJyEADegr4kN2w8gQzj/eM0ZKxwK6FiNFVK+F2A3AjgichiGbsMV9IrIVtCeYaeCuCS15NPR
uy7axeyxAFKuc0+pIir/xPqmEMcgQ3oEFDl5v86TsiQoEu3OBLxv5onDgaOEkYUVfJPMGFpifTo0
+zggWCUNtKjLOJpbr0u1/O+wD9Xu1KRChUn1uaB9OFM8gI4KEoIN+bR/fOeCrIcpBuWqWnvlm34o
BZay2J/tLg45GZQWWXS/QSCR8loGFNrny+vIw0QNDKs8EZe/h0O9KO9TOX3BN7YG84GAs1Og6SRf
6ixm/nlKO2okAU+EZUzwg5Z97jxTVwKRMopq3k70yJZfbgkWgoCL1xl+ojCLIqkuoMyz2WgC+L66
OI5aDACEKIlPDoeQEyMExmJneIVbflbchOy6YvAHoCxQCia8hMz41Zi2/Nuxw4LiOu79X2f011gm
dP4zcmx6boFZGv1Bg3ywK7VKIIQ3GRvqBEU8UuNr+v8i5dNZT0JN7M9qH0rj368SctoChimmk3vR
2mqBKASPWwxEtqqggmjXu+FI+kDGVb5eiuvdvCj8Kt/KeoNt5BSuO6qDp21LvpPoV6DMPF1jSPgi
R/N4pOJMkh5WQ/ui00TPZQ/FI/2AxAis54HA6QXnHUlE90ZkXT+Byb3jN93EfHFu844GDn/vGxM9
tm7FkYm7j0z6MptHI2yAlJuHWelEIXLAYUIxIEy/EiIWi5DloewHlozt6s2SdCRUKvVfs9jPe+Er
ljMkav4ydNzNnZAU3fPCNEmTndc9b3JHGHOygHKVIr0+odeJVpZSnDdBZhG2LiuFrv7Kk/+7gFcH
TZCr0ReDyHPB8GVpNHIjIWF1H4hCV3BU37gMhFX47RWZSrGCIP/J3F1OzugOj8XsNVLtRsOs+T7B
U6y2BHifi6mW6G7Xc80IejMcpF70NtNKn9fwuHiS88zjpAW19Ilhm8hfgNc5HRUSPaEpwCp4Gy6o
q/UPp81286WyPM5WDtDRFYcjuTtrzWlEEjr6UHAMpyAbjP9t8MlhzS+c5JhvBocG/I/uBqNoLECT
K7xxyW90BKPy6z2aYsRoxKqZ/fNxOCTlXYhGuiWiJg3RCL/9nrxhklnMxtK69LmrUL8iAfUg45ao
y4DcprHKZtynXIPsTaQhrm2hlYXfmMkExs/OiSauFRJe+VQQlOcIkApk6mkqf5ToztESvW0CwJp0
m/kaqVkKTWyQwR6jcnZM+ibrZcR/vt80tHaWAuIGjXsE8c7PqbHQoipKPCIRzIn4zkU4Ff4zk088
ijeZmT0cuU+rPqGpzEnkqR1gAtOkvI9GGy0ljhdK3DCVSsXa4Reio7EewC9rcb5DBs2yCbz96HW+
Y8ppCxw+pErwwaECBFp9xbhRvLJCtDYWP0muCoHXIvEYQsmtovlAADLNgVRa5ZIhVnp/5ZdmrH5U
g4n775n+B3nBsTIBnma5Pujf5+2K4/mJQNEwtAIQdebr6hWOdyFZSDjWrTmJ1uX/zUgmn0xsRw/R
w15FCI/wrd/bSsD1lOJOp8TW//a0RXLMPiyxL3PZ8/SLhRjYgt2MRS835tqaZ+mKY1BHglT1nJHX
A5dWojO/0JVKdHiGFA2XzP5KhbNS6LFF+aWleUvS8oO0EZZ1CYVzgVh/flWwJtcYtD+O8w+DEdHb
Ld5r1olG1HrXzEAl+I1OM7XvkSPYGIeo0KI+szNBiTpJf4qYiaMmi6d61ODpJDuyHIhyGy1J/p7s
jwPIosAXx9VfIvfPzguct4prXALl1++8XXZ9wCOPX0Ac7H7/YvWZ5aezcuroEvnVfGFAeh8OrPSf
4AtIztzDH/2sBkA2cmteNLamWxDjMb4ALWHdn4dkUdEAbsdTVfzd6okUPpp+POc6p/aafjE8qzqV
kfi6Jqleuxk0AnQFyxR+H3pTJoSTPvyGYPJy/T74A9NCp3+uxx7DMVpR8wt+AvXXLLx5KhPzpCLs
L9/95dJqCpK7C5tdlsfskAoC6AuQLQhWQcGJQ/1LDttl9FYrCC/yTnzHblUtYwXo65R5fGxI28cZ
JV+YAe8bsAMva7YqE8KUfm90R+1hrtRo7eaeQ5Ln+xZILg3BT8tdEVVgl4F//lnx6YJ3ZPNRWISv
tQ9KQZQZBuC+g9VZwSdHLVca3rx7BKVlocE8ezX+pc8fefwhZwSDGRDEUnRTUNs1lIKV2+Yq4oEx
yAiyhX8CZarNzhi3XARHShddseTHzOUQmSu4sJS4AQc9nwNlc9lJZ/vXhZUdLOifaZCYZyp/odXc
7hbKuB/ehbXbiCecy1VnnXuFu+XzHT33ay+Xal9G5P5VvZo8H1lWIu4Fbc5lvIM8SeLjGdyXZqnr
PxpjNy4WY9oSbLAFWM+udpt9YQHdKbPfFO+p21GyuhaeR4S32qsw+aI6EYTLarTmttQdHqZ/cL90
c0WO2B9/JOIx0m0hcwbO2mhRI24AtoEilhoTNtfnAnfIim24O/VCvKwofATUl9EPolaBODQxhgEl
UXeBO5kWkmHI+FPGkiPwUmfQ7+SY30108XjltEFR9f4dt0wcn1G6ZGd3oexdzZxZX90ujx4PUhKa
jkbvK4EPLkfUD3HcTyi/lRzsYy12iv+JWkhqP7dCiPPRN4z+Re0nmug8ccPqiKqkxfj952AEg9ND
ApW5fimWvrCrcgDgKKGRkYcqCFc6CSqk59ihm9DHgHqNYqM7Fl+2jTJjjqc9chQOXOwEDBkb7oas
RRn/5r3ssX6oSyBVglxDVZDntpa+exI5fi3mK3XIaKU2zn4y9TUjKWK7Q+Qt1F2HKl/t6Ts4Eejc
hHI7d3Dxq0QHaGxTg0E/+mt5KpM+g7dwus16SHqYy6mkjrUz9BBnL2gUcjc5Ys6oLZ47DCPrTVqh
D9gY9tMn0rPmX2oOE1WamZKrQKTKIircFGjfBqV13LHAIcpo6DQI1OihaPAKHXWUj5gPY//CwkSP
l3qwgSKvlTCS5G7G8nvdRffOKI5BJvozWxg2YmcrF4gtrktgcKW5UAgvCA6WZnh3W/Om4FKrdrWa
petOTlQeKn4VUikQYzPEEciGKDMOo4ereW6nAGqbA3bqV7PaFRqhiQ35xZ8qfqlO6ultrmlSi24z
KcSvmyZUowRfW784N7jWn8/Z7UzEdK73prAIikc1UmIcAhWAbfYFYGdA0vUffCYYAgoyeIS7OaRz
UAm4yihMmZQOzQa7V8ovoTRS15fCYbeBeW5VU6XXbhvroHNMKLfdYj8E+LMAR/EC4AnkpZrOlg6r
U/cvc4wb0MQNjjIlg/wC55PwR42RTUto2fRR5Jm/v6C4IbdOlOuIqR/DZPKh/csBLcNupQgGN9Ta
65ui/aviI9fcDaoN+LjAjvfeEPTeT5FJM5H/bnL7YUIng1mEgJjNkHIHY9Gjb8fdawbwIYc4cSWH
IH6W9gqZBuGXbLeuzaCyvzMWjdvOMdN5K2KNj1tLwrOkG6lAe9aQUSN2Br1dtad7yVk1ex4KvcxC
6hkbibXcspHdmE9CMRTt0/FhfMQdbMXvUhTWxdk52nz3IS3sVLoXzLupW7pboa0OcUcGg5mi/1Xj
g8Wgx0yIQrXMt7cg6iV2Sc6ePIN75syMxGLJ8lLNHuf43HCIczascjDOiPaM6X3LXq5zjv7EP5nU
FJaNeAGENSbphA0SWWZXpUThQgvXlS0UTDiR9iP0rmDiewFJNC8s2Q98sfSrws/MH8XGteG9emJt
iwJW9N0Lo0iuoZ4cnwk9d58AhmhKYKT6IlySDw+gkdfGz2a74CvEvBft2uHMV5eiYrxFf2RSPGS0
BlmBRVU49wynqqugQAXr+d5T1OkOhXajPsI8got1eTaZSGapNWxk/jNAxwtiZKvh8cXHKS1cxSUl
D9iw+bl6kXXiLZZroCrjUEr0lXZIv7QmaRH7Yr+eYkxD5eMXZfhUPy+xrz6u9+4wR7PrebN5ijhK
qw4BSc4qA3w8S/QhwK+qby7bwjJsOGrYheOIXSp/1M4eAb27ViXVvSZv6nmcK4W0SfLtTmrrpWIk
7iTMBaF0v/e2zk1Ep1dwq1Xfm2zh+jcDU50EEBimUfrHX/ct6/aVNBOCVQualzxS8JJzDoOVIDbl
LFxFS2+6O+tRXw0l4kAtlH8VOtROoXuPourGJC3jRNjXC3SjlRPKqFaaTlIgAsfoBLNukmQZZuwg
f7LuDULQsN5Op5uhZRLs8e4df45ZlmCpIY6Zxlv1qVDzLaIUo6xEeIKQQYY/lLRlQzOa02leY0p4
FEmuICoF9fTvqkXcOPesvYiJ4Lqb6f6DkR+R1fEtDvH4WWQBX3ICGTQqtDrX4H6/b7+xt6bpos6H
HEhXs2vAHtwizipa+MO66MdnCY81hko1qIEOfeI4j7jWGWGbLf6qebJIS2RWNojHjHECeu1ap5R6
QjASD8ZIaM5NM2AbqJgqup+wBCGVz2/o0+4CP3Pd0bZF1BeXw4SPXjCZBg7higwDUNaPoQ8MB5lf
9kFEtSS/zb7n1wNR3ATtOErJoGIjUN8HXVYw0EvFB1Sh2dm9UA7MglOnKhzm75i/5aHb+MHiIczq
7k3QPmnsntuvksVQ2WvpZBRebK6BD+NbC6MFzgvJmKmhUZYUgXwFP25MJGUYntvSGkC37pFnL0sT
+45hSZjHXluDHsZKD72kai2pl9atqStdiCU4/G5Z4qz93FN96Q1UTVQVYBM8lALn63ntc+jF4DX7
9PtyCY+wHTKJD2yIYaQhqQM26LkJG6i/qyaFMp2SLfHbUahPwOaM8Xan9DVvILkNkry/Nkdt/ev5
SJ1MA/Gdc8sJ5s2nI8YIiW3SKfy501WBOsrdTBxuox3+DF7eSSelDIIwhIso5GzsO/ebVkcVaoL9
GxCfGqMkzWcY2b0/qsvkquBLVCsCgzxCJAUQtTf0lIkv6/lB2aQ+WxJjb/i/p8E0fYiO+Ol/bP90
CSIhEIErZ/lv0XmDZBaMbp2RS6pj0kzBWo+GR4CS2TJD0+r/EyG0ulE+dE7Xq99TypLxYoHGSEsJ
11C5ajbgMegq+uyJYqaLM4DFn2o2iXYO5mdKctNFjuAOjpgCVA6e7nxLZShBtxZ/rD7wq6q8+Sm6
Rdk6ufteh+4Aaj5uLggnX82ZX5aSFWekh2TJMDRiqLbQ/7MTTLvk9TT3fBX0Xf7ZvbLZYlZXmav6
E6r4HDSGe6aMzUH2p7MAqytVky5LxHBtScfOuj3AJxj/zjud0kJdF1ww2glYPwQug5TCrXMk82Ke
z4moz+nq5Nw6MT1Hs+/lGoUsSc8BPhhdWw7MgUx6N310i96iVx1T0tH/FgMypeugka1Uh3c9UDh6
h3mn5pVC+Y0kgEjsx805qesGPj4Xuuv8GmkiER8PqDHV6fQQv87YPd9d8YoOOYhGZd8CzOxAx+nj
SsjLjDA281zSKmN+RMZOwgArgvjx0m+FiXKmb30TvcN2baxovuG8PP2cD2pbtLpj9znxcGUFh6dU
h08KHzfCtjlObU/gup3CNiCuI+G7Q7oY0CMZrSaeoevvs88PAB10TBmNkthD6idVDq0YtBjg7szY
36CQdQSRGGvCvvD91FLa148Qv67CVDHwPjZW91r+UHrjYIyLEdtV+XXJcLWwR4DuyvC9cTt7VPM0
8oM2YUgokkYjO6/JitOnc1s4hztDO9A6cVMmmb+0yM4XTvQ2ZnaCv9YWhvvuL37mmM0pV9QptdbK
01h8pwJoi87S/DQhldaQgU7yIas25pZGmlnAzqffiC23OSF6/W+La0wZD1Skf4ZhAFdaDv9wcxxo
q/MHKSmHmFxlmmrspM6HlyDO+2khm863zHKuBv8s8aT45E4OruPge2XhJBhjDRXdOG/E0wrZ2KpK
r7CxHdXxbC+e/kQbQTEL8Pe8LKQIqmqwHpGtiTn+yOcuoGTff2uB9gdozl0SgfrNxRkgIOIvULwJ
evngN16mPck7xHc9zeWxWUBAkL7NsWNVARFC/axLnsP+bT7z9AvLxHa7sUSGef5hi9Feq3dmrZvt
wblLNCt7ZjBlrXC2wNDPec1F93uA5Vz5q1ofkHuJPwdSnitdQUJhvNIOOXmJR4+3izj7MxNhLW6P
pvlBLY6F5dTorQ99NOarPNxXLZPF1XfhTHRfi74LBNit9N47wQxz/TC5eIBdlXjfKT9MZ+VpS4XU
Cf93r4HISKroNmU8WB7PClm1HfPe5WjGsEun7KlqrbLVaxaO8S7eG0PalKns0EvILuKaVW9Q8SEt
LcA0MH0lweSEtZri8poiN8OYTFKb1phA0XcBy3o9X1OdgwC2kS1Slu6N7dZbH+jeKvsjKALzHLDU
elQAJLJIJWasOb5pcnfqo5o7RJELOWosPiVhnuH61ano4BhOHjzHR5ODAI+9SK+zCOrqJi8ZtiHH
vBXA4voKDP1mJFclt4Ub2Cd/UOOn104NuPtoKDZv/nYu29Uw0WlXbjBOWdkj+SZnOnISm++NjlKe
ZSfyZyoofer9VaeUIu6l1K5uMv+ZLM0pDR/uJFPuHayqt9eGC8X+CeBXswUMMtex8OCtKVcXaSVg
7yFvXg9Vmd+99pb0RJ/uH9Zto+vVESm5RzNxhNKjz7z1JeZCxn40/QJBAYnM2CJpVPk0ZmeSyIxW
aO+KUB52cMGxfnAO5wuyqnFzt/yeLifprqADODVnw6SO+oAOHJnmfyOoEgvMlKjwU7iGHeHN3EVm
NZ8JhbRYgwVEeWPLA0RKnX4xaTizMn0tOJCbdUN/uNznvWOYKwz2jamEvki0F13ee5nUWPQtZbcS
gx6t1VqsC1FUimKV0cLArW7XERDCC14IM5KWefNulz0wD4ZYqlXSDJe0JT9LbDTDn5FR8+j/NVmf
HEvaoPw1hYbFT30Hg7sNzj+G8lEOfV3syVIYzHx/nINGCJD0rNk0MGw2T15U49ny6DJm4A2WgSkp
hqC8N+ANHLF+k31hWKg5xTIVF8nNIhfJlGsm6oAEcUdPWhuZKdOGZ9j5AJxpkAb0WoZBGsasGf/W
/YQ0GUhs/wdFGsaJ9Yse7aHFv5BwGPx0qwoovZ0WQLAp4JyKj6OQz1a6wbxxNLp2A1+r/TrM74pg
7YhpZQQGsNSwJ1xdBuTr2kmJkhKNqlMIkQsrMP3VbvUCM3oQBBDNU5oGRHhQxWFbY5bUvNVKzPSJ
1ikDTLUsttdy9VbydD+qHUBrEWEQpj9+qzhzNIcV3V9C7hNKogj9tMkbzn5IY7PYEDctnghJEpto
duMozTPnKLEIM88CTLdwsBwhtt7BstXUosgbiDjirhoqJZU5YxtEP/Sa3V8FT0GYaxV32EAKTQ8+
hYpK46DL3vr2pIFAdSXOa2lKVolqx3KZ7qH6GwO+wfREXnbbioDMf14CrPsyiY/7qLoGMZcM8rDt
+kGCEyTx34lPYA1v269G7+EYL8K3Wkcjr+RwhUakEDhDDu37wLO6A66skajwqyQynNvF28Ibds2T
N1B3zocYq3q4KmHbKCJ7BXPjQlx0X9Am63+82isbnf+0U9F4s6mfLzKXHQCbiPgF5AsukehObaXd
4GwFweUUY5QyYEiU/AfY0gHAXluMh5mWsBiBuTMDB7HP5yCl7EgSQ3PTwtfsHSolX58DDSTSP9n7
uPzWMtAyfplo2huEK+MRuLtd0sALdgiJpVhK5+nXZn56jZdfIylnTbaezbq9z19eGi6ibsf+uVnc
+sMvHgfqYhVtkAKuoMnlUMmMpAg+JIVJVygZFpIwiJyfnf/QaN5JXPMr4NFFPUoeGGmjZtUi/XLY
74WrsShFpm47pJM+ACBdbV8tPNk3Ve0023L6yJH4WsfBa2eVvcv8534kZOb7WkgVoKluKWx8SubR
lefhDYEwG6jCLvYOueaBsVqbYxi4nSN8rjNQPHfMFqK02mbeAwvzfSpsw7VjWK6vrBNrfsQC6ihd
p9yStCpWAg3unOkUqaO9aATIQXZVUSJiXdwRmnjfzfj43VMxPkgIzHCPwd9tvuO0EMDoy2HuEyuz
08xt+2oKdRbNn9jJrJF7TAkx0mXXhq1+Nw3SqsZAifuNmHswAKSsJQWgGCQPuTjDFTuRFzJi4JPl
0X6uLOzz3jzwtuudPBCSL7M5Lft7jAysLhd78wes7/I7iWaNwxREqASDllSPd/y5OyFMF3Cuvmqh
dwMO6xoeCQaa1fuRrkoZCCYwnhPJnhyXhrGPmEW5MAGypn+PbQs5IUY1JT5k+dOuU9cstb5wZvb3
qgJx3W264y267IUHuX2L+Lh3tt79TKbVcqqP6ql4id1uABhcczLgsByKXsUxVZ0Z82k+dWDWcr2A
/M+2dYy7M3bWTnP+UF2t/UYqSeMs9iYZfz9j78Uq9DlO2tke+d/gsSYlrPgPzt2LBjEVJHsThv16
ZLowOjH/a/7ge+sijd2iHOLaucWZRpa/Hmlzx+A8ZaQs8wbsxeYXyE/JcC9QqwPf3owbema17Rbb
tcLavgRZ3Vis4GgO4qjI/PaWQ5gudiBwRSIXEW+7HjR8WhitdPYUgSY5qROOIV4ptRDRgZbIvDM5
tlT0AKavfEx7jR2yLIwILWmcrgvixxAZF3xJTnzqVrEGSTxB4apQDvMIuEUjHo/rYHPUGQ/6fhwR
NkVQBHGmDm8h+8EeczakWLuLbPCwt3FV3vpMgyigX0fLeg8As8yyLQ682zfy0eWjtYF53qqkNsxu
O6n/IXR0KRAseqU6Xgp6cAJy4o4eviI5dP6QbNnRtL/ojqxlgxh1IJc8/fkav/R67/9+9VovudlE
wyAn9JeDll60nOiyZwn0Ydb4WcgwXipz6F9wUi1GC9grgdIsR+H+ie7cueFyFWcJVvO7yCT35f8K
ltmuk+QnPylWJMJW+YEUE9vb7Ywt3FuZ3UTOIAfiIczfBaei4juuFLbd/Vy/3D30MlWDwj+OU/eT
YDTvDdPVXbg64Qv9f8xpR8VYKj5VZCLGBNA7EE9/QT9U+HQKbTdDNKwfYCCRNCyjc842I3faUCyz
gy7Crhd0ZAM0fDULd1INcM/FMqCFH0EeRD5nT2rSOTkOOyat2OK+82FwvyoTJb/xsKwFh5S5Xoe7
vKJjGVsa4FNOwS0f3pDBX8f1eZ9gYS5vIVir9o3yHZSCkyP2ExsT/Y8gbY/DhOGDiFPVr1yjCN2T
cw2R+JrQXsyIqSyNGTwbd0Q5i+CDiP473JqCBHaJyFtHBIwoH+v+Q+mQKKunftoHDgMGYiGUa0+t
kLCMuVlRrcU7nGvKP/CYN3z+zLxf0mnzqLEKMi5wJyOiCjctrKtjBmc5XXBVOHLMJ6+IlZz73ei/
+PJZxW9cGppC2ElV0ji2hg0reT5RU5Qo25q0D24OlLzTOESpunmwIxTobt2R2NEXxgbJOYT6affU
tyTrHGarBsxAXxxsXvJGm31WBCdW7pHy1+ocoNraVY0tnAsvbOWAwrcPqsODPyh2hjKaNSbDT9N4
urVCgZsLklKgrgiaCX8yXeH6E4oKN/Iiesd4oBsp3muL8I1/2LZtqXisRVZT8VY6QNC7exDwbv2Q
/RhnMQAZKm7MRwuVt3x370y0uuU79/W1yTOSMhsMT3EOi3uyBEweN9otAA7ELDbyO7GRsgDybYoD
V1XNssXCBDihoa3DVjQews77LBTPlLmOE4Ky0+y8k8v27T6ClOc7/yFxH4rKq7WHB/34Dm2DGHCt
3YIQWHxfbZ5m3GfhCu/FIWrXMMHcmQrNCzBwFgCf5dKjOkvAHEReDvSYIBFGvN59FAKbri5o54X4
MC/1LK1KQW14NZyV+w80IYWdSkp8jyWxNu+uEcd1KZbF/ryr2qtkHn4KGM1tVsyp4+bRNY2qijua
y38hZut3nhg7dTcUVCKC44wA3Wdz8Qq1XiVbseYaRV8NqHhIxgcaU7hrLma4wAj2OoYgOjo6AQXw
z/lW61NxYFc2ScyQpb/ecpV7cAEyR9A+FjHix17cG06d/BFja1HWrI8p7xJkm1mIjDtvGoUzM9qG
t9zVyi066gpBJvr7Pq/9CvpObvt+917NXe2QCcmDHDAamVPmM/jd8sXeERSn9BK260mUkmBcIkY/
I19ZhgwyLcJHnW+BxibA0yCmwRkuMXVadi8j9F9Mf5TiXOCgOaeJIUUYgjCmqtbjihNOOPXgKANT
1ykcccoWMS4d2PVD8JbO2IaDrkabHF4WCvaFhr9OUainbjYfT7R1MA2jKWPMhYo60w7f9bK80SxJ
OpmLS5UexljFHGVdT3SacPBY5W+1wXvYXtOzWpIHiJlBsbi5MtXfvv4TJqZh16n5LvsnQkLkc0Hh
jBXWtlJNX2K9SgHfaPWebm5IH5D1n/FycMWqZLjo66iOU7O3WpOwe5MxXQzMEFIwSCtCDHtDASnX
aLkYfo2CVr9YaoYZdSdbZGN33JylOkdQJhNEJvquwnHJvHoyt+3bu2RSdvDoihi/0CD93+oyw0zS
RsuS6G5/Of0KzYp1Z5BneZpZO5d5eXsaS483KpysgybkIuuwsINPTSmAuvyigN8HS/sHFWNPhXMI
WXv2vyOTEBAn7bXMKCE8HZw2Mgwtbszu4kgOKTeSz02LpF2fFP490rjxaP6f+fTqGk5PFlZsrZbq
hDE6MGqbPquEPDa1Ubwlu9tNtaXeoyhxACssOUAP6ewrw8zxvUYjPaEKHH15//Y8k4ztMdsywpvA
WBVW50d8fCrXaRhYhSfeEBJJc+EGenTGzkm0n3l38lCmO4uKAdX6nQw3sNDjxYlEFRt7pW4usgCN
9fEs583eOT9pn5ubL4X25NB3XO1hn1wwuLL4u5niQJahRe04bD/YpkgQyo9k0cWwm7fCn4D7QaAG
XY1qXua1DJuFeUDoe+dkd6nHjusXmo/yOHjGnStYjyWapHTIlX/6lA2cMvQPWlG520IlDybBiMIb
cXOSlkEW3fBGLbbcWwdHIOLCqjNGdAJmCtFCp2AT1Z/SI378Fd0qgqsC/FpEYulLaGbIn/AkEFGM
YXRw3xtrJMJWJUEX1vgtJCC2Bys+XaKiXOGIjMCdtzp8kTqOVdjp6PwjVLRPd50iCHefRyYcdm/e
NbDTnRMm7D/FG/gJGW8+6WlhdNcto7e8u21AoRaBvSoydPgBTa77hlOjvcHI/LqQ3jTpFR2AWd6v
4/K2Trx5pYVptzotKjy4thb8t8CzDdOVh5o6gpi7O69kkxidPerLPGbLDjP1n9DrX3lxgs15bSkc
cklW7fRXpBT/H4VKMqrcvWS7erdtw0O5Ep8DvTgXPEU5rEZKAfZR5WjKIDhfQMg0RxoUYPYSRG7G
bO+94i6Urxf8Nv9R9hgSVF3b6pZaYBfCiQlOfggOHTmL17EjroOx+WZzGsUBCl39IicWvgNqZEOH
qIsQlZXOAghxE7QVYIuxoNcGaR0TI3W/sFEQKhgCcqNVrphRS5RDpDXeZLMAPW01DQlh2RRmeWAh
kf82sAsudiFIgctFLSfy1JbnM+v4yus3TtX7j6tg0RQjsJkXBgYP0765zhBau4njjpEvHKfttDfp
mzPc1sdmTNw0pxNPGCf2q/vSr6Zzzx+c9hOFow+v5q/H9nPIZTIn2V3xnc2oo6w0HvUy47+s6jO1
xYYjfM68uRiYcCIHLK0B2hIJ7u99d85Rbr6rsinmFppLieWwcCfF9BFymJFs8ZwqpdFle1cM0YYh
HmLamQozLMxE2cYkQg+OwzNQKxFki/sE4b+OGe3SiC1QfJm462hgJQrpxIdR7+T2qeQK3rqCDrN1
L53QioFydVMmif9B5Dqg5qR893D03GIZUcwlq1ZbYMAH83LLNtmuB1ZPHW9FAGKnGzPWTOn3zJvM
fXDqjvqUTE7/lWh/bVsKXWklkA63270Zf3ebw+8xe3mv7zKrpgXKKaXOB1xoY8UJAm+Lb4N48mFm
NwachQuBaS+f0YXDpoF+uq3ylsK06OfHrWNXJgShRmCarprVRoTomZV9oAl2U9H4VinyL/Bml0E0
+o+QpLJ5OpFtZQ3fO4eXEja/8/kvuaNWw/PXNjl3x1Qx1CJnPKdpk6Ji+rMeCth/H4OQ3d/iRxLJ
vH1oujqw0RF1zOMk51STqEH4IgcR8n9GhpfuXvKt83fI6ir7H+DC1M5I0nPvuBKk/VxaQOBNlMTc
wdwAF5x9WxHHq9/n4iL+WbNoEXUeV7LAD+5knusdjMoiMSrC4VzgmtUsao8MIjWYxQEcVwn1w6ft
KEVONfEfXySPeliQ17lcqmrSJj8pDtk3dkTScnokNMWoODslq5ol/eZd3a9AA/HvD0Fyk6bSzE+o
owZw8JFAk0LmYFO+mh6si76r5hfMRk7E8Yzl7Ax7PdhubZgR+zw2wwfhJ8lCNIM3k9xVeKRX5EWK
SBKnOGmwHvOZ4ja1S6MIyGqHYHJduzpwgC5tgZ7iR9y0IAD+b2ywASS2NT/d50n01JHNp9TNXobr
PCJGAfdGSKjINgq52hYRg1gxe7WigTEoNLN7sNYJ9xb/3Q2CmFkXPVOgz1V60WfC12k06Ryq7Cad
AJOj5DRsj/xqCTAhN1S9zaCfmyMoC5/P7m1gdh8xI7Qs+cmzqgZ9LgwbAOWU8MqC0Gk9bT6C9RQq
io4MP/kkySEW44CF1Ln558b0stGjCPlmbbtBQwU1yIJlegvx389NTBdG9qje1vRNY9MNUMTYKdhQ
wOUTjCurWeEiepULoxs8ztI2OHQDGYgkRDf7XQ93k2SYi2yy31Q9Fi72A9pK3DeMHMpy/Y2MflDh
XBcH0K0SbVOsrFMbDO3XI2Xl9cRthiUMKR834cj1jB/YNNQCt1x96LboTNpcFS+ht4QkuQnP7IEh
QSl/oXYLefm9WhODvGfFc9A+TWR4NtjuRis6wdEp4W42JsEBob+n2HnDGhH2s2HZsIubHpqnEi9u
sz2r5Yj5NNHAahCikbeadG8yLN2aZNSTwN1fPaM8Ky6MdjWranDeJ+dWRP+yFHxSlceQLcL7DNd7
aR1hE/FOSg4F2KQYFcWb5nqDB1UYsBt+LZIYGidFZp8Cm1JXOLWeUX2AXh6tjj8Rd0h1Umzi7Zry
uI8GhhpnM0vawtVA3oEFeXI9QmfmHIDkHChtgLinJF3LMkZHSaCyp6KI+HpZPhKjFQsJlH12ai6I
rfatmKSPtwtxzFUYnew1uFWXEVasgdSp13lpfyBQd57ZimNn6CB801Ytw+ekzf9AEdp/PFft7btg
0a6nzXt32OZ3UpN2xCfXt4zOLjCHllSjRUnwYEfD0WKOASLWuaXKUGJcpX87Q/PWc2ylsuq95Ych
Yb3VUWqCP7Xiv/Nei0NQootKAKgyR99PmuSl624R2yY6l4d8QSfelaTYI3NEE0txhgRaJnT54T0k
FfS4URvCTfvOUVk0g76fTPzf3K6AEKPyfDLD271/S+SjK/teJBbT+PbPR/nypfVUsLJxbUAsaUM7
6ivqeMYt51IrOMe+Kcd/gPh8c+kdFd1BAFK022z2TrRHztxwGWydStqX2pTALoBW7y5uHRxpYDoY
J5nh5Jt40rM5S95B3XALTG1de8Qu4j1xIa8Ua5MSbYXsjkXJRh1933jnyXNWKzY1fCed5XusQUb7
cB+wvTR0yK8qCueln1QYUnrb8IilVfyjvnOAFXbgtmTqmzSDBgq4smP0Vw7mJSMMlL4RBHk+wfWo
cHV2V/Q/v0R8fSfzlm+y4zMt20jtaqCBYW4Tq3bHbdoUpzZqpGyNvpZ3JV/E1Rj0oDXz6wvvZ6cX
mKdOGtr/+1R3EAQsuYcM3nUnqm8HHjRAVW0Am+bzQw/Ny/IXDRvVHcvOuMwJraUHPzHfoVoO5N2Y
eLMprJ2/ra2m5qaQH/DwWilS39xc99RI58DKki84tS21YXbHDvzacuGgyEA1ZVNrLp5F2jm5yTxv
YxPNmogdMF+fp8sJWgcBW4G0Yo/YuOkLUZ/KE9n0T+Kay8wybU81CfgBU7LtpjcocBPAnohN9qsE
+T3Bk+WhuZYkKSGHZ3eWnSmwKy3jb6+ytOREfTkS/oB6NQ4BVbYpf4gZN0+y8HJqsAcBy6zm/PjG
8u7eK1KmVPZBeM8hE/XK6U1kHw9jH8nZO+fRSeTw1a3+NwhMTKHvPGI6ncrSPX45QL/SWoVy3dEL
JCa0/eerYwdqC6WulONcHlUDb3jgUjw8fvKu/uF+1FsFyFkHTMyK6fqFYtA3rVqqehlyyKDSIZoq
Hlzy5JdPgQQfFWWK7Q7JacqA2c9hfDsygJMxv8UuIFSlosstGtNU02+Thcz5p3beQw/QsrGK7wjP
XbBHk9aomSJy7pp6lojXOYtmSN6CpwFmw4T9qYHmjr7aq6awmwGx/NY0/7tlkF0p/kujzJr8XGu4
qWXyAtLaHJqgVCwoetRy1qZLgSHHiEvYlfk3GGiHJRT4AeucMUpbQFMmu2dvtQuMgmfXylS6u920
lyiAQyD8BuFx9LS8AynHST61GR1TdNzouxu/oiIqejc784+rDjMf9kQL/vSjcswaqNFOBUoRKOXc
ROz8H7k0piEXxtxKqUx/nAE+ZRP5eJSegdm4akgaAW/HpoJGeiGlJ+8P0kOdXILG3WBWj/Z5Nocm
qmldABxyLLvO6eS6+JIAsoLy1Mt6RHJMXBDX/v+jFNi/Gkn/snRqDQ0K0tfXVpJTa0RvFgt8alyC
o/4eAsMOQJ86miZ6oSAdM/txJyyXgzP/ubDbXfekvZfZNlMeEyIbdsYxqbp2P+N8epMm/97+xdbG
yc7/NAXbuZz32tSfbBIu0V7duRdBaj2jkVrekm3j6Wur0lhH0/kAfSizD6km26oeX9ET0zN221VU
E6MlExsWSyrbBmQMuKc1lPrQNTna2voC73M/OB++Jd65fm83wMccZbIN74R8weXLolRoXpf9DM9+
Pl+mU1dXCqt7aAJ8+doOUb2cunYtsaqbpB6s2pbaSzv49Y5aIDMV/BrZjBqZ58hGS2qBuJLYhaoQ
U4lXWYI9QQBU8NKkRv5+XZNQxaAXTd4vy1xZ2G9itbhq01zQiDlQ4aFdhIFxeLssdjd5eMrhVDat
oNEcaW/i7Q69dFAZAqBO5l4ciYTa2u7qjw9moukt1Sycbe9E/EP1xqDrFnE9UFT0+hMj2eDOudOQ
u/cKOWOdtNp3b3k1O5d3i23iP7lf4y6/RKznn8c8rCzxqb+fuDHIXin0vs2ZbAYrx/tjqcptfG/7
HpUUnSUtWD8GOMdfwc5J1GAZWdl1lS0mDq9cxClhicU3LDWiivFX8OIOYk3F+DfqD2WU+zu6iryu
lzlQ9OTKePzSbijs9OLVUQIiINiMkftSuvh1vh10gvKGM1JZGvrqlCUdcL5Hl4tsJ5XyPWT2tdLe
vTiGGWaYsGeAtRoDSTqcs4HwDH0RWGhI4Xut1bWxbQdgvv3ozctwUg8feeC2Ppop/LBrppNRAZNe
Tsi8Wh6ox/Vrt7f0w8/iB/U5kssrY5FP37EvvoQMa9raLMUZmAOi5nsRPSEylEr857ZtmnROiaet
Ga7lspRkwd1wIyraRumpAAM5Jh2DWi7n8olGTuEMYoJ+AV6+3XQ2e1AXVuNUtTEykND03DxJCHas
JCk1rLI+BmSZ5mT0eOk+RYIezvn4ayLlwCohwtrmD4b/KWCU3BmS2IgijpE+QBvbsFZmFksNavD9
adlrdRHFBwlagHFdtIwUBY3BrB74mCveaI77pWSSuShs7cPTqX2QQ83wSqGR0B3fAEIoBo1P7dRz
gW+5P+3D1vEyhkCUDSiE+m9QhpcR41hUT/gcGt1vXsgJiRrgqdGxbYiFMs/LT4ATv1VEmjV61wIc
IscuXtMYyy7Z/vBFRtCkGZZrxxLjbbSyd0QOWSdAsK/Jqa/Trw4LtP1JRmPze8YwqhjMV6536zcr
HPxjsc3yN798bFEQavQJg/IiVXVGO4qUtK0yz5JC6i8nRB9ZvHV13MNo0qRqfXj0sm31OH94T+Rf
DvvFNsZSqWKK0/NhGj04vFqzVS/g8p9kVJrNW0YrFvzSKBtX5SxZMHtAZuBzyB7flB5/a9/SA8VW
elJX7GSrwWJWOQ6uIeK7yKnPG/pMqQCUSNiXYWadjtbRiUvukzNgxmwquODYKW4iKNlvM8U+V/pG
Km9tPPwF90VQvS93csYevvw730TtUuouIn0Id12wutbJ2eb0wEMFHtwbRrLgTfhhR8q767gO32No
aEwHDkMtpSNAQaY1/ybYrsGhvPlNmBNHrjDdp46yDBOXB4Yr8IlWpvAs7P2QXChj60ojDlmtoA5m
Ydk0Qid0U1cp2xBAX6wPOr30s2rhEQGyYEAPpTXN7zuAn21dDD41Jfh866ijodc4apEA/KMyy7eO
0CsebQbn2HnBwEkkSMSfdaOIrz130fAymo+I+L9w+xJFCDp+zQu5XCnt/zltiTXosLUdRZXG8Rd3
FJAwQVXjs7pb2c5b//2OjlQCRK1PzkI+ZWHeN3A16fksNCpE1D/0SDRuQS0+j7+AmVnyr1qpV3rt
4kr2oRxIsO9LpYXm8wtemck1efriW4l6grKA0kwAkia87YLArRwcLtI9aR0HbCAUKH+I4lbjFabi
xz7LaWOx1vOnV2zTSpHrGjxsBjYIV9lztEDTEeSYW7o2b7+M+g7aTZO2kTBjZAQYH3WsJGLbAAO5
prl1G1z0/XETW4jy9LZKVdbAzB1Fcwi/VozRq6Pevq+nTEWDZH21h8prrCK1VEP/abLYi2G9wVBE
0BrFTZzBaograA25MBInvzESgd83Ig9NtlpbmSyCNrDubsxnO3WWg8qwoH+12QNz25PCZ2KoDgYP
ZZlhnnXGui/20ePTwNmWCAdyzMa24ENLla+DVZhP9+8IIq1v9CHdAOOL6Z+UK19HvMgE1zzi2MlJ
rYHjnVVvvSjhmmTvAjOd62AXzaDx16UMqOxYOgQ4evlsoxYmX+nBJvHjxcihyaOxjHsAtYTlc/lS
OolOggkTykY6kjFn4ZqlWS4nQF7R8b/+seik2UASouRG4UHagORyaBGwJL/S0G3T/jscCeM5sbS8
6VHz8CGyU3x009HUeyFQG0I5HJDE8uxZD19lPBrL1JH0wcoH6On4RFzYP1C2Ygl/pPVUPQYKMIS1
GKFBCcNGalyYNkMwgI3WzYSwyBoamH3qIfhu8unBGrtn8bM58rr5Qli1PUu9OmshHo85VljqJqXc
Z0PGWae0qPz+wfC8agOOcuKn6Dp/4rRYQceYWqtUuMXCbr2an7n6KyrDt0yZjq3bw3q5hBUKZSuK
SlOFz5pAw0iIJi6CFXjW6hKA9kDtcEBxzXSTFlkl6H2eriH/sJw5uaeX8TAKh4Ytf+DoSVI2kgqA
jc3iMcWLNLi2r4EAzrTx4offHOH32xWPguEDUj6sTpzSLi7LxSwzB1MIveDCyJeVrxo+11IK3HJd
ehy8/y5xc6gJqeCSPYKx3nUEZVYFXrb8/q+oJHHBNAp60ldZ8PXfZYFqtsCETItvtnqE92Cf5xjf
RMbLfVbaDTEsn6v3RuoG9/WaMjhBnjlqbKVMWkdzQtWCs6af6+Co4XWztdPtHgC7+Xjh5arEttc8
+GJmBEp9Z0CpclEb8rMTUYK2YtkSznB7zWdpXHv29zXh3BfCWEKqF/HHIgTT0J3bnujJd3iAnven
9F+I+CNUU8aGfWoi2EhtbYFpYe8gjavSKeDqdqiXMamWtslRA8LhmOMC97Bnzj3yAfzkTVHChodm
bAw8CmFTW4XETyfxGMf9AP2I5MoDOY3hwz5qgJa1c8YyCDcDNdGmqHFRcKf5BJ1KAV4IDUvDHfEh
izbXHnOAkF+Ha3uYWZ6skCjAvsJBIR9IXhOH2XYJaxKWqe66tbo/bz8muBH7HYdNau23KDMAOwQ8
c+72wzW6TcPOhgaiTNSG3q7bxJ+9X8ylG14lRc9uFAANNYkmGPIXITJHpeBixGkScO8QzfNgJvg4
5HRBs35Jnp6mK5yOfe2IOZQ6xfQGhWZGpRvd9OosJ5DWL7H/srOvJ2VwQ2EuqDeefC/g7rYZjuZS
ogDHlQ0PAI4tR6O/UftmEaweGHnazbZUih7rTlulcRoWtjHH8XxiRxjCLI7AvCwDVYdqGwvRE6EJ
2gvL2yT3+bu6qH3h8z/jLUNijAeurPawvVc2jSD9EkIOd4jy3TOt3F2a2+xJL9l/bbDm2romkl7A
G7+0sGQJe+8jI2goai/p23dTLJnV/k7c2g8NOOJ06KnDlQvBv1GSTQZw8eIOUQEQzIfU2UpDlmoO
3PlXGpdNcdm6DCLme1pJMNOP1+gyZPb7uUOZ86PrO66vHaYI07oBFs4m03JA3MGFVmXSrZVsJ7hD
GFeKIeUl/udMzHgbpAsz2Anh8RSP7ZZKhF3LiGy/2gRSGQotPkxdzMej0zlbIeGUfc2zTVIXKrs2
WKhfcDy5FsM+IZSWw20RXT4xwOQqfTkyI/AeZftG6odGr5666fd4kVVBo57mv8flJK2KjnJMCeoC
DisCUvXhq61SmRqOaTXOC0yel/83Vt6oNFXzZJf3RJ720o/Kwk7qpWeJVUddx1BACZLGBMLuLJej
1F23zRNntXuZnRMH8FV/QxUVYT7qHAB3zChS3QrKi62J735xV3YQcAgw85kRJP9ptWGo2SfnFyxZ
3vCNQyvgct1LPTTfQ12Fe09jyCa+jkSwuKk7W8EDqz3YofUgTWtuVpKPc3mZ8o2uPtzdt098RqpA
1GhLhGFeX2JnTJK3d1ApHIrtIMIe8dM5qllj1ZgibJWZODeqoXyc8CJfOZfhlPwOr1gmmxvcMgGV
pxeyIaWezjSDjvPtOe9L+F46dGoMr3BqPkNZlsXqaZbrstS4aiUQQuzITw//DHA2wZoR0c/3BH3D
vSUSVTnRkBPn08CmRpkN3jG2QvzwDsrVcu9lUNql6kLSyP5oaK4wPuMqU5mWOIcz9M/uuF4G8z9E
HID03fplix64xlsPgkXiyepsAn1bOkZ6DjaGf7TdoK93lujf8lHUXhxXLduH7qsC2DsB4DWbZ+15
BxCWmgIAaXNVkBNFB+w1CKd5Pzl7CFN1Xw/gdZQtfwPxLm4lDgR9OnGYKQFbU7J5iNDa3yMNgYtI
YvWyUp++AcYGXkywNeknhQSNs243+bNnqiFJHO2LrQ3pcCSHckL1dFYjWEcBQi/YlJGL2cDA1i/3
EsJh4hjThwhmAwUg1V741mEcPBRFrzWHi7DSdJcNXjTT5/UZmNCUGrCMujaaNe0pQ6CSGzyExZwZ
D+v8CN+LNzrjoSjtOCVsJ/fKcuuR2VFF6QuTus3gibZ95Zh5NuvZei5OElFgQ0r4mNvYXhbyiXHZ
5u92D7hY1g5fxFAMYKkjcCnMzmjVkViHLyCx1tQsvTbvnU2cMstSFo+tzyj9P+aUcTBqdzJlRwLa
m471vog+EkSBgNN34+PnsTDD7AC9cvNwvUtk7KCjA1ZzwFzkbf/IPgX31BMOIIPIrN1lxtK15ZH+
u4BHheggB0+8T/7hvfkkM+gBIg5xUpRL4VAUBGZiaLVPHMCnXhmd2WDMG+/UyHy+kCiOZFjGB0T7
N9SjzXt5UDxflOm9+5UKtkj+41duotnuZAleGbVd6D0XNm85rK6/1sEezJPErZUpuSBTJcx0gESF
nyFato5A3H2+gfKZQ8oLObN9Kviv+U6C+W8M3o/vn90SpVqjoXMZPeWbQXJ5Ylj00N9T0MI6cvr/
BQZi8mbDTat64vd9oYvPAdC17XlZPd986O7/nlrLGBKpB7iREy2mZZkPXEoOVjTixznOZ/hwyXCQ
eyv4vKm/kySV35d80eyx92URgvG1dKkFtXPyq0HFqfdpR1ghKIwxJMWpI1wvN1aUs5WHIsv0wrxz
ZheomTtx7uSNIQCwQ1LTmdoCIB/tEdvsjh9gYBUK1O9CvWSadzC8AvDrlIya7F89dGALhn7REpqv
CKYoXrIJgTFiHhnhv2AXCXQCvrQdbO607gtJLg7JCEOMv0A1FkStbOpM2hcWOyB+GYg1/xZMvYaQ
pKTu+IvNihemjZyqJFTrztfTOWl/vVOjpn/s0ZxQfxyFCIm0T8i16wI6im0DwUlG6tCmH/vG2r+C
5NQHMN+jGRy3Hw6kGY0XJNf5yoGxWxuajNSqybM7aZuK4P69WaJvJCO3UsgdvUg3+tUdOomRld+W
rVobQDS+iYLSMf7SMewd/4h4KvgUVy2/Wj0AS8zX1FCNRJTyFx02bJbvYUd9B9aIEsj2SrHTz3Kj
Tb3KqCO5sQoBSJyYlx9R3M1QyQdsbn6um2SwZfJ8xpqgGIb3PD2XT/V6V7z95k0GK8cH1aolmImx
73DUaH53/HycgweEcnwkV6WH7LsySdeUYcJYwh6Z3tpDivCF6Ws19XGJ09B2scZ80xIA+/7sF7YT
Pu6oijuznfCh2njOp7cZsjjiVGkPV2NNteRAJAz9HoW4CNBjFx0zxol3+0WPgMclICofQTyo36Gg
okr6uk48+R2lhkedMMpF4+kAndlQajBBJbSJE/kJseQUUuj4o0KrDQmbPlFi8UQfetPiJgT5Oo6L
fsEeBFEYipFGZCoG5dj3+wxGgbn1ffQ8z6J+VGJMruWJ1tJAlfCUOXrdQRIGmGVIBGMEfQY2l5MK
11mrHWsaVRegv4ms677Uw3MzAlc3iD6Nl7LV5r3sKbSl7DfCqd65j2VSMhqmKmp3G4b9qSIAT1xw
dJS7e4u1PJlgMq6sxZIeziru0KDqASYddOywkD0poh48Wy5LnS325sMpC7YpxcQN5tFgRTrQ0khN
oMF8RhpIUfXd2ehHJdZ0U5LkUxG3KsyQr7IBYPm5AEtyG/TF/T6xVAb8F47scq2IAl0ggD/tEYI/
BVufTXWzRlXs0nA9gipDgsOIURaVWBMzibuzGEcTByg1udCgyqj1SsS3OX7JDHcHpqKpEHCEq7uS
wS/iht7S5C8eSA/3Hc68EpEwarAJ0b9CUG5Ndl0EUi0WL6ERJ2FeqgZlQIwMLKcunMFaUwDLjOJm
oAi4GFTSnXbGJMbLlLvj3KmTvlzorQsuJFNlMpZCei/UfmRlNe+hwx8aymU0rZciK7rpRUJixFGx
jCNAZS2ot92T6l17pBk4yAHkNyPyB2quVnTJf/a2Ll4m/zK2gntTD//y9/XBwldemxw2/owaQHz9
Xdlbb2GnheQWmGKgIeedvNGzrT1IIVhi6QHAzNxVJP5Y+/IJzjQRSMDvs6LZD3UczOvQ6ZrqgNmO
aLGiG5IdafiJ3PWhv6LhX/iFe/RL62n4b4NS7XKabkMPPIJevKEXz1FKPVhpQX1wpySblZ34bvLf
flSh/na4PXZg0QEDXGK64aqk0l96ZgXKlTG8QYTmH4DMQ0w/yc6XIL8bBEWp0CKQDyYHgB/H2yWR
QyeeOhMqZfLNP/Pp2nOSgrCzzaq+6XoprmXkkHYiSHXYg0X3wdV0KpL813y9ahDr44SFE4ueg41b
jRGONGkhAbt6redtirJkeed4Uz3eLpiDCFauc6NS46weZ6fKO76Bp9pPK4yMz231fd74D08IqybE
RlFem1/Fp22NF03BZSRFrb3lUkpVf1/jDQgMkmVygcb7aEACItCDEyY7AV0Q0LP6lQwVEv8ZzBQ9
0EPKck/uK81W3YztKhKYbwd2Ep6gSlBlv03RGKDaCCn6PJUeZXlfbvHpBRSJ4Uhvx4QNMQdcwdnt
ZkkoKKgdGs4T4vXRPDELX/4UEc1OgdWebKGp9WOeboaSqVNdyBZcYCtbtz0OFxS4dXOHYveFkj9j
TMxbBWTjhlRuxZAHKdcdKbTnDrB25j+/WFk7GURZWvbu5bSldx8pl2h8V64ZQhA/mT28CzDJocZQ
UO8WMxVA5oEr5P3m1YHTZfN7fYqdh5l6pbfNbe9tKC9AhGttZbPzzHQA3Owhlju9bgr4aBkXDJls
ZpbqvzbJXmBo1WJHO4zHQ7/N3S7SwSuXjLEKL0A+qnimDunoAt2x5XuJ1XVCmXFc/SXQkfV+sj7N
V5yu1x7joLHd6hSa0vAIpZvxGZtc/m4cdAk/Tpb/KnuAndYecTUCnAZOAuPjYIq5jYU4DzLaNPjV
OzYA+ApISZMjxu9kCKcj/AJq2Q5JRHnS+/vyuUxgOD0dnZHg35lEhV2c+tj3HCy8kzzw9eU9IFh7
8argO7PhmHBOtQzKvt2xembNNmcL5aBEVREftwWmYd48TUeYDLp/ioWZ9ib3qPrHXIaTRSdGmJ0M
RgPXtnUJnwyUlk/D2EMdfD1yeA8Dad5fIABfRG4NenwLhung++C5rXCA5JiD5xIXg6V9cQXfOmKU
pq7SfAZtQV9pKXaOCChCglVOGXoDZz1gXfpKdYa7XZKlhMruR9nNfLHTxI2QusvHPJLup0dFL7wv
OLBZ1lbHmzThR7bm5KYpuyBSV4lrfpqfkpKJirXVm162olP27yxlWs2rdr21DBWsRzrCNf3zWL8E
kAP9munraa5ZmgLQTWoPZv0oDnIUHIKdhNj4Ki3WWGUVUXGymdjdcX/9cT6CdxdpqOtnxE5eOzGZ
ca/4cK+2fmnrj2lqtjxpt8BZ019mc0rgvECXyVpKgSYnBTPGemVLhussC6LsYa36lS0Qx5wndW77
lN9EgbWbFg/acbtcvgN0wrb6MS9fe6NDHtlfgjGtXYEIhSHl3oJ9WUAZmyZoSiFsKjROgx/CSUFM
BfDYeph4007lar9NGUK84JBHN1lmyxjgPSg6iZzI3Tn01CggN1eYTCxKYSHPT1NZ7HY6eNKtvDrt
XnrIN2PNNbYR8+rcaMTrXVnCZGCx/F0CbRiNVRBl93olEcWWMOSdWTG+E7IOB6WPBddJ42dCHl9O
oEzLoyi4RkCZZzbU3PGaxe7hC850H8rIHmJ8IJ4aJVtrg2nEu6rnbwvqfhv8SyzKfEhdBgKl+ibb
IsqpfX5KDbtkGmVbhNWtN6pbcTRBIW5bMW0qto9L2OPHQ42JI3RjDKSNYFToxa7lRL1WUxs6elM0
AL1ymvzIa2VyRiRppCPudee6daG43M5Wk48NDs6upj6QrnAXI7/rCfbhAB1hWm5CsiDuo/0PG0/D
kuJ1ug6i2eeZ2Jt5sbunC9SCjAblMnYY2jtpEA4Oo4aAvGIgMlpmweii4zEfgqNFQt6lZMWR9kcx
I6cvzh5/Nf5dRtLPh009I2lQ5xFomiDb2soW6a4Vyq5nMp+4VHbCTIBt3D8cpnDUtsYqXQ8Ejxrd
aXcnN329vxdrDgoDbfE5JPMIsieYwTTIJ5F9N0/m/sCBC14Ows+/vEZU74500LIl9Irz4rpWReAN
inGOFH98Z5p4Yk1K4JtNuJKdBirxqPUom3UKSL7wyAN2xyS3oKyMkdPN6be8uIyo08s4XnQxVpbL
INR76KPOHsmL25A7ad2Be2EUz+F/izRU4ID4STgj4Wgf2uMENL4tikba6MQZYZrVoEqOPvZUJIT/
NmP0J0OvNKVDYs1mBUhdWrZXe9c6Q6VqRUXN8B0Q7sGwRnDD6ML/JLNm95sZ4hTCjiBdp5myFySJ
LhqBCxBsZqiiJ1t8kP+UmYZkLPA5qeMd/NmwB0uz4m090wuSCE7Hz6NKO1kFLcnPD6c2O53wObDb
yMxNjIhvN0+hx0xVNtIEpNBw4XOBpP8l3VtDkrkUVKRRQYSTZXqxzWfWCr8/tS14hKfurB8RbplT
X6Be2baGuyH36RUXE9wtRmsG5lLhHbbvW1xPZYuEZGvHRhBkdlBWSldp0BjKmOtlk7aLreYCzrzK
t3CutxWqupFQCKxoZkKv+3FvXbx2FxUUH3NJ4pWsfj08E5MaxV5jFG4JDz1w9gcFL5LHdISGWdmi
Bs/UllrJoNbISlH+OfKdlLLta3Xr/iTnK9OZ0iVKCQzY16tbL5EhqEW+USh6WTruQCBGRDbcbHgH
AGUYm7/yV+btiQzo3kVUHBnAT1tFOGbNFgrwaTNNoZouZWXOzbU0zqO+KzAhjBB8DR87jRG4oSpI
wfrRrpW9Vm1Kza6etMkgRtO2z2VlpTLQS65mYHzaDmw+Rc2Xd+prscj6fMP2CUd3jtOhTHl/T4br
xxwCGp3yyHXrmuk2KF/EaDZra2aBY+U8cd7NrWmzCuRn/QDr0+qgRTnL97dllXFlfl+WT27djMGZ
pEzOIDDPqyJxnKX5Gqw7U9qhade+CTYcTuedPVF2jxU4I/XbbqY5AjNpLiYzMYHDseYHy44zkLQH
8FJ07jsJaZNwWckBxSFakrNTfmRRy/JtgtrL0bc+qqNF3EysjlKBhPPfwRedtC9pFeaasIPVRoOS
778Q+xHJZjzdkq7AMHvoY3F9JTS0qQfQQ0+3o8jeK1JngNAkvpeDud2hKYBxQUsi7KyUSbnsGYKz
v5F/PE5k8x28n3dgjuco/XSbq4JFETgjH5LOCUHHv1DtXKQpLGuf1x51cFQMx6qjUha0r+1zJFra
rtMqeAskmmTUPsicbhJYentj5wWQUrml2GEYc+Qk9pQyQ4fUa5A1hZfl1LoaLn1MfYL17MkW0cci
sZ/IlMf1kjr5aYc6dNZNbSobLmk0xbZ8SjbCbaXs8aDS6CqH3o/wGAvpXAyQBvswXNJi/RVczTyY
dVgDjmB/8VOqA4+z6UHstd78GtvyJelt653gQI7JL3q1ezoQGh7zyPl/fkdt/lJtj/koonXSoVQS
tL+UARrcQuTqafIRy3aHTM7pNWrVb8gXeU5+20kvKSD6FT1EKaZOuXRPH5iyDFFjU4REj+eBdWw8
XEyt1ZAjSbgEaKLxSe4l9xqw9l7FNRCkDYzhipfIt15Y5Od8gbOT/ylfbxcReGj+MxkyI8BfGuoA
plSKaxmUJnVGpjieGs0RlLofb2NfhQr5eyywwCyqEwR4vQYHRjkm6rxfrrnXmM0Chi70Z7In1HW3
h7DZiKl7Jd54J9BUxYtc4/ejsAwtVwRpSdyJ9PiQavKzzFqZ9DsJTUn8h/ULWyLgAkLoLTJV7nx0
ZjWWXWjxpujWw9+Ee7QSTseW9yOpDWmSSznethM6H6GqwZmRO73xGXzWAewh80RV7yxjkDm5nGvt
jB4ERJkoxCE2S6xqmqNloEE+BTn+9MEC0UQTgBcn5jUxoWtLV3ZDE2y+4820nIXz2BzLyv53YW5G
1o3EBgOtFnt4EnkDz9DarzXcwFB5ZwDx3jrbUxcAy6MECxoNznoS+/PrCuCmEUX85IqglYP4dZSC
3kW4kimYAeEjw+a0Fnlz7ylfYJVVJIUu6elwrpskCIP02GpWpsMNtCWMi/oMQYW7G1jSsPRryaDV
Ra1sAFnnzrSdcNccfVCffrzntdxb5UV8PQ8zT443gzLPzZE0o5NNnzSKsC6ndlx42YzX2eHMXICA
a+ea7Lh5FHEAZ/If4MjmLmRnxub4/RjARfXMXpYAGs0OUoC3d8KNno1xe7ajCf9545rEiTShth9u
svonaVE8ZyjIN4Y8A/CmfEjGxdhyY0Nw0hCj0LEW12p1iUc9xSwrPDwO54dLC2QyxV59qmI7rAfe
jtoWDF8xbJOp0iX00NJQkoGx9zr0XgqUdVFQsM4Vyg+i0WGVuz5zUvs4Op+ToE54O6ewE53rouLb
NpcU4ilOQiSR2XrAX1kgIPecIdPKiNQcqe1T7kjVIy7bS4szNCoi8zzjIAvDNDGNljf3RP0+biM3
TlKS7fm6IKH0FpWrFrgf7r12thXTKwxNuw1Ed9xvv15MdvTa/ad5q9ZUuJjAR/8fMLMaUENKTOHX
+0aUFCQH7pFD0OaeclwglI1R1lGvDN7/DqO0bI96psXquz1E4RLAuTzbV9VhVCeLctc7vwmLBhI5
e/r8TWe/V90iXgfgluCgidsF0ZMFJ4ixY2rxOB3bErelhS3Y5t5FagpI/v3Vdh9PCjZsmN1JuIb3
dZWP4s/T1ZBJYqPz2CPARrvcWMSRpO8gTM2Xke7TL/+evY/e1/wYQMYGBr2+BduO4DpjyH0YgHHs
naRoZimZbgvoWk8CK00gFJUZLw48qJhyq6ifX5FVUA2aX1nTwUVoGMY9N9A3cOqtrLS2ytFESvhm
iR7WRtXng/c5m6NwPg+F2+2K0qmD0Xt1Tx9gVYtCudvdgES5wVCdzY0YMWhz8cmlZ3BLzkbXnJ2H
t3oDYT9TvkUTCk7z78qmoDQIZojO+Ak1xsDSXfT7Yd/SehRmu9b3rqhPknR97XARNl725aZYhzJQ
BlsJ1EdS9OBuyqr2M/a2daQRs6YUg0EcH2HYWlfHpY8ysdtFnLOfVu5kXSJek3Sb3CBG1/4DHYm+
/27Wd1qhGHPMfSN9JkWfjtkuODQ4C4IFfkJ9eurNbDrFdGdsgrE6gJ2CyAYXhv1pwCuWKlucO0iO
hxrnquCVENOCw1OHXx9SJsHVfiFiIMEOzSKpeZKQVWqqmfyPULRBuIWtp695Qr1KX5PJChLcKvBh
S7kqTPxBvYuDHNQvx1AO/vg58zl5WKg7jiOrM4Cjo8DXZR6jo2bdAvhGvzkFteYFmA2odO8xChj3
L2S39lQPwHpOQmnNUmN2i+WQZPB7bzC99naLpqYaHOouV1QH4BnYSIdd2efYU6ZgG7nYcsCY1Olo
3PfpKviIvvCDTSvoVq5pRNVubigBdShE/0c331pEkco8uso4XPE9YMvEScRurVpc/dUC+1l2Z7MG
jPh8d9lMsndpcxQqPIWi++q7QsrGWa+pYm/E4RVtv8a5bGbyCG6pCiDx5FxACyFVeP4P1In5+7ro
eFq+gRRsBvqkbqIenIoRL+O6LdjWxzhpEg8CpNwNuhfBl/IDanP0Sd38NPvQlFR3XVNaSwKHeLgc
h68cvP1Sv+vhbS4i6MVA9+9aR1Udxb94aHF2dI0TGL//8Ma1CAE12VEEJ+zdcOlsTeaWqchE1s7h
8h9c5Nn6WnDOtTnTW9+S/D2BAapWxVxTh6lWBxW8pQhBiWSMzRYIgXZzAAYYk0W66TPwxk/+d9lr
q2DAUuMTpXrsEOd62BdBXlRU2Imj9Cw4nigx+fX1eBXjmESelFffNsiRP48eAaGqJdCqql4pK2Y7
ri3+B3QsQ/DdL2Vq/DVBkJNLEoysexUTVc4p2yiltpM7Tc4Bud7MAGoHixHsuDaC864O2QjrJTMF
iiXe8ysDFg4JrVYFffUN63eoP3tYHNUrPDkRXKPsQ2RNAWdvHrG3u5SbBCnnK3RBZtMqO45VNvs6
LiFl/qDyVt5AzylRs1Df9eLTUV7GbUnSXkmC0YSC65IHdiPiRk5goaVkIgo/a/piUd8IHur/eT+Z
frclTVLYwCcn579wHTIDjK3QQfMpJQvtkibQGhko7Qm9L3ijEjhn2iln1qkeAN53CVgjMbOkZsC5
XUFfhXeOuyGJZorl1Jv/NQnIIeQi2zkYWDXRgRs/QLo/io9+yfaZBXTsIgHQl7ATiV5ElDgrNT99
hNCe7CTF02UWuHC95g5T/ZsIWhW+FEpiezAk/UrumGW+wY1hC5MGrbiN21/OnvROFJcZFGPV8nUl
dyShScQyojPo17qA1Wz0lV8rGSwhDNA7TqFRgNFR9AdKeVs38THmSdeC+UPnAJVwgow2DrHQ3mTH
W6ESQt9Vyvt0BF6EGASLkJQsViF6S6p1VeXmE3n51nuRoo7+y2JxN27eWK8ZRU/m7oK5fLEymEul
nrAcPn9737F4V606Yu1UECsVslSBZi6+HNYocZH2aToaJAYmcVoQb5ycmr1UuvLjGdjhdowGbe25
8KgF9Tu41tdOPOv5W3Q6j8IhMTBWUrl4OeA4VEc4qgcnYn1ZzrVXykNgrFsgyRhDQ25agC3G4p98
Ece/1eTe1m1xJYPR1Zue10SujnL3yI96Ss7agK6vaO38VLsC9baZ2cIm5reUsTKLP5H9zgcyrECu
ORQVFwQyb45KmiJjIutqhyWH7FqpzbSAvS+JOgat34KtAZK0NiGS6fxN12aHZEbCqYap3p1ySr5z
90Ak6gSKZrs6nbdgskZb6ziQPoyajtW+OqTAU834BrC0uvmJ6J1q68swxBMvXvT41zbW3f+Ovdcb
q1ZsrvNpCRHOzPVBv+vhIUfy2/3+4qfY/PrjvYJ3cPjiuphLvFJpR2tksR1vf8XbauTJbLJ6pssj
BezFMm1zcbndswkQLtVRYvEtspurFBIwsr8tSrWBt+V/jz7zOqifXIsqDB4h2nmMZbVLERZCzmxK
ejlD9MTD24FfQ8Swgseu83vyFO/pCMAoWxwqJFgTqvp2YN6iUKHMJD/xQILsRtsgyFfOmd0G1EsN
Fr5sXSk062U+PcPYnVtq08iHIXtodYU/UK9TQ5cFwPmpZp8X5ZAiw7R3b4Eb0gpdVrfB6B/tNPL+
XeA1NU0NmUb4Opskckb+Tzj2G7xosW6CDSOHRMtUDMo+IAco+LMP3mXSRe1A+3yHhsXva6inMKjh
vPSCia8+4ymJLftT00R+RZYNHBk5kPjoN9JAy8FGzyyQQuB943IYxTkqA4bNTJPPyLn2Bjglni+R
gBGgrzHGZ+DAR1744qVeB/WpI5oPTh53wN+IEOoVRWIt037Xe4d/2NojxlecSN/NlOiU9OGnXZ9l
7CWy+X37maPk0Iuz/UXi2V4tOm6FnX2Kfu+4DaEWLZsOAINZB3wyL41dJ7kvrR3TM1wPtBm4soJq
G1EVobKyEWO6gl7dVX8EZBR3jaY26UhYX1dmYFHsIYvrrS8KdaJLVuk6a4AhQCvyzMqvTkDNM1x3
1ra2ZxjSx//n4igpYZvgQ/rXologf7rouz/OTO3PPSZCyDtntRoZ5D/ZYTROZG6bBziNm1QfVHO+
uIIWiKj4rYzhOu/M/VjZm/VzDFfpEnArB4mfIqxa1YtvSWJAh/V7Mwpr5I01vNBhucZVOrWUEts3
P9TVKC8+lOAuLBw1AbmkEKZLDqkGwneU4/Iniil5pr6BPXpn3z/DYlCAjTsyId8kN/7wixXMvyOt
FRgyhjHu8xXowXwcHsE3oM/tjqmMFu1OHHzxQZhJB6/V7874wH/GUo7/gEe1/8IORV5T4u45OQC4
SRw2uFFhnNszbJRLCymso7VlbIFS9HmOKMhzilCoDDJ0E1yYj5KZmgJXWLF7+8Xc84fqX8Bws6JZ
ZhDA5HNOZ7l3DxqPFUcRfdXP1o4SX7P0n3Hq7H7NkiKyC5Eadgd5MF5NKn87xwIzQkZyJpDgcovw
1OgEDPDkqnYGMyiHWPJ1/qL2dn+TpjVwPNN2e6BiV9oYhzHPjX/yHGuUDympC0Jiq5FINLWEbskd
9iUh9MtPGal9GEUOQaGfA1TvWeNGs/SFoBC7QJF/0cyff7r/+IeLc0TNhQZwbmyfbHFYQntgmWZG
AwDzJcW6JvLpehWggY3PSIJ2cVZ4YHLG5GCY7ybESbig5T4t1Ujt9fS3mG/vqoIL/ZDYx5A+8B04
U02DC/hDHB2GE9cGCSE4XP+cCH5gjvFoO7aq4E6vSHbvh652Dg/ziEWh3FUiYCTmlk63Ze3fuvVJ
qfrLi2ZfKAL5HOF5IhKX+WTthz942d3G76JRLXvEIoaOAzQc1NYBzNXyVukjHyc1bTnHdVHZni4M
TRRXbg56O/a9VxfMYiLZBV7TuL+S7cXmPq7phoy0a7w5XgAEwbVWWB588w3gUsvNzc5/N6Y5nO/p
FR/RD27El8+JRl2FtQ+MArPI+AJmqjVPc57Xq/kosya8/EXDdd8MP6jEvxKQ5u5JUuzvWJBFpUlf
m8IY6CXmgmoIg65ujO2O0FWRIIuI3chN7QcmOEPf+mvmUyastMVSas6TY5wSFP6PHqxfRIaDxwWl
yZkXaTmZEPUrvCTDyWMGO16iLldou4jVmQfJ9+O2c+sd/WHplthuhUjxniCs5NRTebVu38xAxcFC
XrNUG8CtFH57M/Sk8l+gKORu7or2Az27sQJviduzeZ3NVl80PS/cfYksh8vNT9t6xzJqClQn714P
IdiUWbAfMOXSjFnqSSG6fJc0nhgTPlxMISxAlvA8w8Re8+H99B0uk8tHs4xmiaK0yM/Z6UTxMAfg
htNhZi5bofom8rObir8npBP0o5rLHYnZK4ivT/oFwiV3gpx1KAMPxIotdSu0SXdUwJrFCx667Bu4
USAZsO4j7EqA5a3VXpBX/bvf+HAD6YulTba4q9F8ZKI9zHNJQtVGph5cfPYVYNBpSJ1j4OlkY3tn
JC63FNuOrFZi1UUFdYZQ6iFDaRhcbv3ti/Wfl4t+WHwaWHFBUEd1JnkKZ7XSNM5FVapTiFgGTFwV
tEysDY8WMDaT3e4V9goInCF60sbTyObUXd/FnkB2SeDfrhBbamhei6phjzpsQgzcoSdYZFAbJIuy
7qRqbSO17h5iXva2g9AgQfu4TTU0YLLHeHYix7D82ZiG+CKz2kok4Yz8mGt/IhtHbmdb2W/KNHdC
eddVi7NQZQ+E53F1q2HjLlJp0GNUiFA28PpRKCbqy49xuwM0suxMAxf14zQbyH17+KBX68ppwABs
mJDjOOs3RuSr3OAR0X+S1qFM8zK94IrStBSWoEbAWgAPYi0RZbVUnLWY9vIjupIElZdiVXE1z2Gx
RpAVkfw7urBaBN1bw5qRIcO7KjqZcgk5X8F3o5TVzvkPnln7KtaRkpGdJuENTWiXfkB0tSvYLFX0
9iFaBFFC3X/DWyYUdaKNbjccPVpS5VNdLhQJ5eI0yh7/fHmVbbcEXuaIyZf/PLUwWhynue4nA5vx
DrdyeyuzN/6nWnMwJhiKuOBNbkEPSTcScVHhj3SrHAx1K1uhgVE4xLnqxUZEsVan+3w+P4tsd8Z6
uiRRfZxKZ2dmodh1lLqtRskoDCbhmagd719GUtalV0+rCLgINvQHrwJcT1oZjevDyaLs/VRBehQP
h2G5NqNKDWMpyBIvdSfE84TOqx+0S8fRBOJtw7dE5ExlEyVLZYY86D/tOrA7+QVROw2mszoQ5zlv
V3hVNSKZyStZNCAFPDZ+F0gUEgNLIV+QxpxzMy9Vql5afC2sxLENhqg/28lfyEvhjhEfuKrjxL5F
9gfjH5AFgqbcBfNAENc+62JikrjGpZ5eZSmGFhxzuduKrky5d4SGjPa2nsJxrctftryoW2faU5AX
LvTBTH82otSyrbSrgUdPYi0wiqCCGH8yEXWkIKAWeeR83q6F5cqzLLHjf2X8JpoCK6qT9saCHVlg
u5PjwRV8dUXGYHa7hTU1kN/eiWvY9ZyD7D5uRGOc+cdNmRd6JVGQ8b9jswX1d6O7f+AFpjlWL6j7
clcR8uOvWPgxZsWCULvN4rvFG18SnSFfKyB+gxtIiPQoN57zYr3/pAz0WpcPygfXhibpbKTrmdix
adU+IJnpeIi1thwEMIoqgqKN31WGVV7dMP0Xeh1zyDuEPqC7goJgqxKw9hcFQbud3HYNlw9k75BB
2mB+L8ePQtrXdpVOcm3Hh90VnUY469mzywWSn04LiDzR4fneCHDpocLoV65bCHDysIq5TQvcTUst
IQRw0ne0EBUi6oqv4NWGeozBKjFsfZNs9UwxOksiyyLzADAzidu76tuWro00vTFO4gDDEMQ6L/12
q8ES7A21iExYAtgxBILruTcW9f6Hi9Szv7gj78fNMFnL6xjZRShGQAU2pfkkQ6ImkCmKgo8z2CEu
O9RswJXN4KJRgJ12WYcOoXUcBti4N+ov7JNPO/oUohHn/0iGgpttQW/5YtSpT+h0oGVFFcXz9e8o
ltHhyPkDeqkr4WHAto7JVLtvF8Yyogcef74zGhH3qjDZxB5nwaBi/uFVaQoieU0h9preWQMTx+8h
F/77Gq+oLfK6q1SmmWFI1OYFA7v7MlqYXzyPn1QXdusMMyKXO01gXgz0Ok+LqcTOCcI+2X/NJIfT
8Rmuc46XHu4ozwcsr99ZcZts6fiEoAO28uJZMeNRFED034uDcg8oBTd6nD7QcKceBypNoxPf68KP
CD9sihv4q+HOjxVaFCTy4ZQu9e1Hsjp4y/13K8RdzMYMsRvxOmKKj/soFIexYNklxvYTW875C1kV
8JAN9hRQsd35zOiJSElqny0gszhwwT2oZL5Z1sL8mMHwwCeQJhFxdVILQbOKMH4sAWtkQ6GXgu66
zuavkx15RnGUU7w+7RHKh8f/RObAKHHa1fyXxQk0R+xDv2h+tY29Q4HuQFmf8h7YcRiCgVzNLydh
11SwrlmO4OA5X3Jt+WN0qoi2h7gXGFzJCFK0d8lVPT5bxLmEVe8ZEzkppEkznowu6cb8eQUnTG6e
148q1ytJ6iA+TP7obPPzlE4T5C28dvchaclRuc46cKmxmo5qu7QIbDNkiOLuUiXSZQkW2v+J4XaT
CPl+y8aS5JCQgzF32c+Mj/iAdDOjhULaxOGDFnb9RUJ2Hze9hORl4V9eynLvkZT3Vvfpj1SHRN7a
iehI4nQbE91/GL0M1g7UTFWJ9dWt09K5tyvyFBWB2VaVZOOKbIfyIbIqLYE2Ba9vCzrjGqIsgThF
jaVYZ1+YKev5N/1OPXoxK0d73WQk3UjntKwSrmrsBQkqvDGXVXn9+keJzN+UTgtgqYJWD1CdGO0z
qlo5zs7heuBm0Ka1Gsp8+D4pe98W2bicN15zG/dbh6bUOP3eeS08ps1MKBGow6kGH0bSZnntjkfa
BLH/pt4mNzXEZUpSKZ3x+X85fQNKAyrEGY7zlm/3dCEFY3oskTkxB0aD1mMizy4gp/oLWvyRT8F1
p6S7ZrO4GYgzjttM9fgYI+QIP5oCsY9Q8c7x0FTwGAqar3cu/drsmxfmkWQN0CyKiYU2LzBhzBZz
PdY5ADaeSo9uThwlvWwOZdKutl3dp1kL+rA9PFLNALDPrx4BfpPvsvn7+8dNuVtMBjelZWozBa7X
u9AM+20cXWiiCn+ShbPv39rCOHxNgm09MsBQdjUyUvvNVUYuH9Vw98ozdfKcqiSyJnH8tD9MBZUz
hBDJdmYtD3DLYMlfQaKasU4oc0dSIngpSx8/KKeLazhU23piKji1YEKi9Ru+Yv4XSsCHtmONmHAw
UiKZnGzrjVxf748vAjIAkN+5Ios/NgZgbdjyKreeL8vKbR9b+UAyTbp+W8AAJWByZ3zs94UbYB+y
DswnTBAMPMHno3bRYH+ty4WpcsiCta28UwT5cHdKA5MA1GB+yTTw8w9s88du35Gzp7gLBZjg8pwv
HtNOmX43bG2yIY/MSfENhvp3iW1hdZKSoQp7ySTQFUGtt39iqQyzPC4fn0CCVw0NiSPoirEAx9Al
yoUpba+zd8dL0QEWCvxcrnQhpCSE0dxJ2Z/ozhxRk/7A0Bi4JZ+3kAId5ty3+B0m3++SATEA6+zM
sk78EOQqeyvIs2hRF77DUvnTw1RLXXAJ79eP9Cmmvu4UzJnH5r03su9t3mBq1f9LvAL9lCdwxQTO
wT6N1vtPSR1jf9nTDUsYGBrOruCU7Iy64lT+w/DAo6WmyKW7st0QZWHfJ4dZPYoDQ0TemPVjH54+
VRNCTDTsJDjhhKryxHi71A8Pp6pxRvPtiNcOS1kWKcM6sBOUooWcQ+5DHhmChOZfU4dqlHzhI+hT
LoBmi/qLKU4DjKD8Uxi0GHb2tI5mwBGeen+9OOJTnqaASDlkE2abAEKPlrXeUgMHiBIaRe7h/VFr
f4xhInf0nfA75u/bbxjbL0y5GFO+koDuLBddi5VNPIyo4Wst0QUH1hrkskoTbmVUTnQ5GrdbNxtl
vqrqEPel+0+arEieMIG4Xk9dIrt74iGllyVLf/g9VSME5L+Bl2VPFk2zx7LQRZWv2HwIbqCNfr8/
U56pbLri/ZmhkL/1NZuzDEIpQerpLrMj8th4IyY9LwdTQ08dSKLOc9HFkrAIRuKC9J7cVBFtC9mD
D8PoA56K45AF8XdKRTvk+XA/58wS7sgQt+3PAKKs6/UEgHWEgGD0JY6kE1i0Kx8LHOMwKFe6MwU2
CMFO8O0L5y6aHaragYL62PEU425kq7bX2+RBroUV0DSKZ/xkShBqLsXOrQGv5x3iQqEoWLvWrKGU
w1I6VvCiF8+FLslkPkvGLqktkx2yHUO7p6yvBV2TUM1/WxzozU9kE9yZaHHZRbju9k2pNQNFzr/7
1wzP33k67pic9VT5Tkn31L4e+Nxx4hvGR2TVY//fW5019VaF+VeEkf44wdMBhKyENj+RaQE7a402
0fCHl2/fzql0SwBkWf3cs7Sm/grLRXH6vHdFLYs3RSaZpuZO+ty8sKdMJbKChV+zWbKrNGtw+RPY
OY7jbiIf3Pks7yGEsj6kIXkCy2KSys3jBXrzHQQWmXo+wbTX1jbH3hjOcLWAXwwjQfW8G/s+jDvt
AsxUKYeOP7w7bhZ3j3ytT4UCr9mQ/1uG1OEhD3wlWoTJSD1Q+W7On3S3mc4rrhtW6YqOjfi+4BeK
DlhbLQv8TU3xyvpr71mfSlwvYJOoYyfHex8mx1sHvcHva+wUCd1BUGdpRQBqBnZZ663ve7UTyXlV
dZe/kltyOJz5euiVILt7eIKXBclgyEXoeF4IKuiIAazeyAi8mME0qpg9IV3REWSt/zjnfz4gsZTo
HUYgEEYiaKcMBfs+vkUqO23w1XGORAZJFb1Jy4tKPljGlPCLpqLL0jvcAhLteKDnaFGQ3FXPtllJ
S/s1ojPnQY6mHVjhyfQQLLSAXdNAcKhXQaLZrz1jGq+XIXRHGc8X7z3ktVTzzaVCpWbjuZWGjwRt
Fba4gz2E5aJpv0uuxeGqa7ztZ7RRdUEEfjwe3lz/1z1EK9cPjMaJB6wOZzcC4JhNBrWfQINgNsWT
8MUKt/DzheDdEevLKyebClZJyjaMDKzMup7GoyayPny3n/R94QreUogkKAe8SuJyA2EdYi1WwiK/
JN5U+aPA8gMrfrL49Zgts8lCpDhNxTHDbYwrCYawd7YgdMbywnVAde92cIBAHlUFEI7GBZMtVP8F
raubQGIvlPAHWScgcuJhAsnkD96vviU/jP139bhZbZsT+TYps8OCdj/WLVBkG0vS8Yj5jmw1YFCO
TeNany6qbNd/QNFp+5M+QkwfH8mOclMg8vrdZ1TiZuh1oqIksF9GjhJdUSFmf8nBS77rpzdFQw+M
c64ZC0QhczrqO88aifVbusSGFTzHVm5p/FaboERcfjYpmwCd5t+MWDb3fnrU5AROABSWjzJWUHEB
C5DgTzQyQUymKKlnWp1/CCdLQyeyWXf6fBEIvjgBNXxMslNP9WLtUL8t8Et29nkl0/r5qe7T88Y5
mQXzc6mgCYkslYYPLip5Jepo6nm3JMxkJ6wjElfSxXYm9K/SpuiXS54uSOVeXbkddg0W8IkaeMhW
rMuYV6MIObXgJfDchMQ0HbSBUn/3snYh6P/dakj+jlJ5VhxK1OYy8/vHcdp/AgorAx1NiOW84dz8
/RGsqYRqGfz8FqLORtAzmiF4g5ClRs3mwpkZF8zdOMtqM3W5v9ujXZ4oZfd06kGmJWSZKejM4V9A
xamkvofcWmktZ7jhDZt48rH8MnO9veL0RbbDWF1P8myP7cLEBtO5Vetj70yE5806R/4L1k/MAo+9
A8pcjWq7NsZQ/US+H1gQHQfXBwJu+mA8A7ibptQ7SP3CrF8WgdV8kHzaN/XljSeU/th3FoAOk/3Y
IxIQN8nJdml/+Ccjnrvhk7VVVlaNp8I3/FaU4ZLq4iK+2/YF4lziUIAcCZaRSHwoPk8fIpn75Fa3
DSj9o9VpU0XpknfoTM+ILHk5uGW7TAbfAIjL/nV/fmR2QhCX2Zb6cfMz9abRwETQQRZRqUnZsTNm
EzwERbMXepRK9DL0vUvHZYlihLDt8BZgdm4UW2g7EHcuvkj3WwF6luXm4G+cKXtK45CoM0WIpnR+
IbvfBBjH15MOl4RbZ1wMc5mdVDX1Z1Ls0gRdMs27CNObHYiGMioBKRlGDcUtckHOa/ZN9XR8o3eo
NIk7FqRnOVO1i8ApumEXkcksJ53XUW1jR/4XEzUPZdFQHEixiGIqf5wF+d4z/f9ttRWenAoQO1Ws
4IlABNsMgdGqYXlPenItfdUdK/WXmk6FdjtkWxdBm55LvKNddtrcbnjjx+9osLrPnZspiSfjHKlD
K+ZZHFAj90yhKxwbxaV8IwuUbxLc02xjJltG0CpZWoJqrsuOlfHHLC42dLiGeA1MXZBdYT0UasB+
F4Vw6Dti6ruHMN7gSpjk3uFpiOCVPhLjWO6Yd01WGX98jTBaWjr3OVD+TRhr5vj262f2PKQViP6M
I/wv54aLPzsHYM68FpTPCY7+xYI68myZR1/wppZe+hZ1Odo6ltEr8EFi0A2GKeQGLUCYpwhF4TuP
zY4vW/ed3FpyeeI7yT+0F62oF5Y6pQfBVu2TQMyYAJd7bB5RlHTy1+cwJWm4dNkjjXo0T+CVlb5p
xxUw+3M8H2GUNSx49/1pkvMaXISb7aMi6QwVI1BK8Y8eJd8A3MUTt8girDFH+BuAyjl1ALBz7aw5
f9GKqGCNtrHrI4ItIddWYFNpRaf5tI+rcRJPDH9tp/TO26Iz8f0BOhW0XYdimed8QZpopZ7HVhCH
VhGQXvUjvsS5gOtBQJmHX9QktjzYqg6wTEyqw78dkYEyAW05QcSaifbGqtDWIZyNHWfL0z6aUwbJ
Xs1NKPb/RGPv/x0GkQhjAQ5qGDH/CE0tpcf5/ru0Ae0581hcE9oOV7Auhn85DPE21ZNAFoWWgMW7
14UFGZ8QREZajdjMIsX1pUafh1ho2A1Hs9G9yvBRSXNv+ipeT7Sd5EzhSF5Ly3k730pe1NXgAJFF
yZZz8B8ybtI2AhjRXcN0k6njDJXpZonpXwlm6+wnMs/gSJ4qbHTuPDPtm2qlNIyddW5XjUVxuz+O
AlYxw4Jvx/ScmaBrdQaOo8HFncY92G2yOngQ69RHemsQcWsnwRXZYFSHkX8QurSU+sHUN/GHGPxQ
1l5EjVHOI14kzPpoDzsw7wfHxK7M7CvUsDEIhk5UgZj9iJQ/P1qGZV2J0W7svsYjSi/+wRWqrqYa
RLC2uIzO687YkTj1XifLH+lmLP0dvHmo1GgVNCx/B/5b4eQYR3GTzk8XrcAEdLQP5A/EKIz+1Scq
1gR4v7iri2LkBhX7/HEHwhRpQbuE5jMBf0LsKJG3Eky34++7XxucoqqaiAXP5wh4y0KvFBQMDasA
I3KokX+9kAAUIotzh7GUHod0lU5fUgxTu3XBiwXVNolJwNTS35Ik4TYrkvDRHmdgLVpHbfXPBd6D
wDkdexK/kU19SHw+OfMlEowa2Hu2rmSgLJgU2trEidRVx5I0Hd0blFJ1atiUzdMldadgDziXdpO6
JAT5gNHjiAMNx9v16WhPG5TgZll7v6WZrG/KEmHtWQDXY6etb/mbhNSZ44Sv2A5Qr9Qlf53HdYeS
2BLKpx+EzM80Mk+G7+SFh3tP7z7WNARTh5ZRS7n6XUqcS7kRGbJT1wA4t8UUryXgHQFbiCmfI2Wn
KONuiG0WH60SLNQilOx2qh9BUPUvj2fG7+hveuGn/aivPgduqI8uqRMt7a0WDpS/rtQey2viJYel
3x+dF+MJGmCNHEcdyShzgbhthTrzFd+9ezar6+Gwnc39SpcIxOoZ+DVhrVJl30s4CGlFBOB0ca46
EsketW75Vi34xy3oodcAA3qNT8BkXQ41miPgrqKcZzVnWhrcQiZ0lM0VTQuNEWf5LxDCRT5zFCtu
2/yiTSC2Qb4kRkMsXRI0qtywlNP1/kBp++L0UhmCkM/cri93eD6nHPhA/shGV96K+gk9NFGbzK8l
OWQm9ZfxXk5VeP9der7H6sDGCRfrWAsWYZ3f3HgrLpe7D3/yJB2OqsXq05AZioxw4jPx+bZMVPF2
aomUjFRGM9SLnWCgJcRf1oURVfXfDGpDdWjKvE5VTOdO2G2VCYSN0KxHfCGZ2O0QxWtA/UWekqOM
6SHlLJTG9F4tjnWMdthcQdgx/Uk7ZvZPfPCOFLLEWSe2TR2wiX7Tmvt8UswayFGB59JT+0bHQCRj
flvgMoDj3zPXYoxD8xHm7936ReuDLYtXiiZFXiigs969kGlbhig4P1dtKUnP9s11PTTbyer1fLSC
L17OLGpJFesw1FAZHBloFjmnJcLKuDpkZvmNlPsvlmiL874KYgxlCC/TXekaUSETSMNUbjwTw3Vz
IsNJXxvYM9ei859Jrn2FHhfFjZzWnpDi0KbpsFmMSd9kcdU6F079BY4EyYo2+qI1OpldKKMooenB
6J0dsRNAzDzqYZmucqrlnHhrSWv4r44TLQATM0HnfDaDbPuwkqjplxy432dCeOrAdwJqb3V8aD7T
DqrSSMOhVWqeWktlT1/bYdROOsHZa125ONxqboE2BHSWvNVwbKl1SLdIh/m+MI7XrwfJxky9EZOp
uQqXZv93VIOUhEQM90Gud03FfavNwf0nKL1aM3Geqva3Uf+6PVWF1btlMxLXDYdj39mHWTyiUpRP
0EuhI69kh3PMHPHDNCUB+EQkH4W5UAwvt3mAn6cNPfZO7JocxbZ3MiQHOh9acc1KBSdq041tquQi
fOu7GJSrmumPNZJCdar4ACcvpBeJZNCNH3k8q9VSv28Ucv+dl3lMN9e9bn0FsO2xgogbaUPiXpED
XmMOz3xYntDPvDyvqcXRlL1dw5+cnVaDJGXvYYlDSXppdONMquVqJ24fyS33zFUcAXstg/70Z5JI
nOfY2spLagACIGaeoCqNRAlMp3R2oDI2NDIE3oaNlEbGHceNc5KfPmy8wFWXD9MpVLIkWYoYeDOj
rUG5AmTfXQP/KSRvQagbMUxPnc+6hfq7kboDRo6sqx5FgemkjUh9LcFkR5PjS74h97Rl0F0ZiHr7
g9FsUC3krT/qffqv7fDnUnDs5w49SLGt2NIzovnazaw4p+/H2kgaO/YSaeio82fPS3gDJFS9yu4y
OH2CNppelxJDMS1QNAn+oHEe13GDBMulgQJr+8iETcMlucrnap4s7fWaDpA4P54kByIGIX0AvcBN
IfdKawIJfCHR7i3OUxwpme/k+FJjlYRUki4VyruHpLGfearQ9M8kRWCw7vxhJJnaJXeoBwUwhYVs
sVLCYklI7TCSJslaAVLeI5JM4stS90BtZwqabJs4HhJtJwoSEat9HKVEJzEMjtrXjfGGbTtqQ4em
FqZnN9JIbsQLhgSLp312JO21/LYlCFrSkiDU3W59E+McoLVOLJ2YalFp1z4008BSl4qka47dlH7X
X8L6zwsQy56DhvlgZFhuftqUWKWS/S9KbuKdsp+ei6y39dIAkmyGUwxbXFrtPItrItbNhiJ4SJt8
atklGRlLwxTg/b0x+EbJ4hq1dlRYf++PYuU6IEsu+SZ4m2DrlUw1o3b9iB9MQ3a1R+VY/L4IvkUg
jEIHgAgM7KwrLPeNJ61lv2ZRVumVpC/fAohpNw0m8nlQcDk/1B3/bwVsPvytwWyO/IKA4tGXWeHz
JbmTDXGMnsjGZV31ZL45EYKpQPKi1IMC/0x6ZbGoaKLoc7ClvhCW/pNylsfgJA/AEdZbx6I+UyaK
VvyH4QRwq60HXEVfjv+1uNYjg6kG49B6HnAjqoBzJKYFPFOCyiHIBP1xHyFpQ2NQ2LJynx0oSP+2
xowHucq3YZaQPZMG8d0W+MgoHrOSH/HzGUzbWEgq28BY94re3AoJWsV90A4UlILAYah4DLDeT0ps
iBHI3h4cxVyo/SzbKL+7fMyzXABtCvX17+VXVBhQopnc1yn61AQh4UinWaDp1jGfG/FIoOacCvCL
oTKHU7OJiozR+9fpq1/hrzoUId6zCRPzhCZ51GUMZbGMKM4uWg2mpMEhUhUzhyjUJAJNxEuLGIu+
DidWz6IayCm12u6HCQ9IHN2UF9S09LsWvUtcT/Auc1TwLQQsxNTBfRpUzdtcRXfB/VWV25911iey
u5wJzBhaX1e1CoiCBlUeyXlIwMSli3JYyos0RVM0D8JmUkadxBm2uzc8weLbgUc9DSrPbtAyJJs6
M0vVCXriczcjtRDG+3EsziDtiRjo0ku+BajadtsmEsBhugFOGj3C19qYl/Mr9qjOGITpXOVj0eXu
H/FoTk7z6m1t1VP10Ui9vLPaQFLkjiwb3FRaP4KEktsk6FuTp0L3DHWX4h//hUSYa9TLtH/QubH7
hZCk3yYR7WFqIRxunHMGvFLz/BhUv19/v9nOnpbvP7p5n4cytUgC4/BOwTidJlLfjuj6cFHZkhtA
vjyzsSs44ZnuM7Rrl1F3nhQiQ1Ay1NoLq2Hbpu1e7M+zXgCqP2Xpx6lq0gl/kFF+ChDPEEoPvZh5
/dENacRtGel/Mp5BKtGk6D6L115Ka2C+9P07XP6aBTr++N/reR7zzydLENoGhtysatVpRaEGK7CU
G26VPKAt5/SqdZZ4sR3w92y4xi3OqNHWmpvI612pByA9z3sb5AIu8AsQhOFeGqakRcxQs/xhp68x
cXAxjZ8II4ab0C7KkepNJGozrMs4FvtoWDe6M2mEjylbW/k8sE9VDCuZ60DgAPl7TlMiofGA1D0X
zGCA3/QX09MWjxQ3F0YFD0gC5HHBb5brvXJ35v2F4QXf3CG65UPLJ4ANrS/j8jeVsEkqcjX6P6vB
tOdjBh1yL5jNo2O7zq1MJa7NpGAJSTnNHR0kwhT9cXpzLdsz3dKT5Hax+5XOwTxHulEi/mRUCYjk
Iq9JPyvLbW2z/Kqj5u73dkLn01IQo93pNH4f5AaaxXkfuRnp4EcKulZs02B2h8VsPPFMYs9Jc5xY
JqJW5RUSuHadTm0vQgIfD/jstGPJ6bM4FPmwxXfV2FU1hk+FFxg4SdWcnfROf6B+OqckN7aWShIB
KYcBCBRy+1JVZlp5fPgbgz5oblv/qcnVJIJUeI4k2M8e0DD/npaD06mgCygzeeaJp87j8DeBP1h+
iMYokIfWcc71x2x2eVsxxSfgrp2YnDNlqWwwyfbb0J4Ezcjlj5rnHKEHlwpzswbx+bxgL/HgCuKC
tOPapo8ZsexMQcurID3RSQkcioyort3Sv7joDAjSIwp46Mvwnlq7qQ8sgtTd+uJhKD2Dzk0wmceS
h7fCvhT0U8ZG0aRgdI6EtDaz+FRxUXFhWC1eLuihWrNxqotuUO4k6EizDxofzE1mnsueE9KYvOrk
7wsfudQe9VGIB7o+w0peH/hS6O+2YiEMymccYT4cxgsKR3ka4AoB+a3HjtEtDXZSEsgXeT27nArq
ZXfmajd4XT4t6estSqpRguatCqdpux+aubBSjWD4dhAiBUQB7Sxdia2DkquibnqIdy1bbStZnRkU
HDA+TVckiILLxvN0iQ78UjgZNKWqD3xrP4KH1qWJoqt+6E2KHCzaZJv2+dUsHBmz7ehRqHWsqKwM
JGtIwDmMfk8bEmyJJtXGhfeOaoOlZyYyPH1vvNfTQp/uu5MEMWSR7dQDaloBPaN87Vr4mWGPvjtc
gMN0KMhZzscSd5lVdCZVdrePbw2GhHD/OIRbbMYKLN6Ehny78KFkvYjPv/m9SGD4qAZ+rpLmipVm
CdaB0h4ny4PY5hX0q42GL18voJiW8a9bqqS9PUMTGmMj41fGEuD+o3sspjqwGR4SLakGZMHQ2i7t
fyTI6l4yBen5VOjSP/0/xRS78CUT1KQ5NnAQesPwppw5WvVIhuIWF97BAewCUxX1BkCpUMBk14CH
AuI2Vd8Ld/LCnHk+eaSSDxC1a7X8XlScO16EGbaiXkm2ejIcR1UX+5QFDz9vjSKJR3kBDLQmzDah
PoQMM1aGq9N80gviHo2IPHc7C6b/1zN10ryMaAArtKezHJICeI8NH59xKePuI6XMU5/c51R5z16K
ko3HpbCcVOMlg862qV+0Ys7z1bRoOOPGa1eAEDHhgV4IXYlbNmifAPk8fSP1Rlh/glzhkDnG27gL
Po/lI2NBHmlpUgn4XwCqhBCJ761bq890R5GtTX9cvQTmDqUMFJ4QAZNt1fk2GPNBAxMIIAzkKy1U
zwmhr3pD8wytZTtCpkWKuaNUEDaXtSclyiuU068RSl0Sn3kquHdF84HOHXa8LDNMstxFU6UyKPAz
AY2ZdvDqoHXYXT3qPrDwlChLNPFuGWpcQFMf0MUkjDJ1Aq9XuF47IsT/TlCagLPo1HpX9wpOR4pp
Wrx+EUHt5g0obBLxKa8BLKr/j5rpXD6Azk8TrRH+o4bIKtRYEo+/ye5ttSsgJh42d6iJAEk2fju6
dxa7sTgHliX0SekpafKV7EcdOvBubwEXaOsnHzV9cZ6gmaf98K+c+BnrhebqHQKBPpp4gXbZTF7L
K1b+ZDdboVF7FO2to+ltoTBhg3MExBw0QKIBtk7RuqkPtVXVs3coq6CTa6fKZBwLgcs5PXrj9b6G
KAfogIn9d7PbOwPmMwOaoKIeZLFr0CF8h/DkdlwqpOhSLMjKhNvWgzZu9mXQa7wGWuFTXrxtPWfx
ZzyB6hWKnsuEWv4qMl4Gcl/4ZV9HEw4XUOSUiQwlO5deI+8ZxrmnpPkpaaoBboq/+PPMet8mQLL0
vuiRTXpmakI+KjW1vj9evnmGj1W8t7KUx/PWL+5L1+O8k/dRNd/QNhKRwvB46a8ckLaz9BaaOruA
/xOZzE0adwBI4z6OTgJLQTFriiEbne1Cvpf42FvOCAWkY01hT/z8h6e7h4XLi4xarSqH5Jn19YTk
LddMfQBWOP9gDMFk33RIw+zjb6T5ArlsI9opIeZ4ev8/UxM+Ea9fRhzubwzQ3Ff0KX7sI0T8zOOe
IKzHJvCwSCQdMQXVgDPoj99R5SWZPXcDV1m3Fy0wfUJl9DGr5UXFO4FCEmoylg4kFmfsiBW9jkfm
NLRMHiRLxPihhBLfUuhRBaoc41Im7ALTihA7L0GoofmzK8igrThB4wrH3ASnOklpCHKO+hw9teJn
bHkZvGmGqGdbECCHF7vHGW92KX6CRqi8sgSmrGQ6Ththv5GSSaMHpqVf7DVSqdXpx53A/iIPcwkk
XxIIntD3Z0Cen/RIL5UAE4aQ+PjoI7cEHOjDWWZ8uHPr6tn19vr6Y6Jwwp4SzL+Wjknk/g6VZFnC
+v+2fIH4kgToQz1ZSzMRDLUagNHsxgZLnUh2xhguwjEwXbfRH0+5zFetUEimteIMdp6ZUoumAiGO
7fKUnVaM5zr1UwLrJ6gNpBF9sHSeZu83qQojNXLQIwQbxPJPzFmneVaf1ChbB0fgF3AxV0FYJsrr
6rzl3e31cxId677WKkLtPYtj+TNS5rBZ5G7CokfFyVE7EwRgfkLwd6QdtPB2Tc8cE3f1ek5Mj7yD
sF+lJx1DGIjuwnf5DfeazpYTQGN1wI7BM4nRg6GyNzWK/e9N4aVu1YW7F2P/LjGYcFlkdwBjwqXK
ZkgDOfT9guNILFBKRzVMJlnq6zOsnOt9WTBEz6a590FxEV8TQJofP8yU89rbk3mpHBZEHkPDYJ8b
N1+okznZxHzj4o6yx2WPqWI5zc6f/jPdFdvmPkGT+wUCsJtdQxbLAY5rR4xR3+WuDlXHcT/XNFsZ
rOxaOY7PvWxOC2+siZQkiwGtofZlNGuIsMAjxWW3ZvDU2Eb3OVQChJJpYQiWwFI3jrpAceTuV1o/
jzqNdbh5ddesnJemwugmnkzmWFeeFAvi1WuKPZdl69SfPObMI+sEitAl746ptWYmgg+8Hw2cozC+
2rPrDYsQWht7A7lZNdm52slWAL5HXTqPPPAs9VZgN1uZKfTbU5CIC8wabLr+8lGEGBOMMsCDClXC
5zKFBN4SAbeKYJFX1bG6l1O88jnVrBVxTxa9Dx/ITiXCvyv4Bfli0Qcxmbr5r8093d/vbjCUFvQt
E4mlO7pfaRtsoh2rZINqdgwLWOhK5w2qrZgWRJPyFsAbxFNa1m0NEqqpA8iIHH+4bwCjpMGCPrP0
CMI0f7myt5plvIuWJVoDwufh2Pt1EPz63fziu5dToN3v8YLph7KVrX5yQHQvT0tvtitsbG7ttl27
euIaT7D1i/IUA75lpfTk6raN0iE8AwqW8SR9Pa8uLyBUNEuYersM8SjktlsUl33WrkICTkR9Lx5M
9WFOhOBvjdbatXyYkkMRC+UjaHXhO/pbyL9murVaHZ4eRj4KKaIoDQ/E1BxpeJi7G+FP22BTV4IM
zR3UJEsmHogvZnDg0AS4s8i0/pDCBLJhisYWUJTIJWZvcg3jJH/Ba0nYo6qG/9E9ScynHhB8XXYp
Gqz5Mbeunh6Iqs5RQVpJEsvO/7TcyofYN6sBjtIjctL/C5q1G/JTW5MiGP0SAsT0zSU8DhMMNFoV
iBV5yWjwWwMH39QirC8iBW8nGNhL5U7hkoA+SGzloXR+vUhN8rCD+Wiu6SMnoavh0EWk2zaeBwN+
9wfq8eBtMKa15PSBXUEQqmu0QY9nA07xbH/ssfVsHK2wCi85Wn4SUd0yUtNdZu5iFDRlrP+iujDk
O/gYvTDPJ/AmbJBp36zATADLKt9oa4W9oeUPXPQvIkYAw8fOamv8Kmsk2pdgv0fR4LEhjU1e9qGW
00ZVflac83nJR8LI31/A6QZoIi9ckgNj27vqdbM+9zbbDHEoeNiXgEWU3WPeKP6oxLMHD6UEeifN
e7oMN1NWCoBjccro+FApaEwR/DWmNA1E2h2mF5Hp6Oo0SGMtH0KlTIoIn/+bvn5ZZhCTQCi2lgKu
grJbyVVUNaXwBwCF7rXyNF6wzcKLbZSY+6Nup6fNdw7PHAdsfk1aMnV/Gh0HdOGZ/Y8Hn4zTrJ1E
DAUntk12nrnrdgOK4LJ/1B2VHUyRBB3tBtfWJ2EHi4KXtBPLLFLeYIevBqvWgKwZ0ssuwPNpTOAy
5oRFQTKTr5qQSOpSBVZGYMT/ZnGRoWogUWKC9Oza0LgeGw2I4sjpdADug9gKLRew02SvVCe+k1cj
rGGpIju94++Cz/MeUJueOroikdVuJ5KXT7xYmcs4Gm8IUingb2ubxuYVGy1K6OKjGeE3csWhoExj
NE4d8QKMtco5N+1EdIP6dlE5ADbVLd6k6+PI9VVerAekzwc/AQ7IoNCV2Eca8he9A0jIQeKEN/tu
ElD09UJD5ZUyvqskVXs7Ejo+jEuxSzljOJ4HyKnlcwpzFUwOIHXSf5GJD+BFJTbhN81dSOAAYkgU
Yzvdtt2c4uktL/6RzdWV7m1Dpr/wqqIFXi1pIuHOeRhHkDIsjaxG+zOj8wSgKfp2xodtq6YwYZJ9
nLvzpD70Gtk3DqMhbRRE8juEHtM1RPV4LrIlJ8O5+8eNoDT6yKyA1FZAvao5FWd1INax3V8XzN14
yRyjw/9NQwA0g3vDLv0GwReFB4q7oHB2Qpf7kkKX9eI6TfbFSBQrXboSLRfnttQj69U3RYVSndoK
96BYH7a5TpS/BiIZGTKoaIiWcRJY4HpeMN46CCjbK1AwDOftKgz2OqEwszQ4v6BxuFilbpyZp1cg
3ERJyMTtJn6dz5kGEtffAV8Am6qssADg/7zkVt5Z+yisB332pFz9R+CH9rTUtu64rJZq/oFmPjuX
p8K/PFwQZMDzc+guvRsBtuhZug8ySlLzbUzdQQvFsYzzX6yE0/rarZOf2UQj+xCDYn54znnsK/XF
pg6xie2tT9qq+XItTje/BiLI5j5GYV/L7OGnx3gDT3es5ZcMgaA1OQpS+cgFdNsqj7yMWRLTuxr2
YJ8Iz9ofNKhLj4DJtkC1wBx6XA2bYxumnmfLwMQMyjhecwdditTOg333l+sWsHcUF/7/X+QkrCk5
RcsNpWVGK/vn7x0wsTFgrfRXyU0JVJ50G9/4ZvG+nEtuZSNz/OQqQu5M6etBSAamQuHFQ0VlhI8I
4auCR3if8VIb+MT/TQs/LyfRmefz7ST/CLdnlAP/rHrH9nog1M1mBh9pzpJ8Wvn1cQhwaHQVgLmt
UyegHbOiHFLEnGd1t31CqnuAPw67DK9lv3NPJlA76IYdDuxF/OfmIq+SeQRoJXVcI33H+3JLz709
ZCrx1jrziKHV2Wgu4EckS2/JgIIbIor+OfHMFZ9V4O8LeM6jxdWDLlhLBt/jQIxB1TpFccsfDbDo
IfwNhnUqjBs+SBYlQLBaZxfM5EgNyVHJcSTou6K+HgpdxMaVA0BykgylWr7+7CDbPxP4YOl+257l
+rBRP5s9YV+mCm+nN1fak5XDL0gKTpJAPZpAgGRvtZSxF2We29RDbVfC91RIeu1m0+7b20aSH8hk
UgozJbFsWHYd4ZKhMNFCMfUpgXrKaHsm9JEpQC5BHnDGhWETbHu+GXzzZh98tBkzh/11NzZixQTD
/Iba/96eEZ/I/V9q4q+DkXP4VC8UH0pWYvpfbpO522i+8+KRfHIrDWCplBZSQoglWmTz5dO/sDjr
/+OSQoAOyoyY/NA4z7shZ+qKgNCnZo28n4mSLIMCIcXFok2ZpQbCuLwC/lcrfeuERehS6bbzZlLT
mAJHRo5ddK/siQ89dYMNcoCstwsv4L0hiY3tTVHc4n1aFfcxtDxmr+gf5QJOx3611qXRA1v52b4g
Fq38eDwypjTtkA6g2N+CJwd9+ccGZCH42ffxzGYNrvfPCbrroY0XkcYxjrdpt22eXZLgzKZkUuZV
nm9ReTphQKS2LvWK2c9s3F5T1pcUj8lKe7mMEM9Y5UVMW8RlVtePwyUODgc8vZBeiMqH9NiInBfJ
UcjLjg92lMccfvpKaI7ZZGsIBA5YIiH16xRdiyBcAJ91/YK05KMQm5v6o/qYq83+wRWI887065AR
W2/e/FBaSmerB1rvAfxXKVMxqqppFXjORc1/uKZziQiKZfa9v27giCWjibR2i6oYklacpieAGO7n
yaEkGsTVkaMgqt6wTI05z3LFSFyTVdEKd9qH+Gor0TaJJZOvAKxjPlERTt/PV9NcWcPPfZZSYIFW
9/oDCa6blSEP/l9M+9I1iUeKBb3BrSLgqLgmt76gpFbQTyyxrY1srhU50DRhDGSXpDgz92IxX+SX
e/HQASl77VBwprdliBATiX24EOPBcPqk6ifx76c26OsP4hYPcDIGMAr43V67tt1I5Oj/XEjGdx62
uYOyc0aMFusAUpIiRTRIaNjiyGzOTKXeYIg39eB/cmbbI7BZP15763rzO81XP/MJewE67BxY6SqB
hoIpUOiiQ/668Iv98KFlFxMOpKa5We9b71IBHnAz5y6Dy+mLYyU7BweqQt360hzkYM6yEbUqqb3x
jDiSGKyk+4dBstD8k8Z2guod/kFPjS4dS8NGiaR0NXWbddX1Vri+OkIBtoZOnzTmn9DqtcDEtjol
cVMhG+Jol4IVto8rEC8po86ti6QoKTOOKi6Li8ojmeQyXqk9DCGrvcI+xSJBvsGAwS8G1kvSsV0I
PdxCk8ffFQ9K4SO6Flv/L3DFKx3oKOrV7aj07XMfgI9ckAZ10sKAigC8qnZ/0euZtiQD/Gn3Ubeo
/vEgmHY9tq2Hy2Iuf0OIuqrvnHiVZL1izzQPwcA/4KRxZ+THkmlE72CD3G2hi66oTbRnZQ+trdSa
ik68dpobxgKGXHCe5Gp+BSwzq3Yi4Pd6opLb7mnMYkYTpv5JjzzfhaT0ojhJNUYWbJDHxy4Z+70e
WJMjU4hbpYt/2BCqVWOUu1pWOCGF0hMC9HUNFoN/8AVO8ckfN4ZOv1HCqDv26gumZDQpC2gyzEfx
qJKum3tvTvYxkp8VDmY9fZKek737dmJitTOdSXMB5Vld7fRe/TXEYi4f01gJ43HVlkj6MWj/WL3h
f36C/DRGXRQVfyDo7s9X3ayemZLtRN73NOsjHwtXZl8R47oVprpGVpYkaEWFGBz3byq/JdWtYGca
SW0dJhTHHs/O8sCTeX7seWyEkJS6RHIOov+yshbJFnD0dAcLFVFjQ1x96oJ4pzjJSNTXTv/UP9La
rhLsLbobCGO0w2xZLZ1Vn/lvnhOC5rLeZPQw5kyxaFOr5hIk/LngTIIPHDoHkubov8dWx+27+6Zo
RBKpQzjsxC2xzfUD562drem/WlcqPPNf6auSu8ty4NjLuxq1Nn0OJO+Xn9fdnM3MPsWNfpZ2dFBT
1B2BsBUy8ajXlw30DeNryc4L5y1dU7AlMr6a7lWiSaO89iMC1cJogcKkSNSiqqWbGWOEwm8wXvZ3
I7V4RZwwtV748YHUtTgSfz2dfchE3pOTAFnzkrw+0APlOFj6WUfvqAx9Rf67yO0TyfAbyNNx6L/M
pRuV2c/nE5AcFF5tZeixcEzpx19JgkBpGmd0JCstROMHXYLR1ndlewd2lYQmm+QaF8nLZTh2xieR
LzhXYGqMiMbtqpHsOuDFhQRBJyTdaJFeySkJDEw9D9kHkseZw5BiCxCdAlKExUxYjb0phaZFtx6M
dEgidX++9Dh2dqBc/s7/v/nk747hkA2KuFW2rYbqKKHtvsOOQcib7+mrd3ZkDtlYNQkrDHKTCwPm
Ne8yycY+KG17UZwmPAUoGAHysQmpDu2x2NAEo/L6SMwzaCeb3Jxi5ckWOGRpYuELfNaRubtXKQYh
Sn9+ARCPdrN1Jr2R5f1WKXBFW153uKfNQTHEoTFrWqpN7gzF1/7n486Cy77wQ+pwRAzggV5XNGTA
OXrwPqqrZfCdyFM1vP9tskqsnSY5XXNocR4xsZ9lJ2o31YCb7J36kd1MQTJtqeRA+dAiD3dW623x
JOc0U2WUeESJg8JPGRm3QpEzvN6VHF7s5uWq9bQw2TagL0jdLHhylXtEX0kYuf3TnufpQb6BBe7v
PbdN8c19qyjMjC6kebKZCdoi/wTQ5ncg9OEHYSC5H7H6FhcDXXWKLMJPZHmMOab8JenSXZViLRc9
KvNFnE9xHsYpeg1YLRA/t9QhnJbAAjUEs+HRkFyLK6mucRnEgH15vdksrilQV9DqFe66pNz6daNL
Xtt3k6J+crLsYEkQcXxB0gc3L6LNyK+wAnBxUbuo0knq5WP8x9IVnTi3iC973Tgi2SRR83xP//+i
j5+bkxMJFxu+u6nTrnH2DbAo4QjJEsaRHSatetVnymJhEQFWoICcA2htuwHLIul3gsyp4Tt6n85Q
Zn+4WonmOMuYQwfCTzHU+O2BZaKbiUDbosfWSQg0t+vernV7otKdEChg/NZ+9jn8AdXWpXRfqUcW
EYNM5dr78sVH34R9OqdMlF/XmD2zKf52n9hgrB/eXdENv7eP9O0UjYRW2QCsbUJuLe3reppQiua6
aOVai5l+5uaHKTxgpu/10icNVFxY0u0zABdPNQjuYQ0ntcEQgSmVM0kjbhRW/0gX54gwLU8H9vua
ZIQNeLcXa132WybNcxkpD8I3sR30ON48/hDwIhAA6etnxFWWT4mV/XMUeT3mdGUuFDccFenWU1uT
mqUpX5eBa6u4TUR36RCu2Rq0s+6j5dtYIdoN2gcZ6ZE0b21VZ5NGmX1VPZObRVhnh1rYFYkLFcEL
gwu8LfQKAlBhXLIb6tU6AFDU1szn11lbIfp3avDbqiZSVUeEmepKpdQRa2bF2QADut7eckRoTbA7
EvbIz+Q2FdJsCjClntU7Q2hjJWXadU0xiB7qzUb+FqYB6U4NzMSPnjaQMMhSjhRndwGXmRm7YiLu
VmtqlzaK9Dn+u708diXQG9skQDqOMqo+d/0tzhtaARYYFzJQ4I05UmP3n3nYJjexbQeB5I+a8yRc
xYbV3lslQq5+JsvglfVElnHigaPqv4qWVha5Dm2gcmdnygLr4pPrHhpjVMHR4LvZuP3/hznR3jO9
A8NlIxKkVAdxTaKdg3OHKckjgpEcNUe2QLfJ7cz8B7o8Yy92H0eB/Gw4x9dQ3DNUJGnrP+zjQ4/f
CtoKTK6lJ00INH7qwiZeCITRIL6vf9TpQ+mhBOUVbVOQG2w4D24R4gUXrEOoPMWffWUzDWH7s9Z7
TkEfltIMXfMh1tsuW6kJRIx7DneZZwag1FQJf7t5xTrP0zXQnSsI/Wlq1kjy/V+x23lin/NRrndf
sqy8JEXAX4k4gjt0Jd7ssQpT+MyXvGEd+BaMQiz/JJ5saMgmx0VvWt41Pg1DPO8MrkSmDdyXSgL/
7+2wEF/OKqt+n1h/jIPr8PWwLaRsxRYCnhtLhI1jR4nAuEqFQBX6vsZ5P1KDXwPYKA1z2e3hyRE1
kCqbXG2MTFZRWq2ywudP1lErldvxFzoi/EdMrnkEv7/pp7fBzCHL0sM/Nt5f5eUNDJpEQk2huD21
rxcr7Ld9yehXTpb04hAI7WZnjYQSu+G6/czvRYU1RGr6/xbp9V3sDiIExp6HkrDP8GrOcMpddmcG
FdaCQ3OCJr4mLChjfb2YS/KzBqjlpyaJynmoohslV3R7jMleTQHgoEAwyU5CSzk0Sbd1Gjw+O9S+
PyIwUKniYtCTvteE9G74igkcq+z0BGPFHyrFOXm+VG+fcKv0sr/Qa4TywnaNaNE6m4C295l7uru1
vzNqVTWP9YeNN2F85u93EDd/28eGYx5KqivAr2hIPnQFu05/ORqX5bmjefVUCEd8wiBJup2LWBJ8
cPlA2ex90OzUGZ9gUNjsdhqTJ/ADLptpGdBzG8GGZAap1iGoJn55/nGNVA8cnwoKfQJ0d5UVJ2Yn
I4fFPTPyJAlBhnDhZ2FXrTTI5BEHmDz74bgJUewXWxYQVioAWS274JARvPnjXcPLfMG8kVE8530x
7hExNaIl9SDTpxLYYr7oxztAJN8UPlP7j8FC0+7F7vuO7/zx87xfDNJyuXZgkeyrGhcfBo29INTJ
0CHmrTpA9zfKvOEHd+Q7/hzMxF2cUi2JwRVoXZCNMM2CrLINA8ndexwGfDDfL8zUU3WK7CfBUsOT
yxqO5QkdxwIjZx/mvntr5TWgoHi2FklG/sXgX4xcl/aicW7ppsIlCE2Cju595A5LPYdk/ELnKcdv
1PikxW0Nrr66wQRZrkSBQtu1UZzF1y7dR/KT31kPySMga+7w97gbAmw3zFX1IJHI83mybJQjiomX
TG1SBPaEsw+3v+waSAe71d7J12gAW6fO22oywVIIoK/q9N63Ha9YHmwdJPdzk7NqROoddxGPvk4k
5/tc1XdAAO0LbdeZMA3+0RS923imlJst83/X0GE4wsRkeLkbq+7LSvkkhjGvpycPSBesrY15K0CU
yd3A1QRyoIU5RjXL+9DHjWdUHV/Q95b1l8ZMrRLBz6IzY+jO8ZU+3IIEUn/gVA57tcKvmIM27pme
TV+ncw/+knYFW5vmJJ1qqC3Fyy+Fs08EkL2QbiQeRTSvGVwreDlGfzSRTTGWe9TZ15bMshOV9rRT
hT0h8C+aG3nrv0eqHG3kU7t96paKvQQFbANBoaBM/ulNFxsFqC4+iLnmRGKhXlSoaNLEF1q6frrZ
OddZLlAAZx9l0Tzm7u/De71itAYoyUF5O1A5tdYFlJv3JWUOzyYeL0c9fsCcJNToznQyYvknN1eH
qO5DjfIFADv50WAOl3lCadR3YeCX3QUBF69twZusJXd2n0AXk0nRCgS1yE9i5Q1MChvW9r9d5KWJ
9fb9j59efsmxNC0YZE1hjYLiVaK+uudiy88kEoA70gOEN0ySpO+IUnBKTdCN82e+w3oXD5zDsYlu
tYIMYVxdUNceLbqZEPy/qKp9+YIIK2Y3UaFPuUViKGW5gTyJpeD9xaD27WTZ2/dpcWnqWVucvrWs
E746MfvSVnSHlG0P1aodMxOBb0xcREe1cBSCeacnD602RYOZNKfpbkoY1yMOXGEcEp/99HWm6uTj
n1xjrsW2gQ4tyXmdNbpx6ebg56fHISn7NcMUIXPBwgg8f4vtA1YqsDx7HQ3qCWjqYfjQTP9+ccjk
+FcWMiZy623ng+lFI99uYmkMaAXPkdqXAFcTAdCQW18VmdS7erQwciKjwnrT1WKRdep5QtIRWJJx
zav0xzMxsJSvf/0nydqTmQ99WB/thqMPsQJxJO0JShZDmG5SZybAqabEaBx8aapkomxGjwGt/t0h
NJkm8QaxyEYS8jL1Xb/M5RBiVr/d5YBHA6KPLmL5AlpaTFfX1XBV8Mx4lJcs/KnCP+qZ/3/w9ibo
fQKr54iIlPT8IWSKOAHnzM835cGx5Z3YOwVl/k1+MmdoqOxy+rN2HU/Bn+WCGOLlWX0723xgSYlx
QWjOvBn4OD2TsXi+PCkCeRZkzqc2kdQkV5A5jfSeNHDj00WWd56kOoD0rxZKGTurEwtzZZat+l8+
+SsdbCsNKTkmFFMmwPHxqCpNn+n3nDUiVU90q7zgeQ6UM5kikIr7xIDCFUfi+cjpLkMS/hY7esvI
rlYyigdLxksBRZzYsuNaob1qNk0uWmlB7YvLCvJnE7EcPOnAabX/Z6iOyts9jXPY/kaE8Io25hZQ
lbx1jzx+jZvpo9F9q7PVjaOMobeARH8m6GIX9LavUychAbuSA93t8mSOQt3JqmZV4LEFto7yinaM
VjF9pIHwPnUlLLwdO6MtqTT+cLgRFHw4tAgh6Ji5NvKI0UHqyqsP7wXp8RqkkbSrus7WIVOiSyj9
dTWXA+D2Gy8HI17o80CzOWQIETbHrIKJytw3RHr0vlvzX6r2Wu9deLhYH/37L+fuGk9MB/7veUh1
cwOGVRKjkeMwgKTx5b8MtYbCvK3SSrL2awOwYqLjrJFXaVK4kGFgD4/nkmEg+MuWvzIigHWgBPxT
qEJ+hCifaSVb2t6mND76evjrxP++no/k0rVkkdbVoUKy6rzEOLDkLpK0hycVNuUzi8cZ6uNZsNWa
gc2/wDt3yJtbFaxeRU2N6q/ioY0HhWFfuV+OzQ/XHsNVYEJBe5j3r2W61d1cAh87ZOk9J9Hsl8FK
duqxdSoCeRHdQ7qUtJWCSrgOzRTNMHXykMXrH+NTbhpMHvXNtz9PvbIu2Ted+ma5ExHeFyMmn9+D
HsxCTpKfFXHUss/0xXRWyDI3gLJzdbRnTn57qS0Ftl6LLCeY05eVTECKkxYG5KpQ6lnA9CpqLkd5
Gl6n7YiM0fcaSBIQNc6p5W9DFgKuV0tZzD745tNs5rUyqRWB80FDVPoADZzYQUUKqdmUlDSrp5v/
P2itWJfg88c60c7+Wi82guRI9dx4FNELefcrNsK+7dvXaSO7v4lwm5oPejsJzmaJaX7v0ZRDIsp9
9OR/PnMvx1JIJTgoTU2RKHSF/ztYw+/ClbEd6d0leDNxY19ltwKWOkYfxAmIclqfRDymvJSmEACT
OVJOusviB1HC7qBSq8gwn4uIs1vOaYOoXF10lhPW7VmT6og92CyBX8MMlefEGRDnaqOZWXrtfxoW
9m/OYNrVNfBap1H/SUrtvBMqlxV77hlsbtCZcT4K2DJENfrT/lVMRyrxHhGG0zv78N9O8w1i8vaX
X5on1Ue1ne4S3IpKPkw842Dxtdw4Ga0nmxODfEpnrfkLS9/9tHd1DYsA0qR9QGbzJFUHz2wD2NKB
Huc4EVAiGkvB2NnfpITgNcs74ciXHjKFQdZmWjfyno+2DtemsvJUSFe3ygZ1onkjnNPW4/aV320K
HK9R5y/YP35kdJqeblm/sioKCDG3zInELAO6nhzRHGLBak60aTQR14IahqJzhz/+L+zHeUTyM/ho
4BIU3vVGtI95zOG7lQoPxRNoKsxGdM+F5zCkSrg3VkU1+foOLDtGX6CV50dUzo3cKrP1LHkuRPgo
pJSDTNg/9xarFhkO4RIj4SmJlnoNwX+iWp7DfnA3aUEQVl1CKQWgUGuvSGo7kK2J7ug+5zto+N14
9NThx5f7OfDZiSmck9/mwjl4Wl/N9zbrpmxJOdByOAsFQ5XMWHCHxSUvpzIPXnhJUTAGdKSUDzGi
o1lBKYvpdYnA8kIAZRBXPUP61CXMVEHE6gDFV2dPL2JmDrUNRhkIzXOhQ7UZPFC4doHsEGIlAdFe
ID+zIeEHlI464wqntHJ+TCAv0bNKq+GPm0i5Q80f/kBniinlg5sXP3VQVAw6mJ8GbBv/+XVW/K8l
lWjNtrT23Of4+KyTmjnwUl3+iIhKGnf3o+DZZvDMjzi5er04Tal9Kmn4ADYw6OwjCF8u5kgDa5LK
aR06/HFRGJPGLBD98zK4PUi+/XHGvETQ0pBkqlD7Q37zZYMvrJIsNf5WNj96NzXVmSIUtK1e66Vp
m02DNbGgGyWnHhm1C2JMsPpfkWjKKB9ykbQ8CI5/3/sWHlElK+ewnBbia53h5H6a6bVcAI1DV/5y
zeceLTLmhuitQQgXc/J6jF7okVs0mKuEsNC6jFDr75xte6YNHqMXnFiqWoBrV1ywnfsjoxCyvCbV
wMAeRZ8fn8r0wtD2tndaBFP6Lf+ufBj2VI5f5q9B3e8D0+fyKRBdZZt4h32eq1nthFLI64MbZhtL
sOE7vjQMSWGJrNDE3lF/lYD+To5zEfDlH9QGa6UWagGrkbUURJp+SJ6Fqv91Io8fpW0TYH2zAzC2
TczSJNs5qTM+vIxUBCRmHKcKqdDbDgJhRURiX9I9hk8NXrhV9B3IKvq1Ez2kHgAwAwt11DqCX3yL
pVLFulC2xbcUfnrAszoaVU6iuLQAObB+mzG/52W8oUrzLnD4H9uX500f0y3v+guHf+xIpAkMMMtO
kXVXXlrDyHFQhBaUTYZ/NYsugaB0HoZMqaJqvPwvDIh90YDvRWMeVkOB98W/zkTKEkXSFoBtOIRt
XyWKPkjvuHVvsoevGyCZcHib7COZduFPZ3VRwDs8a32LJXztkbZj+EkcLZO6nT0iol6za+1E1LsI
QzFiZdk7hsL6W07TjGRuTfZGPntEHQ8UJkPhyowx/iEooiR7TxMzVEq1lhbBLoPvOMDH92YMeEun
XNQ7lOfux+967K7y8lVs5wMZcRR7QBw1ulhIeofL+yaZLSCo5S0L1mk3G2zcBjOXZDZ+FHdB/STX
UbxJNfM+GNgbABINE1j3PunY/ZCe1tCM+2dAo0WsG9xwL51Sk1PtpDY8/Jme6KsAVXQmBt9NRFCN
bh/8D6IM8EBM2QJURkRazeEb12XlRpk4OkGXc4rNhq4ri3MtjFdWCL6o5CmdfTM/LAmke5s2xjnM
PSSJlqF3Q1/2dKPDdsju+RhaF2Kwbo+9e5wfoBCzxaGc0+gXzOZ2afKDJxRzwLWhFbB/gLhIvd5I
3zoCR6elP6kovxZgXf98uQhfIjfj4UGr++EOhtSKC/qkPgF54IOK8Hzs/YBvQkHs7HXBtpyighaF
TZzspBkv0SpmWdgB9NxcaHa/OSdEwtjSm9s/yAEraX5sDtzhSh17eR+31V7A3R85jbhD3Jr+4mRI
g1/mhmlDVrmjiQLXde2oSqYxLnpuJ0o1J74Ds8qdNYj1AUGIkXVI9q3IgzxWDK7CU/0tsZ9Ca67Z
d9ECmRbRjOpX5HyaFjbddRafDrO14dCRd1p/BWbtoTcraMkfMgOit00OPvhI0hMoSfpmM+ZD3tBX
Y3gUQSp54k/nVLUMzG9/+bKSkUEMIDuWtfYvlEm/zcOx5lWeHw04mVHEnVCDXS7og2Aa1wBUhPyR
wq4WDZt3+G+tpVqHbONGh+plSwcESTl/Gpx1kB+l7udFyvafqOZ8a+sN2vVDBHf9zX5mqBtL14Ul
VXJ2UAyfm6J9LpogR9jrx44omxcwJkDbH8e2jm94cmm94vrSUa5PNNnLTfA3NMncMYQGadgrCcsY
hTMCG/BaqvWUMKiNW8WXy00qQJwUSxej/rkp3MbEb1bQYidR7LqvNHqjWtcmWhlztxLNHcPhhOIS
VyA0ZhQIBr2ugsl9LTVb78WfOqYG6SfYYwx6vJGXoXAed8Mu8+yYPXD5+L/cij1U9zhZQ39QQnc7
IF9xGxJrvOQiYgE0bOLJNtW6H7UFXRbASWCuusrT4j2lVZsL3vah9uNgzwtB484vbVmd6WrRANps
GcNTCrwiRaKiTv/anXeYCw8ZhN9JzSWE3GY103Llte0afkJ5hPY3BTZjEHiTRxm+2ra9SyDIF0jZ
gQgsJRGpg8f+lMdgCqj2sKnsLFGU0RUlzgn0uyo1nCjDFcSUUiPQIr2HBsUfQveH/0fGZXOk8XXJ
/I7QFH8VJ3JkxB4cx56Li3wVxAheSaBkDF9UYG3g58H8luwvfDWTvRCN28WQw3Q6Prkts4zqW92U
D9GDmeYomHyG8uoD4sVh5IzQCVa+j04zleJ9yR2hwUAEk5NbM/sBWFAwRhgR+gnul1rTDz4/yVwo
1LaKTbR0IqQvwP/T+YZdSTbPA2WjeG0Wy/Gtu2Dvqht2AT0V23r3+kpaOV5Y2FW2KGMTG5YYzXtN
2ev2J2nD22ePVF1jRG6YE9/OvoIeCfDZiT+xezRCrvDKUtswqxz5jJ0NIOGt6xB7JhOkeRp+5XEL
guSAtXEDD1CmxAF93dENcT3UEEWHfcbIASB2MCGkqyeN1nsa/9U3ZuUhuJKGeKkNptqAHwz9z7Qa
9WTZP7kLZDhw058k1iscmm/6KextsdZ5nFCaEsQMKuoeAOAfSg2dA4B5FUf7EFXaQSHSLCzDQcVL
6olcY9k8jktcmsyPpQLkXli6sOGIuI5NfesfOT9W11WuDE1jmxOyUAqwnv/1P1fxRzTmMrP6UX3B
Fx/J+j5YUJo+/vQsQELeMvYVoGvj2M4IJ6AuYnCVQcDs31qqCN9ka1jzziJD5oNtZ5VzeGM2zMC6
q2AwPOcIq1bjbKgECjdODsN0q1NNKc2YFZkBoJDGMz7mu01CLISolDMXyBxQpd6T9NPb17BUouOc
jxeap/6F3yJlSf3XkqYn7ioDzPs+aDStd6ONK1M0HUzt2N5a5R37/7q8QbBp0JyHymA9EOpXRi8q
JSfuQHwFCnAm6tY/jzsLilpfYGTV938TwrOUL2wvlq+ZD0REGkKCrERqNHlFQW76x1nnCFJxEXYc
/8JrslQ26fvu7EiLqqmC/HpNuZnDMsSeQJ6sU8HtZRNOV9N+JXz05zI/wvQz/fYArLcx4OgAH8Qb
dTy9g0o5eVVqu4Jp9vcx5ixAI8+RtXA8KXGUUnbcKGZhOtKYAywP77xMqk+H7Wy0H5R4FIKoxKLd
bDBR1OG2tMxly2ajD9xlSwvJ9o6i7FN8ZPVZET1p540qYevK5EPjEGvlcjIbUA2ezlZaKeq/YXE3
yvJfZnxILclky/8KJuoxMaNqZvb1bra+LUpevhEIf46FmwHjJjgDO6FZT9j0DGyYDq6F7m9mEI3y
yVXuB1fPK93CnpXWNMfGfSUhKFtAJTEYRx8DwaNaUmxV0jwp6J0jzwqeNHp2En+FiNbLAEwWoz/d
b1mbuVPbFNaY/tI8GqQv000Ew3I5Smmx4F88jW4mQdabwnCwO3me+a7qCZLhxC/nMulzdxdKMpTQ
JSW9d9zJQDKViya3n1HIw6BN01Z1bXumRtUn4/vafK2sst15NMVFMrmzar8V8ZqD8s5PbiWYyAYH
lDVry8naL7QJi7aXQeukVcHWJNJxbXfe0TTtmKP1SqjRFzmzMrL/WBS3gu3WjjPLVs4Oy0oZvy5B
c9olU7tGV+FquNDJC0YRpt+ephSICojBcq6HNaXqo24yIn8YnKjgQZVO27l0IKkKsZE3pE3cEd5C
8oLf66fA5RBeps1LgqD2F5hY6KCgXHbB6+qhQBuVKYQFXP6qHX7x49TpLVHflvuDgtmgzCxcBQw9
mogZqxfrH+B6oElrBBgywT8XU+p2e/cIAH58wiVN41beDBT/md+YWbEr0qVBxK5ZNrZzBfLGZ2oS
s3c6ba6ZqYduh0nrNCie8wK7iHkjxNvDFOBySBxR9GbytYiuPzPXDp1G9N9W5WLoPW+DVcG3PqNd
A3DeCFWlghqxatXo0JabQwQHthCgDMP4KIMVp9pJN99GYsthCFpjD+bUZKZjUzep8j8NKWs5eLQg
lH+lBT69Jc3tpRc554Qsla4unbiahoj1yZyftiYefXDqsLVOfZwxXjym1GGyUMNVSlnXvw4NAoIT
vyzCczjC803ZqpZy15rFxAJqo6+eLcB82Cfv9STIeZVzl7XV39rM3fS6Kz7sFflXlXTsIV0OogjW
NaL44l30PbfLvf/2arF050LiSGedLGxRvsGT3enln2E6w6H5WC2DKS45KHtcfxCstXVYYFNuD/DQ
7WDE4tlo72Koj+JJ3LksP/wSiFp4QzXT6W9zMVr++R3wHzlxZEhD+kn14Z4UNB+oH61/AZLnwiJG
EM/gVMa9mfdlrxQRzz2HorUH22Omiha0rdh92PWjs2UAYqJ6IgdKJ9EkGlQPjpP2bk+OJBvZggH3
BPHcQrm1E0+2vUsOoT9VSoV7AhIOuAORI5YGZ+ongA4WyWEHbhD3p+3YYd7QI5zh2KTb6O5EeRFa
6iaOZRY84yJ5kq0sfKbvNYrFeeadN6qKNd8UFQpAAMzxvrQ6ixa0sCZoqqlRGt+OilMTCOqpdYBp
v8Q/JRRToM8oP9G1O5Q497zgRvp5rhhIg6bigdavscHAc0w645J8Nb6gwcD0foBfNW3eANNQkIMP
98MK1rTBd/rxNElB4saEZCyJ8Hs9TlzB8G+gpM96rzmGGbR7HLfZypEyTYsRqgYPfjzqrZcJsp/R
BfvAqUQ76VxnCiC9AcpcwKXo2yJJGxDgLHxGi19hcsjBOBkXaZ9Q1T1R13MVJ+NtyYfzqi4mlL4C
MmKg6Xkh1cweAKKjQyICT4NK352ubFBdCnInTPSebSLRyavOi5k8rddECyc7gOkXfUmC/NzM2mvZ
KsmRv/1pk5K7dnjSTonqF0kQNAkyUg/Cn1msvYs55At2DmPNfsgVHVU5Mk3ha/L3ataURTKVRnK5
sSakl2oDqthFhS6rH+EAHKKNK2Pi0lGLay0j9uPeAttEVl7VEne1ow2x2tmA30nZtRKo/YWNGFky
acJZ6IGdB1Lt4BxjD2WJpJWvTHTEHzqEcO3SXmdHiPKZYSxQ0/8mB3lPBmThZWVXhpH8zbWel52c
iByToj0N9Vo7qgjNsir5VHtGkO5U5EQtTOEJaPuX/DZ0Uxt0mr8PVHl+D0oD4fxJE6bQySN7s2kq
3R8TpfAumE3+g5WXdN456HkaHCBX3grHk5otaxUuj36pfWCuoT6OESIoj2Tru9bz2zp53b6nrZ6J
Ek5oc7aV1188xB3x0v+tQVZAy0oLmEL29qgnE2gy+LOyKRiBoEuzQTceDsvOxQmMuE/n4rXpz0ZH
aypOKalR0WbX5DfQw5fbPN/dQ3BSR6Om/96067WfaycRDn0ejRcYrFp+PXL6ZeM4Q7+tFv4L68vu
odzYGrKzxEQrbhgsAuUePp590XhqRxmhbTpmPVtG10tS3jz3nSe3FTRUYPF11lHgj//OXi7LMoGc
Sl7We+w8bGG13aKhKTkkeP98JAqtRTtYcju+g//8tSQvYlyZibsGUFCQCGDFt1l0Q4eblr/j32Bt
x8s4IhduUQKTByv6wKpGx+3eO0IncY8Aj/eeDbDf9xJOGdZ39b/BrQsayblgW3CVNAJ8HZQ0mMpk
zzqOkzglTHh7c9aEgeJM0MhQkCaWxwVbKMUMUeAkkNntyEqc8cjAHHkWoB6eRlhz73/CMGYk0lvV
0L+s20HLq2zPPkPy6fNZrfLtEF0k9Ih+PbqSa67ruFNYr2YlmIwPJ7cKuCN7OCjA+eKckQCztOsw
tcAVhYYcVzoB2wFpvh9DP0JH31QFwsoUvd5sWhdeLjPLMyv0h1JQb1S5ZyKtCcB8PWNOFHzSGhkz
0Q4vHnbS1+aIcWz/ihCKvv8G22tnbaMLhNKGx+JcaQFh6+n8meKMpEDQXq40g3cfV6KkqTF3ohIt
QbAfZn8SvKRlYwd16VFzdJQCnYrFoC/AXgUmyfdCwhJFxgsEcn9te505DTIe3guCAaPy5f3DjxBF
e9bVj/us1FQ2rthHFoV/3rJm5J1Qfr9F8bJcBWA8rQrdeaB5UHZOYCgvTiO5uZe30NvWZfD3ZzIf
ZDj770rj68mG/iwk2UnGtRvp00JeX/rY8XDnblbwvL1tBHh2IJgpcpU2vkZNIPezjGTdqVwkNrNE
9gliJN+CIUh3XAcKxEIEfB2s7fwu/ffaYMNRtf6esZ/9szGKTjmbNtL2fGXEOljq2AlYnkiJ2371
8f3kr4ObzoEj8J1RJHa3vzxSJD4mQj5WfLNHneiDxzFmMFEJugzzXpXSBGRYvojHd5x+33sPDyHP
Rwc7EZV/1Bx61RPsDYqimZKmRQOvjXQjezCfaAtVFNlbvN06JGl95uTuPSrd1AXSTSxBspNGf8I4
xNRQIkvhbgWTQYXA7jrY9IaK4GCFO3AkF7M1T9NaUoUGcNTLg2eEF1aWl8U9cxajRvf6HLzKxCZb
h/QNDrq9o3j4E3ExAQxdNZ2waqaU++rcuzWO+ai2+z09pYDkHyIeCeUDe7KApr4+qSljVb4P13Cf
9d7BWLHC0+B7JYgKaTfo/BeZuDnPCQHDAKMmNssWbgP/vhUXb4odwkeBGrVKbEIZY/uZhBKVsYuA
4JUvwgASIAuEZJjAqITRO/DGCCz3UpKlxXC94ADrbYUZhVVQ2IeYnMbkrllW2On2v70In1ivIe+b
pm0LCpbLn77e36ByVwapOoLGbT+dMkn0tDXJIaQapdOry3HCBzzgUWzAezJGY3kfrGulMk+VtTCu
XjUiKz5KzZnTydKxh8/I8c3npTY0JElkz2W2naRPLaTeYo8PdivJgBL4SJvRDEVMIK7LUX8qBpKd
gjZS1iPcxCEtZhLlgBt3g4zSAyl4L/ocOswIrnJtTD8I8fXsgPuQb+CjDdtCgst6Kxfo9cpm0G0J
xV5tBtupl9WyblS8kldJM/p0wRlF+cgCn7nB76IXxuVXpw5irq3FlbpaAwukjVeS5wqwH76XNCyU
BFW9AnXrDLrcGGm8i21Rkq3NKc55z5y3Hi0gU7HFafGzOXNo7Nw961v9Smfg96nezNmIwOOYJI3t
NXfXBQP8B5HsAPCgf88539OYTCn2gmpfzpWUNhOtCSzm3EBE/mDLguksXxeXq4hG64w+zLivAhE5
2ShHcwvfan6o8hhgegqAXQmg/P0mgkb1ntg0rylEP5d1d4ZlJI5b4RRM9TmjFKg+VgU9vE6AUYcs
D8MLvLPd1zRWS/aAiBqNjMo+Qg8jhfAuiCPBOYEVg6tPi3RWNsDCgXEiFk83Estmm3lTHT8lCFXP
xIV8LL2w0iD2QRhP5mHz1j+Y2u/dqGj4tjbZAprWcTL0L84rpBogpcgyDCHKt0busXWlxlfwtB7b
JYqzIh3+JXZMhxe7yGIhqvQdjSdpW0LBVjc+JvpD02emyk4v1GZXXqpmYaPIf9FXWVGngNrf6Hcs
f/avNcJl86K8Up6k8mklQe5PGgNNBmAZLqSw7c4k0h6/MDtcwuyFN5ORsAgaG2gj2xGNBi/GaBoY
ZGDBCt/vaJyOAbbfAWjBRr0DtQMckadtfctWI7JEVN5/P0hGltC7mTtrrq6EHftZWtPAjav55y/x
uptQesAtjkPCSHrkhNuBVpvakiASiu4JYisUTpMmENfncCp3ffOVtkWBLWYocoy2ynLWK7ndnEBU
B7mMAloxo01rLtaExmabyE1Sz92/e3ocXaIqd7K2EFlrt+acf1dRFqsz+UdkFvRiwDSY5bGGoXAy
N6j5G5biVYh7j6WRiR5N7alh/UuraeNMfubWT1sonLNnSStXxcmUubN0KNZag1mwzyVe0KG4+a4m
MwSCSTrZ9CHjMdZpBAfYHMZIQjQPMP99+QDw54egNk0cf8ckGXPmBhkDSCUZCHiM7ijrW9lRzlnN
4sElWG8xx+Pv/VYbhJAQWunMV9Y4NLtYEMUoeqRt2QkeeLRuzIEVC9hlLH8rctQJLgxqVp2FrG4V
78/7xUoTTJjZll7JxuRIbZTLxwwhXC5R/Q/9bzWAT2u3I4fDeHdYO4PaEiWRLxli8K/g3niPawKL
04DNF5LKMB9922Hzlxel1V39igra5p/SFTygjKSG50kXFOqZXZr+NxbhPGbsjGEuWr+4ONV8xfYs
qvr2QlY3q7D6v8CiMDB23xEC4t88pU+CX//sIG4m5ZPFFxxGlL1f1sWo53ppVpXOmOoyLjXUE7M3
/aoWVKPXZ9F3q2QYMfewEAJlKvDLWdtv5eaa6tSuaPYifOA0s14LCp92tMjwbG3FyB9e6panNI0n
kdiiYP4gfGzzKtNz4Oa0Rm9cAhtSAz5qTnt5kngYlmV2BrRtTiukFOESKudsgDzx9clNY6Y/X3pr
GIm/WfgFqiIvSkRkx1OExtoDVAEF8gT3rdfbyiKvnBbCToyQrKqboB73HGhaeBV4PO31BpzLdbp1
AExXkDQkbJIWRjuxB6/vTi4Iw7XvX72Byf/9Yp6bd08N0iZ6BiHNHqthH+KnZSeYhI665rLgmh5g
Fuw88BkElu3b8viRPeZe8ERSUhNENc5XVm6OsrBBUCZe6T4P0ZhcVve6gum07u5111FXi8V0SGnr
8u+rS74bwcPWb1aJqTWWPftZYjsces8icVwSGTzhMT0VdZskZ7NsGR5ub5U0sY48ZxjSXeipkEdN
hsJJKlWiejyWXDjGOu9zR+ulzF+qvjUWxhADHRF1l9Roc5P4lGGd0apSgKjPwplVTway730aXZYJ
lTbNut7MnNJHHckaHkcj2MeBplBEbZSGxXWh03uSHXgUilwNGofYVa9fuyZGPW0QcFgjvOkTf2cj
TdQYAylr/HlnJprTC7+ltK1O7U4b0TjIYd0ITKrwWbPV7UoMwL6A/xWDvBl7qHOTTbaAKNS9FwhV
A/XjKMXQGWIzxBi+imB37gbMQBi7zsc8OaIiBFLdqODD0Z1qgGO2oTfVdwGIy0OnvLKtQkCDY6I4
KPBtzo9R58I/x4sSy1+s2qYDfvj/byF/Ht7UzP/CwqvXo0mouGMDRAuPbvz5hgPSNizIRnALF/oN
tyrQh+Pr02IoOGQAj5VjWDXiAZPVzXz+7vD20ybcrrS/+AygTEcO2kEasoKHkt0nZj/3yn36600a
BgHdu0Palpk+UJwGTY1vMDxETnQtEHLBydKYKTVoLIen2utZozeWs3d66cyxydoUancG4IAOHu7l
26FmXBqXzfqjJRMqwVh+YAIH1X8hLADjS4o1Fg85KRSNYsBpWMJp/25ExpczyqQ/jcjtVK04oUin
kfMesbGSJnXu8XsWjX8rWimjUBPwZ/UXqT/PB7t4PEw5yqBb5Mu8H/4MQgHTe/f/hymE+Ge27gog
xEanwy3on13sw5bxS+KPShQFg+l8mZ3dVG2ZcXYyLPk5dsiIPdYTlkfvgnKhF38b+cKbWGSNvkZ5
lYmSdQ0cTNqy8ojE9RXmg9JVni78z7yXGfLJKy1zSxdemd1LhkITFDhq7nNf15fDzX+i7/Zs/kbW
obbw+9NU0oRXpAz+K3JF047d6Ei4zdNXvQCdJd/mC9Z58mQRKqpthYtHSXmXSKn3A3yR44Ouw1Fh
VNcV8PV8CtBouTo9zMi6FhxHwrTZq7lT/gwI8huQVABcPNr4A0JRnfUo6NjbybGMYi+oJ/ZuPGPw
kzPUgMSNjd2fwApNqMJUQUUXcV2meJDiPn8+HDjHiSvElhG0spU1IJYjQ7axeF+5JGRHusAIuB7O
U3IsDBf9JD/tIHqMs0mr0T4rWcU2+N2t9mmgAHj6tROHNBNXPkL9/9MiB5mE9JysR26Mh+XjJ3Yy
8HrzKhQTlvnBGoBIGx0szolhZz8+UUW6cQxtuws1L75gE7Yvf/ZVM50UDtu5DXZB8GYsyk/new7/
DYeLnut84HoQ8DO1NwODjaIm4giBF45IXJxuy7oawZHFqY3iBfGwd+ZPc1ScQoLg/ZWi1ByRctZt
b0pbkuU+gsNLVCv4Qz8qzTil3lVkaRIo5Pgk5duu/FT1sDxTPQadgExres/5m/omskW/lo0HSPE5
LL9E7QhhT4LtvjGOyTGdqdtAZM+fAlSpMjHruX6BRAZ8YWUEq9rIBfl7qHvHHtxjcc2ibs4jWJUF
CDZvgKNZ7hEENIEQm9L0+Wtgj4aB6AsOwU/jhuMKaqUaH4ouSfS7flbd/KTYkjL3SlvE7aaOhU5u
owKcITc9xJr43OmFY+TIinMhVMSW8axpyWtn/jeJucJWOHzpOkVaUJtj1BrmbVURTUoNXZgkykN5
eUb60xFgODwPHJN/UNeRU4ycS+tWR/DfcNVgNyzTsnNw1/XN0Sq8gu1bQGLEjezpsDGkq0LPa5Ga
NIp/Q4r5HnAEtxZcZ6ION/HIC/1iI34OFrvF7M9eGyMhUfeS3FlQSfGU0PJD6SLYfsXMOO6oGJck
l7rya02zcSbb91lelLQGFgnAfWWVgUQ6KFhe0tJaE8Fpfj26z3g21vscj+FOdNpUItebf+3WggJm
0g1S8F0cF08v9kiWJmS3wLL8IETCBHlHqTtiMmLlSqIJHDbDZo9XRJ5jirlAU3gxIHWL8FqY9E0f
oYOQcIUj73B7WEBuwehT0hgplTteulLlI8KDz5y12KsMxhPi7wPm61O/rUxIHz9oAyi3BArXahL4
YAqor+MZHMZpcPYgxvBCMBRMsUT9SUBC9lkJL5c3VHzcPzMWnH8zEpyhxD8Gw7cCGDD69wy2wZqW
e9AKh4roCGfgaGxe3wyZllXqflZuRDzFYFd45p0n+DnWiDUrb0EUMCj5RzSiRjjn/A1ALz5vyH9z
5uixuQ3wIM94NmQU1et4HZXfEMLjJF1FUZ5XqMvXytEGDtbMWLKZuOx4NCv9JE8ROcwNjOrJtMoX
FW6MvkMaYwtVCyux+6X2cUOHKnIEY6zVqTKuimf3YPFu7fPQwS9ByogitLw8qAxSztDqLWlXvt3s
3fvoLSmbbZkB33l/6DlRbFJutJzml3zCE2yp4FlNat/Vz4U/xGk42Cd+lEZkFjqTLyUXf4jslJdF
f65qfIHfNq9khvfI0qLJD+Rfy0koup2VZ6GVAAva8Ka1wsCUQDUqlUwVRVZVLwBMwFG7/AFBijto
2nZ2E30YSHbdT4bwXMKnk39aARzzZg1SGrKcp6h3IJVgGJCxyrRlEh5DF0XTQ+rGfdwt/aDexGw7
mTseQ5CbMujos3xBlME6Zk0cqgUw8+4MaU+057/EWk5LggRJOIsbBphmJWTwQ5PWxCxCPLtTTqbf
5r2TbXyKdjm+7/q55m7sBX6EObe/DAGC2t4itfx/Ayb1uVYzI+N7T9MEA2FcNDBK3MPbfSPSwyLs
boiNBRm1GDbEp95kf4fRDLos2Zs3HCoIkAR5VLd9UuT7copFAU2vaAgSCirzbn4Ol6Jsw80NqPJS
vWH4j0/kRdBWYFRTt0oTCkkWer/uieU+H5qBON85F3m3YsbwbeSVkHYjTBJM2ZpcEGIAnuo4VCId
IVRH+b0cjoWlS1eA1xGBEfBKNUeXzPadKBmc0NcSQyZCYhMbGCW9pHi+FVvxSdqNLQY8GtN5j5kv
wbsBlhAFwtT8bPvcJFKsSNbfh5oVblXRlESeCG+howKZCzQ0dzTPVEv58eEcoVZiwspjDGAoAqAO
bq4gjPZ1O11WE1QRpUfwhdmCEYj/0zq0JMdoKR1hs7nrL9Mf3TQGQfUYWqYumRuuLBgcGvpHfbID
f3ph/qlQjqjja4mNMS7UAo88fDQmiJer9aNoGGiES0BedWAMkoJPqLOxAR29wSj3r8ND63RQY+8s
Xg4vhzcVg/R5OOUtw9ddCHWS6p9b+QOLoY/TKKI96Flnuc1PVEnoybdH9W/BggpgxDmLBPFjRpye
6LvWJT7tLgcjTV9pXXDlZUJ9dLnwG31NbS3FAVllO4ga2IZtLvBOC/wlKDuIpuFAGf9A2+HxhJ0c
b24VVYqlZNpaFpir+9cbarm/ZtlT5cQW0efeEZ0HmUJZlfVAHLfEbKY+/BM3W6EIxPrBGDaBAuHB
cvluAWI8Y0Tb6tctMKI/A3Oj4DhIPSKdFzvbCPOQCG5AG8YP/sZWp5FqtIVhbRry2OBhGvL8pCYx
OmIXIy/BfQRDM3Djgf+wOxojJKfpn9bRqSuHD1XA2qlAuNc1j/hPgXgborJwbySt4pXrm40sSRKO
zcgfNDwHtCFw49HCUDzYsaNahG9WtGyzwVQVh8o/3ALvkgu2qIV2Q1Qvwoc+nGjWCTB8SlAP6WaE
M24g4f62iNcoKBGtAcouL1vmU9GaRZxNNcq62delYo3ndZjGJ12NgC2vxCh7Y38DBxVU5t5g9vdy
e96P0USzG85qyJLShtqAAwAQogPbedAcNWdPFGh0IoxMC06+apBF8qsBTU/1XExjdiSJ0FehJ1uc
6aGois6cZe5MosqJtn3P3FwOnfaz97H0nOobfAJ8TTFiPZGNnW3Shi0ZBE/DXbMGtsav3kIiEinp
CHKce8zlV+mnmFlx6xrLMNJsjlEYBIv8imvmOramxBrzChMPt2bBI/khLFJvRqgjPcDr2eXfm3J3
yEBgSfiY1wRM+KvD/S3JQYKzIHO1Qa2m6PXq3Hy5qxMhWUhKzfbIU8pJtieqqX+zzPQUO6TzSJDW
yRRulgnSqzYdXBplWjwx5JpTZg7eNBmcsjwv4MMl5qvttAD/KPLiFvJSQ2DFf7NTrvW8+QCXALgQ
F2tPDzLpdpx/ZW7JZBvSDBwD+rPHEA52YgM1zkMn/GpLEcsBmgdIwhKQEzjg6Qq5j4vzgYu0OV2u
QQnjyi0/jDEpIovVQbzfPCh7tkBJ7zBSlJXljF0OQAFe8phDVdDIJoFKlEfW0WQNidGLaP69NwAZ
dBlTdX431ju7/7nrHQq1uD5t9wfJaSwqRAFhkCHfQa3Cp87gsUGygDBhGHQBWwSSBm+C39Sh6WoT
EqwBH/w8/j5kAREEDB4HScdyMqG53zlcxJFMAoH+KHAZmcWE//qibak3NsSBYI/P/MZSFjFKS8s2
noPSv/thOlFgqPw9QoCytWCKSqH2O9PYdevaV6AH3qCGXhaaBc/Mme0R0TE2WvN5UYtbDSjU52PU
IXHhIjBCS6Bt00cPLJeKFVa/vnXOBsbNFq1EqTLAShKpB7Y9ESWTgaJ6vgO9rfMLq2pUQpuo/WFB
VDaSHJRgE/wuzDj9+dBlrECenNY+1YUx0B6SuwdsKt0itDCot9iZdFJqU55jXEvmF5NJYxgHXi6x
+J8HHLavYuptG6dGVaqFiqgLRSOhEn0kqqo6n5JH77HN1SIExXaxrjLs9RcMtusgZjWYafiP6AUV
tOMZfKGJ4IdAv9LrO/BwKbkxTiBtNwc5R6Sspo7Xew+wMHZGw3urN8xtaOOf4tnNvkkFWiIY/wV5
JLz6rwMeHhSQOXUBjteTHAPZbztCkYbBQtJ13JR1kRVQXOCfvRd9EKvBEvmJrc7TjLY67RhCYvKk
41DIKSCxHUVnR4EukSfjwmanQUdNqMCstdqPT8Nl4Hf4FtRIQIb70D98NRed1dwmeZ8K6M30p4k5
7oeJTTQWFao14Tp8beaij9VGe6OFvzshzQFXaCm8LG0tqxbTfcirF1cUklHzVld0VF2y+47FrZew
ES6bqNtIoDKnIM+1pjp3bfwYHmtRrcVO/WUz5p/mVYHJPTFijbo0N3Ij/tKAVHSu+7YueEc0MHGV
siSo1l3yp9nL0bxK2sW/VPJ0iUa9A3w65Je5Ol6F2iLUE3tsbn8ZPliQTnFQjdTchwjZ86bxxLAo
p3M13YadfnCHaPEOhiaxPP1VPkwqsI0LuBkOzbmdQAANSReWsIWNlhvZIuRYW5Rk6BLODvGOFf0F
sRfDv71PGl4ye7zEDxZqT40z/Lw58getKX8NnIvqAOfOexoUCnP2MZX/KmYwwGvTm7nAhkR/RaE1
Vbz1JJO4lONbVMcmgqEOyL8FKpKbSQ/ZazwzN84uGkbFPV6nCWleuFblbgfzxI16QumE5PV37J93
ap8uglAmtxCYlxy5lBfhfjBjIWAVSO66ps9c0gPEN8H27X4s3ozimZUyBN1DcX0bhIVoL/bo5313
c0J5ViUOsJJDd2L8toQPWhoWQhDbL3xv8ES2dQRY7/YwrwB8JyGXuOMjjaWI66cm0LAu9ujXPjbE
YqYkA3qnAWSoNEisigUqXjwNpqlSVwBKFHc+et/cLDopHsOptyoVPMr3ARwAln2hRUWiuwPo4GeH
RkABrbc6aSynrm2oDx9e96sOMfcCXdwZpXkL3c/kaOry6Jgmtp3ar62c6Db6PQAC2FsdhONqf9dP
8uSF3UZ7z/W5Qw==
`protect end_protected

