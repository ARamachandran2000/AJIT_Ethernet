

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hYn4T1Tz8lmB8loeGYuHmgEJp5TdMkRKn5tdK0Pxo3wkkBR/aG2es4RXT0Kx9IkGgy2jVWVPoeKB
usRl+M6Pxw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZOTsELKZdXMGraSgAw9rgqxvSLbW0aT2lTeYBbmmRdIiILVX40Q3XF89sXvrmWq2q7dAJSXvpsX
1JIpxbCUMi40Nuru7hdg9WkNNMs1Q8UJCou9g/GNLxJnh56Wx2JqOiplBqlgeaLjd0T16sGmIYm4
kTNGsNPOASR/dWaldsE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o6ehD67QiTZFs1auOjL5nkbDEbn3neiXmbyTqqoQKK+v0TaPL6hSxGHE/Fz3NtmR3RIza9+Y9rVH
Je7RNuyq8vsgofAGK5Qpf28P/9kF6eDh0JgLJHOonk7lnG+gufS3pMHIfioCEe/2wyoIxzbwUPNl
TCIJtbzDvWpcCIKBgiQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cASOe3RHelXhU6s/jEEqAnadTjmj4ihjbMuYb8YjKT8lAROht6xaHEt/3WXUlUPXIpDwtJlexClV
csQVUSlNShzZmxBI5epxH/HJqLhQYwkRDFK2BUAagxn++cS1iWJGlow9Gha0EU+PfllVje3OWy4O
LbiqHgQlEG6sIGo0ZCj6KPC87SBAytHtAiVRpovpGAxLS/DLeXSJaavSSwOc7nmWFDaNEi9dJS9i
qixZxDI5QNaDp3uaBFLzKqo9oSPgNj1mYKRZp6XL0ganfqQCHh/snCyymi+o0DC5vSM/+RtCZHXA
A1u3UsiXv/IfegAneXJ/yU2Rpj4P9iaLKgmtjQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kAlIhoAHksCGo5mF85FXcP0dM1NExLuDn6ZkyfgoWH09b5qcw8bLJnQMlkLvdLRrczznUPKBLrRR
nUHSMi9UTzRZ0rrnazgGnHFEV1vyoRgDQDOpkZbrkgl/VynbkoMBhCQXYT59yyHhqjI6WeIYVipR
zyn+NdmUB+/GwlsSYygywX31rotvUxb4RZmCqg+UCemw+N0tS43QuIzJuG1JM+3+SVbU3LuVcClf
rOwWqAFHsOXBSrXNoPX6QeNlYUKy8gcjiaQqPSrbrSJWdgvqshdNnvLWuzkREOLY43TCoAFwM8p5
73h2VUHmwffIqzCELbp3Tee5sQXgMbvJ+Mbfpg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CFQ8408huN9E8h2/r246qkePkogHtf4rd5gf8GO4NiUzetOQ2my8cbvxYBjZy3yQSw0/LrN95Drj
cc3uAe9r+wOvBQ3aM7AKnKpRkAvmqyCRt8lkW5NRi37udLv8jQJ5gVByTJ76KIn8s2kfj/iHou8+
VyK641fcvp2Fk/dmC13HALsHzGvO1m9Kg3zHT1aJxtdh2FDGLhOy/TtcAEbSWUhNkclp4pw4r97T
urhhIiarPZZDEkAXG1Ezi9I9ebmvdHMRRa/e9P95Xg7vwS04EHfmVTpFKF7UHncoI46I8za8vjyZ
8MCKLS5zKbgCU1OCJ9lQ6mJX1roD79pJrnKYpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
1n/5t2pelRZWsUdvtJv6lChe2nX2wPcRXZ5S2/N51Ud6r+47LHmlMJKInVOJwL6fXpfWoB8W6VHr
2osqNgq07mjgq8Ug8hYpGPbbI51vzHPQNp5BfNcf8p95X2RknhE70ZDuJxy0568OF8NNyLmfzRux
bxc7CDIQpve74anAaXaHDqBoda8XPzTRfvO3ISLm478RK3laC1EuwLGjOn6RPcApfrXlxBtsIOVK
qRVo2NDY+BtpNp0Jyp8sjRmMrYhP8Da/tUZzYvlG9Z0fX/jP6jDDS3DSnu6LMkaUnwPizJ57WLF6
hYlFyRQRpKB5iGrNXhUfoyBvFacA1ltDHihcAZbOh8Vm+fh9yhc4oiw30Yz0WBKZcQpuGo/FeUAd
Kj2YIJyxYOcVinR1UxtrFyObwmzVhkVTVJ8eBF5yie1XFSHhjDzla/GeVdY59uRcuZII9Nc5s5Pf
0ZKHMIavt5D4x9RF8+WB2j1OpvZF2VFbd1hlnySUhq5UHp+beDg6llAWkPfEyQjn/7SlGVHhFM5z
UPwiDRiSOW2c6DKEOy/nhsZnufCF3wYmv0Y1YWO+ImUDyN9Lrgs2dEVpVUjSl/BobzcB1FB77MwL
HU2fWJG4ZCpQUlhhs4lMhiS62G0pjMjuq1otwRhX4BjFIx3PxUYy7fwblrt9rF6K4kslTRr0mk7k
UabF/6rqpiTX7yGxUKkxqr20QzW/PQaHCnrdU2GGc4lnlgEsHgEqdt5egOfuZjAA/hZhnLLAhe1X
NMlGvYpEMp5ttw5nK/KiqNME31llmMmFdrQ8sOgh+L/sdhkbsMc0tpiiKhgqkidxLJxX6TMY5cif
XcvdoXS7xTSGg187CL89pi2g2KywkpVLu6ltTMq53hMy2JDg9Yu6uf84aSLLfRDIcsqBtCGMdh/E
UgBZv4tti8psDLFFKXZwmgGiZH6tmLzC2obCHty7aK25yF76dNst/JQ7pgk1kho35mPk5XB8ELzh
Qp49HXIk40hHhKdFgtkqBSbO2P3DXhOD0skBnaiCeXY4Z2zT1eLUgl0d8OG1SQA8z8bjWmdEPrjV
G9N4LMo+X1FwRi9kjWFNtPegQByQWcrGy74pNoEyGP/3EwSzsHYexJTtPyEWViV2moZ4dpFl/74C
vAijqNhLwY6erhg8ztMZnYK2HWfzZFMFq//iB0zMAkpFVv4PgVKD3EjbBn7LaeDQWYYcnaWEbYBI
gvyu0aJJfsX+qUs59QBZwvmfK6zHNC77b9ApLlUifZpAA4gEwLHJ9Teb3BpsMtPZaaw0aaVmWbQ9
z8A9RZNElzLe9Y+8li7Jo+jm45ayxZustB/1Kk0M8EoJ4JuK4cfEa8JyJJKVFo0PmkLp7X6hAL0Q
ouiLYP5KaZX1M+/R/fAL+eVJw8nsXimOZ7vQTtryLBYNNw6vaa1zGVi5Bajsl0wmz3EM9BSIqqzN
clDObAANI3xNvzHW8wy7Y7pUZc2olN9gMUrBlyUIMcf2Yi/LBZ7I83kNdXzxbz+Dyc68ku0aOsIK
Rs2BXqPMEU1G8d6JqG3c4LLb0aXxROd5Ch/1ql7LX1j8KMLHsQenzuMtuE8F2I0p1Z+nlDgR7XJw
3ORgIIVcFXRCgHCW+lVbEQHcQRvYPwk5lVWw67iIkDZMbvSj1RLh2AHVtAjJtiViIq28RNZ7B1re
bl7pHFGx8p0L4YP/PbLS+JONwEBunoflk4SHWrqjVa7iP5wOIGW6dTiJtmdzyJ7BiBXGHellZcyz
ORJ5XTgH0iltAATRN/ebnST00KjnLByEx8U29K/nVYjI7Ezzs+S/ctH6pfoUMzT6u7mfG7yC8bAE
NDRyncx7FNVtlOV2qcK+s4Hsp/Qtg7soi1B2WxOUIYnp+yGG1R6VlFlYbkkoa9JtdrEbBYdGqeno
59KMDojatEG0moLO2qCqJap5jt9/x1fFJ/UCM+4tCGaurECj+wDG7VxieaE8W5e3OBEQqTTpp8ft
3J4f+JT880PtUr8Vqv051Zs/E5cPHodcs3weA6B6vbm1bAm0uxCTAQzp47NV34HAGcew3QVYcOZ5
7LbH7qI4AGZRDYZRCoYp623WCG83qhTmzojAm56ImekzuimvJoqg9xuOMXzJbzinexhjVFQH8/KT
ZFU4rWG940C33eHcZQql43xN9CiNtyH7aA5FwSjHxtiQhSBcm8SyGFIuXaSjRk31MGGw2lUBqxzB
kDd/+rEGNwutzoa9qU4HnuWuihd9nyfVLVaAEyiUlJ3fBrl0fao8qXYrzpsoSn1fAdp/4tlRVMHW
Y2RvpK2XPfTBq+9b2Q3ZILUYyCB/SUQ3BJjFvRWQ54azNSijf6haFvyp5air5Z5q6W5Ems7F0Tof
O4aE3v7x0JxDbrT6G8f+AfEFCq7C8bqt01z3gd/k4EYmNfHOGK7yMvkC/V4wPDIYsKKcoPLoTiV1
z67i8MyZpWvLty4h8hUx/HPauUzslQDOclOitY32/5nXVzSuXU54nsEJ8acIEUAJHrxDpRIy2AMt
uC+wY8xBd9WZyYiS/LOa/uQ67GgHWOZtKUAp60lYq4NuE6KTnxHtW6YytFJ+1kwiIAjigIX5Ukyx
4jo3vfvomjz/MnjT2hAr0sWDsnHgwF0qAxjgUKikFZ+/Ct9a1kv2N1u7qUEsNzi3DAidujSWdG5E
eTGgF7xvSyDhD+DWo4drMUjdt5Ev73AyAHnuAYY2Js7Bhq+npdmBvDuIYzVZCu4CksQEFnXMKHWN
LdaTWrCrByHrZ5e7RN1b6tEC2vxHh+xCzCvzVSvN6uQRxwOHgqj1A6QhrAFgur3l0NA883GzMJKu
fAcRqh/42Ra+LJbwSAfX0e41YVe9P9WR8XUK3S/T1svvpcLzgssnS9kewTMyws8JIKzqG/wpovlg
ctlixOqyD5Ps7e4R3dgryIEMjBG+ZnoZikUKdUz3Kc4zq3okGwFnbvIRJKbdhdw5ALGGSRJ+J/xS
fAiMCohgcd+Ro5Eg1BiuUtRfXqu4xfCSHcNujbWyho82TY89TaEcEK0fgNId7z/M5j7koCbtPcHp
liWbOQtaHJ64htj4/Dr2xVPBmIwDjLbt5NKqpevjT1XF4nPiYsg5DRWDrkIP5Pl8lLdpfwJGhLHh
GDWdS6CYnRytQWjYZ2cNh2gDMRIh4DPrwQv7QxWFrfVQqotcLEExPdbFLYZf1gVDtI9CooBOsNMU
Kjm56/Bwiyit4JGMIOyTyQ+CePVkfbfaxfOq2N/5Mc2GDnrKm9vY4FuCePSWGck+ZVUEWNVhYls/
Nl57NhVVNpzDO+GOHTwQEGWUPbCFKVLGSbcyuCLxub3IijnadLxAw1d5mNsSQ06UH37FDDocxOb6
SYxbyQ6S3BFzR95nZTaNajvUYFf+3eZv8MfIyRYefOyY3YfEjS62iNOcAmY//cd8F24NQnpAonKB
w/T8LXsMTgJRZSTKZ3ohhtrp1LY1bg3BDd3CV8QN7Fu0Ahz9kOmy8l8HCoIyYUGh2Tseg8tYKxSF
tONpLdlJvEfWMpjgiilFCbDGelBMDcO3LkfOUUHuXYa27dTw1p4wC4jnPVHfpolkL2xTW9fPeB8G
WGbhLb3UFrDr+uHkX6tEsDTdS+B3hLGlGJkFpyXVQrUUklH3QK0BWkNCHBrdjPeoUvKB5L0FlKJi
+w8vQT7aqyv77AnwcPFvmrtYhIGMJ4XfKA38XXtqnBI7OcLRGWfsPTeXr49KUX9FxP1jSE+XvKmI
MRBsdlr10yh/pAJgmdxrm35Y3Do44BpSc79Ey+cbBz9py0p+Z+SUPq4Ox0QQExPSBpeGuHihXWzb
LODAgW3Ibjc4AnIhQoaD8NmQnY3i1cv6b4pMp5y63nuUqPyRuXYrD+/UXlMDBU31T2FiV7i4flAb
VXleuH1xhfh/Z5AoTnF43oWoAbRHSCh00bbNhx3VC8XPtSCxWW1Kr/T9Hel3pHRM+KICldir1Udb
+p/zlcwiH9zNosdah5MCuvpQ4LEFh8LLIAX5M/NmwF0Apt2x8miZp48WWpDquku48mxMMCevX5z8
YRnEkFvcuttxvD+oInoXC1yYASFf67S9BSWZJY6U9ceMIEghFtIAuXmt7zgKqsQuF7ZFo8aMlVhp
CaQJCw7bOyR9SYw1YHGAYzxx3Na/PNqZ/NhGelKaQ3nza2btXW/feV7SZJ15INoOobyTaFTmgWr4
W1cXpxs0aLKtZGbzcimOJSw9wbhVZdcqwk9sw70pWbRfwmraJBkAn2J42J/BFfh5CKRF+rP1DABd
ZVps+odvm50XrddYNH2kYSu+Mh68/iwk+sa+JW0+gmkm/MepQK7dfJJWh/XCusRuSpeqRzTEfQhy
8mahOnuFHcVAyFT3lXu1RIkOCKAwMO2md3R6dLoCBRul0XnIyREKiCI4U62PWAM6u+4KnKbrKwtC
c5m/VsR1LfELOWUT4r7ti1sggecy+xWVI0lCePgq4sRfoUoTcsAJJNmSDBxpmi4tc3uUQf++LhL8
sxhF/m8YRQByoy9HytYZ0c8nar6diAHlxTj/i24KiRDXQ9NvOfBWYjvnj6kjvcS58khOeek7hPQD
yWBlK1lgGwPrnfKFrFpxxxajNonoPlVIdMHsl+lwDbRJKpYCgSLecHK2aSbEGZQP65fQI4HvCpNl
XbzR6AEcRHOSsVh7fmRHUn8dYwxAoBFDSpUW7kih9RRBEAiLREMsAXs1n51PuFayghmjUWYCM6tr
1c7NuI2uTvLa9EEJUkf+XzxV7BAY0QmciWBS+jjpEqhHBMGCM0+ubHsOXzQJXiMdwDnBPSxjAKbv
QasGrnhVb+6aQg5rTfD1rp7wsaEQJJP8gks9hq/3MEvk2S8FunSVJpUjF+p/PlX95Dxj5/WIT6Dj
vaDGOMdfPo2HKKKGNSqz6AKPzJ2BwSpcsxHFk+2mF+kQivLHJ0G8xNaSpScgcMcScIOSa3dCH2na
fweb3FDiHMBgDKggy45YhCcmYL0P16QclcdHahTfuqJ4xNquVlM5StJ/NuNEIl1ZBxWzV4PM0N+P
bOJtnT46b04DxGtkSqTZEmWlAjpiFL9B9NRPSRSqFxKxj/ExLZ7bGh7WS9w0iGKdTO7tFNG+DL3U
a4FHucSNqGAHpkqxPnayLfdBk1scOG/KPqdcJZvgG2efx2/lMUsu1dc2bCtNii0WlHEboyNzeGgi
LHEsa71A/U9TtGwP5CYL7GAsGlco48Jvf5b/1yJyRbm6aPqBX36RD+gpPnwJmKlMiPzEn4y6K+To
pMHOtZCWRtPYnr8n99U2qv3kDqTd4iebKyr2PbfxH0LrSJwOA6cfx5YBJI1FbFjkLYRzXA+pOJ7I
DsY0w9s5L4PEUPrJ7GRzb2UezkT0UfVb6Zb/GlO5kZ1FmO5M7ht9ebDKGoC+AJICU+UHyNYufSPI
h8j32oYPb+6ulVBwTSEGbvB53IQ9oSUf5bwrPUpZhCI+hhaz2XmCZw0pKYX+e0zTv8A/BwKJ8nHd
L4tbhHj8qNuqCRjVgUCGlwOyAW/yKmfO7gOJsvj4T/0xxCEboTWluLCA/5pSyOYAzamLuP5vqkxx
IoXSfF3d+IvC9OkhYaqXBRrmubb9sIzgSoOdGlLRe9ARmEplGG54R5FjG65KKt5Io35cxWggNucR
ieS0MhqTfWZVZ2tHIWLF0t7lrrrxrkiljB9DjXoGEuPovC7SBCl/+YpXQ3gO9ky8/ca9mULU+JUn
r0Ph2agM7C/I66u6DKawprqk8H3eYsd0hgiX5QQCsGsFU+mrZ5YpnAGKPHgM5L4SsH6moZTedNpc
7EbDcrupNCFEbb0N+cV1xMFKXCoD47a2fr6hG71brrByfL0bu59ZyN921kAx1uSuh4U+hZithMa+
Lnnq6TR2m3g9IOxjfKif5M8FjloWuBkyOKMsTVZ5Hmr49IrFcvb70vbrTmqgIxoWN2nwy11QEtXu
4mZEQOwGdL11Gdw2X/TyCkUHMWi5/4ztPg4atPx+JTWtA/oMYXKshTSo06W2JADfk82f6Sc0rtzu
qUO5j3bMd17+AJAfSZaR4G5ce3ta5sURXAHDAu25G6AOZY36uCrgfTyFET2QkMGnSxGC3KOg7Fpp
pzGs+JE3+o0mVRD4yJ2fDsfq7mJAPsxCInf7/jvbISTzYQR9X+rXfNWjNBKT47sC8hfB64UzuIx8
t7ttT9al8xZv0h5Hqzb0wv2s0DD4Agf+FaE/pqy69kKJzepElSkt5APvwLjJxUHw9bx9kV85ig+4
XoNkP/w6hEvOSZlB+bhOe/UG7Xum2QDaoK7FOSGPJpb+6cTCFf+bRLFEohwLe1fHEAYUotLNeRnu
9BB7YKagDsvr2NbwwdzgZUKxCoNPWxW6nXGwnbXyEl+qChEhsGUVEiwadMu2XITDW4mG/iJVYduT
UO+ltSdnrFTOdYJo+1EC06tvf6M9wHEBtWwB53X1nY3qAxONRbbQy1GY8BkjnlbOdRIc6m1GR2DH
c6QUezRpv5YmBv+kIiSc6DvcwB+pOvOSob2gLJ3xW9CpNPmHFnKHOeojGb6KLKOSzPPGz6Trfa+A
iYD4jmW9MfzVD7aQ7HeRKH7P4KO1TYpZyHdqEv/di3Qf2mJPifZFVQdbdsn+UhbXYVJHJp5nmkUe
lvK/qrG5ELHYHNOglrHAuJf4MIOimJYyc5hyNmPtEvpOEv9upUmPWisZ1FfN4oNowF6cuWaDuhxM
46LP6ccGNQiCWeUBJ7iSuVcbZSmrcmHOeTgjV8VuGDGxDXdw90Iqh+P36p/AcptRFoxoiNgAZJAc
eWZSuHjqUyk8kQo9TTv+llLq75CBpg2guVdlMH5/wBmtTaZ7vaODuPtmtDcuNm2FpSxmUywqWoUF
RoLWHEm9tUD+4u2hHontss/b/TfHO5Wkr/ZbJ0HTRC69HOaWvvgugVqL0uEsH7IgFh5dsW8w9aAp
yV6bHIenT5eoTIbuONtiQbWD52dlCK94GY17ZGVgq9R/avKhxxl1esUEEnQUl0lzNb7BCIL9cnY4
I//xDRSGevy2I2KooHRWT29m03xWVH72WzVEh8Ig9a+nbNNqMKOxxONfO9ScUcomvwRnyHOwk2g0
h7U22Rn67yBE8pbrLie6QCMQhYjXCFPJkNpQNjZnybqU8Mkh2XqmpJ2yV5uf8TPIChUj2Xa2IzIB
D7Q1sOZUhs6syDxlogqAN/mWY0Wqjz0B8a5SMwa/kqCcnpphRa5P08nZSWMJygWhKY/UrF7iUPXq
kUKchMc9CjAx82X0gDR7qtvmdOtZpJVsnIFWn0TV8UrKQ6hkFhZxRLMswOhbFuXcKCMUa9RKhB3q
QdfMFVYL9e5RhnssgATx16wTKZPeJDt0zz1jjNfO+2EqoTC2R+21yCy8cvolGdeqyIxncxcdRBAl
NwuvH5WHOxqSt9/j0ZWFJ0qBmmzGbheSKeno2OosG8OKpnNgeL7g14aQ3YlK7IPGuLHWpEy8fvkn
vUTz4hQvN6csTebGVYUEE5iEJ6ZylJPzQgRqyouLqYV5SrnsFJ+4zhpHii8RMqmsJA29OtFKQEWn
FLi4HVTKAci95sBJihFDBZPsmngLISZPfhqkhQ1HFPhx+4Dps8LImhtkfq22g1OMMqHMC0eJqHXJ
rjuXcvYNVOx5rZLxGx795SwERmNaoT+hQP9uJXSeM7JGbf+e5fdXddU924/H/qGTrlQmOcXPaocY
K6WiLlb0Dk/RvA8U2+eO9Wg4lEQDfF73PD3zFVSAkDUjz7bPAMhMtD5Bq4hfgVrjH5AWUZ/gJiOd
L9pGMxHggn7J9hq8jml9CJrBGAyK6LBPqkgc6E8jiKiqvTtWMjCgJVEIxebkVhuMwpcjXCB9To7H
gmVmV7OZ8127SflfGO/NgvnTBaqKlBv/dNKurUkx3uNNByQtdi6QjkbpPHHCbNsPxjHd9P28Vm6e
vbIxAzZSlaaeFqVeGRScF9y6FoEEfqY7uQcT2CCYO6X20gsaCc0INXUSqQ578462BJpf4hX5Y9xe
Q4RCWVIhCJIdKneroa3ooLqiyHHiJdGZX5ff1/P+8ZYhKzmvjV5Rg3I3hh/p8fKEYPOqcaXGziuA
KTnC5Po5wlU+xj6PcgsbDC60fIkBjDiXwPBCrJyA/5E4NWMgte7a1L2EX3Y3Klx3q8xoGh1vCKNG
XG5GSozZwE4HBjQ778H2LJyFXSZBgeQ3PFx7Rh3hicUqU2Z35QOqCiZ9YNSGpXKrHflbncFQOYG6
ZDIfYTSp4vW3lpW30w78ujQ3cM4eXeig6kQsbJ8kFu6jzvHTtPhSZd/5DDB8vHTVQ3/5QwcoQXLT
79OQFr3xLqnIvDl3q5F1M6WEucvcdFcsPKqv1X1mOjn59oCPU7Bq/eps3Pa8gYOOegEo3+maJRti
mKcQ9QMiqcwDtgVvW1p/58xFtuMfBTUJXKsEOKx2mEWCGoE5PJNotVP+yhPgxwlFGtuW1ro2I8ek
tNi0QYhBNznNy5IY921Upumer1qYPA6z+UJXpUt37+cqDfe7vE/Ot+ZiPzjIAogg+JKQgHn1aFnk
Jnjc9xhmRG4xt9DNT3B809ApL+uKys74tj2ztS+ttjnPhb6pSlrnXt02TQUW88/sqK+TMh3ODQlD
+IctV7TQa0fsf5xn64ePzzsrgpZsMhK4Ts39CuJgiAF0ZjK38NFdu862ekNMVEnzc0W1gHayo4Kz
xVSmEp4twm/0BlKbDsMjpwrQ8qXJOSHOQ6u9auSToxo5td1zBB8G+Qx9wI4Nl+tA371Y3cnSfP1p
MYzosjw0ddwM7FFMVGddZj8u286P9hPEF6vwy42wE+ELLimufZdPf1QFI2jevkV2Uq99+VPwKhEu
/1sdVkdNu5mttFMXyH1YSzOEUgOFHf5BRwgkvXIJ6B4lMwNgR0yvHZ4FrXcPrq3wmYtknzCC3wUL
Wg1SqSzWC6BmarO/wbzc0c9XYi8++gvcDIsM5KnhZHRUov57SJ+kRS18nMcNBeh+H7hWj4RKrgOM
A7BoSKSDv7xeWDZAH8ZaP2ZGOtrVmfaQoMYzTb5czxtbB6KM2kD0Y/VT86hGwSb9ELfTZz7PPJBe
l3q3b71bSJH5gAjiYKNh/CoGf1KpFC4m1cRyTW07zZmAbVk2ZQJHiTUct0U572A6FXQOMOB/BGtI
WjbpvMKo9G2oQR2bHBsmLQY4CxFCqSBMqTez/e25pQDBmDwbLmE+7rkS5OySsrZjusbae7U3seC5
WX9Ra085nmGdktqRLyGmq2vl4562ByJZgHXhXXDDyrEZEFhT0RfcN7UbsYzWwL0JIV6rQpi90yN3
v3VSbZKyY1e3dV2jlJXmUFXvYS8hN5/X8CeFovDLii9ch+8LMDoTMH60KI0uaqQOAsLTnjTFbs+c
785ld9b4vUvw+dsw23inLjhkJsT4T/LExbPit4+81gAavupURw/wLnkVJb7/B2ghi3bt3yNgS1is
NG3VTLpD84Q1852aieFZ+ebVzEoWWr595qgz58aVLOIUM85foPG/MJkm/663TkTzCmgR0pMK1sD8
EK86E9qphfCs6ERjWjCI/huz37chn8RSqy8zJADVdM0e2Qcy8qvxXI3vokrZntRrxh125yKUdTb8
LWMI3NvCyLTwzfvQs4S7PHBIo6o8Cpy599A5wd1gAAMTFKOxkffNHNjhv/aW/gpeLS9W6P8zqID2
BCmuBnkognLyhCzZqzgra3ZZj0ktkt+qThJM5iI9e1NUMg1r/WoElsxVcnWzhIT2BNJ8Hi8K/QhE
MncHDrZsrjAeDm4WzZ/nrZIPZWHAyA9EnOYrbuboLKjb926nLobf9Wh21LITktevO6S+sTT31YcI
9e7vqeflYnbvzQCrIMUNo85j1CQlnOH5MwiUULHhRm1PhXOl+li90egZW2YCXkx2W1yRn25+jGbo
RBw6f695rFIodmGXt9tZexXho+8B56buuNiDd0GMvcQ+V6MS1uGm1PK7kZYufPcOYoMI59O9BFS6
2zRBpIPckTtOVGOWHwgNm098eLVl+i3aIMYlIkVU0YLfzB7L2RAwyCU3Q1ktp6hv44P+LUxt3pQp
5utRnXFE1KH1h5ExYp3MLCMcv8KwcmGClCCHywtARFz7wjFLnXeoqUmr0imCEcipjbRNdZ2qYe+r
Rstr6AuVAvNKB6j/NM2g7kT+nT24aB0slqw/2BgOnFrOlQ0CFebGmAx4gEf33OKvVgyMHZMNQg3x
hY/JGykUJTs25C2FAsMOAAhllWFJUWPxa6LVfVR0b3nDYoF3gPYl9iLEKj3Pq9sGfBNunGCG4UMp
0p5d+hmY9mtp+y+HGzvWjQzXFaYD1uMUsMniFCEkxi3La2oQ4SESVjS4c2dQu6V6tnoeyuM07Ke1
2tWCm6uoPKW0v4VMR44ZsGeQr5sA4KXeSQGUz1yC4PT3rNvZkyOdca3vVUCXsnUhymoPtuOnuvjT
K4I1qOn6vbpSlJBXP2KvyBHIg72tCFV+LtWcPvxUpznzMbyc1aQaKLk7Sf9zj0mlwLCgWY5TVcpV
PQxu+Idaw3Jxu9MObJadrRjEWHSD8y5RvfYbhHvfdYbr/4Em91lcGD3UcepOOOFirYiaxdFTVMAk
fAiVvBu8FV7VCyc1GV6QkO9qNCELMf5robpekf4Wu70bNQfzqnSEQ9h9qGShR8slF0oX1v0hAGg9
BkRxlOT62VL1xwmJ+YJ6i3L3Qy1DBQs0u3QPKQNsOsjZW86/ZpmwzOyaGoNtSt0mMU0+GnUSQMpP
gmOih2nQID/TdjHbYTYUh1v1n4PGqIKZY9P0lPmY5ATrbOJL/e9/dwynbYRLL/ksfu4Q64e6Q3vY
edvpnu/uc3dOzRlxBI/89Qn2ENAJ6dkVE6WttKhvylroUvmgacBtmH4lXxFuvGoEGRLPrTRGY/Ra
gbTi24SKak4xivCY5FFA0x7YKaOlICBzcRDZL2Lrk+onTQr5PAfGUgfKHZbnjyu6b5HUAPLyS+qa
AWt3i0+BIaIo2JpJLp5hZnRjyM4eAFKSOkLXNopWkG0qhS9AqepZUDe0NbFOc7xh1n093d8XLgia
ECoTlgEfthGJTRNwSy5YHA4CGFnITZ2p3YeDgvFPIgszuZuSNPz0zTOywal4RNtzTMubgryozPrR
TN7bnTuFuxYIl+i/YsP23WyMue90Spd4QkIkMqxDbwN/q2A8lmOKFV+GthR1mrV/hEOSNqFUMiRS
tc8Q8LyOuON//xT9zzD70O/qlAAWCpbo7P+3nwAnlGcub8sJ9DnH0UeEUpAOt0SLTfa1mD3Q9ESa
evoCcOsj8jDmLnSH7ZKaxtjXjaCl8r3OKwsBJH/+0ZXNk6TWh1uJ3W82WYujif6S4BQwvQXdI4LA
tTcxzzFvcqkVnIykF1h0lnHE6hqsXWxXlv5jbz7Y9AuRb9CKfRGK0hWy4GtRVhQMvGNKbCk9IhC/
/cDM1iR5R1GuT28Zc0t9xMS7eAvEF+XA06drJ4gPFLXBg4IrUwNyaD9QOfvyf6Wd8MpuOCKJFza6
z9K/7J0pZkzlyrGxnpY9jnaQBJAUstdxcvbGsL94XnBOU6tFJ9Dfx2FoB4BF1LCJ4eoKxBVcF0jP
M8fIeXx0H+HQCQsOJ7lQmkLmAQmbV1it+eeUSIMr/GO/XSV7zNBR2Ug/QWeuguW29bhfEaogb+5t
pgH1OKIxneKtmAYNcjjqGmHrNGFZSIKHv+vcVrVfYSsHVHEVmJ+Noy8TqD9IazocY5LvC0dwENPi
O1EW8aLHe/b5O+XdOZJqKnWcdeqr051XF/BVnew2RnXh6+hbf5RLofImeuETVpyfbDZuwIIPpFID
FnBGzSsECCR3VfPwDa1Ll4uJ8/voe8TkF47NyYrFh0l4yYn8k0OwbHl6BT/5wxVmtWJuyW3n3kkA
VFY7DdV10QLRvU4xw7dWCN00HOacWFn6VtmJnmrkfya4sUyqAFG/mG9hRmo30Uz1jjcrjYdif3vl
eKaYwhLmW6CvHwlMMdSDTMQtsqXz7Zp/u4scsfJ9CcCL2XA/aco+FvWT3hLSk/+/LuDi0EkZYP9p
JUc5afQ2J19nrbH2nv2t2I7EgR03gZCGsHjs9uivJzVaeFW9E57eFdmDWmiRlQugBPZr395LM2ma
WX92bIEYyf3+x2DufjklvCcvjK+oqyhTNVWPzDIcx/1RN5KEgPc1zZcelmz5o2yFyVyqxKEwA3g9
7O+Y/l/hFXOKN6llQnPCwawgve/42cdRVnTWzNxQAWsTFkFz2IY5LDUbMFp8LFXfVWppUAmsmxxL
+pFhoVWG0SGsvLqW+kOdzMAaM5wgewJdGRbIzgPgKu88i1CID9HH9qMKUa1XfyPQ/F9l5uH01RyE
UaU8TlnP+yHl90Vs1OEgLjlgisRlt7Lcr9dF3z/xIi4CIom+4rQKu35X6g7+BwRmTXZLfp4YeQQN
58dlDprxoBuq6La0UqVpLefaUuuW0FTbn+42UNY9uaJaPjNo3Rp8fgn6Cib1ySQvCmZuKAv3ygUM
11h1NFCA9bi4YUcQqNCQPN0vdpNDxFa2FN5c1PBv9noxnrMjeQd21w2DFWMwaQPAZkS32tb2gh+l
u8Uhuz/UEd4EVC3rvQqwP95Kl0cg1dXR6AZIkA/SjNMtjS7W32yS2aGw2shjNOpEEcUTMZiWe6kZ
wB85CNGTAoANGsYk4wEcvJwfHJiwNWcWSxRdUGMz8RTA8WqShgzdB4xIZsZG0gTrmAWO7CspEOCS
dIzWC3z+1/2US88VLFCnb6uXaejOLV6qxwyxKdLoRvZ3V/OUjkb0bGk4wozBtXoigDOmk9UMLEf4
Bk1kYXteuSkoPQLwpw42pCVAeSkKnchvD18P0uYKWIBLt7lLlpYPyHaWpJIih3z61vOv6Jtq0YM/
2PtqnngnTgVlEVZq7cuKDN3SzajqR/CviONucSSaaRRSOY/ssPJEI8i5vZtLRNms0AFvvbhTctLz
Pgk22T4Rihi1bjHXAG3nH6vRGSdjBd8Hucp/CdbhCwkydsVI4ELkl6+/vSGxx5HE2P0L4667nVbT
v5e0zuSu+0gv0NI506gB89ryLDJE3qL44BpdgN34CnkJkPo0N93NprJOR5ZQv+8G4oZ34dEvky/H
5tTg68z/4pgwu76NgAdrlGukXtUY1DAA1dd24Nw1LYvu4ux/SkcIksgFOysZyvxUA2tkAWX35oiv
Hn63msXXVhpzFMtl7nON18uht9n9peEe16L/RubQFsuOXETzdCetuk2OBLzsSiGfLuaGohZzt2cQ
9y2ciC8PJCEMTiaXoV/S+zey84rWw/1AH3EC/swJwODdBPEYmre794/5njzYlyu2kzfRNijo7DXj
hNQDiceuFf63hxh8rckxauZyDSgKxnIXtInl8e8FvGmibkFlxjdQF0br5gH1+u3TqFnkYkfWlVmh
hlXHnTq7s/FMBJHfPZ/aurqWDQ2a1lL8cx/fgM4C8d2Fxlim88nkTOaXFC+e/0Gd4ZbqHBrunaX2
T6OpeK7cVVy2OtLxQUdRIuD5moNx6Lo+WqCbA0zOkEjDL/hey5RovPcJoKvAZ/9IjyyWtBw0ozj8
3WN249VSzk2xStgVhiWNIB9mYXZcdic3FGmuEbG/Ej1AfVIE4WFmXQpa2Rfu9NgUMZ73i2J4Rt/t
AY7Q+OMsBsL2o7UpPKvcNXFu1U28NhfA/zUnBSy1ayeM1kKXWcS7s/YbiazeByfw5sT7vfHIBa6S
mjrhT6gNv22oKhX5IrH3Jk2xY8jfqhFjFMKAKnHKQe/QQQPr5ALuUZ+JYNCxsYzV1fHCGsIP5SyI
xon9RzOM8X0CSuS/DZ1UnTi0dJ9/P4FVxxLSNHPc8+ijC6xgIAt8zek4hEj7ZjFc2A+VBApyh6MG
0DMF2JGkUWN4shFa6/wiEuA8OBpjVjzW7pA/TGzkwID01BFamjcNurLX7n/6AFBU050bwXOQoeFb
p4t+L0Tw2//lTJGXZQd1OG0vRuh8x4lowSwzdEeChZSytN5xWJ1eSNSwmihp5opk5NWbkVPH+VTh
u5r1hLZy1fukGAHE9Iv524gVuXxGqxx2pgvS2ysRP39QB11nujoH7pv8P8VfuPOUNjH/wi280e7F
0DA5+eqd0Ko7USh3w/acQ1zzSZ0zgMIplGlEKXVS+mG0WLmv3r0eCKKenAz3D2Tb7c5Hm+xAfdwb
U55RpqpCdObhVeiIqorwWDALU+oRZ/zpFMHthSYqn2fm2yLmZMejHawP8Kvt9dGS/Y/s5Nab3txj
+TCQ5nLV+NTtrIYaSzH7EvOzmp/AsXkW4GVFmncT5zMmcZHcPwVXEzEggmWnpesOe5w8OWJtB/js
NkcFomyUeGkSrJGEp2JS/V+tqK7FTroIeGCj44S7jN5+gPlfPGFYwRCE9dPP0HQxinInPA9MDiq8
evr6dKE4DyZZlqikAJ7Npgt5Xd9rJiF1XTVFKIYAlnXHwvdylfxqUT+wYy4TEtA794jxzj46Bmmz
wE/i7tiargnaxxxQZmlPsRD7ppqIzqhhlG6Ijn61pz+IOYyAmnf+NpvHIrPDIpF6nZVaM3LeYAUq
jiyn0AeqtGfUzSSxVKVt5z3JNrQVMgNWuQHrPCmdoCZVBdlRNaAvF+OUEiAF6QTeGwqxlZr/oEly
aJymgOnoEA0oj/jG1sF1LhH+eSl+5ydaYukBWccDGFvy4BLzVpOrFNw0YVoO0N1k+bXJ+YjMjN6V
trvabdoZqjxBcIg6UZVEGNm3kaw2FYkaJB1KDOMFKjGvf0xiq543MQ0KzIHTXX745orAJN+1y1rV
yLkUhzYUnLUzhDOux9VLTL0VGMMWzlS1v0eaX4S0GpWcAssTfTuj/2+8oO7KMDwfXxPhhKSeauDw
Sd74g5jrDJqJw0CGs3uE5g7IhCc6X/hhdTHZIAT2uZGEwYDG/WbuHL0PSKXF19zuAkYFY07QmMth
uwiG3EAANzKtSwLEv5FS6Q+vDdDKvV2OIkKVp19liShZB0HmbtIAP0oih+12CB04VmUAT9NgTVe/
I2tj2Ejelt5WwiD1sOeCWCxaPCzGFAutl8vomoYRkVtTB54/W5FurE8GoLeHGmBZ5nOc07fbedEs
/VdufQtVhWXeN6XPf1FZZu0jtRhihL3qupVXtLG9UEtkP2hIwXXRUZ8ibj4cQl4qBGqwE0787NNN
z9GD7vqD6WbxIexbBKy7Q+CtftgEciaSc/wKJd8U7Xyu5GlOU/tqxdcL9cDErzW9jmhuf9/uRzTL
j4+GRgcwIT4nILQFQur4odZSebd7DjEkyCpa/yWC2FRSWoG82vhsKoFWUJn91ImkyYFftcCt90H4
dSza7B0MOuYrx4DVQsDCpqzpUzmWv88ICQFA+qUo9+GoGQASrkK0JxKlVYghuNcLEYMvA8nSGMAL
M2SwhXgwqHb92GQEYJZ0b8ynWFKm+ame3owmumPyhXSlcJMcItC2Mtu/MvX3MCtpdE7HtpuK645x
FRBWPIFpicWgenc7cIjItz8p3+v+TNkKWmtZ+3534I08R4m27C1l+NQjIY2ZBIsJW1grcYm+6O/y
pYLPt/wffOfUqnDIbUYlZC8AdD5bvfr6+EzgKIaSZ2kU8gON9VgvwEIQLmAgIq96igZBhSxp0XCv
GRjUi39eP5kO+Lxn+HMleGYtj/eSI1+C40k7gk3vOYpfy734/c9cvbzXFP9hFfwXtgGG/NyNrZxt
siAmBJEEyrmKlL8sWXhRCyJPf0UEVeIkKubc1VWtunxQ0dlFyZmMU1ZVye0KM0btrDv73wEldbEL
/dS5ZJBpAg4pL6vrLKY9FwAgXqXjU7z2zI2ondxJiGTsTTnMd8QXgxeLKt1hHr/RBMP5qbPCKywj
V8rL/cafyFZBgCKGZAFGVN2LwQjfRupFBUrmU6QqkuNXZyNwo6rv8BKY2PGFz0auWvGLwqO4EprM
oz7O8aUY4EeElfBTf1ovNuZG9KiTMskOVP9yI2w9b1QXH6w0jwFnDG9Djr/Ms1lS/9iD/OFpQDY/
GnaPGMDFe1NRcKpzEt4LcZVQt7XvkC7/iBUruuMi6ReWjCEdVffJfMbKml+obDUC9k0lNyuxOIto
pELGOuUhTJt166x0HPNodAmlXlucKehVvIE2SRTzbi658zeHTT8Ag8kgHRFph4GtruGAdfY43YGZ
J2c5Px6RGUYbusbjSoVNdwTchZLZt9GFLI2lLJQ7qz0cIoJMYuJl+sJmNcySnWfUTJYTBQ1UL/Sm
sdg5Lgrjv8gGAb0R2tNOzADoblSwEFyJgXEAZXVsb9vhR483ZSRtxUBh9KvXpL2kffdHjD+Les+1
YfAG13Y7Sjit+lVEOnl5urn8H3JXISkiSM2GbjYt3GKU4MzwoWXBnUm/oETZCugv8l0rvY4goaFc
F12+nvFk99cgrE7mtI7egrLDn5uUBboO/nNFmzBxhPM1uG45Br9YdoWQRRQvYlO4W3TSxRA576rt
3nhZUMRKmGx72u0iBXushMKqVZ7/CSaFHVEUKrm/Foqr4XEH7vCSW+RvyRnm6NPIhN3OMr0/yk6q
UPlVpk6a+BO8iZJf4ZT7x6eICEsVfDZEr0xqioj13VE7S/QW2cXK37tcZRIOJdyQ23bungi4OLXs
U6/UH5u8ilkKmeVwHK4BCFEvxtrzRtvKBnaRx94J86aPSAVzKHve6rx56eu7YrsEkdrx3IYsLujB
8dzShcj3p2dLNbYOb0EP2rzPE91ngQPdszl7/MHvoQ7EEg1UxGAxQBAZte2Lvfgy6uC/b8Bb+KP4
2jObi7TwSwqJq/qh5m8HyKC1M+OU86mR2rDXdOL+a6y5wGEgvmIxX/NOS0eRmNnxMjxINxIMeNo0
GdmuLL2m/UttKfFDlNnqK6XTnOw5Be1PD1sUDespUs+2gyIRa7Atv3ClFSjasRnbOxLzPxkdyuZQ
xzPoyV5s/uxL2GZ+1KPkhRXAo/fePfRkj6xrzVqtVCPp11Q9dJBcZW/XOdAvJGJgOE4jALt968Ry
B5S+kXW67qIeMjxfmWuPWVZisMjiRBaHwdIQtijl9qTET5qYtAd3GJTFSJF3DHpkCBhHLWyl9h2Z
3kgoT4RMRztypvaWQ4Ds1uZmxmZcnzlECskU2WJbexOm7YX04LgC3peNR2JzQT2uVvi94Ql7AZDz
irbrk42/DL19IJrkqZSz4AnrAnIep9ShwGbFm2dfPw5Hf5dZc4Q0+o+bibKAuOwJnLwkH+B2ri9T
oH0CboilbEFm/SES+wqYYA/Jd948OJa0ycRvbStrrwMFYQgZO43/STCCNd0rk7a8WZNVOfoKTN6T
aFzyaXmtLsflEStQfbJiSAEZSk/2nPRz56bF49bhtIvMDYaRGPDxKGqO+P+2sJPBfwoHOyV4QyYf
pCCNy1Q8CjzHRQSgq+63HAvm9L1gT5P2PzRPy42tj8snK69BhNe/uOVfRWiazHLxD1cUhIk+Pong
C32oUrdY3cDVcW0OoOAlYKvwD3Tv87m+zl0ZMwI9c6CEPY34nKCWUhYKM8uDcKcjXSNrqnSZpjbi
CveF9CmGPCHMD2g/tk+sr6eLM4Pi7P58T0gmdo9oeEI7XsMfNI7iIdm/bq34f4ZEsmKAJJjCHB4X
RBOyVJlQXPqhcA117aXaXqYzTx+9kqxqOhS3hoESyKcdJ4y9sD69whheGHxCKB9IDdqWLlkFSUau
OtOLcAjngsTq3Ku1CIk6+6HFRSLb7lcCyBl2ACbuPSSR4b3/0493xWfkmpmGqG/sQWvuubzFVuJw
CjF44gOQoGMjQ1ypUjbJwu8Xf8FCjnf1/HBlUpvfNjsn+wQPcQfgml71McelSa3rR1xzFcMgBxxE
8ZtwPr7pNc7c6bs/bYJyUcGIx9pvQ58b2KntRML/XOWuED6ZklA9UrFF5eHXflVlWMl1od90g27t
llBiQiJ+CHHf52hDg50x2p/us5zYgdkLRsMnleme26QiFOsZdoU8kuecnx/hnXlxpV9IW0tLNckz
ot6g83+i6jeT3E3xnzWi+b2ZxBrxzSqi0VbnWJ8AVbli2Xko+MQKzmB2qhxULSmojvbGfRlP9Cxv
jwuCdWr/a0UtwQg/JQ37tn8TnWTj19QTHAl8BcFRbSKwwiKz/zX0Y3YXPAWFJ9ndwgIxOm8sFeu+
oEAW81WvH/4s0xOzSDgs9iSYK47FASYq3ksFRtBcOD/ff2TqUQ/4L0zoXQvk1lZo08P5rT2tCmN1
XyXoBwv81yotJqf60A/aTAsnwc5cgaaGG62rmIzuJqOj/JJhkaaHZT62DL2prZHKkHpIhldd4Ud/
OB6lmL1I0Uc6J8kOtF2CN/kzSQwKi94S/jclS+unovN6s1SRUhaEBeSDhgHy8NHjCfn9Ee8SC/tC
+6zq4tEwERcwyz1eP3QRXwd9DkN/jSIWLVz/U5VKh0OQhhn1KlPBU0rf4CuCrhnax+U7kK6v/FH9
Qx6oQU12lxxQ5Ys18jMRiExN1OtYi0x5RLvvSYf/yh7I9i2EQl0GuLpxGCgTfXw6qmvXKRxVGpH3
J0f587UI5X3Yo0d0dv0XDWjZ9NOgP6VA+uJG24kgqbK7JldCWB76BM0kIJq3KZvy5icZEuspcTry
hPWFQUju0soLgO8YBGY+mS6fAWfsRfBJwh3G9KsU6ruVuiIHMw38OEZdlFNpnr8a6eTGGJxhg6JN
3CZmVCs+rL6+IVpUQyUB11PslJHPD8re8s/xve5pMpcTlVSq2/FifTbzffVnY8PZvddEAOF/Eikn
alsAEKVtARsUe7N1tzzLpyFCe8is1qaTa6hMNid/Fm4aN1xHHScAgX9jCvwMoWPhSicNEdvXWGI2
H6QpXc4s6Y8HRC+5CyflOvsZxC+GhQhWPJGATdjXqVHQwUPT3Gm6RYRB7+FTrNxnIab0j7pOUErT
19VMtgzjDQ0vOrkKiEdDRqS7ZR5xaLIhGQdi0YZfnJNtbmXVPlNyIVAm8hWuA5IHkpG+gtNRY2wT
GKqRXayEpJ2+vVB7YMyFGwgeWoG2iMvRTNnKax1i0AlW1viZzTg+o8zLji7a08vNzGBtoncCO1oF
DfPl65/K/uYPcq3nWwb0T9c9dkR5ztLABrSP7mxooy1j0bjiZ46zmf+ZcUszbw2XN10O9bHMWeng
ZbPg3UytUUWTyXwZMqUYnRjEzLX8vRfimgPhg1sP+VOM65+H8IQCu9WfAZzbg3/aBC230VtPQSw+
er6kr2hWQ/CtfiMH7Z/mu99m9vUMD/lBCmUnZVCO82Bp1y8WKq07bCLGaqMRDYDZuAkh2Qrrs1Dt
johYqiTh7nUS+0dZBeKGwy7lTxtj/cXVm6RoQcIOEFGxu3TwMfmugERFrJXXsSAd9i5efmk60XhR
BLACtQAWTpGjGHcP5KjYhbnSLWFPYMVqtzyVxWO0/fJbYtJdnmtfudydgGnLLnevHXv1QTnGc7Xa
vPTxi16xJfDMi+eVcsFrH4gRDxtnop+kBmC77jNwlWFfIWOL0bSBNo2h8f3uLmz4Ana+9Wyg/0kD
37cGLjK6pmXdsblCWMuPMaRAumhXFdx8lhUPQ4yA17cwduk7bzFUHK3EGtXWnvXkSmtm37InteDJ
N4L2fGckPYY0YKaIubkbN0mDAhvRL8DC8N7H9QcqwDQRUPqCKaUbpcKbf6b1+eeNkFR41fFixdcQ
u3BssVaAiu9VAiZBMok08pcnGf4pwkB3RfduTe9He4cyYIQbrzdcsSPG9fIhZrAwA4X4X5jTbWX+
2wVrPOk5c5bfMViLyEM4iAffjYiyUXLOMT198STGLZQKifNlPeTpGaE5lr82Zx5Btp3FD64yQoQo
4LLuOSCDtnn0Yx0PaTMgxP6lTu1kFHQIgCzHcQ8n+f+aMkMk1ie+js2oD5rr/C9TiIQX0zXazZIh
/utqEcpXECCRdC/Ii/QlEjqnL+o/oldaRR3uFbsbG4eoZIF9n1rRCVqLJ8g+1GvEfwGAXeuZ3seq
AtnnG/2jhZGAkzRNeMa5dLaKsw6mS2MFYxTEhRT9eqiYqcvXdExKZ8wRYv8bTG5vgMbYAXvlrDEm
v6c+rr773e26bePeDMFLmEEVhojL46gpOSMI04vboLnchg7LFyR5+3fdz0LKLu0uvR5X62250yyy
zeYT28y1Hh6kEbBqVfPp05N6DunhfGsjNkWCa34iUQ6WGVZReeEbRW0RaRxVorQvvG1jpCIiIaLJ
1nr+8pN0DjxWTqFapsbLhbQ/MIQ2/eN/EAw2ZmD78i+UZSWD+UL+K2w1gZLASV3fYPU9EKz4+6i2
i9Hjrd8vhI4cvU+UTQAf1eQBANw6K8gAWuP+Riff2OTvs3c0w3YJWx4K9AOJa0k3/V6cKuQjPrti
S0IIf4lN1XJZOgeKM1g03JCieG0hjqEyBog0jTFtUEkldNz+5HYg9aCEDyRreqvjyRCAfcLTjlhA
e/5z74Xnm5QP3YJghsOL9uQqjdrB8cM/i3re5ryTJW2RnnSxIrzIVPizxcMzMnzU2C1SUdpbcvmy
ut9avXvPzUvE+d/Nrydg13+Ki6dUglAo3hEdJ7jj4qcny3IWygsXs1jD8NxUFH9nDgtWTvRPVc2b
uevqIy6KLoNosR0lW7jln5pvMjL41XU3zNygHfL/mdgdVHNePjYHinEvuG4/K6yHtYkwu7+xAhRH
pJknnPLRJf8vcJYRGN7jX7iQDIq7pzsMxeHpMaPq6mzwfH03QCVK09RJDXMM+ejP8tHYkAxU3F5n
CP69ZSFJZcRfiyLl7R6YiSZk3ysZ+tUoKQ/CH3PCksjk5hDA1f+nJ67AQP3wc7orv74hx8Bju1E7
rBC6HcxScGn3yVtEbnfggb7Bd/iVmTO3Ymsyxi9KOt0lpuRjXZgg3yTVdwScLUtCO7wIDC1x+4/i
yVPzMV32geIydHQVOUKGpDwhUGX/jX35FfnBPBuHPcKASbJwuRgZpPWc0vCKbAjkbHORLFuSBsux
JSpEMiacaOZuK/TRtgDVamR2Pm/od5LY9vW6qBKZsaD+03k12S0NBzZgkCyqAn9bKMfdI/czT7rT
SV+E/ont3/XjgBi9aR0KrASsoR4bWAiB/CxW4fj+RqUByDVpb8Vr0IDn/gGpIncsxmaixwTKzJaw
wC1KFN2pjXTckGr4WJ27Yn8YLH1/dWHSt9yTiq4dEJPac1l6j9aJ4TgXURXDH8CGYlVc/8qaHFIC
X+IoyIbds1IS7PbMhatVC0WrIW+1UAGv1DkhvTMp+cFLUTkhP2ukCypizjwg94djWdk3ECa1eQDm
BNy7SbvSIrcr++mD8y2AGwgwaRGFuGNub185ExnvpEQAvybqgqsyu4S3bDVOy5ZL45bZ4hx+qr7b
HJEpKf0Qyi09iLvKiB9Ad672SB8WdDjoSbOltCUBodgtntoQw0LJadB9egR1zYMoZsJyhjxUW5RJ
E+Swzo1AHlw01+CDEFhtV4hTaErAjbgW6oZnv5cUB9xZfHBfEp0GB066cY3cEgXk3TUtbEwSWP6H
ZIQBtvA9fhrC7XOj9EzMvHlKVKuny+2IaiOhJzCCnMJndENuK78NTt/04M4Doax9m2jJ6JaEoRid
7FzJO8Jp+13KupF6aE719f6ZQNvmJjjMql+DwzJPQviKXizY4abdr3HKGr4AtDFxO/XDXhJk98Xb
9XoDakeTFaybsuAW6Sq0tLdmFyup6bjvVCz8cGozNcA/hb9cZOoL19beU8CaKQduuvGiKvGywTn7
Gw3aqoYzDCFU7g08HJLPaircglFrK7Sarvk/f0PmixbC7rHaMzHW7XJGMeF5VrvGfRQTEBhNOKhh
5CKpBNwpYeh0/vc9nh7XCR87EbI7+duFCSGOADAPLVylFjC2Qcfb21eVTQZA0SMMTyNtO0HvzQDf
SpU5IVcijdHebfxlELRMdyzu/Bxy2r1/7WdRq4pLQW/8lkp9QL9gQ4jZDq4Qp116vsIRoKe4o5Al
Bd2eRg1Uxj//fr1N9pRI9qM14Mro8hfLJiz/pb7i88fmuuZUuk//J1Z3S7wZZeoPOX1GFwoAdfXQ
Ju1QdSdusvIRIzAvtx46Xf5SZd9EHCbAen75aAnSqPp5XISk/gykhdaxFYJ0IbrytSdc8TBAT4hD
BoDDEL9eVd0HgPHXUZuFAbuu6Oo7sCzL1ItqAmfgKFTrr0qH3ccnW8dEr3PVIsME7/J+y6I/nIhu
gZaEPd0sFAZ0iV0RQjlqvHDFqC2m08063qKJvyFPRo6NYzBG6MEzo+8aLeMOY2o6EsXPkJ7RIl/Z
746FFwYwOWJHWlUckjO70IYQeY58NXYBZwfneKppG5P793p71VHaHaQyYh6Cuwp1nFTDiTfUKUlp
QPHrvD6dWAvQwDrqGzRNH3Od/R6DLgLJgb/s+Q5Yltfbnsk/1RIWovHz2++xJmATtwgEPXx2XdSk
N01Il3H1WC2sNuZHI2pGw03PW8BfdeWCVtTpG4yY/Q2vrVhIF/V02ZqbtVNBgM0PAQlZTM4WJy8O
DJiCqM24pA9aO95LANFrFGS5Hmr7d7uRdWibrTnbL7YXIyx25kEk7ar3Vo4262DrCJkQdtzUrzAE
4Tv4ujwLusMKDVeEacy3Q7HQpEHgHe+8pUJzYWiHTGW1laq/RGuoFg5sirAL58VDmhZteCCpuWDp
SNwihzEB7yfkDBdT/K0MgZ+ViQDJBwjHJMhcXyJPTcwenD1itohxIa2D3DO+RrJ8GFTRiI3909x9
WePQJPEqv2TAjFFER8Cece1/vBHRuXl+4V+7t1gBRQa8dHvLoDEbgj0x7L2hL8WziGIRlqjDZBhu
o6R72kLPGHnDxo438t5m10UqKxLlm1qHrnaAJTDU0racjLMdYBCETIll0enujyMMcFmBS9wdutBZ
NLNUoYsTad90sGUmBLcyDD8SwDYcKUBDhRs4YWUY65/Jp6wL81uSrs6x23481WyFpFwfz7y6UR3A
j0wU9+RO4e6tGt0mXn2dC6MgX5eGaDC7dnPirvrXV7nEs6zjUQHmpY25PhUBSSaXS5Pyudsv1eu6
JJE/dva58UGrlH1qKandpw4/q2+0tKTAYhhWjmhUpsqSStm/hS/v/Q4rPO6qzAsQ69oDExLpGD+s
nvBmw54AetzDNK864CPCVuCGhIr6sfRXG4rKqyTGoliKO824CorltzIl55zgh3xMm2HCgmHtlt8h
A8b4DBcvTNgYeE0YqmyhFD1CFFIn9W+xnjDFCc5CkLKbEl6uCNnor56yRCB9oIWbtU+M6XrPnBaV
g8h05ZOY++vZmZQb8ju3Ta9P5rkLZwLDqhTFdBOOW6VmuUFo5eLLe71oLpuoQhJQmNUTn/lQgtwY
A2ksrn9jbSH6xx/+GJjGwb5Nrw0ixnlxguQWf6kFfqA6uJe7SCUjR8AfHEiFW2j8walY/BzCPjqp
nVtK835vjklShM+SRQAxm2FqgIyctbJR/mHfb3KfAVJWqFQKjLcz+dp3ZysHOLJRMaXZXRUse1Fb
uu792/Aj57ZkS21KipWLCqFM6Eo69mefMVRxIMh2Iyk6f9mUGev/Ao+xSimETGH/uplL9m8Yjn/Y
XgNAHsQZwyfAGo5YkyEKNxW7Uk5NLigWMOC6Vn44AVaret2KVLLxzA3LJyxaJVFApQUJOt8EYID2
3mvKgnxnMlCykIx6ttKGI1UwG0TicO4YGsBr/YIReQGHToUo3MMoLglJMqnWwU4gp0bbhkj3e7Ae
jEWfocVDBkPK1JC8J3OWwonP1E67h7NE+5chliI8dGniETvShv5ftNgahszL4HhBC09nDnPrzVbg
ii0Q5lgI1NKXLcXBIfcYyYLj/M5iHE3cyZSxKYmiS+xwTzLYOUVRedeghERTug/Tz0G7ELnhC7VK
96v38MNKkTGMjE8UrmVA9gfXXzR8w87V2xnkZQ0qkv3px31gWYrgVp9CkJIXKXzP3p0JM/pwzAZ4
2bb560aZ6a4dYfQMKy3FLHkt7WzHzPEMt7QSNlMURjIG0uuFte3l1agE0vvjpJDE/h4N/xV0FCMB
5283KjlbZWhiexz1RAeeH48yqsAKyZo6WvSD5EoQRtYCJRNzG2kB7SGSpVOLNIVNopgWbOgG4m55
3ijCiZdaaDBvibw8VkwcvTtVXMcfofjkDsebKpATzMZxoD43lUV2Jky3N/ZI3LJNP+76L1LI24XW
4T1tM5/wraB7VrhG62bCwcTMmvOZcqimHiUH1rJBhJjtrmJXJTVIE0DACbMLGKinxFTVcACJhPpq
y5lqSUEDVAXy1E4n8uzJM/ldxxiYhwW6FxlVpEenE4sM3jxSweNwvynyo+NXPIsGBGR0hT6xn3JL
ZkhQEdm6y6qSXResai00f/35kCUXQ/Cl8W6mpXJXjMGAJgUm6i1kS61WNnmUQxEe0Nhtu0UO/Tgi
UHbYzmQEDuoXHqiKI3nPKApX8BTYdI9LEuoLob1OiA0Og21ITcBFEWi7cZ50n3BcmLlQdxI87NUe
etXPJQbeShHKq0wzWYWO1XHhrVGc73uXr7xaOfVNQcbBWRQGzLgeopP1Ck2C83LVN7TF7DJ/RhAC
FpPTsJospfPJHBKf+5bSBGEUw/o884o2M87MvBUsnlHood8z95BrWwYImOONVz8S/dhvalTvqJaR
q/ckNbQx92AJmuF7qbDYkLqvKcoPeOSyISSVTSlNH7OB++crVOf9T2rxVFjA0ebdoDShoswcC3zN
e80iKFQ/terZRohjoPQ6PlKrA0YyRpJMr9Upjwx22+p6P2l+V9FnO7o/IhuJbzlwN5nSaxXQxt9K
/A7LtncD4Ar5sbFBUt5MDhwqOP9tAA8XxqH1YvTt6q2jqUTuAY4SqEuP1B3i9pjjLxqTGdCC4jry
ddPJ4UB+bpeC9GNgtVxJZ0FVHod9ALYfXCXSUsePYkxL6UF8Pajp5dPkpHXz+OVXzfF9YDtgp30b
XBqGnDmSmkpMKBaZLVtRJuZUozQ9z2l4TX+aRodvsepRk56hlNQRguVGyc8RKbLd0R6mlS5ogeTR
iz7+LPtG6G1I3lB9lzbMqF8lADFpdwU1gf4mcl4lqsNBl/aGpdKp04dzZRiL4YH3UWYB1dMkbu/Q
OEKsvY02BKEavPfXP9dYXICQpQBu10Vb4LjI81Uv/RdpwFT65k8NXewPPwW/awg8ipGuqLrhjp1z
kaIsd1xyqnwJfqlXO98hTGMiiToJEiXp0ja52GBnUbaoyYpRld5hHX4rQWXvvmnz18SiYeKJhNwc
ZuYGgWAk0sWcqYq7Gg9HPuXdju7FPq2eK64qhljVV9QK9d7AS9GsWsd/6v/s6gGyNj/rvCalirLh
QCi+Dr1GPGHTfWCQqvEaG8yawfjDPIDwjIXXp+6EF+a6Ei8ZgQWGHL0ewBT1ACbpgQkLb1lhP1fg
Bb/Qo5rKqpEGTGZEmP4RIYogtE9JXKWarjW9Ka/l+M8g11JrzqQwjbWuKe8Yv44LDaXcr2pz/1so
aPN4WwzkqFwri8GSm5/RKWhf8W2b1SuzVDf69Ze8oEK6ZCalMpUquDUFE0NlYnprGdKORbtUM8MQ
cxGsT/YgyzHgQHGNajHQHrGCkBzm9heSOXjpezjbV1pz/JYqjwivfW4Um++PqZzH2xnT/EVu+X4n
33eNq/PR70it9/cbq8vZMJSZsJaUEMdUy6QobfJ32XvYu0z1Vk2NO9HDO6wigMJseN9dV8uvRoDJ
0fcQOihNt7/3wFnk4aDpUjeLwfGpjFXPym5knTcTdxDsGeUqc6e1NOvnyiYTDDd+xeUwcOJXIn94
OIEIAIuNj2wvfOCEsEU52e2REHTBL0ZMUv1HbKMVowNu95jtafno1OF0Gm0E+yY2qDzEymraNnD1
p6LLlUnERSRwZlnP/hFfycp/Tr8eWmWTrOROUZHe+1m3g7btV3i2MCp9Fhg2WPasHlfE6d3ZQD4S
PUbPFBDR/9mGyOLlZ8NeKKDQxCvke0iLVquc+aRX9NVPDijtORosbOF6xGpoR5dYKzvVzgUH6K3m
/D+JnInUutHUtJnAU4hJU62Z1iYToxo/lXwCnBnXC039FglAxR+q9BncvJMK9Efj5yDhIpPnXMH/
rN0e3ZqF0JTNlGN1f4BtxN2E+mA64PTi2+be9FNRNzsELlIjmBjasLjgy3v50m8iqHLgXya/YTuO
7Rm1QXx4dIK9j2jZ/2GMLargj7kQQOZHHxgmBJmiBwBY5u7ZsaMx5BOLGOFehdthkaRHc0plrhaB
eLFmRMhz1xlbXxnfFRT/DmYGXB5NRYwEm7ltEAeXdckIFFL7RDf2XDdGYwKz3HGfZ1KgqtQHgy4t
LNZLGFXNaacAokWt4BMbU4b1eRfj+ycECjrC3C+LBp2zDnI4VHpYABleCLqnzhpVY7GTvE8toj4j
5WNhnfJW9PuWjm/lzRm8ZOaixiTc+CAMm7Fx6dfZzuwkxmIIGZGGcKofnn8dB6JYL5qiPKKGQEZa
xNjgxd2WOmWpZcjolg9zIRD+sCxSJBXBdGReQVy6iTky8Il39Ulul8IDWWB+nU5jkJ7DYdVoBg1J
cV6Fs2zW0XN/21Xdl6klBnWfaOftPHG6hpavEPMii+VYaRXl27dUhxZTxlSh9Bt/ccYp5jWIxcGJ
Fg2D9PSviaj2Y1t9va2bamANziVBseVBC4xMkGrufAFsdYOF1bVrQ/AKzFaJFKBuMcUXvL9PPfqd
HoJudf2L6Tup6yPuamlQv+N4Kcv+IS0JRwNCqitq213DCTBpA7BBmUfiP9iOF6xWlXGuWmlTB1vu
5OaNEdzh6eFAiGm9QRzn1FkUqWmrSn3RGA7CSlTKfBd5R7Hw57s50hnifXI1mW0XMgvMZK9y0uRp
/87VtW4rW8zghhBWYpPHvdq0ewMG2A6IExVpAmKHmJo5M5DNh43Nna93pMxPD8VjK599eaXZGNxA
3crhYMR8MC53f11RNM96X9cxyBhl7D0Xe60YOLCWYag6qAFjVYbaevzIzBVjM6Tm9Psu1GniRLoE
4Ax9epcWlElBfT2p/KA5ZqlYFTbp6bwR60z4qwSRGtYJZuittBDSX5E+FcvNA5HNTel8Om/sYGrj
4Po9OCtrTe0Fn1kjsWpLMKiBCK7w0RCNwusxb9kXMp9o+VfriPCWctiftnepaRRl6ZYaLOdXajD6
QEbD3rJv955duzfstSNO6FXM7d8rGFJkapDJK8nITqcV4EKwHEodmgS5LZE+N1kgxT3atUEinl+e
e5sHn3L4B5LptJyhcEEysMLcObPgNA89wsY5Ntk4rmKMu0hZx4E7gMApFsb5lRwgyCxFQ9MldFS+
u1aXKob2iRTl8SpxAKumUQEWAf5+qjDIWY0YEl4lU7h6+tf0bolkgjQ+rUao3EeSb3Tf3TR5AKh/
l0xudi1aTBh025f6/bCIBZxVNdW7rtyWlGT4SPkL5S8rkFiXGse0mGmBv0kCmDILE9m4EokySWPx
pdx+FhAI5i6+DtiDnSu40c5/0kUstX+V3vGdzkLnhSkklOP9xkXuSBOve7WdCD6NQ6H4PkSF59Nr
nlyi4cTOkSp3vPl3qY5snJU1jsh+42CiohyuGbJsm4hYEcAY4BtoeogDvqtJpHAjp5r3dDErASkQ
K+vcbXxUH1G0fByPLRxPEl7kCH+OsRmrJYAvPbv7mThOxc1I4+heaPvc9s9cIGq3yrz9DOHE5VIw
IR29K8OIE1jahyEzkHlrbUu8WQSjLt6saPWGauN++rA+Gih4lh3kIeDSAsuhpKZRGVSaN9tFBiDC
zteYLdFG2CVqrGd7MS6tjFwWF0e+EejP9IgchvXZ5BsgygV7aVTbdax6cKE84YL3W57tIwKqS/iw
flU1miwe0F4bGBmxzNFm+SnwEb2oF5EIPNMsfmEJjhKOEbD3pzjB7uAlsPUwVf5OgwZgee36YDCs
F9PUhk5DsWXBoZ7jmO8uv2tPE1588pOyGPukpPvBhqZKJkrwPWnWibvla+KMYO9ZsAZkipa7uIO5
O4eIav/G6yQoGT1empJsUwk9v+uaSHxDem2yTjWUq7BZJ7AKC0VOxan4VxhfZ6qzupuWH7KwxY7C
jtED8ZG1pjPzab3Y6aGPF1bxuy9vvfkHvedQACRlvV5eYHtznGfqXw9I550N0yqk9iz2vjKaE9Io
c3rgNaxYYwl52cMG4PBSyyMZJD1+YwniqdvP9H5bvpF3nUamvQkEVXV30AJfBRfsD9rCRIKcr/b/
z9JhByLn27i3VgMtjGvjVyilB/w3YxltlCdsM0lU306RZJQYFpSDh7sybjMvWKSORQ/Pi2B5rgEG
/ggw6/bqEpMH1IYE8+Tol7HKl6QDxgTW8eRC/S/kQPOSnV1g8BEH0hlPyxrDaRky7e1TSyIXGmvr
RUEZEFk0vE8BVk2aHV4ZB0gpGCftu4wAvq3KNnmbB9xtGmtEk4pVf6jdPpzBqtpFPdSp2sB+BETG
x5s+t9SCtXP8S7H71LpVOAMEDz4W2THA3X75U7xSEaAPc4MZlRLD6VPG2qwP7Jo2C4GLkLVk3oEy
zRDNZdkxHZ5b1TcXsftk0k4Vg7p50Qh5Yi8yjYJojF5oNt2RAx5FMvBslxPblyVkNkh9C5dCwuIg
dWX7zYkXlyrBC+PI3SVhyhZqoC8hHYGcc4IE2QwyaErq8Nz33wDElOL+Pws3zM0PgYFadqb0PP/D
p+6/HS2D9cNg7L66XM/qNYt42wrbXEqnVwKUjeLzL26ytU1QJa+zUEAT2x/zL2d6N4Ncpx0vJm46
f/uVr0pFJWU8k47eKZh5Wf82JVXUWrs2cYeDGq+V90s46BCH8Xf4m++oDWOK+6fAPFJP8eH97IFi
XNb9nR1KGYEY92bcKfKdYYRrrwCJnS/9ZOokem/p12CDDD7qaq/LrXpmYpGOtU03gWm0jSAYi8Lb
TSSUoUfFFi9t8ptsHCkLtVN9qSr0gU7ga3vTl21Z1PILcnX99M6RSmMiOINGD7QxnVSqWwjn7daA
yPG8BXxfsXwmJ2hzA86VVDPeTPn9ZeCvo64xQDGIX6S8bFj6TznTgNK0LrlKUMlt0WpUWmAlWNOc
cilqmO8uNBAs45CF2sVm8ghgeuAhtY4zHNuCb//QXRZoWjSX4d1dyUBfy7ljGE/+3lNbglRsoql6
vmLrqWPzzyOeOd+L6NUq9IvKQ1dE944S+2tKk5hhsyai0dvl6HeDEWKGCX0yR6eITvxFAlMB1FDe
/kG2XY+tXrY1mJiwGTAQk+Vwv3xiBjoMT7XnBgXSjG/u0VfrYlF+IbRpSM6iDF70mFTqoQk4O9Gp
mJbmFWU6OKTImybS5WJvwyIrCU5/zCk6f+lP5Yms516xWICBItEPs2N9pxCTACKfHOMhFAXgJvDt
K4cY6/rwqw+i464ZaI77XbTuqqvzJyvuCWm/IhdkJFfghQvUxNzYj4n53AL+jiKJViakzJbNAqZJ
Ac41ht4Hh2khyRKhJe/xbLINm6isG+cX2YlPAzUsS9wMZBGqawm99wmimriCAkfqwEP5c+QdCGv7
Wtx3G41wAEBF1orjQS2prdqp3GO5lUh8HVjZ4d7EMk9p4PRNBZYu+IleBKqVAnH27xiB9fBaZAJ3
8aorNK1XeqmOXIJNQBU983pzxHVguRSu0MSg2LTvrNwZD7+BbHv9cxPc5PWvSjJNHY2QVIGwbQB4
c8jUS3Lv3OpJLAWdtaevcIQjlF0SZ4z3/0HwMdyGL9qUsvGmpbEJBLgGrHCyaFtD0wSw5WUcbuV1
4uYfkZWACA0BOHp5VaOwAcBHNVsUW0i0cKaVOmCUTNN9y/dYiu1T7JOluwAdR1+lhYKeFCXOmePL
OyMpGu8vYAOXJO0lhU3NddlcOC/CUIASH8IPzbFQKpum7IN1xPaHc/TL2p6JxJS9T/QiSWOEJhjf
VblqiOK2fD5+BaJkMvK7IiRs4MBO6/RcN2F1WYrYj8eJFrTqax39/c5nbmVWnhqGj4oYhjwH/SDG
1f0ttz/1j6nl2xKfFP3hzXAyoH+STxhfBGKV3p9KQhz56qw44WSYPFha+6Wov1XqSiHYeRch1W72
4nY7hqF0XXchbM6yGOW/pGlhg5t+9WCFsm3LviugPSXFxS0Lbl7kQ4gPYgNj06Elq0cI3qKtfW+l
djBfT8qXDAsFEA7zEVSiUmPcaU4SFcsa1NMLoDrWIEtrOQIXE4fi/U5N/bAPA1UNhlCd579Ue6Cp
GLCd7gUh5lfucVxoSvpXBQFQkYRGo0XwYxIuNvC/eNBGodgrmwcK2byoM++PMwEQb5/6DRIsVuJ2
3BzM18DvXuoS1ez0YUEANkk4RXQ307ucdNRRIaJgoiUKytaMdOCP/1VREueOAfJjdhAau5Nxsoeq
Ojrmv7GHTFis0a5Ox0Om9WVm9VwYCqvDtnkGTloSIoQyB+ne4zGy2WWc5lFkKMOvLyl5R1KFewoI
Coj2CPZmV0BNwzIlgz7Brub4MfB+8jyfGei58c/Zi5Gaic3kPLFdERWHKSdfqqBEcKLPuZW0NE2P
hKG0cHWDS2jn2/uzbr1rVI2lOPmj6I/Fq5dx359gMI3KcajUItnMUjOGdvf4VGcvqYZ/Z8SDlMTx
cRF7uAtyVpdvUDvb0PRP/xRGA2GykP0B0RmxiesgO5E4ds9+e1mcYswoNz8E8OC14y8yZQlSivtA
IMY/WUZ86AIteL9rjNdr7qfK3evRg6nntknrtCbaYC2bE27BKW5Yq6ueOx6Knc5Qol904+840Idx
zrroWk4OWLBh4bhBmGBph2piihzkvf3bu7F+VbBl6PFFthiiDoWdLITFBkt41feyBa3PkCx3ZH4l
7Fu7Gla2n1AXdTz3bPrNCgnagz2s5KI1lCEKmqDzghUoapgMqJl8KUfzQ9+nYbF26sjmEPCP8SdL
cIRBc17XH2uXZqbf5NcLECHa7rWaOMTYsyITeTidjTgl6OYDWiR6saPiSkm4ddITOLECVCXETBVf
ArQemUakjMF+cjtHRdYfGkLdJkpHOZNCQ7chmjL8kRJgpjOLAlACymm0abbaqZJWToP/Cs6/x6Is
ph3cYiK6K/Bpsc6xUaNaavgVJphRxsUe/bze6BiypCNDrkiGlSwBqCnEmVbsZSL4f7M3RmbGoizP
qkPSTgRFyNyvFUrXwJYl+JKEKMmgnjaRIMMS2/ZD76BJVspiSNsqvxuDmwj6p1a0VMi6QRrR+n3n
/YffTNplmmLXcBgWJ1ZTAHAg/O5t8OxAtWVFxYkARZ8wAaTksPWxJJUL2XTMuXTGQ1oCr5n+qZUK
vsHvHM2cJrxZVOd0Wj6hCOOTRypbLYt1qksZeCN1mNK+iTrljEk7vfdvCxGD+Lv/QgivSqtGeXw6
azGJa1s0EFELGqIMlCG1g5564Lz9/YKwS/Ai/n5imQBkvrJhW7sjT7fLEvseZBrZo2YZDm9n5baS
+l29PdRgpNRZueM4EwXceGnZ/RA0s4zENE+Kw+vYkkDPGx4mOjjdNVoBd6nL4RAd4DRpTDMVNm8f
mERloUnqSlbpcpl+8TEsgeb/YMJLbsWAkv2Am8rTH+j/KOKsSMXwBM387wwMDTVQKXzcioNhF/sz
gzFWQ1q1anIaNmmDYPHhHXsQPyThGo0SH1lrtoXCKURwArAdyrjwBVVqgpRenETvgN2Zh15WRtZy
H9VLcDqkNDE/Fhl5iCcTq+gJ95q9AkIhjN0nz9zIMbDHh2oEijlyXqvIBRqIqXtMBztZEIez9Bg7
NY19n1hPwlz84jTO3jVnY3pxc5+7ykq1Axy/04V2WNHvpg3KpUlMdeICMkNbhR8Q5LmogTZa03et
fP07laOhgT6jsUPnozmu2Fcsh3bxNiyw42Xg9zS3wOQZqm72hzlsTILFrhHx4smZM56Fmjd+aHqc
OkP+5TDBOQ4kLyWMjrZu50dk2/4QHbZAqbWfDRopbfly9DVfbwv2GvRmwwDA2HKlQpJjU9kVydaH
suFCmQPTJ1bNj5jkv0fIPxGNzd4SivQzuEcT0TKYNYaYue5d+ZHneAZY7SvC6F5gwf4bTRt4y5Eb
ipWhsr9A+3o7hnikAi3Z/iAKPiWMY+0jtRCl4ujUTVCY4+8+Rdf+w5uRBgMgGi6aEfX2jIVN7J2+
DfpE1yeR63lE/t96Y4J3oXYcG2h/VYzj9eOsnNQGhiiWaqkxze4lo8yb0teR8uIvLrOjiZU1Mnwu
2aicvLoDIDSbv6YP4oyY5B1FO39+z29GxDGli5T75Ulfa3BzKsslq5kaGTZ5Ys6JfEcUaXHP6hDE
Wk16V9xnp1qs/S/6IVoGhnPLbRgf6boU+vRW7IDZIpQSSQhflJ0Uf4kDA/0J9lWlk5IVAIZMkAp3
keXwAUr4ckc2wcfvB5wli82KiY8nds+kpzcsJvro5DX1GBmsIAnuGDNa/7NbmcOch//C64L4G2HY
KB86tBai+L2Gu4hTDuq9x0SlsokaHlT8/5cslHHqZiLcAkZepQ1xUi+0yjuEyPeR+1e84Sp3lTpX
k6n4DQWmbG8+0BlEtX4cwZHlngdJNej7QesUcyyPcxDRRbCq+P4koplTX3TlVEeHgj4eiTa8Fwn2
bL1sjbYJNOD35Ms71LGB6ebzdnfVg4OVg/fmsVrXQGDa6VyZRpou7L+YqrEeEtXDnEskW4B6HPHv
uhQE1V+hRJnE95k+lvLYBUnpLiOihpUg/48vkcVRoMkg5ao1E2v2WyYjK8+TvtCCAqiC2bZCUnjX
Q4Rvqo/ElzpM3n6CM3dIOGXFYd5GpiLT6CgoSJ6l73mBLScgJABMH6Kd4DAY7sDovHsifN9ABBF4
sTSMAPt04IukfxHrCMhWmKrGrnScyXAqvcuLbwKGQGCp0PJHGzMIZShwwbks93n3nVDVfDA4uEm5
sm2pcEcEJNiuSpTWmSjkrv/P4nXElVROjyEgf5oGKlU2kqR+cDlPk8NUdAxpacOAP3FuGukpnspj
8X7G/0zxBtLA1WhKKLDqCRGkukxKD20tyQaDX6vA8Kml1h3DdEyrDuiQXcS0dJPs1iXYMxFzQJVn
vOj8X1SeVrNDw8xpu/Qrk+lzwtIrthXXwf1kWpI6HUAOdmhfT37a1QJ0ixir8BvA8+NLJsOCkDUA
vqgstNFMzqsCyB+IUiIm1etbVTw6IAD2LbhThn2FweIJ5TwmMKIZhC+6LK5E6aQJ5FFJZuXBCWx8
U88IBOBZ4hFVfQi5rme6ySTAkUeNXUcnMO7N/9PYl1dDtyumougKdZp6mCAOy5eSU23nZuMp+oWW
OhjcI9hHUoxN1Q2RZdiRbz5t8eEOa8H8cE3IrUOBqLMh3Hp2EU+J+NJ8CcoQXfLdlh2aY3sTzkqv
57Oa3S9MQuNfwymSoxqc29xfGSnrApGKMWQd3HFhehQQruBV/rMRwRPXpGOihnQtTl+uwPw1YfQT
1TC2w4yI5XqiBCvT9AZSB1agvhM72IyL5eURFuMgIbm/YIQWuWwl2bNN/M79f1Qj39j+QXfpT8dr
b9fhDmGpE7jwQABMBt/AOQwjXWw8dQ9wJw3fItbvQfxpzOvkawcOkqKi08jb0E7qbV8dJjpnILvw
RUQ94KgLGBO7veG35Kc4lhwxpWIuvzeI+/hmIE8lAKUGLpGjORs/GyQasiRuF6RW8WYE00MaNQvp
/c1qjmn8FxSHWD1xjRrf3KIbAkK1rJ+wTxusVNmGrt3BCmffvMcigsjRRM+hX4TrQ27XkrX1nSzM
GKIOAb9L/9b3fUhB4lJzGS/WbqhqE4UVxPVeMRc5Yxb7QWeYMoN7GEccCms8FOJnSzjhWLl0MP4V
uPMEdbnlOLRLHduSqSHtLLTCNpExUQEeqBtA+JEIRFUQfppnM9qEhvLNg826mKo4UQG/QWxup5PL
s6Es/tYclhiS73MlXBXNZDwGx56IAxxP0gczprvxKf074elnOGdZEAMV2925K89Uur5AGtV9Cw1+
hw7y6nFprv32aC7M6aCVCXvjgRcho07myT8j8CyED3j4MgBILd5NTuqSS51ViY3uCZS9TI7E4lgG
hDC5pY3ddG5vdvXdhqj0heQQh9usOeyN9Oo2m4C0WTWH0y8bxNXxV1UWUsV4cjJN1uNH6QWovyG6
67hqBxIBIKL7Ox/vT2Y37QHyIUp3Raau9v6L+W3z7Q0eVSDS18h/l4peMJiM3OYSvE0Y/dGzbj7H
ZNbsEor/kYu/wSIXgSWzOogksaTX2hetbZT0AbhOWuc69pnwuLxH8HD1OxvuNfef1ppCufhZBkbo
G6IU//c1m6Zmke4RX7PPAKtpFS96Q4m+lAN819ae705uUAWUewnRt8eD9C+NENvcL0N0euVeG5Qi
yEDzfPlqEYiH7MteBdVD31x5itBbFem27wRnbl3o8TYlKi17pGw2P3Eqn/ioo6RC2azxleQstTJe
GhEKkYjA9ncWI+bY+TGPIuAiZNvpgGs1HKvS6KfMalZrQjswpjd7mxxKifpedgh+qO1hSPzCDwmL
QuHmNQ0pRWFdnBZgJm74JClN9HVDolymQsSmo/FCagV5NWlXl1FgwVn4oxiXg4qDEdgXyVi0gJF7
OPnDx2cTFqjRDp0LsNUU2f/U9urtC9KD2wCf63J+83HcWScuUfxBpf5dMakC+4LgeyaTf4cty3sS
vwUDQH8VxLB3KsnU4Tp2qxhYPnZytZcIxmFLPexjlYL2JO6xTJy2AKx9JxhNTz84ww6cX2xgjxdM
HxqdFTcANioV0NvDNByuxsqoBykAOeFXBg/GtjpmiDDtlDL4n3b5AZy8A8T7r7V6h0j97kjUujSL
qSsST5H8qi5oFOObxVFgb2JYwNbjWJc55SL107rOwvLiyeHNR5FukGu2hD2ZpowZ676zHI32jpFe
6WA39JXDkUA5dnij++rohEnm4iENYcv/fi4inzTUTrulyJ9FY7jb2lJku8795mf545rr3/YX371I
8hT52S0a8r+PlkYk/gyObDuiiUlmW+RCrPALGx6tGKSRq3nYoVsxIUWxh62oitsp9x/EL5rJRYAE
OaQJhnj/bGmmQFpUthLqhjAAjstXZMk8y/6IHhbjCHbaQ0xdh6/LpM9BBgG4Bjny601lFVAB80fU
k2VTN51LK914siDEFQUlaSgE3tLK8liPZlmcjCwHF6rp/NGmkE0na7qsZjh88ZfZKm22dXo4F0Cl
8exyj5X4jAykesU55vpCmdSoib+6RT8CjcMQ2rEtZ8F9FMGNaeS8x9WhSpxZ6WSBZrKP/uSzWZ71
FwRBft7V8ExTO8E2yXfhUMmaVNdN3M/ShpEsoKPrz5j9zYErX/QsbR3D/d9jhDdka0I16z5dARgA
YNzXbFmWTjw8+xNac+AawlAxsX4NYw5+TVNdpWHrl+qDtxo0vw0RtlB0APC9oiAzkjJ/ZLQCXoiS
5olG3A9XYEmcIUA+3cOTCTXxJtrPfRxS2WogQDNvTEuxlN3vX0f21otPK2WDZdp8EXvdpORQFICB
OwFBXK25y3ZfFLWWgE93dWXN5NfViR4w8ZXonIfwbSzRNuqaIS7BON07Y0IE0eViqLfzGMggBv01
P2vbaNJ6CoUYWPcDCtC8govLJ8cXvnDwddWxU9WfLjgakFK+Gp4hi9TQ3DcK3EdVz79PEDaYSvhQ
sb+t4SShUPhKSpFqEqxGtlmzNgEFzlXfOyJMR9GGocuWUGxpp6HF+UofnCTlD2vS9kgnMjjy0fvB
fXNWH66Avr7j7mby6qyVJg877ojKvsDx5MFjteanFIpx01XymWhmZ2pUG1ePZr3k5nI+83GJqeKO
wN86ME85hXLaI8SiHDTbcwUuhIN85OOWGDVjUarJbsi6JyCsY4ygndYOvqQgoeJdTETZarJSIKHJ
FOLw8A3qKjZbojAH/zrfPWERAWsEwUeAustMRLMPEO6ENvR/yek92loKu0uQ9qyRAu3YTWBOvnEE
B5t1tO6vMBgkkOfMWuivZdPYKxBSlADB5bBF8pwptjK0pUx9cIfPkDLYbk+yGXsrS0PrY/BKzsA6
Q/YS0RRHLoiwoYGTmFvCzU1+EkXW222qV8iR2meArIE/lpgYtHDUo5XEFAHwnGLacDoksCTJoDga
xVbMmn++GykP/GeER1eRidUY+E8HnOw65YgLhMHYCRSRYDFDhNwj92sssR+/DF0GZTWakk15ifqg
FBLd6LVBvvoPn3oUG1FBviSYDq/farGBPPES3Bk5RGCTiYrHQ5+s3zZ+sw3IhYPOaqYtBg1ASoac
NjFh7Kr/02QdJj6fc2X13tE4b4GKX9t6R7ZKSgLGFLTRnNiAbOnK3D17p6xH/HE75GSBk/QE5NeK
1r8YiCoUJ+FRw6J4w6vfSb4JjtYNWXkeci1w3ijYoPzcb/R51XAEBrc/gdLZkeblK0AGZ6PJqj4J
Pl0/9hm7qe4Q92h7zfCvwxxvAFsxqEX9f9E9WBsGWwYTYiyYhDkbgAqemZLL3E3Kq0fcoWd/oM49
NjwFiKoX7nl0LMQhHunHXCmRW9nozs1kyIRltr+IDHNfzw3wYyQR7c4F+O8C4uxJpkF1bqPmU/y+
9KXYZEbWQpgDB+vl6bJ+5KMq2PJtoyAknl4XSX7B4HfKKRT/gMPt4jseyS23vZ5DXnVBhTtdOf5L
iGdeuda5Yvv4GKRJDR8Dbjv6JHnHBkYE7B+zSXZ64FEhup39IPsBZqSpWnLY0D5GHcH/GYVyb2N9
vCiDltXCg1Aun3+JIoPllhfJOSXv8iHtDHPZx2PtUTbBzZzl0SZ5UVzaYnB/cXyV9rG5hyHN2hnY
gjUzubgkOI+fYwX08sGLSURclrWn2is+xIEpmn+NCIIqFz4qcTWNL8qPYZxAGB7UXb7bETrIfKwv
7obu5XvhwJ0PB2DwArTXDrKj2ffihEmJnjaMZs/u3B3r5dbs8udQhyO29pTudgs+ai1BvM9sYqp5
1fujtlS2OJG42yhFvXubiQpAAJyjdlWrylAxlSmPKvNRqgBlhsZxZ/nq7SwkZXQ65ykeS8D2a8u4
47+aLww7RHopFXQ/x7ixVB7WvMW+ngleqkpEQBsTNCCJWYXp8HX0TMLI+qr78CLR/I/0wx1ZINWe
DVpFjSurPPxRq4sK3HOZrEXYj24pxZ+qK32U7l4whjfroSs5RpXCW2iRDc/pbOF1sXMZuPV3KNuD
JADOv4q17giDgWjPNGx6S25npSKgsxL3TFoP2i+9+fsh8IJQYpEAHR6HEPFtGd8nYxcXHIdMpD9N
perQQGnTKr3xQl+JwVRNkxmd1N4iayq0ViIOl9GMXNjr6L7nuzIfjHykhb3VUFOzq4lRzZRq3JEV
EoajPKQo2pzaLnmZLpPR3Dpxo6z+KkrGOwVtlA3XMyXdwfTf7NH9nfpUULAsE5esXYfAMhFBMkcD
BV6FUbo0HovfE6U9DkwAogUPGWonFCJgZHtFInCHUQooCr4WSOq9/erv6O3Q2IMQUFDvcrbqRern
oOq4I2yQZTtLbmCX5I75Pn1D4KfI7CUhDkgDtrNazgWwuTM6XmvQ+mrUaISNkeOUjEYRT8Jmkqm1
yip0yGRw7XGvLroVLRFITf4Yafzaj7A6Pv3ORvPJZMcMkU6so5O6/3kjBymbQqqCLv/nr1J8Vbdr
eqltvvLWUkzL4SoHvIK7XVqLN2dS8AF7xv+Y/jsSyGXZhd4IEU8pe+utMBmiFxW9b+dATJE5tx6T
iFsoyhawRmWHd2TvqAW4YqCWP9z9IgmHkOdVqliYPjQL4UFU3oM0hK9KsHM0kWrLFNOXa0a7QHwO
y8zLQ+141zO9ZzfMNdCZQ7q8qsjv3IDpGg+CF+SKEZ5oPaEhDD/C3WBwgY48tqU73ES3WxsVdtC8
VRp6daG/6qE2LiLP4hlTfQgVMX27r9+Te2WXVKKeIVZoSqkvfxIiojvD+uYE2wh4PAjqo296Qxm3
btWlTR9Zj9TuyyuxSa/233xEk6NP8x52APJC2MaJcQS4njMKGj2XD7gjeyBG/8SawLLtInx7qiy0
e/GNV8MtVwJIAbhONTUTxA9jEq+92nS9jaKBUGdoBS7rIdIIlE4NB3bc40qsYDKqgeSYIJaP4ymN
kftEPyxH9DxeH3+XjyCQvm5y/Am15bt1z2SkQBZ+eVhq6gkkXuEwAtLbjOz+YHLhOeFk0gqI6bRK
P8AFepRCzfHGfvSXe6P70oUTJXQKmtn24VaGqnBSEzVDdE1r3lRvZXYYPd0Igyjon6JOu4BXrLfG
+zK+d3+tLoqotgZXZj6+D3G7+55Yf7CNMWHK+jMBR0pBX3kj31ReZJO/3qzlj8dsPxNi7NCF8thJ
NotfppqYfKM75LFnqqyOH32+9BbLnwOSbRChjUarwL0T+M1DAQWcTQoy7o90JzcEb0WIUq+/Dj63
JPu5Tp5cK6X94ejx6xy6J9AnC2QYYtIoYxFxzd2wkoYwgy8nPID2/2LuRzTTG6F/Ixp/MjuoaJri
o4/KDahS9WT6RYdXE4/Atjk4VSyhsBndzLkO8r1OlRjp4kYSCDsmrtR9DYUb7lbcyZoCTEmrte6Q
8wxlS7Fm5gu3oAOsN5oK5kCz8nzwrlZ8vlZN/2FGYyZsEIw091x4uPP2yjd0Ykac57PRwIc8NYOt
RMXL0lErZ0I0YsQChN1tsUEaceadGMgKRmsPyMFRYpbiv2y+fwAqLHU6JBQncgmDRSCCEEjWorjf
gK/bXP68kfWQGBFZRPo9+dhNYZL3fI3xsJYH8onYlVMWbrTn7i2Ykc6EF7amWeNET8U59OX4kdf6
36X6d3La3Id/n+G28dRj5+IWTgXDnIEG4t0kOoDe7hiZwIBaTLESGoAfE9o2KesFSb9dW9y1ePe8
9auVCvOYzKuHnnLbrJON+RIQGwkjz3PV1wXJNiBTWjbDl+znEB4o/a6Gn76wykk/jk6wdsM/boQb
CTmPE5BCTHXzzXfRJqsPSY6BWBflUyW9vfPiQb1dFRHQ8b9gFrUWxzTFdYpy9tqWs2TUSMYaGuB7
f2Y7KPNsAcAHt1BLepMSYFEnQZrylx3LVsV9rgM8Uu+4cUxXuif7lvhN+p27D2xJYTXsfafUyw+T
niHUEuuz9dzUxda43K9watj8yUbVYTqtSmuMla0ZabWm6RqsIlYzGYOkXDFhS79D1RMIhG+TWZT6
Ze5tDNinJjNIzQ9k881ambbEtJLdmZMP6H4J6M2V8hXXtWV5Dci4ygIZ2TUAhUYX5/sbq+0UjIU5
7wQoh/g93mDyOs3vRF1vtcduI4ro8D/rxwiEdGj/cAl8nXkwz25eoCXgs0KNmobxBPopsTM0xlzr
pjuZRXiZyx/0fQ98Rxhgz7bkAKINAQk9DOoske3BRtQ6B8+73yZofl3gEjmyUWfKqPDD9ufJvM71
h6zBlzTZtp45phDcaLPhEl+JwQtK+UPMrmrKSGStEHbODIqIG4P/nRtWIAnO/S0Qa2WeKXVgcvBD
QcjfxgqdjcLNjToa+vnev24787/F0TAVtS4C05IvzBAoNu2d1dgwBrlQyK/00z3xAx7sNI9cSeEU
Wl6uvcPo+OmBR2eNbrUk1BX74+O4XVCuUwdSz0MK/WLSDM1+QWplx771sNj6IDjoRrBf4EpyruoD
QEoXNU0JI7Y/XQHu3WwNNdl27Sp8qIGEP5eHdoX0SfkseU4zqoJeEMGDZsieWohi9eewvbV9tEeW
S1scyqKL8DlWI/PAVrTGS8EnC2tRHgWl4Ia/lWAxIen23u3ofARjRcTBTaSjuzSh3q6BjvO+YvvQ
47K4eKCt01wPogAXfnV1HJrU9j57Xav1YA967cIDVEx5+hwhrT5xtgjfSsM9j/CSpd6vPOaykyYs
L9ZeiV7+wRZFEKO2nTwMWCPvKoRFbWwQkzPu0fx2ToFQfAScPDg+13Uld7TfVr9bEe68XQKn1uS9
FkuPUN2c/QrAwmNIhkZu/rtbENwnW/KlFsD9y1bMQytyGU06lAmDbfguv9ZBAWYJ4KKrKaiHsUf6
6DicB1k/Rkf8wRmHzecbk0t5TRO3aBF3C0IsFkVyYsKw3a1e89gyagRvijxCtpaLlVf0cA9inTcf
9p8Rwj+t/46awUCjlyzjWrEzJ28XmNnABNiC9gzdE1oIjTLnJ9h/mjd1G4VMTZn51FYYYxUMJnZi
tMZkQfTO45rDaNaJFdNlp4ChqUf9+kigCCB7YW1FkmtjMYgDAY7RlAMcR2hZDHLre4xIntu7zc56
zeEsUCEke37XdfrLPu7FIRwvD1dauS35bpoSkz7oVZ0vY//l5N//3YceETdQ9AkaIkM9ilv21fi4
NOb4xU+UmSprQYqsaZHSz6tLSCFRosalbIACnM5ilWW2xGx7xsxgAevcjtGwGsTSASkqEDIqR4vW
hz0IQK/xvqUWYMDpjjyWd0A3BsiQ8RVAr8c8DYz7Pst/gomDVCNVA3yiW4JGAUggbkmWp6ly2nij
i0eVfgOc6MjzPgg+M7LNJA4oP0XKkkZ9g2ovIfyupdQuB+E5v0HjySqVztDh3MlsX6KMCIP37Vg6
TQz8kBxs48p1kIcZ5rXmO2ZCKy37dleHtyHQs2S0kGLcSIM51BCMD9Yxxat/ZPNGqKhvwRBs+/t+
1FrlWCyo6YW1HfFNT+maBmzYfWdFtSzaw/kTdgBtzFoKzRGWkzzwrjMtfzU/InDAFZibhBE9VK14
njmMVbvvp2rEjjUohVYI6RG7wQMHD68qfY9KpS2xmpzQMQDgum1HypA3FK6bYePS6xkG7ud35HwR
NSspZjLf9VrkZkAK4stbC0Web6GnqSwgy4Go+A5HkpWhD7eIGk2MdDMGXo3lN822zi2aUHi3vuEf
fuYR4huPoDO5hBsb379t5p1o5yFhc6bskif2Gx+vzTt6x7wNw7DYp2mdrFEvtabJRtW2X3mNpDf3
DRw7nArU7GjFxn2M8Cs3rC1mqd5LitdEq+oRlJ7HqLioDh9WYWzZNj5yKl1xktiGT+yymPrG99Gp
K/1NpybzePAdiJMaYKOSnTBAtwvhCTllKTvE+lU6RUuC5+oGhXAXK7kklCXlRYBEs0bS5n44ckiE
RvgQOEeeU8EcFa/5DyEU6w4pq85QIKSW8ZEax5eMvVrxt82CtrNyAqb6Iucd2t4jJE2YRLb1nWqk
wg4hcp8l8H25+1IRLeyNIXUYFNLDRiWIeJp5i/SYOWfgO5GvolVSzVMN87bqcxiMhUBzdJFuLVdq
aWjfrIQEEWaHnHAzApeP6z+CAE1BqyjN7xBZHT7mha8klNt5WyLRQmd3NC5kStiEpzxWkVpmvQG4
djq5Uuak46Ks5IGaCJZJP4sDYbTNBb8q7oSAfTK6XHYBKAvlWJSpPZa3fPlj3UXq4hPQqldqwkjO
YNBYIT++p3E9Ltrqqx2j7TI4LD8tFG+gi/ZNLMjNt/yGalJ2R/hkLZox55qeFfUNGZOgFMBPcwQS
MbGtBxEGURSk48KWPDUWMKYJlvuNHASy/l2VLR2aH3OgNNtFGIRtbwx3EMnxm0nl0sxXwwejZhrk
R/h3UfPe3rLHRHhdN4YTUmmh98MggMe1RrmeYSU0NwccJCUthKzahAaFQVx7PSmrWBoajpidNwmo
lAaL/WZwURjo9Yn78+EJJcJABPInWh4mPxfAlSGO3WdWlAmQpionc37wjPfvYHkrQ2VWbNEMpOVY
A5fnmnKMihyAKZUECUtCXQNBerzJgY9NRtD8U62YezgTV1EtwMUfauUhArn8JHO3BX2lv8dfaPwO
uGDsJSt7TDZc5g/P8rQFp6tLthipIiY9BBjP/UazZdVDtr5CcZButwMhHS/I8KJlsluWwb4g4mHz
8jcSgO1Shm9zmfVQ5OEJ1TlaED6GWW2CKXbqpC/UF1syPUSpLMm5+i+FUEgOtHNUBu2+EmZ/Ae2S
970ds39xH5jNQYSKM/Pyc2UjAAxP5dLS/Mno14Zhe8DmD0hvf+VjJcs2EktxH2soK1toY7ruHmHJ
xP3tqd6+Msqu5qEfAlCRlWTxVQaH+FTnX3KOPI8YA/9KgRrpq6hwDrLpJcNl88ZAmC6bBXpz5s7h
UGpyrp4vyk9c0ZElvGDXNqnicechJ+u4q7YXSd78cjVNRDO8fOKRRCt8nGqJxSxVgIA0gzMlURt8
oGcbLTOohJAO8CRWr12g9h29o7s8WzH0tLHuOAL4LnIQ32zpPKg04o8lBqoGmGhi6ykhiH0CmuZR
EQV0+QEWd76D+lR3BeDCPBKeeRCi1W/wh/+uQsZz65jdUuFBktAXiMq+p+yvZU67wepNT5ysbH6+
oz3zsKrOPqyZWpeDY76gEVPZ+INGfLKXbXivQQ4nWF15bLqdCgyYePCCkASGXdmlafyc9DmaA59o
m5FgMYmxK770xPR7dvn7rQFjY5ZKRr47c6i5rx9NVV0AiEiCnsIAVRx4XIhURvieyihSvGT22aGz
lAe7Dakl9f9llGVhpXJW2BgVhEe/b6jWpYgsLDY+0omySfRXOmjurgtEh3kfcBHTcqQGdtbd4QIV
UrKV3nBRiaZaiTwEHcGEZL+o49t6GmD+d9Nh0Qp4M+iG9DKWxAkNb4aL3J7vh3A1ZJKNqqMMY7dT
GNJVOG1muPI/+4XiM2kVlX1dSDBJ7DF0tja0FYqms7b3NaafYDAvtJclzSmlpcLrSOdA917tH6uD
FJ3OPk3Qi0Pvn4RfpqzaRi9LbpxLoQcKuj18Q7tP2mRWyOCYAAms7lLV82TpnbLlJZWA6/1RjTTR
+sY/Voo6vxD2UyU2mV2dX+2P8iUwikhJ4QwvhQA/42ACuYbMhwVF6cWpx+xW8IAcbucTU4CqD9+4
P8PFDUGEOtqUylqVCtEItn8Awiky5Zdftqs42KRXEocw823thp8VjRpLRsUvK5GhN0zqRzYk2ctg
yhmXkpS3SHtPfbrRTFELiiqsYp6Nl1H1VggH5MkpNe6u/Lfiq/bQBUm2h7JFYMK5f4sOEaPL89II
28FdfSDG0ZRPnTeQQU1JE3LCXGiDbWtzAM1FXjSsprtiEkh85SpNFDzLK4a8Rw6yVG/S2fPzzKTe
5PwNXtgSXxg+KsTkHkxUEEc4R/3d/yfuPd+up+FTexNd9ncpi5TLBJWlcInjKpkT80BVkwNuMkP4
EJojZrr5ifbePA8szmuvt4XflGG9Bjc96oOo0rxVlJVX+y7AHqSONfds4ePU0Ly1I4nlhqhsK24U
B22EQtpziK3wV1bO9ior9pb7tTFLxJH4IXDosK2NNBfc6b/kb4zXqnASrGOAP0alSo3FA1LHFi4v
97B/DigPxXHe28HNp66EyRPtXk/qFT5USFhHDc081he/zDKPXpE1OAhWx904yhkSoBog2yCQRukn
ryGIV2WsOexLw82bk1xMT1CwDdMVnhoZgkWPjsRJx/N21cmGwG2MdgWWzNNvcEbvyNfsYz6UHK0t
EMWPjrnOQmjNAy10+LdXc+z3OzJmtHyf6icrvr/yhjJSFHSzEnKbTw7g870HfjMZ+nbSEuSXYggt
qrmQ2DnfL2rZN/7wy9HYTiS1jyvtd0ig1ByTwmiYxWuI/D/iaO318c4b+NhMCByQJ9klwlrUL0S2
3pr7AGV0SWtXWLXZCXZz3MsMtt0ieOS0fq3u9so+0doa3UnztFTpn+H/cTw5yOAIp8ox+1jpk+6o
bS0WxsGVTMFXRqMio1fgJmlIy2OtlluZzaUiqoRiJzVjQnYt9Vrczu481PdZ+mZBK8tnigkaPLKW
O+eEBP9OSPy58yDZwUWj+ZbwHHqxxzANr3AyaHKF8xkzAknJp/t8tlWh4r6v0HRl0Wq9dP+DSbfo
rYdkmfKb2PdKF5bUeHFm7Fy7irLyIsKlXEaGgxWHqj1ZBYPg5cBvcJ5UtjlfqPELK0CFyOMJgTbt
6brhOBTmfMySxtHulNbjOXuuCmfoxDnZYRsd9izRI9oF13plW0/yV82Zk7UTGOsAgDXHQOV0+EMW
bDsBTZJhEb7b+gMKZAqcEgA2fmAXTS90gVJAEH5h5bUfD58LFU/tDgX0JRV2zhUTKl6wYu3nTt14
5jPSRWTqIWRNwXerOE+qgAxR/X7m8Gcs/vIRciNMNrI9glrdipchXLhlEkgadZFrBp1m9hvYT574
tSBxh9MXJa93P9Y7WZvJf9TUiWNZP5IcTQxXYIkhOpjdRnBIONftGjnAP6URCHUld4gkcxLjcK3e
E0bRFc3je6qe8LychytllNq2zioEwyxGuorAnJ2DCuSQ3dUfR34fCFoJuNGyidpBHYXp33HmVilv
OA+ddT2OK/9GMcQbCW0sjCDNjLYloq2s65LGCxgCl5cFHyK6EbNES+hQ0wQb7mm6/OTEzi9Iu7TG
BD7ToYeSTfOg9steja+Dx3J+nXPRnPW7ps/HEdJO+3xWLZZwulxKKgLr/bQ+sAQ8Sct17sevH/Vc
Oora8MDZHuxOz6Bz8YBHPsSz+khaw5bB60ZK1Neg3dM8UjkUdfxcxnwnYuPHX3dCgGGgOBeumsTL
8m6Rf7rfh3wOjS+f1bqm/er4dCoq+I9bVsD1LiNs6Rn0wORuYPUlVWCpMwlykJvvqlHkYVU0xG+a
bTodp6xqAaATS7JZ7JHOZpqE4Sgo1ruCjDa4lmICHaSGE9dkkAQ+yJ9S1W1KtEAFNfP69FZVjyw4
IhpB0RAjI/tLDgneC6AUHaZjnmf/GtGBlNmdWbNBpuTxNTnTqyecqzKKqaIgEKSATlwykdlgXMwn
oKhaDlQ/WTNEsJGPv3ePvG4kx0B/bQ9LiwgSADh4As+7ehFObQSTMHEsnd0t2wVI5YWWmVo8FlBW
ekzKzhJYfRyWL3jxDYhkdk0aoRtUH7G1FYHxI2HbGh/GnjazIAbBlZzun8TycguMFF0D8rBGWcwf
T/QX0Kt8OYt0xIzPdfkYGCYYjWsaoweNtVrsga0saFq/4E9cCgjL7WNNdPTzqA9EP0AJBUYWnJIS
flNN7W4/mXUmLqdrSdevvaNUQmwJa0OGTcz5nVigM9rDxEb4H2hMJHoRoF8Ld3gxC5xIHR6ur5wf
BzrRCafXrCVkRIDU8TlOntvHmD7ItZe0nfznEuLFNNKZxNhWTki1Pog4bsiHTu/dTWpGK+l/Vg6x
iBr0V0f6skHOeBXvXE9CyEuAQoUJV4EvQNl+iraqFOpHcru06aWONhR+stZIjg+RArdQrrEwC+id
oB8k1ESMTSJQDgBUPyxOSN2n04yVeZBegK16ysBFgbmY8z9kfQG0v4UsXB/5/hANcFwdjs/iJVnj
vdyrl1uJrDoZAdC+mu2Lxm3sPebxMmmer5D7sXmKsvXCU2he3cXAaYfa33NUPMqiHjaRPjR/JtZx
cLu8TpothKDCkRT3fOkrVK2OAx5btGjVGBh+UO/FpCsTlSCjLC9P8FLjyKfhVymyYm5FrmcY9EQf
xrC1nmY101e4EnNomKj1n64smW7nHlNSCnLgFt1J7fzCzcKaGRXSr0F3YNcPOEPcIIoUrFmrkyS8
aTqi6ZV0mayEgRtgiAY6KtKyTRB0JVS6wOVjP+fSrJDiwRbvX6NNNGBi2fgrl/pK8CVcIQG1i28H
J6YwQ7Vxi58PcU0oiKqWSHCXKW+x4sFn/erj3RVytDvHJQz9on+T0waHB1L0BnSvlD+3h6LRLE3P
eWJR1JjSpZ3L5SkjnZJfVEctqGRDiikmrNAebNEd+hRmzjmbn1eZJUiJYbvOWfyNO20G1Sno6pcJ
cUAGAeYjhjEz4q1fdGyccW8Cpypf745ta+nXBNc3yQ1F/ff3Ly9t289jvy++MVzq64ptrGqMtJhV
4dJlR0/CH7LfYos1/gPj+/LCXrqjQi7OOudq5+idkfpX5e+Qzf2gxd1GF0q1Vq3WGCy1TJC0pqk/
YTYPHc+9ReNyDfRVzq/ohtHu+w8lSsLepORrpvVxnkFgBGSpaOC1OOb/3dXieHdjl/dGfLQLyATL
beTVP+00ZhjoMQLLe2q0s8DAoZXA4KNo9eJ1ke58U8P9jVKT0NfF1DFpOgf32qmPnNtmHp6fviIv
ZUCqVwgh75XBWWSYB5ZMWQkOdyBdsTzvJIZvqc9RuymjP6vSnxtfOdQi+1Pd7gQCZ2L/x5PU8HUX
axrRKipt6VBA2a0QZHOHes3jYWD7RHy9cD/qUvxlUHQsyBMuErnrOtTZLS67BVSLqGeHBV8U8EgI
ZVNHucl8YgtZidHWWsI0cgZo3p4ESElveywPvmzeo95q898e+cnfq48701+2JxbsoBdULQycF0h8
g/cxfDeQguH45No9EeEI0YazpviMKTVO8TpQ2IFsRbHw0Pawr9k/yyZdQHfA9CpVxz9eDiNSxr37
qlDKqrtitK/89NEhtU7rgrvMUpA0b5Ru6ACoe97O5Nzd6bMdYHHeP5T7VUeLQVSJRtkIg852A7td
NVap68oQ28AKjGzclIdZtAtPGjtSb1mJrxSoBXfxm3fl7sG1j0iqRUyPO1ILgkf+nrXfsrwp99Qc
WVceUkkrGzfGNQiS+GhMZFt+P0gLvoUqCQvWNpV+N7pJOPFJjJ6F9IvHIWcq0xBOrSpreXHW5Rd0
FguRSGlY9UsBj6MJGGFgZchiW0AL7RMCJghjNo8UOWPaG60YAtxwH7spFHTQve3WasF+s4Yxbg+Q
A5Itt5zzpyfZ7aB7GUig2FIVJuXiWuHwuO8lotYS33ZWEUrF3KGSgqE7EEoso24XcHFzrybmitZR
wIoy3DbQXYmsi4oxVY92dJiUrBWxxKSgDCujeu29xPlqYkieoRBRvH0bQ0miqeqNUCSKF7IuhPjs
FNKYCnb+WR64HEXmWQ7pTvQtw2KyFt4g/7z+HGvdH2mpBjTkTqNV2SCAES8Lrr0Ii3RGCcd8NCLr
WOnQSlkFct28BIQZ/yCale12F4cPYUHAYexxGt3n4ll7cGMfk9E3LPnnvFM/GP5n+3E7DZ+ujImR
cDn/dDfFxgNu8wppruwRJTgoTQpc2fGkYNXhzDyRzBM8xZOHVnTgQPL/z015KVh251hy9YSsv+59
4J9Q99bf4FaJaUQ/a8jn1vthkQDSr6xF7Q1+aLjlPGtr/DkHGS6nymuLrX1GBLo4f4XO0Dnt3AE8
oU2k2XwiWp4DkTtBwkgVWJXokbmlZn7FyZWZ1JKNPOdZi3nnj4EVa5N3IiL9wbcQR1WdJrXxtW+l
AvtZaocXBTd5BCaDAOjd//WAEi/vF9FF/YRYfB61ZsXVzEEIJTa7OJvWIJhbeZkj9+vEwhePL9s+
j0wDwS09c9Ttm1ec+VFNuxrgxKtEscF+mwc/rdAakfZH6WhmqYwF/sGeop0vTj/vMxskuLxfFLEB
hRYRb9QE0sCkj4EK1QVmIBkzXamHmuj6DJJ5wqdRrLNLP3T1IrzzBLoNOgkCkGDD/IE4UbcPeNXk
qDdd2rOk5fDZrulwJog5ilnJhl+iDgWbEFORMTTyobTicC2lqNC97/crk83DaMxWOPlUcY+H8LoX
/NSKwKA7+yjoA+HFWke0L624ntnECRQ3uAqb9+nhvWpauoDN28Xw2LIZ/gAa3Spo5co02ihl1Hrb
KDw8VKJSo02XOa9OY0gKHJ2PyGD0/sMSAvaQXvEO2Kp5bzPUpL26pvxVPMf2fQBVUPU17AH/BpyN
r+L9mMgmvrRqyMTBMmhCS8ZBTAv0hq8DGxCTuB1GBg3inECjFZ7G0MsgbfPV0HmSQgYnFcjYQHc8
phT+9w9DPNLwEIWPba44zxjIQL8iYy+JXV4FbCZgd60CLIpdi2KWrDeWmkHlvvY0uyagt7hZD1tT
PjltKVs5Ma580aS7Vy89hNj3t+L3itxpVfyoj3k3QYYaFa5sD74w+UGezldZauDy52uRdbw8JaGd
Np8dwVY3a1UiQOkky+ngfX7PwNBB5hGnoooKrLLQYGDOKJfyNMFbB/pUtUDWod9KLO/g7uC3iAVX
Bg1OQmCKSYwKCFTY8OSiZTuVr/MfNr0I0qeU6ayJDfQODKOZ1kUoInCIlw55g/tEHeoFbRf1/VPd
imNXhoS+I6GhZEEpDSxq5TiWl4otAwpIu4eQDGyjIS3nh4vZUxHocbxXq+1Jwb4Frc4vCuVnxubv
gr/jFZVjtZNzbfcWnotBDkRaqgmCSskL/0T8Gas+QQ+ry70y85+CWlvSo77H5uqCo556OYYAF7uq
lXT+vR9SumRdjqhHNMe5c8/96VzgcbAOuYEfpG8+GsGSdpblfenAlPVmnS7G3zRBWWBYhUPZU+0L
5f85w7hGEcGJvmqQGfBEEWYgahNU/f0nE6DU7e6NU/u/V1r3HR9YCG9YisuHT5baeZmAZ/+EpiTZ
eUnuGqEBe1Zq79dIIehjHpzr2Iwz5QfmsFa0RTJbJWL0tFzPCSTc2yomE/bNBXJHaF+PaRB5P0cP
tXyIRpZo/UDbINM2cAvU7507W/VpxouLTZVR1C733o4pw4+Ms8o6oQcb4KomIKe+GI1CAyiqNbfj
EQjQwQ5DrxNpvwpt+fJxJpxaIYH9vJU6Q1HxL6N7KF0rYE6q+Z2uB566zuXltCsb7qjvqXGG4Equ
+hmIDQrwayTxF6UxWMM76mAk04DhbRbKDdIE7nu2/OoAaIRTunIZKMxeJBpUGBF5n4mRceYN7n+K
TRXvJUKmt5piU6OFSJvP3yZMZJYFpjJyiVF7DUu0nCi9vB2vwl7C2UvPIZheFTmac8uC6OdtkWQA
WPDsO22NhVndGYxxHZb9z+8TNUXwx6v6HID9g9W7qZSniZyqooAufukY6YbvAqDjxTTVujNQmKLG
84SnZ/Ce0XC97mr3aatfHJzSa36AZWhO/xd+K3mnxcg9ULidgZ9vXrCMc1TUHi5k8mWlnsgPv/48
AsKNJxLpT7c7It4SB7LicCVjj7Mtp5D7FGetWR2qCywqxrKnfIpz9ggyvPaLGrhUWHvtJDYOtGiC
zu7wh66un5TfSxfN2mpYip3WpSu5DqDYsIeyhddhUrwKzEFbk71Ayj+HanKCnnFBTb28VrjEQ++b
VkZSfEThTusaLCZdQ6JSv4j9nitU+XSpnXPkTC1ERQ7RAX6ik7OUdkrcDj3iC0aQgGv3F/LFdLWI
glCKeavbhQFCauDdSU69ph5HhS4gjWszliA1sqNFZ4kkDyM0R2Ruecxu1KU/qIEudLOupl7IsiPU
3G5hnYg644sj8WTyexxH/XG3svwuV+OshUWGIhZE/dCMTKMepDlUnS+vMBK8X5/DWPCIbA5mjkPR
FbzwcZhZFFRoDGqkfbmV3QZ+gtQwcyTyjCocx8Io3UUVsGh/FbW2abPvcnEnds4A2w9DhdsP2tWE
ezhm9Vv4+BpaxAdB3FUiEzgO4bL0VQ6k8VQ2Jt4PakFKfFnnLWRDFOk0NWujkXCPJfX514KGiwkg
Bn846H2QWpak//MzIV6DNYQk40jkI9LlXOnJRVAJiZPO+w4y1yp80H/W00QuosDEhLiAeep4fnsP
o+l1rojSv3ClyUqlF2qM5LjSmgtGPJ/W1zPwg5b/5t9IYMFXGO7w/LrV6baPjYvuf/NhxI7Bs4ZX
y/92QiVsMVLMRgTk+LksEd6awE5CbqS+4d+E0EtCFLnkXzHaWZ7+hmNszvqDBc5/8sh+yBYWh1/t
VSm8KbdepSxiZgtXUJu5v0lPDwlItqU7fCXViKDUR/am3+Ba+1gHOeYir9emarojk9YDcQZ97da7
hFBYvEOeodub48NSlJrdLfSlMjWdiHEZ2qNykDoxThsa20gMjO0+zYyJUfUZnSyiLJhyHAFWSrg6
3uDQjZqYGZo6Y8Jd+ZuIjG8XjomQ6EVyPOLjmAxf/ZVgTyhaLUOiDA6rkmmNxtHCo3jb5A5gDss7
aGGG/ILv+Nhz6ouK7amicn5vTHg8ItJsRcqwC/0CTbBEHJsfHIYL7VtVuUitlQ3G8b7e96BmjXNP
A2ulGpaLaPSL1JVyN8aQNlinwPu7YZ8zgcf3W6kgM8KFqbYCOYz5qPytmYYjTpItPdaFSGoc/G//
YapZ0G9YJ6q/pxX6HPSMSyXuxdpNmzPmC0JPtveggSaA4jBeycI8cn8r/XRxDq1q+7bTLZyTEEXk
IyAbsXa6f3VzlsDW6Nhg7uP9h45oSBkyjDkYvcG/oHtHjYHOFYpGmSySvZg/mu6Hfatiy4mWLuoL
byNZwLUNw3zvplSaaR2Kui3mwLZcpGnKOYJPApSf3FzaDVwFFaoBQNNkK+dfBgFpL/JNnsRBayzs
l9IpHtWuiv1IyQLMRp9fZFXvsdHRHrTauWswRvY4z0HR6+gBEQnR4G2IFBNv8jECQDBh4/MVyots
6CiPiZFx9RZL4Z250j8WF6ugAzEdylhw5Mv4/9qMP15m1kXm+iikz9v9+8o1bIbk79a637wBFdie
EVWIO+cu7eqPr9tYioLounAc9QRXKIYfRCq43OYwX4xkL4hjU0yKNrUwaMDtQz+202MvRGE9EqqV
ouVf3mdRRxr9OjJTZ8wDuBXLaR4NMRUwJGK+Nx2dN/wPfmmtoO4+QtLmS0lfif2FZM/i3MQtpgt1
jPrMd/JvzFEmG6hWNjgwxdFoVwljfPl7mXwfCZVj4CygNxI0n16iaGCBCZBI9NbE+/1i8Z39B3sb
qyz2DA4SFbUR/vBdSyXEphgs5jAmAjNv9rImEI/0yHv4q/ZI/aGmQqTTOqeYA5JYrSEf3zRRdnxM
vpxFWhJlgdxNMqUqjoE5q1hWLF24muXp9RDjpoyRjo8XPA5qpTRz5WTZz2YQPm+1YqSv61qAjKH5
dQBF9p/sC05XetNbLlwxw2tTVROEgVKZYajqVVWzZGNNMOjbps4V7an4NriOA0YMtniPM5ZYS6MM
Ovmss7zaf7RKnQ6hjQJNm8v+nVvDArxCtdMMVgZkRoWLETxyvw7OII/Jb7aa98Yn0BT+iw5jR8Zz
wFBRBBJ42PQgz9P9kHRdvCth8ecsY9pv5B/ALssSCiTDplAPg8KW8pTDhLkxtruI+fCa2oaDOI1v
CH5NX1BjB+51TItsxXbCPzxgZV1jK311Ni39ZuVUVGvyUgzlTsLDevA/SK7cQfBCEBCM8ZuZTeYg
xusXS3wt2XqkrA7Pcg5E2Bv3IWOGbFmgVLZurMgrg3WDn2STmzuf3ASrUw/KgnsG9yPu/lqCPixG
IFgdlZ2PKdYY/hgE09z7sKVexpi2S6GkHLEiIDOlRl8+ttHBFH501dPUldJu9LRgDesPpuj/7rga
yjxh9doXQmi49dllEU+Bs1Ghf/TExGo7NIf4fTa/SKnWU1nzfjtjo6Sfta5jkFcTJNipUtE5TJel
WkuJbQkppAphIOXuPCW2PhWW/O50t4YzXXSNukgStumibz3052e+BpFYQerhuxHDGr15urw6ep0J
/PTSTChEkb0WHsRjq9SBzgbLZJRN1CPQ96HcuwaXRg20Kp5Enws8MAVxK/Uz7JXwSWxvUfuO2L2i
AlWCGIa3VQ2ZhlRI2IK8Kq88NL3+wMxbi/aPyjvU2SSs0a7VOW258pD2c0eNlmS/w8CZzM7nY/Xc
H6sW1jx7fxBlcEjzIA4k8kgn0WYV68bhfW6OsMrNz63amRHN1oWVQlcI9SfqVzHts9XXXNPPSf+o
kEFU4fCuRyzAPdKaYOGbF4pg/AL2rsmiCWJufl5M0ejjkeQN/qO2ZRUqWeIwzMxh/CXEHfICpvhh
TijAthUzKI0YfGhaEswPakJOoMw0L+WZmM2/RfY4cj9X2q/wRDBTkpffM/nNseB/BLx9/pNsh5rq
FtAcUCtRaVmDVXCSA+eO7sKi2N8xdTSLQQXfD+hLtgsGO9/tKbDtJfE+x3XOMiCe9NWtc441cH8n
JppVlEco1n0az45BV6D+OBnUKtZMnlzD8OsiOjiXsPE7+YoVp/wHpOM75h+eWGqssmDmVvtep1gp
Zs4G00yWlNwqFZAGdmqv6ocLr9+fumUWx/tUq5S7D2BPJdw5wsR1cSdbbc71i1rGd0yUqkI/2fZ7
r2o+heB2KfEBDoeo2FVQGlrOZAx2x0VJDAuvzX5WUGyrPJ8ri7Nq9GXESJLEwS4U/rczPBXolvWb
LU7m+GanV4jn88dhMSkqiSiGJdXXCTym5BZAisnuq8Gc58wyh1FEuRZ9zrLZRCW6pA0xFLV6Jq7N
LYB+d0UNj4gIOaKVALzk8ZhoVZP760nWhmbOSMYO+LcTA+9EQ+EhwT3vNn5d5onZ1mCbpmmmsf0l
QnOB9vq/glSHLADStXeshXVX6c68WZHA/fmGv2tHThALsHVOnV/6p1UiFmppOrQAUCGhFgA8evXD
qLbUGBcrsp223hxvKfAN1iOFacpMW7OnHXdYXmYX8j2e1lmWq4e3PrQEXEct5vpWNWUT1N6FC0Pt
in/IZDW4l/qBqDE5SckKo+fiM46DLtTSkapsxyFXCZxQqCldGCWvfsO1r3Gk3i9DDOqZIRuEWA8A
Np+vPnNu3HMlRHG0Jnia8m8WXyFq/okADx8Xxbh5TVJ0DRsuN8HOj/UMvRCpI1Z5VUEB0ySWQfYC
K6wQ2vdXWUS0XRP2mHNj/AkvRGQbd1RYG0biMbTS47BOb3DYx8ATIwpHrDZ0aeDcqvQ5/iwP8Cac
jwiD8yJwxVC6VkYgTOf69Th5R6FvA9VXp41JH5fydrEvqag5VmWhhZDOeZJjS6SBwgNRhqWrgPER
YDORqn+8smvGpcWeL/5cEJZ09v4u2Yw79RahbBjVDzNPl9FZlzv33oQjoMJifGZ2kYRW6AqjiERP
4tfKz1f54otpY+IDebKyra41knPRpAXmM3yCnQedw6bLgcHqGVKNHbMa/a2DiGE07TyitOBvn7HY
WQUNepX6YprS1ja2V3MpICX2p8ImjpDjJLCF6cwbES5XRgkEEdR/NRCdAFSXpwM4y4YoSnBHC1GJ
bmEro0FEHYUw/WnI7K4o0Y4wNjqZvMOuhR4njDQOWI47EK4XRLEXTMu9nImjx2DX2Bfw9/bv5CgJ
5qLsvZhF6sfmU9LV30ow+EUGTOIY8ftnEHkrsPnwCrAomyGMLUivY6TSsZw22F/5EBWLGi2F0RUQ
1Vkmf0g+Sj+AKtGAHEoqSAMOOXC0636szWmlmqlXpVvQk+S1qXPEOYe385zbMRbDTQlVb2ZgSdvk
MWPiRQaMaFHPPrj79MOVmfiCiMkPr/zOWje6NU7wVIjWddCgNeHYWNbDPaUC5srAUl3o7xWh1gkL
BRR1P/HwpWGbswgA3N2EEWBzQAHcjlQyIEECZ4q+ZeH10xJNWZWbCkVLW/k2S2KKz5ZR3t+Vo0iN
nNofky08EhXvBYfNTNlBZQLE1/vW9vCduB8OqKJQ1UESWRIWuownwaR32FdLuGjFTZcM7NgDdoS5
t1etkLHuU3kb5NHx3N7Ed3IulZNpXd41IvkRc+jAbzomcdOmcM69NaTqSAIumGhzWY7LkzK0ZGMD
e0DTIJND8amj54f2OklaM1qM5KAJt2bX6DB7xyX//IUbYgp5V1IEg9athCTnKYkSWiH76ocLnqRY
+rVAfgAmtJ8Qyr6d37ZSCE7pasbdV8IPg3dk6R5Xxi4559Rulla6UHrj3swMUq08fy7Uvo4RmYxD
NfDqjxT6ttqsejueAGQqQGAx3F5U/m6GAnNCjCHxQOM1oI+Ao0rts0c63PXmzxa68E5Y353Ar5eF
iN437uRQlO9zKoTCAk7e0ICI6f5ow32iaOdnrUg9q1ffqQv2i1WAckcKJpGPZ/03Nt6pt+iMP+LU
18pwlJk67Kow25yXxMAOFARJt/pyrZ9dYqdqaXmsK9OryXC7oLYYR3x2QHHSqxANdwMpi9d22JSv
9Sz2Kf7SqS8YIYc25aZY+pZ8mSyMNRquGMTZiW/353B9a6TVtl5rP4+KnEvo9T6/MuNp85elGGlf
oIuqb2xzCXAWnICUWfBzyEXPRLITvbN2m8zHR9kqEvW69A9INxfb2OoHYs9Cn0/CcWjxDxilKwjZ
4lGyP1h3zmz8lRabjPe5bTjMVo0b6rGrCTSGXMt+u1IvkSMPTN/5QxARwkw9wtlvfYb7KvWjwVeU
PcnTCvpTxBCsNiHwuiMB4ExnLZaUAjZFPU6ahhQcEDvobd6QgrhnA0FWCOMyJCbLUFmbkhIJBVkh
XirYAdxB1G4sc7ppv/9bBP+XgdpVTXNhjx9tDGSIzRk0TnFeadm3OU60B0zFwJg/bjV7ik39guY2
NdxROTysKIXwE4AND0ZGCGGMRuv6g2SHhRFmzTlefhOr+q9FiT+DW2DUG4/s9k7jCBUx2WnvHikQ
DLMvDRglIk8any6G9JL5Bx8lgBErNMpWKLN3sI53s1+zAXYegQ9KbLDvkfR2XXZcMNr8nXdPEwRl
uQb3EZxFXuE0ZOTAtwJNNbPWRl6fQxbuSw2kRsoDR3s2wrsePYCkOs5vY/KvTkhNnj5wl4iJPMBd
+fsAjoH48WLtw3/mLU7xUOtaOr1XlzhPSXqXtKp5CQfKaID7zlq3YOTqEc7vDf1sxMj+Z8NRgY5Y
x+n/2HKzHqd4Yab4OjpDvAzJuEHMUQ9ZIy9JmngB/ow+IXgiFb08IOQXBr/lpLeKd2YiRiAilJMJ
JVxGspR8/wWsGl4cteZ1OrEovog5Mmq/tzbU2hxVRsRj9p1MsyAyQdF8WJmDgTNuQqvJbX8v6qN0
p+QKSOggX28UvlS7oJB8qdIqdQmDfxZsJUC+PWYrLDRPtXMGyytOPmVYrjIcDUHrILzAy8oMHNuS
56RCE5w1WzKb1hWtgaU3R/HqG2GcfQmPmKxxAp1JFK1WxiFTzKY+iu5oh3pQMyo4ZCe4A9RYfhwo
yeCg+LUg7I1L6N/XTVqLRAEGkemnub7X5+jYcO/Yxh02f/ZnZcQE2IF92x92kD0Qg/vuBMVPSTgD
65hA5y2Jkiiz+Il6y8DV8XI/95fX+rZLnAS93H1C1D4MvR342OKB1fmDD9wOL+0EJtm/ifIxkcGP
SpDY9CFR16lazlAWFpzcdQIjSSmqhSRLqa8l4ui9UcZNIbPKk1Fv9AP5kUChPnIOf3CcGjNV2OKo
s0OeawIvfnc5sD4+TUERZ1Kagr0/N8YP+D03Oe8rD81GBGqCZQhpPQK9dMmK2XPPOrg8H2wc9A4q
srSngNOtg1mmgUfidN2bMxiMhaw27I5h9psYs+5NDFHFYEIk+QRs3D7KOoqfFiRV08zm4SVwCuDP
6FOpz5ubmIgWDryKEyyiRbxVmKBtWKiP4EBI/TkdcpELqC9GdMTMVQ0XW/ApnLE/bVlusg3ASCR0
JXdPi1IyIMlJVNsDydSzCrRUGgt9yT1fdBCbMpx1/HW1lPEXKsFe+kp7f0p4tSDteiKYNiIWFwJl
VKlwH4mHOmSUVN9/88X2uvjIh+8dLWKuGfJcCoJ8bI3gLda0gRxV+BWwFMh8QI299aZ5PKYR5Y9B
DIrdwJHnlmM3AC4wpMUF1j9XjAWER2pSWngIXClEB2FUIPXbgQhSh/8KhoPdsa+epvkWfeYExEeI
+jnQhZXhU25oqONfpdathJag2VuYhPOK0NHzzITsCmC9RATtfZlDquRBZh1eQhAvfj/4DMHV4voQ
opsZdBwxOoEhS1zHDTcmsEkjaCj4VxeKZTlbFvr2Eex/kS2D9MuTXavGYFfhIrpUhV0TSjYSuKMB
GSbBrGoFJGAu6Xvaix8SldOjjnlOV9fj8mMjJoIa0x0mPronx8VSu0sceiF5vrhgA6ppF582faSk
H/4eWX5oYEnSCqWevCT2NgD5dyAW8qYsGLomwdf11aJK4R/+SxV8BtH9jrFGzBhDnBvWh/b4rw4o
GUYpZzTFSftQ0HsvZbaa5eqAl10Jc+rLb8gX7SeE/B6/8om9PHZhB/dpT2ZJLMLg23yN8nRjA9vQ
K6uDN1O/fEyH7oiza0jeP+MjailQ8iF8msVRW3vADcqG397aqobG3SRO/+kYYTARj8oUw6DEvSvZ
MxTLUt1iHTS+wjwPV2kAgUsZ7ly5nbVi65+6shcWOFGWNgrgRCwBE1MR3M67xTX35nVbXRoxDCYV
q7RcKS3lofCc3uXmqw6Ld0Vf7jX/tu0gHv6kbv7B71/H+YcUaOAodpJIWrzEd4DfNrI7qMCzbown
l4SaGg1YO6JUfd4tsLw/8V3nUul+TTlpuvF/b/2pV/LGADjQpWBHIXNEax8VWyklvs848GGShBR9
v/zy2mY2dHdgrBF3IMfQImQTldd9S4WaPgjYQIA+wfE9Gjcsa1bEPGyu0z9FwRVwLYi5DONqM2IP
H8ryl9V6xiW0Pq61mPuVbnSz0YysuXg6BUke5wY5A+8XfmKiw9O1qzvWfahLobStofjzrAmW0UuL
mi2Q7/B20WzuKkCUNGGNe3P6iM6FcMi8UsqBT4HodIj9YMkFPulLYodET3wJJggorTvDN4Yn7KGe
mmYTbsZBMawpRF//fR5u4o5Uu536WaTdKfeffy25D+AAepS/fd2+Gg5d5E/JASerrp0rN0ydWdMp
vg+z8NOpzs37wbGrBJWjcVMeDHS0VSgWWlvsGErhibZV9q4ImD3l4VxF5tMzb18nEyRD1FCAsc7x
vxvoWEOCEm/rzR5tbKa5z9JoWrHfJ8V/mZLfkYNXhomNVkcAHgYoemZFTizo5L7z76YRmdK5mC2d
c2hoMlQfVWPMz4zU2qZPMYhlVQOzTKt8K1xrHYUjb1lSe6F2+qGCOnYi0NgTe1Say6OrmiaL1i40
EBX2bejK7CEbXvdGMJ3ZulHLKRY5Ckb77m/GFsRa28mUb3lFGWsAlCuoSla9OI94RQdLNLOqcnX6
aCFHBCSTGJyAilnynFVtJhuSCQ8PyH4lx7KZPqhyu6bDO/Ut/HK01/2umbsI1riS2ywgoIcYvF0y
OAffJ+lOLS01myXRaT3MtZeT2c7pMLa0c90jjNzJWFnb5nUO7tXmOazHNiEoPUezhopCLwXkG9eu
rg7J09dqbsXPVTgzNF4adVkuzk2H7TD7iwmc/XOpMD2xLYaLuCulBy4J9Y+b8+Jlpkfn8qXUoI2V
hn8UL3lP4/zWgAL6iS0P1WYNB68rEGrPP6A5uE8mCYYr9e1rULCJEJX6jgofj4trEXv9bJ04T77L
5LARQrdPUnk09z7ihoRi/ny2Gk3RYsPkND3ZkpmjRGNqpRG+Q0pk5zOrnyJPYAmnrk1OS4zOjdUg
OJuO5jGCzBMK5qXcYheUAJCSxi8HR66jWc3Phe0oV5MJoviK6gkIWwVW1rx0vhTZyEnir4+w/CQt
uhra3NMRnbWovho6egHOaAv1Nw5I8MYGsdSwDuVpgLx9APuY3/Msr0J8a0m3WDaMAT2QsZD7gMi3
+/VAXz4aWxtuznMoHpKvYzos0UfeDL9q0hFxpDJ//gB1t6DGY/EnsbD9SeKwlGeADeSHhn38uWnu
JaMdvWOvLJKuuCvxBWk7+dPOtEv+4DwNb2MEbxEsbw0dz2U2UsZcv4B6FQ4JlOTKz1sr9pwzFcl/
7JFwN6FXG7mgttNs3cPdZYnf9rtI1jMM3rXlJ9zxkT8zDGRzBtYu6c5fs0VK55CW3NL9LfQquQr/
kTpau271asOYAg2y6L1zWr75iYaV0ojAJaggGTlI6xtjy60+K0IMvGrvA4YCEDpHQKGpNYJo90CH
TO0f0mYHZg8jB39fqu/qWw7QKBSTILDv9Xiyhti0JFQNEuFXlmzO1TP4o7hTaJoZZsWY4rbYY6ER
cn3H6yrkAJ1GDmsWQNIsOCUVt+d7nLPYKq5aOhxUv0Y2poBMBrBjLXyLPYqc2rbkNcoU2+Szg/5T
AVdEO9o6EfsI6tlJKyQc5vrdiALoo9kr0ZVJbp2UYBqTn/BfAPZxcaeQPDO1puEj4k947Owpp7HZ
AGsGsFqz9WGeoaAVm6xVibBfXuQSm3D5J+L/g7NTLX+N90S7rpLbgSgXgRg7rBVDxzUH07umLMem
h+LssWcq1O40nAQucdvcYBPbuOuAEfrTFNjfA+Hp44exee+ehVcQQuR8d8+fkIRoageRPrVxKdfr
uMddp5875deVQwqP5zZcUkmgFdNxSrpMb5uK3AXlbzvpHQsdYv9UCOtE90QU7R+cmnyFPKhGAW22
CvmqW4keoF/k3qTnYTmrGqvGAJJmnkDdRirnZTB/tGYw8Tj7j9mtBxnZ2ED3Gijffb3IiLoAA0PZ
kCTxO95jmJxNUx8MkRlDtsgjbBekV4/e02MBj3kiHs7bEoCEwpLWR9DQncdWKEbDqmjs+OpOTcTF
wK1bKrrOr0usrC0ien8Y2dN6IpZMO4ZLIKoEj6pZpnLaRpeZ/E52eqQ84Bno3cOkRYymaPU+8bf3
/HHP6VNZdpDLTaVNvflwB+SsbeVD7hNIsglhfDvgYj1UmewmthveHhiJNgdQ956ZxZgS01jjW9aX
q9r2lxroxBau5hMrFS/Ntncw4UYdgNE+IccQz8hNwttDEicPgKuA/Af7BiCRfM39zsXL5dEp1jmD
ZCweWGjaFT2j6XuG2DCwW8q/oKo1kl7+ofAQstnWB5eSroKvxQGENCtgtXo9o/L1U4vqbcmkBszY
P2PazuIhiqAq/bNqNQe3bLp0sOfvVBrOMRadlZUlKgMXvp8okiCn7mchylwfULVaNy5PIpW8N9TJ
iP5mAxGaPXdOToSbz2HgsLn9eJii7w36z/7TMwxY4CrcqOLayAGnygzWsldImM9B8DuRJ4SWtQag
aIm/joH7jal131ryuEd2h7RJhp5OX06yIiEOzTSzJMRkzRI6/BzR47CBNsoLQJ/IDbFwy9ArGfaJ
XXi1xk08wp9YjzW2ymnEJR7vDmXdspaXHQURKIrh+Mzfi4TTVvlEB7PD9btr9qhv+RgWRsl36bBU
QNznP4NrcXyplB0ods6g7xFVjRQPG7XZJGHiFZ6vhKT7GC+acbDAHB5XUowzjODM+KcUHlTqTcmz
YmLpsKzp8qa13tL9jX+e76tpeZDt4LNXeFljMo1rOsccrfDMwthF0Q1Dv+ZohTNZJrwvLOywfHqK
M5ssC/vTBKVpCxjlF4Ja7b1HN1aqsa96rVZoZ9u0ZuhaMaa8U5F0hENk2NcZTZZpeM3OKhKg15ja
BEp9LN6Qdwy19d82TCdXCQ9DIdB9BUUzZLBcdHzJXhMIsMwHd4Kfe+V4+J9jQPVqytw1BVOf8RjF
3sxwFmpFrbQA0OAk8orOZSx98e7N4Gyjvz0OS5QFlHhKpYsyTRAOvYmUdy19GvPXgvgXXfuizFI8
5fdE0X6+O6Ygh5vBusXJjN9Lp2AvqNSVZWYVxKOs9NRcvXMIUsOyjBu0AaKEodxG0Ml9bwLBNiOw
lLy+YlibOp75J8GjlB0QXcz2kAonEgzN4FOts1OjWiL3g0gSJieMsoWYS9w3u6MS3IVi90jCkHj2
/EbIvkN+hTLaSoNRwvsBEs9nwHznsVa7bZo4cz7mNFlKTCMI3dhnaO6GrXoA5vIwcU4k7gtR9C3M
dMsBAhmVu4Z59Ohr1UV+D+SZpb5eSW0tuyuyhKCBkpylCHvCbCcsQM/ra0lrf3kywnwS0/eNWTd/
bZ2NOD3u+jVQMssN0FXxKV3cXAESrJLJ5+/ZySz3GgzoSmhsu16f9bKVHCGz0G+DRiOfSv6Smzxz
xbyWW4i/a1wF6Jkd2RncWbVPKkT1AyT8OiKnEu1L8+WBHTx1qv+ohCdwaemVugN8xQ9mURC67oEG
gMwr4qeprHyCnvaNtdfRNZTcdP/bqguDYmgCL0a3D/cLikRRrs/Y0JbStJy8CYOE3T5N0eh5qL2u
zC/loRjt2TQclHjzFoIb0RGytWepbxZn9L1Z8+w/G1j6ot0/SqA7OO7aQwbvibhCgIzL8YCGWBpf
w1EEeCcvVt8/W4v/xd/95H8oCnZD/e71EKmSw/4jlPCeddSp2Ln3daD6QUF+5JIImcrYGkRDXGYP
vejAu2IgTvQ4+yqG9GjRGKV4O3LsNjeGj5t/Oj47Py80BfAuKTCWGHsG75HbyV51ZXCNFY9DSBhZ
VUa/mfeXrGGZSFS73p2Y7pHRuEt8UglVlP46NBCaxbYSWe9DauvYbX+LcGHtXcrk6XKF+eu9IMbA
ro4doRLngBe0unCIqqJFte1dr/YFJODCxJBD6YRZ3ZjEvLsPtEFfWwWiS7tqhJvwBJeVe247CGOc
p7vypdbN/BinAUvtFxBgcyNriQGrFYxGK6iJGMfPgCFXqHdE4u6NnKYIh4O4zPXWAt+iD1y7I056
mmPuy3Kksq4hyMvrObBVBC9YzRiK2DOCYacSpEHmxPDaIZqtugOF3l+AvZhDjlE+VskxVJg4qvu8
BffWbFnA7PXSz/00rQM+zINbWbvl2qOrvqJEXFUG6TqY3ZxXUSY/rRcJwy37QlO1bzliGmJGthGy
tc4S3nP8qfiPknD7TJxAoiJEChAobv/d6mjuT52b89hssWA6I/5jcCYLNA+712t7S6/FmU4j+Xz9
m3DYBfiN+K+TFDyPy2CkEPncvroxMjYBFhGYRoV2GYDT6RtC67APPy/c0M2/ayyJ70DHLC0e3KSD
IoXXuBaDcvTlYPXHdbtr9QH1vrhwMegOgBytxpa+gqhHlGJUsII733X5LgL+fsowzRtP3kT8Y/IO
ntrtMq/9wVjbDxuf4P++62qIyBZkHDYaMibhki886/JM/AEcu/IB6heAUdEQvhuZlFUgsOdY1tsQ
N6t23PgPegEoEId+jrNO/TnSZF3RuG1vXIvGodsencfsO0xouGwOfSGaX1v1vWBaJoxlT0AHx/q/
1uR7n3HGBJfeS51JA7T4RvmruXlBx6QyweUt6LIm24//w9Um0Wjei5lNx4/p3MDnxv0GC9xeG9KF
Trmc++fgbcuRs6W1/CtoyuDdXbFVAbdJJBP84+PdQAYhqcK1schTnY0DFP2rx5a1IgTA1xiinUd3
n0scOrlHAs2OUJNvMqYV0/ETjc/lKuTIEk7AmhR5pfxVcnpTg1XE0cJRO5zgksckw1V+GQBAxtoe
gnEcZ/eHN9jqNfQRJCMtPwNbL3Hsj4SntWftrRV+21E5t+TJ41KPC44hRK23Evf9l77VFdXZpCSp
iYVl57DAOoyGm6i6zfhXmebrxZLfk0xP1zuEQ8KwbWNKSPxNYBoovpkLAqiUuZQym7k7zSe4VAkj
Oo71cIgXqyiukpkitmFTCHe+cnmYDniiCgEnRqoghK4hwlweZ6hsDq6xFNaBhYfId9OAENVSFNbd
PIymmMSAs3sklgDBKljOZwYpZ4gRc9+XvvjmZe/oPoGfNJNxlsl+an33tCK6fXREXS/xDUJ3jnpP
WBYC0MnqM1a/9sJ9Fo+eQ8Gi6pb5fb8Hxd3t313fpa91JwM3iGVbk81JEw29IkMB85yqp/UTCyYU
8MJXzjthuArXi5m1mNodGJ05/ZpyR1LnjaBXSdnXA+5RIJeacgJab1eZVnHqrLrnKXXADGfzda68
Ag+MewXzuVShB90vkKdnd4udc5p88+1JPd/DcjSyvy7dhM4BKa3r70n5h0Nqassrwxh4CYy/owMw
1OZO3p+sRtW1/fY9ZWbxqYtAdM2XsnFu7fP3cMx1vmfvLZpdTKoV6jq0Umh2xvSHxuU/ZPYKvON+
brzUewY+IlGt+9hLgcQqaSJW3E4NbVCD1e/pisorc6EGBJzADjS5JSaSa5YEkYpNO4F5UU+1yzdo
V6CzAPP5bSZUpMCHKXrBUiDPsolqrGAgsfTh+5QO+nbA3skTVbD5cbtnXoWyiQl6kZzIKhdL7Tqq
f6iz1alfWI/VGsGkDbVFEbaW5cTNksXzaXk6GuhBCD3okb1QeakX3fJi2kIhIQhhIEIUcGGvqFNj
Zswu+0xgRrbDRLp+tlKDHewWyVd3tL3Gr9qLjA0HIRekcwdVzKmBA1JhaIFLsjR84QgNf8RbKqsf
gG1geUPscSH5CkMs1B0jAEQbPIDU776sd/8X+fGzOQudkrEcqgdNUSZ/aRAbT/0ff8IRYBn/2FYT
J91WTyCA4anA8+FPNAcXZd6M3Doua4To5tFgVqwrCtFQ6F6W2rkWF+Jjgcd8iNiJ9RUbi8ht942G
Q3VwUjp+uusL44bc/NGQpIjcuZPWl/zS/0+GMWbMVmnb+HyzFF21tHo0qaRIL4TAaDfP5Lw/LGpo
NJSSBchaMV0o1Bok3R6w6YkxMnsnBF/ftR0YU4grQsws9CWVbTYg9kaRGbzWPmT/S495Ap9KK8Yp
mxacpBgj/AduZ10JQ0cx7XV031MSYnno5aubVr0QQUTdVd6J1VSGLcJch6R/mkt7j1+IZyMPC7Qt
gMWE607biXeC68nuqV8MD33HmLvSEvWiXuNbjPSRjLiTLHU37f4EVibII1JyipW4NzHckqO3Ca0d
Cxua/MlnNbvbaPMyNwppkjz5QDEALUmKWkBBIpIBw11Vm7RaUFctDosNFfVlKnZC6xmzVIHUI8yJ
r+uQzXmvaq9QF+xmVhD6UNefrlVe6/Bny/Nj3PaY15/GKB7Nlr37Rqd8+hn0O1SlIfk81SL+KCRX
zgWEAi4SQx1vFwDS6gF44FLweLZF/VSfZZO83wdgR4O8IyZWNIVGmc3fpw5U+aOeDw21dra34la1
EIpMfYUpl4eArFdl5FqYkw1X5fZHOMKgNH7M9Yq/Zk3Kisa2oh42dah0qdw0AVyaOb4XbUAYx07T
WqeE87v9Tsri5XXmMGr4Mkb1uDzSReJbdIOR0ClqLcsOYAUesCoGkXnbEmTSmYsJyS0VauR0YhH3
Lcnm5158kqjHqfJsTo7yMYyMqQnzvgYmFUnx4XO4A3lmLcYk0jCQvqWpx4o7ofXf+0aeOz61WzYS
mvZjQR/sRYNCmN6GuQJ0FcXmnOLV5N5o/j9Qdma6kb0Gtuk7L7lAhbQa7Tm1agKLiRbLAPa0ooGv
pkFy8+Oto7oc8ySS8kpI00rf/5ly4wQEcKq9ynWocCJ9bVrASmx1CxTqle+ywRJ1+NTNDMuVVPk/
vGeU0SOCJ5jwdwhYeSkQYCw8PszlM+TMgewoqiDCDMeRschcuhiFSulWc07b2N/VwLpK3F+MzvOE
X3k9sTfqqDZdiJdd7hMwIwfbYQ6kmt/2UuWBw6ErerL1FgU9p2nmaKeBhhTyukh1nQu4yY68jttU
HEkUBWNqeGn1zYHFf9eNO8tW9+SgXeZXlKDFra6c3Sw5GJS04A1alCIHRAwvMpcSKQR6r4oTZfyO
wgX6NnysXEmb0s9ZioZY18LUPtSzB3CqMU+pnBxuVbkQe4whDIysQKIpkIFOd2FTViapFwaiPxWe
8ILNsZhyX3bN2V5vwwiMCHs0NYO+rK0diTA354H0TBIo3AzOOQ7UKK4p0UYkgIMGs/Yi6CY9Kbp5
51Q9nKjfpOaOSNZwpUvytOEjhV8HEdVGeOCiEsYTkjuzn+QFqC9UyLdprJeSsw9UDXEyRRdhE4Jd
PybnGlB+oGEY0R5OKY3Mv4LbFfh4MK+ra/nPNbHW1Bas2Hg0OjnbMnIkKkWkGMrXsBr8+dOTOQTE
YSQwC2/58MvztDIcXjpA6D7nN0JtDnUgXyMObkpS9tqKIQFbCsYrhcdGxGo/KlY2GPaXxOm9FRKp
q3h+gJCBJVeu0JDEBfQRRBKuC0LMrhJt5kV0T4y6ur4PYAkx+6L5lhD9/MajP0jVK0y1spknXY04
hU4yjZ98Tz2FAiOJfIF9E0d1a201qnW0qt0o/Pd+vsKMV3khUUQ7qJQ/YJhrhqrHa5RT4Wk+pjZP
RGj69B/2hf4Fb6zBii7xqlNKMZt1TWJ9sHdcC3Js5VdH/6DHkkCmT/kzwwTRAsALJHvJ5cbogBDW
PsM9OVw2aYcoofZ6K/i+ztRR5mAGvIVlVlFtMePAu1NfeRwZpaq6aa6omku0txSpJSb56w0/GcTB
2r825NTTddaNpINynXs8sqeZ5snqtdW9fRz0GhzzPvSjUOOLLfeNaCwqtn+fgboqcZVYYV8RRshm
pOCWVDvkG1/uhxPTGJXnoGFHMqUM8q/LRhB16M/4JL6TXLyY0GEeIRc9w6OLv4e3E9csBgWmJpqh
yxNNl5GN+VFM+YMfnLvup72LQan7yJ5R/b1/i4EN1etSKC5VGaCpsJ3wgMBWXblgeg/RHLx24pnx
wGsVRU+/2ZDB6BWkTw/cLZ9R1cl46eV34tUjgSYV1Q4wGXAfyeBvNO4TbsuncKtlJpvInU97I+4Y
kIRO1lOs2WKVg62DJH4dOJcCx8n6etON/YZ8CSRi1wMoZdthIPvL3Gc4w72lAtBlofN6aNQh2LCP
k4nlFi7SZ0ElsigD3jyL9Ttvc78B3y7lXjqrA2FQPyU90Fh5VEbiNazeAr7B6VcelBCHVXnBsWOp
8B2hMEDLCBxa5jcSwyIwP+O55BkyvBBnwO72PWkyY9ymPpBvwQlv1bYu5QqGSxrlF73qNpyXxb9/
/Zw9rQkdzlMAHj+IxJJ/YJRjEw7bwYYy9gJEtWsb941k7XEM6nLKoS/Z0Np4VsIaut4Yxj7einFj
7t7iVLSEMhdxme1Ffq9EIeAIta46iHtXT6dWlvkqxi1kmFSu5HFfHn8K7y7VAvJEtYKiqaAsPZ1z
m2JQM6pe4aYNZjetPUl6V4/U1MY/KtZ6mC7Ks8/0OA0i/slIhYIhnRQve/LQKRlCQglYef44U+3f
qaybvFHcekaraiY/9nhDourDZs9ZJ9IKxoJtgMxYZinsPo3nsp+s10tmmKVmMuu0/a0t7hOXgs7n
/wyQJa+BKTEUiJuwhRC2diSonqq7tVoVqXX410gA0TG1lYa91o0fxlCNc7cv/T96vH8VrNg3YAES
Pgcah1LyJpvPDB1FCLNLO/os9qijtAkowc6NOnOnqRdvFq3XkYw+45p6OB7uUmQc0y4+DaPkig6F
rOFNhBtBfTvxvga9zCS6B2dzGVmD/dyCHcllRCUMhnzpDCnFmZkGx0TTNEMf+f3mykE5o9W7kd7Z
x7G+j57ti8lT0R/ngYtGlxtkPXcu4sMcpI4CloPWEQEbhmJnUKW/3jIA7c6GoIIJUG6QG4/XjPmC
JRl4DldMafY5Upg1H3KbZahXL6nYG8owNn1Lgr0SqTh5fvG5pZhBkWSSjio9ECnbbN5ogQPqwAWI
ApBW8uIt6UZg/4cHtHswp6Qc55CKvHdUFOAYWqEJd1S30KQsMTrri20hLQXliPIeU8YgSmAnVXx3
JbfdD+k3UJghOMzgQ66QRghuK3ctd2mUR99rZGzzP5QkwuvefdNStiluGfF/chidGoaaEo4B5opK
IaEp3QgJFdR1xQPbeRJsMmcwHyTkftdiT8pubB/sgTYSGNLOde/uJsFJhGzk7u78QF+noKT+JW/R
Z3frKQ0/GsCisNSiRpDRO05An5euAwDw7JG0R8JAVZ3xxrE5RA7jP4SNy0xA2BnPtM5UD4cMzqQU
EujyCXV4ae9bu0lUNBzz76T2KHitNA3kNivXo+oJrMD3TmYQfSUa74jjXkmLZF1AI8LL1wYzuRrz
84nL291caMhXBIbwcGqdETjp80+2TlkEr8X279nitTvbUMpvYPIDgswr4hDPoxmyyf7nPD7BLl14
j+8UKESBZA6cvP/1FJL4g9iKKzlfT2ZyTraEwc4JzhDhC2kI0+0G6utoEoWgSUQu6N+9dnGbGNOC
dqmUjRGHFlX3Qh6NS6+pzA7m0/X1tHC4HNL2VxpLhMjiuVPBVMoMrAfwOwpffhZHcrWa3iqeO5ey
0IVbJcS+VuTBzjmu4hNrkNweN0b0J6nLbikYrw07fwwhxXTKNKUoJw6bbHzJMmP80knmPb9gEhTT
noaabHpqTvQha/0IZtrNArx1VJc69uMKXyscfXpzh4go90y6MDwh6aWelFvNBVpVkNUTv4qvXcq1
daocZ64z4YPabbQJ8n8Rwis768aaLKdmTjQxszLH3zRBHtYpKMeprD2nfAPYYXxd7DE72c+7ZxKP
LaMj5+PIQyPlA7A5gp9fkd+HugKdipoEmmraDc+q5+W4TExpulDQTrBNzWel7yVuB6KobKQ/qd7N
6AACUOCe0kP9R72IaWal3kimEXyK+24tZCN61ASKS9dT6L7J97sO8W4Qd2OkePk67laO8YJp2SqE
ldPJ4bvM6giOn7eA6xEfVfkt1K+/S7aXUdDNhbKDOHJ52pFnwsFeV+j/QYByiw4HMa0GoWB1uqkH
z9MDzvx3iCbBipy5yrMF6Drjdp0foscfXK8251B1d1PQVDPVBNHDNuu099wimgfIQ9iU/hPT2u2m
ZDXD5PBSitSIs5XCDP4yx9doF7RY1OPQmYpmxPU8c3t8IcwKV5JdMB2AJi+TOQypO/HjMKpw2H3t
l8DaYm94nLPoTN0oNNnM9HwATGgeTzME1kU9L6dFpku7hATG+LXFEnmabfBT9RTlitVxIy0DJCes
GBkdJSqVlWZIblBpJl98/y2KbArNw4NAJRHZJJ8iQma6lmGEmst38DFT2jv8HHJJiax/PUj9Upfn
08tojKBJ/IHgrfJHr5YsIa/DFYlB3r1Egjy+zA7O7y1uykBPWvJkFOg9Rd702TFK5KRutsPrlPiB
osXTqm76xz63GIF6Sg1YSRDRzzIoLzl2SbcY8mEfwmuNQe/Uq/2TkfypBWHkSgTyn19EtGIfzJEd
qrlpYErn4fDbjrjKAgBx7qqN6QlFU3yQfOh5BEV+slBauZZ4G5C6PNZI234MsBQklQ8XhgIoshKd
LO8OMTfuVaFZ8NiNsh3zIZCZf87Z1kdXQoKXUWVCMrEiwUcH13Lnlrj5MiUZM3t1bIrUzewBa/y5
c+3fbJcfLgmKTb9Ekd6mZgqWyPwBeeDK5nQBpTcBwcw4PSxT2ZVT/Mew8Q/83IEY6HJ+KzFtbr3X
KcZjf/4J7GFdcgepdLGG4lqfIiHXazy/JFtnex5Pxnr6pq/XSwUUmo1da5lKXEhmw3VNwFZuxpWD
RPfNQAkJKMAiym47D5RMhw6Xc5izljslgOvxjFBNylhlW28fUqdXQrW4oyiWl/eOyzrn3waRm3sK
FWjkEshp4LRASvFQAljsc7I8uUSh4P6xqEsf8+/kqbqWrhrgOPh2QTpFdogdGqKaq2cmkoeuJK4M
AEPEAVooTMEp12afE5Ron3fIUjVWwmo9p3RC8P+XxtfdU05nCtpaTg5ga+phdUJOeiZxubjYipav
/k3qVnF3upT7qh1DephqoM2/sMLoa3moxAcPiQ3yxm5F4xaOlUKeWSLPV8UdtdYw/K1OR586iLAu
KBfuuXj2PuULPAM4Ygm18/yOHgQh1S1Wr82wwcWh46fV7oD+eRsE58kAX+pxtcmA4fp/qU9IEySp
em54QZi2xY2o0aprGGkWwzN4sybvNoFYIiUBNj2kdGLLYIELO/jT7aH3USCXZgu7cKAEHt3xQD/F
Y8s6hLPXmEvXR9oILGox4iB1oXnpNRtAFRDdR8PDdLKK8OCU+IbXc5dhRWxQF4xCosEcI45UGa68
TJZhZIYywW9aPrF4+iGcOXFbAD8orSvnkW/x7tuhhe28d4so0nZULnWlkZF/A4gXIHyy90nJXpHe
FdLRRRDpLKuc0mJYhUp0+fkPWRXn4niMXYJCa6qB1LskFeRWc+CeBL3xOjkuW7TDW94UcwBcGbZr
qHonVVHL6yCnQOAWwVrMLPymGfJ1SRCpjZMJ5pQZjW7vT5F+zCdb26gJp63Rrv/+1iq3ypHNp4Rg
ICyqf1/+tJoFoq9eQ9H2AhydfOPggsUkO8nNOScjRnnIaRuSxXeW2lNQsEDfnT2rfnrcbUmIB4s0
l8cLPDwCU9+FWx8U/LTv80I6Mih+wAr7lkMd210S90lvJ0el5MnSolBjenxZ7Y9k/SI7391ccZbR
MRma7a44MJpQ1yNInRiNUarPIpNnUU0YhL3wzUEeOPjfu+FiR9eYoMa2+0DVnoComqaY6p05j8yt
ief6SQBQPBKposUp4RW0eu30VwPThD4yidOOEr7iW7Ecd1USAoNMM7zd55b2X9yFRJUCNvhztLxP
Pi2Zrfd65q8PQeqSitUAjtjixa173Jhnd4S8oKlHaodtO0ydkJ4TsuT+WJxbtlatr/37wt6tKtWP
Ouet1OMb5mqSQhkPMq1IvKnVsAI4NUvLhAJ5KuU1n4a630h6X1iyWNUZJdz5tvZcKn2P3OwEkUgB
BVDbkFQuwo+rVvWXJX5GY4XF9lIQhp7vdXfUYTCEdIyNTvQErGA6veTEEfsS3CCh6ZtF6aCgoX/+
AiU9TUuLpFLLCZD6SY0Szkj6lmmNdlPSn16BA2w75E63VFh20ccoXI6LAGmJ91TBdYIjzjwjSqc0
2KKf4BgcewrL/F1nqOoyV5D5H8QWdWEUNIgWuMcBrDNyONR6qKGbJ/9cWXlDckEl6O/gX6TN7gpS
LjexB/Tkc/TCer4wDUxm9YWpaVl8AIyuKnsHed2W5A8T7mw0j30rAwshOWNwZy3OJ/IjizbTLvVZ
pO2RJDhEaVCxsMP08HzXEO3pM2N+xf3HOa2/VgP/SKHXRIvZ0U5j05D8Jm5lu8Ew7JKh4Xq/5pCk
HAqUsB3aQubwPFnqhcdYIl9lFSWC820vGzrBEgFyeH7OoO0xlmcC4cFPWdqv4t7P9nV4CwV7CA+w
a4dAcXoUwheUbc21LS30d+VoBEs5FhrJO8AC8TWwNLNAK1q9PTHQxwvkq8pl56sfx3U+zdx2gEvi
Op1yJHcLbuzH5gSC4oPbGwcAmoAaLSmuttyL40ZCOAYzegEkdwlOawDIGyWRJ43p/VsxLNFai1vj
12QSrw3pJD5dpE3TtV4KRXdJuoSuOLYhCztDbQuhFOEquzuMSNmZWMOiAp/vEqoxr2+W67CSBf2k
V53SIDMDhBTyjONAKLedfmSvo0l5b8rzEAYV2+iL+wGTH5n/LeU+8egEIaFO8weTzKwgwOK/6XOW
meIx1fGRBwzmzIV3u01Np26Xb5JsXMXEOjlFOatDrcCjtBx8hl+Z3bwzu8cuzrVQrdUqBnz2Ufmu
Mx4D7ZNwJqx34gk/uzV6MuQvlkZX1Np86AJZx5/HcXBCoCII81NNy7rsIZQ0eJcZC42QHH8jPaFx
k5d7pO+u5TeYGU7SnWEWUHraA5N3FOf/g+XJtyf58HfE66jMEzWuAgglqjgLq/sSCECBBTTYXAVu
Le7iNfQhgD78UVWrTSG7IhzAzMwWry9MKWJxnXjFd/rxOrLNqQBZ+4ls3VLcoM1JEeVGhM2wFIDa
MJq9knTekKeFUk5qwJn16Wq4QN6XWmm1STqvrBtVbHOQXp9/tBtQyP60LkGcnLusVBMfNtMdUsD4
AN1cVjNpGImR7yeGQHLZ0D+x2LSkblfiFt6QC0T6EV7fTGFQqBcTzs4xJDjKFp3ZsbvM3UFjH40b
S1gXRv++URV5FepWensmkg7OmP3pXBeTcNfLcPrTG7FBBVoGeGre+3QhUF/ds8Jme1J0PFgupKbo
TtrKs5Za77/9ITQc4s3e4BvoaCh1r3GNj+HL/ZebVBA/huSULWl+mOc3hrvQ0PjpWqs5KiEOKMKf
YpeoltGyc7gJ3D4S3Ec75IH1N7WckHyf50ri6Z9x9X/+GuzJsNgXmjjPVA0WKg9YMw7CbWEiiAj0
MbIaa2q2IXOmakfhztlddNUrhJ9KvaUJVmnhKpKjBVTDjKs8Dh4J/ple44skymdjLIIN7/0Lek/x
jW7P0MfeIfDlTzjyI8YulBgMZAlYe3YFKoo3yO0bDh9AeqQ53fh4JAWYc9CEKlHZnu7Yc9Xe3bq8
dF2aQHH7JihJC5iSE4jc9Ue8eVLbWhn4Ege5lgbE9kZmEoD2CdASKxv0LIfeevXICtTHa24fWqAl
FkMp+x0B7C1OtD3BQin+0ukSo1Qt9JQwGcJE5CfFO7Ptk38jDF02wqAjgv/Ghm9uMyUDPXLAuTCM
V0orXlsSGYpiyPwIa+mfg/5cWFfqBHuLZnv0AHvueHr//IhUpK+liNJ8r6GQdmPOYVUwK+3xCGhb
KDMGgi9T2hqb5jM3eCWkcF2Nw9kgRy+62PGitrJxQAsRWzRwy4oqsDUit3NRdWHPa4dSfo8Xy1m0
Gdw/G1tKPZvqdxWgraTXw1rf7m/TGSC9b4yvYainedbfVv9v9ljFJIlhmwZSqf2qKxEleDguuJQ2
u9wGsGtFahRWOyoxMgZWxi9LC7TyyufP3wytJK2/lWUnU+dhZE74YaL0nO+AfutjlA7Ih5x2UtTE
usg+XKA7qNYLeE3QG/C44hpO0XRCWTmQaLT5VVmSXQcAlMIu99l4KwkvGJ6qWidLi7WGXG8We7zP
Uk3ofERlfkY6Yaz/II+R9zmZarGswRcCYTiMRqeK+33+IcQDZ7mMGIqiToYSW5zHnvwz61alfqKv
GWt00PzXY9d7sMuIJG/kdQqG+iqzxmilbEbLHCmP19fxfJyKtfLtfge8a/J1mO2G87Sd1YLCkxjq
/3spMOwWRa6ZXJnApt6sg0EIK5tbzcO3tFSU3EQ/cEwSSjPDkFG5C1keBJpBtSCIKdn8bnhC3c/R
sPByodXhbwDhtl26midwjtkT9zknDD8WVxeZ6b74/GgzHNY09X4qT7jUe7hEfrHPigA2RhIJjXu/
YjxkwRSUt+OCGzBD9GF5JQthBbAAjqcUG9eAing0AzLs1/82pPPjgL8RqbEWOxC/xWTz22O12D05
G2Yk2WETvW0qea0glyQch57QAx4Zb3iUdIWNsxxmwbTGyXlvheXez6mBXn8gcuhuQ/CDEDj4i7qo
Ojg4jfKAll8XBUXSo4QWKMB3jjrrAf+tzwjVOyT4oI06l4rP0hn8AU9KI/taczqXJJHJt0qCqiQY
OythA4RQXLGylVPFpmQzTfNd5Pmyu647k90aMMLztpJVK7MTq/sohHwV/Kcic2IdfQg14/cvSuck
GoN5w1RH04WbGgHM2Gk4whlM5sAD1frj60eLNWhAowiC0cA72/rf4nCsmxhnAj/KPji2mRVrxY8h
eCt6sqS94/jBSXDpKZrG7SlCN3snpwILOHuQiYoEXiBuIvEZBHQHfZcHHK59Yb8Eaw6P/JB6t3xI
HKO+CTWDyLdES+0B45f08HrwyUqRqDJ4ilM4qqO2gEKG5wXVkaQPmTLNp/0SsLxLd5Z2mJOlhLNq
8QcDtvbhAXGyXJX3nvYyPflUnd5pWMo+k96nultLINU3Asac4PFb9Lkb0hgvjsZzo2Z1DysiH5Gw
toD/B6awTo5d0A/iIk8VXgDAUEcUIHXkyYVes7FLxDTlGgC/l+wZa/94bYW+Uusmz2EMbiYrNUsy
086eJzrfihoFEhxhGxloNUHjnoiM6gQldiMAta099Wvt78LD/I23Opr+eJpPDANW6j8IppnAHuhT
0yfPCOYKapUU83cDg4Mhc8n8fFrVVsoE/0PWvM310Nt5UytgEQIgOTPeMjovaPGdZvV3MkPhAnq+
MJcR9BssNzlBbBBMvwFIe6ugZFYBj10mHd8bow0KCAELD1eolDUg6/9PWYmTURbJmgR2I6X+upAo
rKNqt9ICeEbpR6v1FfNdt0VkTP8Jrn2+dHB1SbaKMIxgadjzvFn7UI3tisZQ1vEg/YFTyFBqJJnX
2xlL+3UOgKlD+/xoXCLgJPc/X9x54KoxPpSDR2dW7sFPGEfwoe7iAx7YcopqqWQIDWoDoYTt3aT4
4JP89b/zK9zyzp23m7T9ADXeQva+2dB8kRDBy2DNY7pOuzVmu9/tCw5XfSpTLxG5LMYx3eKESkfU
aZnFnYg1O2UF6CV4cCvhRnIaSuGo912bO2pxxUtuOoZnW8VxadVpie7V8jLkpf4Jw7dU7GTf6+zY
NfvqGjIBvFxj9AWzRlvcVW0QjtYI4OMheRZa3Zfuoai/FwogHHbwAqPpz/ttRhov0gDA7nyaiQEZ
X6h2nWA1b5s8k+XUnIoA3WMectqryr9YwUb386oqjq9lEJNRBEjOYim/hHy26IopWXD/GgeuC2xt
h5Csj85QEQSH+jxwboidWuoxvcKQZfvNHxg0vR8YwC6xbnkk7DE/x4DBcPVc4teu0O63TIyKm47o
xItHF5iSjWBhDHeGkAlWHR1AJUc1PXeSCYbWWUWx8TJw9FAw/M95GcNbcpiLu7DHe9zSjwH+GHpB
x6gGQAgdw8dVvVHilwoHPBbSf1NO0SnLh48+Ct5oUhtVDRXYSnDqkALA+IS4SO+hsSFrTZhAq/P5
kxmNkMMFbu/qhToKvMh6+BwaNy3vsHYE0O0ztrGaQh4VI9p+hJp4oC5VfBRxA9g6eFgtUMtaEtRy
rr1fLkAowQxOgP+SVppBp2CerSSzvq9OgBuRMdOcYVlQBlsERXTGf6j+ifwIjqqeSX5TdGBkx/3B
8g/jAnltuOH7EXmmVbz9SF1GgC+jWzZQsWDtfYYqxUdLEVmbzyJLNThRYnXE5u3olWbBe6VV7Hc1
CShCXQ5xfiqjQWWLSBpEXeTKasIYXutZhwKyImK40sOWw07ZBacxkozR1N/P9fAIg/3vMhBssCOJ
e5tiL6KND1KzKb0/8VY/6rIXDcOsYyfwc2suDf9oSsjlnXeb/8TPzwhqJeZdOztrOrnoles1O4iF
FDCOrEXKcVY4BsDo+gjEwI+BQXhNIheC6DdOVb5ojnkjgH2eVJL4Ftd9OAnfSvZW/CGCGT9YVMye
a+fEuvuRdaOPeDBDozgAuJcOekUBDm+G3q9QA6XkpoD5j4aIo122KVqGhDjs6gnme9XothZva1pV
lysQZuABma1XPzvK8l73GjqWK/wKsm8bhlSeUJkppxamnQS6n5YOkPfFnI6TdQk09eLb9kGnRn9E
9W/bvAMhiXqJffqAd6KtCPbO7TJHdpZyTIKqnagrEP4+LMaXRZkUyE1oDE6Gxw7g/+9x1Q2P/5SR
cknsi8VxtT76ITA1dXkmtfNp+/X25y80lm3pTGDh3mv9/S9RVNN7mnv9vBwfchztr3+jyCZc24kx
lBHA0kkLcmoLRpaIfshxWCPjXCtGvkvQMmF1tVXP/K8g0LKPtBAgV4kcLEc42KEUvmrVIw2DHTJl
RHGMgofQJUsQ2Nd1XlSWSpO/va4LgHKKK4Uhtfh5vDqlXKmoLK6QPkTaH2zmB2Jdig9S5dr9yuWA
iQGWYzD7TlgQIv+path6YsZoDcgR5mFlMWHL6eZA3R0mu00BftfaAd4VOE7rl4dhwm4XD8c64tL8
1QSNAD7U2PzF5Ra4XdBYp5hf3deDeQOZaw3Gebwlm8vSCKVGFgxbdY0roPCwkdpHxI/RWquAGEmP
QKTqU8OiczBpwATOzYtQfuqDd1+4mrxLcx5hLaWhDcWr4kzvqmNdMl4v6td0lJI2nMZF/MfqGlaJ
kJdi3ORyK31vVxKN3jSWd93gFufPFYI+cNRnyj+hPgW0NaTnwwEGNAwmDT5NGGO5LeqH68v0qZJk
5UU1cxdxEBbMNoP1iaf8Cs0LFDGNiLLUnmaeFrb47ujFzDehDTJeRcZCH9RDO22YxgPPxSawP8SX
FL5SVpJmd6IpvNaNhSYlH4lyeQVusDIs6ABHBLSony2NBOVw+ibshPFFD9mbUd04J35AbwVzsCmZ
v75FNVzIfyD3bDf2t9X3+Pqp14nj0YHQM2TWOZHQ2ehOzzeGyZea7aC37e4OpPcHkZhU/DpM9koF
39u1om/pER6vx8ME8RVt2P/6ecis2axfvqzsC3mLbPifFfC4Z14kow98QlnlwZoGeSKLeKP0jETa
dYme9sOqHrvPpRtj+nnMf4IToeCjRo8m2ub3A2f6yNX7YDmM2Bms+3JCfXto36QJ8nU3RQIZgtQm
QCEuX7jAmmdOusyDBYPOwLwE0HZup+gPF+KIiZ0QzzIdd9wjAu8w3RdLgw5ZYy/AgTynK5tSgbJ2
+Gp5T/cBm3v00sh83cyVnda/Lq8EHOcHEVQvoVMZHDsvOXcVGdOWsXTQ8ZvCl2NBj7hHoc+KqIec
ucmAS0VSBKr/ipAd+HajMYTEqufsc/CSHQDxg+HrVxZedntMy99FHHan/4GakW//d9JdyVypjH3e
rRExGo2wnT4x6bBmGA8Bi1mMQZXKJSeHT6B1/FkJR9Nu2P81U7+IDChLp/0d9jdIe9LiTEDnrSOz
2IbQMhGXmOsege5N4qILjXEEhdG07hTFe6E3MN9x+iMXUnCY/igWh9TxfMz3VxbfoLxIcZhq+uV+
xp8x/QrLi/9DC8fhDevOgPIZVSCAuyCB0+8tidPMdFB6W/KzLYAe5eO9hR723b6pQES/Id2ROAg1
7oONSJHYWt4Gv5BwOd0WrADbVfUVDE9sklRYIWhCqrHVPGs6pXv88fZQ11I2wYzrjXl7bsTtt6/3
H5GoA/i0orHRvjkdjvsJrvorjIt/ICxrPM99pZVmPgUAJok3gHGMaJniYoitqx1wBNUgdGqD8DJ1
fAvAyMgAzQovFYwPxuXMJRZ9UKAAe9IJw5If6MaehuNJGGLREUUM0Xp0lrvhpn93YkIaIJ6AfJYK
Gf91ip+syHcFY3j0Ouw7vnA8ErhHesMsHUrrO3pQCY9iJYtM40nOpH8RryKyrex7xsfS95wo08U1
6uTlZ5i6S1lAko65Jfb7hhktbht/aJ2Yw4iOJQotc8M9K7mFJY+KiFnllQf/HQO3MbE0qpMqfz4s
4A06CUhktSPa0Msf+iw2IFwI7qgk963R2EEeaU+GQzD/5WVqB2bVNykNt8EaN9aFG3tEBRjQijG+
WEetkbpnr7bTIa0jw7FnKi4qGMGlKusetm72mHoKR15m1LwzhoMtuGy3JtKzF00yMBYdnI39V0eg
xSNebHgD0KUXZKY6+ToVynBPS2tiHeN6xvxCHCNbPkZ+n4cxMHM2jUppQoqLT59YWKZuedYAA0mT
Eb6qFVcFJ66pLpkrflDxsst+vpSYOk/qKL6shCTLQ6PFs9q5o4HHhZ2Eb54CXiUyvC2o4xzald1Z
a259SkajrG+UeU2CLJuzFi8o7ZMIZJ3yXmm95KpUchEPGbQW6A7zy8ztI/gi+sCIbI0fsUvqekbT
lAFH9say765rM74IHtbypVhv8WY6lcI7ZqTbL3n+GBd5rAIdq17bAJ4c0elqJACrOfCoCMu49s3F
AqKkA5CAsqskCKWAYaB3kA+SVTfc+8XdQ1tOmFd97itIej0N/SE4r9WQDrNsyWZsrpVg8X6MU7OX
KKM4IlOE7Wr1XCs9bSLqJpI1NSGXIqyZ+t45HJAoRxzA9DTDdU1zsIgTAaz37OdB7BN9Yq3ONotS
rPotXgU1g2bsgrLFtAsXancbtCJQOPh0OfdKqO5Gd9T5UWFvHSH0vqbH1eIt4jsMLowOYFaEXhOB
qnhMbU5FneGNBbrnjY2Ft50J07rGzR/bgwkQKgwYz1XvSEYyQOrbh+tu6iMEds1Mvxy8EmPOA9t3
VedUCN2SPRXj56rPPtSAVTCsANYtft3tzSD3obwJiNs9/rLUOZiu3sZDnd2+cc9jVZqh5CDZus3p
srNEiW1sY3GFK72x0S/Pxgk02safoVJCCX/Nv/eeUQHf+e0kc+gpVHZ5GWcnukV89bRPPX3xZPqc
OkvmmMp+OJ8cbrGEZ4fz4LRWYmC88SwsBP/O3qMpuVJoo9fMuYTYOdBQb8LyLTY/tbhqxzeTOeUV
cwRiJayQN5Vb3CniOW65PBdO9z1y8Pfb/fMXvHMylpgnDCN4s56qUWiDNdMh+qty2cHs7r1xSsMg
SRzWdCjDlsfKo6tGxce7WDgP6EX1wlz7yXmqTq3MpVX540jR7eV0q8RGb3MUdHdFilKI4lbxAHj+
OfJiFGN8do/SdTeG6dieCAsDjps7L9s9/A7/yT6JGUizFK72/B1fInmXjrwLC/AGikFA7wR8c9OS
0astzqXeEOJqC2er/BHyPXpQnnGuo8AZA1QR4PqaQ5HK/EwoOb2VBED8hMah6XMXOLW2fY01CW1I
6lbTK1qe5B6mHztSQKmYUhPNQoVc3Pg14heVRHKLephQkIRYikNABoVcjXSxob0bKuRixaW/thVC
fyckRYygEN8MG0S2t+aq8rDAEIh5703R4Zj9JVcrXufPZ/1iNt0LQsPcOP98gxcSvPf2lsqfRyCG
NuGPXNblKA5Kc0d0G5srneQcO/z7g+BaTgmMp+PvWO6YVIHRDM6YGS9l7PjOuhDNtkMwDkE+xWf6
trKg3qqeA6MXvLI8jWaePbUUcAuMsvTMspNhHxev2YEpATi4AieHco8Tt+sRPM9y+c94Pnom+Fyp
huhw4aBactHt9q76yPQxtq7W5VklS3wHeVdyQIkkjdLuno1o+9rkwCDMMCE0DOwJ1mo++Kzx+Kjh
8HmTf5UEXP3p17bZ4RP9QNgViC2SxdSyLC5HEjqOcTW5WGaNrBR/tBtZOsPHYKVTh/tCvh7dnacL
YVtGbLJauFbuRlGNM0nBNtTTahf7L9e9hgDw4SPJtAJ0f2V9bu+u3SscVq2paoCwmllb+9cVh9A0
OzcuyalRFTZZiw2g/dfrGojm3y96GAWEGdq/cchpaLMqbPgLNeRO83W8SwkS9Owj8YEL38B9Bq8k
GFIHO7rrQtPelXQE227a3EviINrlNeN234qgL9cGXzVU/wUc4ecGv0pluZRRkhQKESfQBpyYf41x
vIxAfbaPH1NYGVTP3EK18mJhFnsv0e/yNddGTiXE0tQirBmqIB+vWHewPFzzkpFGDn2rMIL2dY7n
iZOBKd6dXdfzXjtxpgGwmgHkCwrXrSPn8Jb9v19p4isFii0tixlzvkS9UJpC0iDmsgtftnRUSN9Q
M7xPrTesMsj7JP2IW24orLZM9pEySxLBMjowNjUfmeiE+jvw02QjiA+Qi2P4sbyjZg3eXt41NF5m
KJVUWFFINaIWL3ZxST9YWWLCpJPaBcvsCIFJqQGvYxHSjYg4lrOhEWKDH5pX30x6EYXvR9YNk2fV
3nplqOh/mnpUD+63oEDj9hoAcnsncseqxCdGpf7eEJ1XoRpQVa4RGD9shFr8x+Jqv0x64E/1fXV1
hOEmxSqjnjCKT3y/cDDsoIIgdZtMK4mLBpZGgcbM3QnkM5Pq3BUuhGb0bkvaODHwbvBXGtPE9PjY
8Qmynpinh9cotV9B7QaefFOXxN2csobnqpD/odeEgsys1kxwaXi3QmDU7bzHO4tdD9sYWeGEve6/
VQJ8B1MPLbTzirq5utIgvL/iaJj1IYldoU2+q1mxwHPnGLk/dWO3Rp1bYNNsMtUQkD2LWMfiOHX9
ojllgj1awE6PprMw9msTRcb1SX5wo2vATJxMipGsMdx2QDlWkB61oRYpzH3oRVS1V5AFrj1EPg06
lLFNBm7m1RUbp7ZV58SUSwL1tRZgtv2o9Q82+hVLDHZGJufhmYAtyIFzhqBqrrPp/zZtn/AGLbKL
fRjtRWeEgZco3hFWP/IcJCss8rJOmGfVUeVmwN/RlQetiOADescuF8572Zj1jKzxCgrS/E1MzL49
XmrxbzRyAZu80HZPBDOE3JgmaxaQTjLZTEXLn7X7ytD/K74EcuRkNPpqeiZBk4LV59e541R5piX1
fxVr9206Tf3byX6AhEhXv0L5wgD2Obv7ViShQrOmRIL+4G1GAmNqExqNeTGR7ykmMnanJzQYH3/I
u0No801YmYYsGJXYxQa673TC78CKtBOwH4nXYyfckAeXToJvLGalJVc3At9KQdS/YChR9pHc8BkT
GwmHOCjEbiAh9kdKwwfjwimc/5I2bxuBBpv08smgXf6SkAM3A9jPhSXFCPQhiaIHClkXJGNtQpsr
OhJiF3m+fOJbZe6ly8xdLs4x4XGAlMquslBAgW+MXA6you3n3ludtGsqW05vGPZcqee6Jt4QYRbO
FVVtGQAFXte1hUGfxdRsb97fS0oaV+EAHpY3PRBgEgRQWxechYXycGydjRQX2D4TqNiy6kboPOn+
vQxxnGofccLyOm34p6culuqlDR7UGxaqVW44+dkGfbeeAarGwPBMAQfrjl/yHrgJfUINDUP95SMZ
llDYG8+DTWbOgKR/zAAbnOl/JnKH4lfoHXa0iskfwuLwXFVR+m4mLyG+oYRcL9N4345pnHwuBbZ5
fjr7pMD5Vu5Ahxa25WIg+0b6uAVWeqrTSnIx8jzjN4W3MJhgigkYn58BjnZnTFvqo/KqNntOSCuY
B6cI0wwEqj+sk4ldnphYEVXML6wWWxkM4Ce45KJRN/Tz3J7pmPuSMELTqgHip93Hfy4zUEHnCcpO
k9FCzmgo15bMeHZPERntvqshR0Y2FeWBV5Hs2gJDRDHcg1uaSSSFHN9ARkPn+seGY7490fwNQfDQ
2DSMR1LM3N2V8lkXCT6f6KwIgcUj18YTWY0ZSSrbMLT2A5PG1HwNn6v1VfaazXlaiGWorjB+hgVg
5PxWSG1lEx1dcm9QzNoL38XrL/es0WUZEabp8BSEROTLwQ8A56dRWD8AEEanyhqFVytTf21kFxUM
Ee8WuzjvzdgCAqn3a+VjrgDd6XZG/OEZIA02bnsiXFoDyj+YYNVcK6Pn4tkrMVCP0PUnGIA0xOUS
k+PyHBSGF+BdfT8rhR9HZITDjrj9bwGGEr+S//r5EyjCMCUsrZwvAsjeue2/Mwz5ou/75YyHkytk
oJ5RKTR7sup4RP40AIKt4oHmi6gs7bUtcvR8SAzxhTKg5Kd9iNR8G97Nm4aK59YjZ+1z/BN8gNly
JQP3wl+vZpMtEF70JeOIs4BqVsgAAA/kzvrvf3k66JPMHJXxz0E98Id8sCRMcf985KQzdg1Oy/FJ
YwYCH49Fr9p8R5TvGD8DzLuK/i2plGwSiq7MY70uIk68faL652WWGLz11gr8D+U8e8VXtNcVwwmF
8F7RUdD/YyCqERMLQW+m4jNu3JOZKjcxFngq2CaZwHW3HIEW8T9BBv96Ved2/FxSIjaUVCdBD5G6
p6eO+SOXN19TsLadvKZRz3TPU8c22BQQ49mWkjyAc0DVutVZ1k17LG0saUfMON/4HcywuBjAViVi
LVCjDu1LOCjkvONkSc5u9o+Wq61yosRNI9jtWc/7RNy2MyvcV6gpeWnPG/1f22xv1QdoVP7y46AV
mKaRRxvZuCY9IhwpXLB/Uz6eOTBfky7UKgYv0sopsu3an7+411zznPdt7WYq1Ugt4++jFpGVF/n7
/D+iTyasMRKtqosJbIyXaZdf38xrBBA+yk19q8BCJEm1JAfTX4yh2+71NV8dAPG1Hr3y9wCrvDrz
NBX62OQYJ8rKDqEkz/Q2OxYYPSDKdRqpxax7RfQTH8CzhYjsHKaWQmmqw5cZendDf2esxCcA6Zug
pv9n8SpwY2hYuisfrxOr1t2+k7y3UJiKBBVD5adK41zlyByyV9WkvJ3LqS8g6+krVpZ8olx1x6A7
yl1bacmoj3uqJ/IBjnnfmIGErkLtXmTNVtCFSwasuFBHhsWEXm+IU9FhnjCkU/wqwjTf2LyJJxzX
kD3FO5SEGRFLeqG5XRjETzq0J6AIGgGjAYOHlPfym3SmMKiFHEIYEDnozzSh7oTSzRFjrEGi4Ngm
tw8TPTrzLcQg2dm+uAZbAyI4koiKzeF3BCs7RLBMwAHP+XGB5Yu6atTYP8S7RWBkHCIhIF35gmQt
1vbS1Z7CUwUtxEJCiJWKbZQU9RSfi3IWgzOgLxQ30NHzbmo5kIMj/ve9gyKYz/AJpLW6mRc+5BI5
eIFtxczvHsMbJZz8+8F+xhgKG8X0G6Mu59vG2wnCR0khvdpmdrve7WG6L1PQCAI4EKNI5pBMUTna
Gtfj4X1nDgNA/ruk7SlzcCHl9Xdq8wl/MjJILHaRQm38PdyfLDL2PNZD5mpYLrLTgd231cV7dtcW
UB9xd8cx7aZeHaUfzl9ZGT5kPBNgUCnbLhR8jlkGlSfkU+Q3hkyNXdy7aaIIxxQgtTLMwsjGn3dI
+7oIOO9jVT/QyPiNo/9u6bIrn4I0h2sZR7UIyeveCN/9rmhzi610Bh1qupSnD/rmZNBFVz841Cac
LK1JpN49IgaYh5JoetqxqUkWtMsyshCV9n7lNQTwsX9kNiwlsf8Eb+of70qJrsuez0lYNlTvSgAg
rBqshNC5t5bm9fDLIkwnFtCGtBEQDLaPP2kUUsZgpwaiG8yPZOok1nkkW45hPKko605RNzHVwRNG
/Kgj91NafY410sCHOh/q76muhAhFc2KnaWkIiXUPxbLxbp7B3vXfWqAOgCTYR0+rJxKG41Tu8UtG
mPzPNpOo0fXy/jJ3YhS83KrV9/ANxnSUrpQjT+1Jz7R/zKPFod2x4o0xXlho9DV0nqU8O1bdKoRT
L4jj0Plpoq2BdzfPveQGzqNRfFHjuc9svmpHXRrTJXhbf7Y4DgBpnSc2yBh0+GO3El4IAaqdJ5dB
o45hNPZumWJwhsLwdsr48sQ8Af2AeuHtqRWLNUhjMXj9Sob6P0/g0ZfmvuBfOhvrtpESWValsQ1k
xp4UaZ9XIeYqPXcXkzkP8jGI+1LSQUW/wrhHWqmGc4JDyyXgf5zZxf+DcqQ0wz08acpkKEh8ZBkj
UaYCV7g8lkOi8B6MEg27giFpBKMxkKEkNCgcSNV6aidyGHFeRF5+omREz1OmslpuvYyFIzigesS5
XKTUWFOFmY+QLSQhowJVS+pJQ2WWb3uSikWn9GsJ6z32jq+2DPUJVUD+JjVaOaJsqYHyPp1Qi40H
/V22CxmOOP+KNOHpqIRSDeQj5+PCSYDnIApfmggGVxfB1+n13pPgY4XziyAV4uo3jW98IfAmSHnF
68zyx67WASAMGlhzUV+IoFHfftoEy50899/cvxZ07VbGHiJpWijUNgetaMGzC+ZtY/WJYzk1klON
/lvMVS6aMS+kREU6CmDNC9N6VyWK6rZRtzv6Ot4gjmlQvV63foRsPMu2vhfe3aPB1pcMOLBdjxx1
+Pz4coXY7frbEzmOGfRQmna/E3ipst9a7omOFLf1L4e2rUKKwJn1yZQymDYps4Ihhhlh6aMT/+ff
7CrOaYwERElpQmPqGyRSTZQs/0tUDkuXdA0JyKxOgF3i8kkSUuPG+YYBDZnE//EszC/XJQXx20tw
ChO+/NyopwlAV4SvshaMs/Pam7qbnWsZYZ0OH8taReMh6jKveHZgmzv/c9NHGXiqxkj5ThgkYJ90
l+eB+xjgyLnBqoyxED1LW2OUpL691ZQwQ34xPyXr+tmyQk2sU3v4fIKaKzvErPppTGkyeCM1txmk
TFbogU3CzLfyzhhgDjrrImTuQm4dfsuan3fjFdMLbJ1ifDGDQ8wXmBuxp48ZOQdczeeZjnEWP575
/7Al2/bwzehIdIbmyvCloKDkHoXjNunQjwj5Np0svuwP1t052KbwgDihi3sHY7ZOZ6KWf4fMscLr
I5LdKM/Gj8DTqM/omrzMTK08k04ZMhQANDSN/daXsMSV3f9jpgttMYUw7DmpSC1W/IPXHhaQzxwV
J4zxrw4YVQPfixsoT2iu8y/IJ4hq/loMcrvholEGihFGEOEbCbBE2mPzpZQGMS2nFD6Y0+eb6H1T
ActpVJ50A2+F7IgnXedbDVudCECbB56KtXmhSL4q/R09NC2xM9+/yyNm2BATYGscQwOosBdApR2u
qQGUhV14xwBSUI7WoBvBh1hCozCYfBDnc09FSIJWNmPXGq6cD42NZx3RA1KmKsg0nSkAehP9Id4g
5dB4DwfMBGxUJI6YeAfylFUu/iuCQwghyFnv85AZBAx6pd5jckIjh92eB1Ng2i0Ewg1X8/64UpeD
rVW7sCgz9vGJPm3Aq688xqYdBx27Ykb/e8Gr6RpWm+mNMwuxkj5IRaEkUV1RTuhB8Iya4bvpcjES
3JLIUvu+9vFQYsnPsKpuWHYSDqfJX95280xytIzwdLNY+NQSaRScOYGeXtmAB17t0PwENwt4yf2q
ccnwtYcQUbA8k1MZL+qnspwv44+uIrcxCm4Y13LMo06T0A4beVBsN+/MN7focN00KQf+pAngVBQE
teUUpZaxGBc/7LMhkDmCWE5joaFJJ6jKXhsUsFlBYd7lLLZlFsXy6fpKyzo1L5VnqaBVyy7IBvuY
rhTuIPpvEoYw1hge9OT5/xVRxptvTqp3kymAQ6d6kkKUMZNeIEmB9BxRnklHn0v32twnntG/hzvC
DFaw7UXrvGljthNmK0hckw9QgrQIjPWhzG/QItJejtRADrEzsLQiYibaDOw7dO8HRk2CjeLdlTQn
2q235F3wrRsaJ7vCFsUaaAxZQij/CiFoKxdD94/5OucEPhd4OP2tAigWVAFn4Zwr9e30C6+LUyUv
u9gvtz8cLfg5YAylTwfUMAnR3+IxlI2guTqLz7UiT96JqmdKifiBL9IJyLq7j+egBASTTn4yXKkB
e6/S8m4+bGGAcr4VOdaYpjv30SVEe4MoUljDXFZfsWFBw0u2F+zPaUguzE++M6bfmaZpAuOH+SSY
anVGurQdRjbIDLvzuPPZUqhuU7X2MB3EYfsiRYCCidPvF923ZR9eeJK+ivDpHy+Z9D5B94fxjBdq
X7AFg5sX2ayJhvzlp4RPW/7ZqVsX4vEyDrgNXTXVSIazn4Z3bD9EWJexNfjQq+JYeQW071r+yYh2
SqHAm3z1rBbdyW1E4zaXlDwTvYMXVGUiH8nki8kZ091tqZyrKAMpxRex79lQqWwYZsNdbbu8XgZY
DkAxFUzT+/DYBwtuDi8jJqORBUvGIDwXI9iX+y2DxXJMNC2btOoAn9s8q2hLhKRtrBfvxRiEoKje
Ju2+JyCgb+CTmY35xvdqzWYEpr9Arxprw7lJW38z0MrfzOOTm51UezmUHNx9hpf+t1ffpqQCMGoa
gsLjOgsgC/p0J8sGZw+M7sn2Ery3S/hpc5Y+Aa/39nuxxn5MLkJHb95kdxgMZ2eJYdDgaKu69QYU
RR/rR8m40lpefTPyibpvHodOWn59TQvSRsUS4jrBam5Z2dLVLF/cfcoVkNcJCkpBOWrbtqkqo0Id
/jl5k+pgi9Imeft6V3Zj2m1UDnOiE5dW3OWDJtXi0Nw7P4lMv+D3GMEyshkfIPFeQ2LeRXK9BdQ1
a5ZRKoMWd3ux2phbUKHkOBpLF3uplncLg8X5cObA/WvxBctlM0VS8LYN3vAxxOD76M5SEIV2Uj3Y
0ncGJXty9vsZ47pXwwvSVuDTMHEHO9LnIgr1T+Zs6o1mCoOqgSUsJrP42bgciLbTi/H36rs85AS4
q0YBcwFR+N5wgktg2IgIAQnSsYA4CS5Xwa6npLOI1w6jHJNg3pB9QOamAptBDpPlyLWKvIiAIVBI
HvWBerbqdUxgeUnGJanNDSeBITKK5pOFXvavKcJqJ5aKJkRBqQ0wxA4/3CKGGAZdcOhIV97CXQbr
6Kd1dVurYz2C2DSknpm+r8sBnNZr/U5h3FHJl27I2YIj9FFlf5EHwK4ohCZx0tW53cctg+q8kEUD
2kkZFIUdRrgoIJ61rZn+7Mjbx53sLl+VihBUzy8kMcZZvA/yZvHWrf3DjIfZ/OK7omx76w+PAZ4D
930qcmcnOPWjUolZbFcXXGUSQ1vqyTYDfgTZMGDNKZ/7BRagi6GQ+uisNwtH+nyutI8zHdjKRV4N
g5oYuMH0rWjvoIPDwCOwyFrCW4wfe3QNjrTbX4EuX65g/Qp9zat+Xk/Gop51sqhWYbZYYTe06lw0
HjjnWu1OXZrTkSXdDamMLuwxqKc3EKJSZ/WOVdAADybHyKRDUtFWk/MyzZxmGw5/loEv2zcYpXKX
IL8MQytIc0LUDXUYTvlTh14Q9ICVWrgIBjWLjwOZybVs3YWVGvgm78IEi1Rjh30th5ojh3ZWSJ3f
wzt/YHDlBH71wGfi8KgQ5H2PPsyxujnHlzg1RiRuFhcmlzqknPFRCHjxc1aUQKGHkFxy+rJs8aHa
4UAhaFCnV4WxGqm2ZRzpRpG0fhm07wW0UmEnIOvvZ4cnrz6XpCpRgdeIq3/e5ybD/eLdy3qPDszj
5gJRcPHTyNAwisz2/p+7m8sepYfs3l/yEdJVqOAKcqd+fTQB9JR2RIAvDttkeuCDoz2qzp0l3pEB
oLmHdvou1aZcnb4oCLEaTDFMOTdqbFtQC0Hca5uHOvHw2xryb3PoMmNRy7cJL3sCSgLAINe0B/Xt
BAG5yKh1xCtAvO1D+wEzV+R03BGO//aXONy+OoMbOrFJFmAu5p2yhK0gev/9wdnf6rZxjQoo1ZF7
3DFY3aW1jE14mSfSH1tL/qGHLjBd3D1ktHaUR2AHJ/psVndfy7YcQhC98kweQBaMbXm86GMtwzgV
2K7cQFlj6Hj4ee3oXYosXe4uyb5cdjC2AHWMZHL1NiImTZxhV3ZH8JU7zcbKQmCGOd5uQBCoHlrX
tIJrCJyn/Y0VvpBqTfLkPHr7J0dwpp9rCbZvcStzzDtv2fldhCoKEKHnV3bgmM3ujn0kWcQKuphD
S3rwWHXGTRzSdMmGmVA5hLjoJf2Pu6RuS+egK1P3OLzBcMecEudhPfmVy+zmvSwoQTQBviGodCFq
MjZMBk6bnMvaPL5TB0qo11iLUnATkGMT2l7OQbRBhjxg38ijfHx0MQysMkq871hrMa1WPp0apsKB
UU7o/URF7J5iBS1vCkKk8ez91FoYxQfVVmK7niynsaVWMONv+1gGZtFa8ZEUjHDRAzDxa8tmj6sY
3qfVh1YZTBpEAfrYVIjdhDHe1fqg0dGmT+K+KWVHJBfIlaHEjjR0h6s3zy0acXUu+K1MIETdELYP
wTbmLy7Lfg2RL0B4wMlswJzpcfaUyyyXBwyfOgMrTJVj1f+wAYz682scbJ+H1W7sMmyufbQlgH6L
bjcj21C53Y/VhXNkwlz4gSzR5OcAVzgEYAcwhsLTtZt/wQO/8+88PLtVAAOvRZZEi/C0CN7YbrhH
4zzkAxsrDTd623I1sCEwtJgPqsdJMu0ZRULWuC4/Wf4WnlxpprGDMmDdUVzxsG8E58+ibmYG4Or8
hxzmU/b9pRdg9DB3mGgDzDOpKY/O3J02OJSVNpZxWBsdT6rEt4D5hHkPm+g1Et9x0a2HjjVLyBs5
cc0GZUwAuazmWgF8UBZpT6jFnwFHNgUHEa5dXg4v/No3Adk+US2ssFZ/Q1muL6NVsfFCDgMP1HYr
TD596yoCEvoerlx9gWore0yU2oxv8buzFcILfQRhFTquDoVDnHaMkPk8WK56N08zkFoF08ugCLxP
UToBmfAsGSIqYn198mUTTpKYe+L3g9/Epz85bv5MWbcbFuwARJMCfjxCobST6TB6JPFo2BVujIrS
KOzDdwIwFVgrVbfdhUKB+zM/E3x+SGHS+YmNYFl0UU9zcPx6qSwF7TDZBTgsqrumk7LpDm25/ai/
7q8BeALKDi4J2Vlh1PAJhI3RCNFcUC7vUJiuw8nwXL5bVlUuCk4ogKoKc1PQKjCshKmNrhFMJr9L
Y9AJ4dGelXRf1VLzYwj2FAz2C4zvufHKHGq0fb9mEsnunBhJgFBm64n0dEUpctC2s/zvFTYs6Fne
tVrLPM0OGI8PP3pkBiDjYT8hztQ4J4jk/GAldORivg3pEi52Ri+n4bGT4rpm0pSZ5t3Rms19cOJE
4ABwRr3tra08a06fr7ifcspPBLpONcipEpcZa9Hu20ws0MnAvYfAktMRZdxfO/+HgB6h3TFswwLi
X1tOHRrq+TAPNpoxByiDg3cvjQJVrfBeSlgCfEI1vUhbRpUhzh8whkTsOTWyVhLeWRu8XyobfINy
aLeYuRnFhwZwQH9m23GP7DLFj693VoRrqLcY3/l0Di1iJmACkfabFTFcJ1o+AlN2CS4sSQxsf7hw
oJFTkerfqVj+fYwOc6YfL49Gpa7Fq0POXkgxvJcczyBiywjkbhUEj5TVCNVawwcYGZmYgD5ZuiQb
5LyhxWDC8cJpsyq6wxUGUI+hN7kFgU+GL/84duyDsuGXZ8oficyDkD9OLUZv9ylu2+ChI1M1zO+J
QS4yzEPvOCx2TBjRgIRVCT2bNU69hPk0hmCNWAMeYLzEH1GmE8kmq/cR+pvXOIikFA+daQlAW8qN
2svlU/DYCIvDQ5gAMUx12jN0ds02C6fmRngLlQJLfrBfCJfwtFrYjLlTb+zYX4K5/gfWZOlePVq2
ewDlyJd9LLhsBqQuOXAQWkdi4X/r2j5YiX/qaHIWgKhkp6OGGnKvE8sMqCjmm9GHj5rdm4wk3NFi
NNclyvXiUPcqzM4ceN+jBQRQgd1r8PTt3CtZw/EHauPhf4SEEFv8ByFBfKQgkb4nVdT/YAKtzMHN
ZElqxw7nHiEdHPz3S28Dkbdy62QxwBzjPDdXSJ5/TYkS7Xy6fBp0OxYkeBBAHBg5C2G2K/aFMBBR
CQ8oIQCZSSBDScnq0qAjwjJX+DhCL9lJRwu6AbOqKWWhcyHBj6NfBj21afjz5knrRi9rL17ejuoT
izoO71J7yVii0FQ4mAAm3FPJXRXAbTRiKNGLCLRTyvFD/W0B1h111VX7qSiEPK1aV3QpjWCJgGFC
pHhn6CieX+y9JQF/vtBs9O/EY/BTLMtSXzBwsqOY3CQ49y04OQrfNHbiQMSUw+wXgs/W21FjMJB4
0NOTb6pEGowEzyBj13hlrqJLACCDq58TBMxR8zCtYCyRA3u2DzZeLLs1Xj/ciXtj2i3UboJfXwYg
k1zq2oPtPIl3OKinUQv2VtNtFCjBoyiWqKyLT3CT0UB6oibEw2Qui+c6eE5cR3ZJx+4lkIjV38f3
uJGZCJxq5eNYIjAZX06Hwmo8+5dtiwX9yx28gFtv0Lp1ABcBx50vAqbkZ8UMvttQHyUnm2uYacpF
KkTHs8ixkhGhj3Aa8EOPEz3y1hMdzSvIIe2+AGNks8tZk4fHjKlC3pZW41QFIzc6RoLJH45dgO8n
N1cY6YImJ7xbhXxWFjPGIxCueguz6M0JOS+6XABPnehW5b8V755w5kCHY/d5f29MPDOQSXl1jcrG
lQ1mdWs721IPzIMVDeuAwq++IdFYU4ttUdO0caGvcFPENjJfzmdcvQCUY0x/6WCyLp0NyOqbSjUU
kUWpX01XHrHK6Ehz8zp31W4LHNqAtNxkb3rZhrl1o+z/nBhC21bkIPX8+1cdfs9NU1E2dufuxr1K
y1cvJEc2s7urOg+Zs5YXj9Nl9MUM3UAjWuLpeRRxqyQP90btO77GSfjcA24M4saJNQnRij4Hp0pl
Gqy+DLn6Yyu0ygaKLv9uIT6N52eXzu+eHIEPKN1nWzhjLjwClXH2XifJRuYrhvoYl11+nMcigOdW
j9Alv+CavU1PZSrQPeS8PklTHID3m/1Kc1j5jfg+TIAvBhf7UfT9rW2GqUlmJ3LQK6qni+PfGqOX
j3JjrGmuD1GJaNVq8fivoELizixs72LIfzK+jHvTOwxQ+D5ARKYDSbso8Fdy6AEL2GYnlN7/bBUX
j0ULv2dXuAIqapv44gSUmZKjEcqnyw91dMnnj4TYml6E6A6YAU3O4hSSJze4R7To0g8EpPld1heE
f15AxCupPIbfT8+SvI0P8PrH5KOE6vvx1YexGRCTlsIGc5cZI3rK01mBlg2OvmLMFIJJLrZSnaJn
M/15SkoGjssmPC6PMTeP3xwuJMI5tfbA9LubAgA/2GQpdDTgGCq0zzpji7tvQY2skmAMlv/4Vduz
Qo52UoQ8kMN8Q+aOOzrwFlQrzMQszn7pYLjMLp5qaeCcCzqzf2VTGPKoXI3ltuIDjY7HfcBypcnu
Mly2MfAwTP5uKv26zlhmXchhbO2PoV2Aq1RMGqSnNdK2w9T4bQHOrT9UzTxu3j81xPwyezZ9vPXt
wrGVyDs0k7IFpgX+e9upHdRrpHXBDHffAQ1Us5LSU/C+6NS1P6DBF4rhvQ4MzcfRBkhavNtsdZxp
Pic5KJrz6NKpkMATRUfl5g3yCPDuk97n2iX7+Zxd89a6YBtUiILKgcGQRY+5X/GJMfUWk3HE5lvr
BwSld5R3ie7B7np1jv9gAN/ceFAI6PdW6WIJ9pC6lwbYWD3ZYAScLMPiawsq+QJIEcowm7HGK40I
25A9aKZtuBeZ5pMUl+QbhMQo8KA6FM0IgunNf+RWtMyIlGVqjb/ihtLxIyEDn0KSdTjtSIi58Tft
fAsJTNIyLbaP9VGmE7iPKDTN9ATLu4WjjFPFHgIOmVIN1o8mJjkP8Z2hH8Z49Kp5Dss1W6gYBF/p
y0JTB/6tViEtF3wXdo3J+lmekxceU2E2xlE4YPcf8VGyC+qyeX5HkGuh3L52Zx6rAwlhZTQoh/Uz
mOvWG6HjAHD51mdBEq01XjAEsjsL8Km/QsSjlLb1Pg7FDnGjMfwFQBPk+bDsX+LkNWihNMMO3ULC
Ht/gC4CuUo/mJCuVFki0tlm9HKNGwNUVB02mdNtzrrqp6E2XSfu7R6wRXaJ7UE7jDPQXKqeMAz/f
Xl80Qzvi7YWO7lFSeQFTN0vM/ofij4nKwc9tPvwt8RoVbI8NdUHMLvPqxHjfG3Rnkt1/DTvdvjHz
F1PR5R1trcEaD1DBIxZ+xsUywl7t19ohlSbOVw6n9IA+86kJCwhyqZJLGszCP93KytIqzWZNrvJE
yKo6MQutvs9jjAYowDk2/FYSO2nwu7qWBNICSl2xc59AOhHLROCWXYFj+i5Qhz+5sKO+pzus91X9
7S8QzJR9DNvNsvw+gxAXWw0F/6wNrVffIsr2O8hkH8Sed9uAA6u2rVNktRwPPnVQBklOrSn06WN+
qLzh8JvOYuj/9kkUtqqpdQhnC2ibWLhwzUUQCTZkruooGnTQ2385zFnhHn10B/58yyy0Sp+OUYcj
ii8rzdf15gzKHV5ugTLnuw+g7fetDmGLLAZ1xBpO6qRJoWVmw+Ib9zX4f03KKZZe5DZyLegsxkJU
oqlC7yRqyIw1CHL8Oj4ooxyzg0RF/HPY4NnZvs0i4tjsys4Ofm5ZYrSHB8k/ROCmpUWZJpo67vTK
B/g4xKGNAqNy8JjZmzQyRjSYm2Xply/Kniz6+n8XjTXxOgztMByKeefclLBk8sf9Aqvk+A2d2K3u
+0RFmkDeUorVrhU/StNhLD2x2IfsiHKtw+iod6pIR70fUPqtl8ITOyfp/HLTQUOQIUn5D24Tc9M7
mB50mkbTmBAGUOvNnxGKyKGUMAiwB+hc/ZY6AGfcQxRE9xxYG0J0irZaSRIPE6nMYN2BHMbmUjKp
BEXYML6LTqfpYiv/icdkmhM6Xqo+5vvs5eDnLF53aXSUuAk/WBAiWGxHYoOTo0bx3Jp7PtZUSw3k
n2vxzDoA1C81Dgqb921nmWplsDuYVTlH15doafHFYWJhMFhrqpzk3lmWUsa02Xsz8mSTi+ABF8Z9
8gFEAMNkMx7XPKRQ2fwSDchRm5SXgzkzT7+eNd+SxBPbJNxj6mfG8tJqz3S9/3q9blcSHZ2EUHjX
eWb3pYp64WzccdrSGPrjL5LCmgRP+b98sa+RUOQB7HOw5U8cY2JRHWFeE9ZtLA8v/bs9fwu1Y+WA
XCER9uuGjOjXK3UZSc3uhi3O0HMpjEwc4bUTOHxPjiPjUkYOEoX8++jjUkEvDB8lHirSXFuEuwp2
eJPX9n7l9nFX9uIjZRurvm/L2cqvoVsBM3c1kR7kCPRLdXz49vQQrCOfvCGwoOdHBk5V/ZcNppGZ
6ZGdSLPoVe9ta9wuKMm/y1RUCzrdijvxoaIe0nf4jQ3xdqPdaGmfg1YHr/POQOVGy0LtWTaU05rB
ZAmrzeSIG1JvVjG05lPveT1ljUYOQgS44nW3lwwk2UzJjWzaUuS5eegBsnXysI7MkILDxpDiaKch
QE+DWekhIL0FjwuY9LnhIZDppD1cec/D73QHFWL6CIP9dxjjubfGVYHB9o8HaerYx3+hOjlkJg22
kGnMJI5ITUKvlhfhFeIYghKd1N11BLX5TrlxYMs2znaLtBGvqf29mPLSR7Yt27ALRYD0jCJQE2+H
7fuqVSftxNEFxe3atpOKXYF5XYTXU/eJ9yqnPBVpJSTN4VzIKC11xCAelzhJWLZIQPeTcHZQt7gk
2hi8aZZcbElf9bATapH3fScTu1bWHvqh3gc/BeBekJhhWmub0UCuQqzTW0G2DduFidyWUP8T7T8Q
g51Z3CbD4sShTkifWlEtCDut1ApA5d5bIw/NzhjqyRTWm6dU9lUUw/h42+V7+T468gc007j07Fb0
u2d/DO1FDa/z3zNtHsyOoMELTP4aw/10beooHkeGU6ZRFv+IIlsZ1c+0F4+eHvsCd124BkE7xuR+
33uW/vSDO7WNMR25AcPxZzJe6zszC9C9pk7jPJyxQiJbpd6SnvcgrGz87eqnU908IAngbz4Yn8DZ
+p6kWkBqudR719cPo9tiXnJjr/bjvmLOja0Lwvi4uQFvcozEqf76ez/kNBYSF1s0Bp8pQr7AFEFn
aWdik3C6Rib6ipl8Cx15naxeoFpU2bh+aqDv1fWNVWIAMl8WOkPGYqt5plOSVDWBdMKLMbmrg7b7
lHB9/pEx+ZGqoIPWepSFswthB9sRbc/frS4PenOPtu5AFKfrhRGK0Le931HK+Xkicc/kPobcHU8s
ZXfJk5AcstsoimQbTCDJs3xdv6Y/yII7VRBoiGa+JEvy+uSAsqtKkA3JOZCiifkEYs9zW4JwYL16
NQZZUsA8upUFkiiHvKjZMBAuOYrfcoyoK5LzWDDCZ1X48UTCgMHN+C3H3InzupB5izGMsqykGWJD
jNRqRXjgHL1UFKuzIrlB1nDkNXiiIBmhKmdBKayAryy+f2kmYPUbBKPNWUxSIN7IfHgqPMkGZ/zK
yvVJ4Gv4/bRwwoFA0JjjT7JkdjQih94PYcsUgL0EIOYThj5Xtj3FUW04meaCyuL70qnqOfKQCycu
UbY9+ls0VcUDihHvMrGzRonMTai3m+PhG5gLUpFlHkFp/+9HN7YUOak6f0QM+4rP4d3+Pb+KCvam
aKOZQGFH1EF0RgnFqOVp0qf/w3J7R+3L7+Gl8nvfUAFOMGfbBCgx9+GB/NwXFYF0v1XZWhvnFyMb
M6EybgcyL4dDCaQjLL6Q3uHQEITrppoP3XYY0Z15neXgQu1fu+Xs6pxAtp8LlS+8lLO2LD1TRUfK
jFWOo5OAqWXt9F4p+nKQdf1CHXsP3fIdDP4On61g9DJ4yGPM2hX3GBW/wQGsA/3jHOyGn2GTUqX0
d2sobuuVSLpzarMQmSAZu0nhkDWBFVzfN6cHyV2ElfwOo3vNeaa3tUCLXqJ8XZAQb/y7WTJKtkQL
xjbYgifkp6LjDaFkN9LjGfSiQUqqCrt78U0IWEGy2yihfSrnmiwQbj7NwSqJEWaI71S0s5mu0oVZ
HfmO+rWNZt/UhFhLTrfBWVnbusYlEsS02uziGoXIe9Jl2QOZ+3VedSV76XfWZhC0GPFmVUE3vCYv
8sw8ah68kaNy8j80/Jb//qtzsX2uqY+OS7s4Kb6Ud03xYNdTA8u2xF3koY40KCU/b1/9OZ/BgyaZ
NLOXr6ID+0XgIPFR3c+/AU28i74xbLg9Q0hzqcDljLbvz/TCmTIQLrBx/ehquaVrQMmTbxL8ze4K
xZBWkfYOlA1cY2R+fdE1usu3hTvRU/DklxS9vtnGrb2Br6CarGQ8r3n+gIZsj/26OqjayY8/GdbA
0+NGaaZRt8XZbVUZ1dEqisHX5nvJ9qtV9kMsv/WDkOdp2J7YpDGGVzsWpc4lWRHkfgjj/BJSbS9a
0ACOCamdyaGCPsrbaJAU7MT4+KzEPznmJq8Zo6zwUFhK/1K7mIb0yLMfK9ND7uXXoKcqPd1lNZBd
OrzPjARm/bbldoR0E4ibH/ueULRxEHpGQJ7TchsQmfjposOXQoPTFR1VGiC5KyqrhC9hr4Fxj17c
E7/q+TH3WjjiBjyU5UizLv71h37K+RNiQBIKz3y35UJXMaIAAADVwdQC1mIdRSpT1CCy4por7s+8
qAYoJinZwkhA9ON+4/UKUOVeugBXOUMCyqPRkC0SiaKUK4PB7KEHD6kpVzkY/okKTqXsXuUBeocZ
uptcctuHcof89R/b7T3J/uOPIaAr6DEu7oyEXGXK97rQ6JwydyeDqe5TR1Idea9OW/raUm4n/p0w
QKSTycjGXKwtEd3XvtOQCX8NoX0aFjXADF22TxIy+GyFoftPWr6lwXgU/dvjV8sn7E1sdubwXqbk
a1banfnTSFWJbVFGjcJysatRFMxQEZ27UcYPwpJNAbJ92MLHvqTgTwJUn8NmFxNerpNoyN7bctGx
GuLEIpJ5cVP56So1Tl1btmLWGQ0CXQog0i3rQw/3dxqDQJ/wHgXPsTuAUPj1JwOypRI2Za+MLc45
/OXFPHFC+/SBHcO1gEKPNtLcaTpZ+/1DMRodcae32CPtUd+OMogh2aZk8W7lIk+vLpWoRe3qDVKL
hrp0AB4GEf9GIsNhuFC4tnTF2BWn8xUpcZ9AaQu/7WqzVMd7HXYJqS9gYRJ3rWXABZikXq244/BI
HQ/6pC1SeDUfcn86mI3gEoX48KmE8UVWhvmaP7rUiCP1lEtKlcsJ4I6kQakuEh9jsNXqtl0SHfOy
wQ4l4rGk6I2w5AqLBXxDQQRkFWuG1sV1PPStFwBC4ZMLBdXf/lbWkopwO1NUNGWlHSdUAkV5eW5P
EJehr8K6fYC31gDkWjQdUpXbnPDgeH6Z0a06T6asclZOa8dG75E2yPH7VvKXugRttg8jQ8rrtuTB
KMhrk9vNsSXxmN5ZgdYKRiFfP7V+lbKgi/H/dw74Yx/hG5JUVIfPSKKohbpDb/VjtcQ3RpblOWCk
esqTu/FvxSkPKTKCMrJe5A2UlD9UbXvB/clfV35GNLseVJMGPnVCRpWigLvHVj4xLaL1QXjQe5dB
LAdA9B3jhvf5GHiFddLrbHh8iVqiiEN0r7XBcoIUWqprxpjPZ0eZ752N51fsd3NAYl7UccCtO1Z3
bsqI3lgppqtTRZVqKccVPjHPtciQpOVd8WuPlwfY4lA5NlHgVeWX72YtqmTR1EN9/Ui5LanIKnEV
PITiuQqzieA1KTUen4C3WAyJitpt867hcT2Z18RJg4xIS8sj7HUPwH6hPuLz41BHmwv+G38w3BQx
NZCWc3S7z1gM/RJU/t+HtJHnpybUAZ+A6wKz+b3kDyHzYginp/vMFAZ/Co2M0dRgji3Q230ai469
7sDSm2EVoR549gk1ZP7OB4MTtAVKXrrUaIsPybH0qMmoYhw/GOlFj9F/wxmKxdm+XnEirqEJL0NT
UrftFI5QPfd64dtVrQ1YkTVU+rvHesiFrLt17MhjGDM3xt7rhNSoXXz7Z7orsdGumBp1gMJ7Z1e+
cAmaVYNh12d8HBV/opEp+kRgNj9Ikaj+cepFvql10ashtHU2I9HG1dB92N396ndgJE/4fIMxuMaw
sH/FU/bGSSXKVJH0bvBu9bhQhxX3btyLbtw0iA5t8vnpYTHft7hc5af/BovlytnIRHqHHJjvqGdP
fZ11j0nwtyrHqyTP8jnIEOMT88pJ6ZtlmSnLAW8BEgkKUp4sxKeeBzex4D+NlJy5Liv89KTJbj13
nZoTzr8SCPijmuxzqDFqUq58zP3j2sQEW7V01AjHNL9z0WIzl1fMscv1LcDxSbbbyzpUmci5dogP
QjPs0eE0l+chz7XWtom4qs4jEiFmm4/a2/8FubAzfxZWPpPPJdyMVgigw8Fo9w/osl2z8EGmLWe3
gHcyj6/kRBWeQBMpjYlhzTBv3f6o27mvJFxpDFF+HQ1zUgW/4iGsHpepnq2YRoyPvQmPfUuIdJis
oOtN8Wgnx1XO5ITrIBryEL6OFd456s6ohoXiy2Lq5gAJywal3IpiBTqCTHzDxYLLT9qzFYU+MsJ9
HC8+tEOHWCL5ZyUcqJXzkEa4q8x8isYgKdDiblp99lqAtbuLvatz95gmY5DTFH/8pHMdi/T+BWEw
dgMdnprm2NKr+XW8SeDcDLfMCpXJqlozBLKv/b6I1n6ITIuoQE0Ada9fIyx/bv3Pblx1R0pmtBb7
o+3wWkvKN8jxZhGKMdwNI8Btm2EnXsQY8cZPVirQsjEIlTDShP3d2W44Fddr3TpqKo9OWP8nqSQb
ofoJ6PBnAwcU0QXjRU5z6XBZHUpd65h4QBTFUHbfmG1lpDM9tplkSXsIc2vBWnucFiQRTdHm0l7T
vhMbA+GMd7TbwyZGLA5KU4pc5sNPU23m2DgU3w7ZP9nCvSUdXBvY4gWno0NNOoaMGG72dueaD6XF
NzLvZpsZVg2eDj1lbq7/j7P5taixEjOekz7nwm0Hbij8U1zu2vrEVQt2Mhvw4sXIKpiZFkictFdN
rhxfjFSg1Q1wW1NOADLJPJsYw7Eh3xskGQIKLMUhB4XLooMTbzdo4T2YCQrfAxywqPL4r8B7UUNM
wUZi9ch/+37XCoyQRr4dJPJBr8SCDPWld0kKRHis3hD9JCviomRhKo/ZM4jzCv5VMKvWODlvBDSm
BvG7ArlSZ7fF8x/XuTRMgFJ34RooK3KZiRj0sE2ePaPWmbHsQFWSTQP7BcfvkE6wRfIiMSoxMcVi
4dCu2gJnmwmw+64wApGsAuwKJMbbrg96t2kl5Bz766nSaXJuP+adeT/4fPJOD3hc3+BlqJMZSqQi
t1epoLnHRRxxmfVD3r2sSx3KxgFcnkSf90dCeIl0a/NgiMAOktUWSGpu0/MUD/uJc+nRq3eGQoEc
Vfe0R6nyu5s4WcB3Wy5kasiP1IzwEz+yvE1+CVqcVXeFqDXCfeOP4edspaDL0jlSt75qd9FpnDoK
kLpxKhBccM2xz0Wwh4z0y3drwWaVIMO2ui9oWxYBWObM7aPzSr9KL0WpdwG24RTNwyup+c1OJkdL
z6wio6/ufEpD+OiEFOUV92QEtTLozY3e8l4zZ07K4Je+5rjSLDR8U+CBu7hgMxfswjjbyejid3HN
JvZ2wX3TsS7RXv6NyWhcV8grtVSL9mCwDw41obhbEpgUBNMZtNyU9/ropTcuFJihcmnbw8w8gKPQ
6sNLVBV8ZjgKtuohxveAeEjK5IGHolIvrXA1OwAFld8wGcoY5mt8OMwp35ooXo/F48jVlpKTJz2F
zz+UFQAl9bK+PRqHcedTUvZbRVeQdzUigtG67eRRfeyn7vbt5kLaaXKtoUCyE0/rZ+KOWq2rSxZb
H+oTVvkosAELf68GQolGbO2xe8WbuY5qf+RDrpEYCdmVwS8J8FI+nmV2nnt7+AquTN+9J7dDEHsk
BNnZR6qSpHO5bJ3mSWwbtJ39CTiBrGhuoEYhWzhUGvb4jpbm5oBXlWaHxbbPLeTc/N7h8DL+TDiC
HLeH1lIaFwUmyOTUE3XLq6pPKTBnAyFiIgrRghMSocjejaLCt6LQUlf4UmtFVZQ6skYeyB6TBJz3
AKl3u+IKODgqSTBZkOeXB34ZB7Ji8LCPlLPWG08IIbfBjmL3yv4b5jQHsTxlSY8TAg42vk6/mJje
nswn9GOx5S0hbQfEeC97tzoWkpZF8TrA8YbrpXPFjn+p/UzyLY+XHCT5GIsrcnyGXtzq2mMQKOV9
vDm9VlyGvFt9cXq7x+lixI0IhQgJQqSiDrUFvYKPux7EES07cUnot0MACagRVNEDP2Z5QxtYpHM7
JwOM0e2U6NWGWA5YFC+tWy3WKYlEi8mPj8BLCFEdkEknQZmA6ZLrlvr/N24SXx1Tm7crYOExDo1U
whcWlLUELvg2gp+r6mkmqK7fqhDYeTuSipyHd5mMAAxzO8Jbs8JKj2bBDcqfXy92+HP2zGeMefKl
3xcrtm9vvDq0R2ZpQEPaE9wdzsaZ49dypQu8DBb7P/8gfv6NsHTk1Lb+Ot+MMPE61D7SrUDdiROK
5oVsstwhzLpIuyFIdN4psl6PAGuDhboGqRmtCBmllJxatuBbG3kWzSMAJQQE90yJFr6R15iqMg0/
2UwUusHt8mNjhwk58Bqhlb9fOaIqaqfAWtxXSbbwcVyrdj/8jANWXUI+j8m9hNS3BTU64toJ52f3
cWJ8Eh4m6ZTrPUFs40hCeOTDOj2LzPfJAGEch/la/KaZC4lRgIiBAb2l3t1ojRU//fLTR8cgtZ9z
1gxB9tU+hjCZYO7IbDoIZ2Jv7+0+eWjzV8VJg+JpcLTqLBw0QyGmiGASuX0qpj4E6TXEFgQz9LL4
l5bdcXEy941HlGceIC5eylJn15L3QQz2Wjp7fiTGqQw/uzdWWPfdpRsfw48ACstdol0HwJJSJWLG
PfGbNT7IeE0NQz361DUGG493gicCNgCRV+GwjmW+nTJURF0gBytjEql2oXFvFhEm4h0CMjhZA/qB
fVHNaer2iBRH9Xp8/fKJPxg5is/eAb4Vfd4llE8DeldIRR1s5lxxGDr56QG9+SSCcS5tACD2Ye7i
9+TPlBN/25bElWlhdGGfBccyi5YTIdqVPzJandCcJbdzXSvejo2i/CYmM23VHtMJ+ds0UypkuGYH
yjgpsQLXQn2wQbu0+4osgsnoI8AwT9DgNh5VhNvPX0/sXhrnWcAVlQ22v/pGK8aRgxT2ToAyKG2e
hYQJGNVsA7ZqvCCIGGSgf9TDuQ2kiWPP+Nwuvm4APP6Zs8kKE4XJv4D01akgGOuldQV7GYCtC1KJ
7+PyajWg4GU9nft+MrT4Pf4QmKYKt6yOmtAjW+q+chVorYuG4t6zfIyxbY01f+npkSe0Q/AFb5xL
I11PLxd3pw+d50AGSz5DH4JJc9KIElrqkhjjPxnNH1hQFVmdPYrgOLUaR1DzLokucrkL42/Th7X9
Y/l6po6YhDaVhRZtt/YP/17mIw4qKOAzM/Aht0DWS2MAVmbjVOPoyw1mMDzTH42yrgPjg9v6Q09d
avQEkNY6XFaG89mp9933j6XGFD/OGfVtBlNPjRrgZnBhlTQstX0OJAn0Psa7jtHOzK+dMHe/DQ+l
MZK1KI5AmnRqHGnajQMpRH+0lh0t+LQggfSmgMv+nD6VznXoUrLEOUbgfSkG2miRUe2FxzFl+gR6
F2fkZFLtUQhyflWLMFn16ou6OM+d+jfIGwz5SnHIT5X4EekubYAeW2NjU9aofe9XnAHe7e3bIQUp
1A9nfLsr4p0VQcbN+ZcDSAlsiNzHKDe4qPYQ2BODV8keEUea4NXwlL4Cdd2PX02/NWYz6Qwhhi8F
5IqzOryRTaXDWxY1U8NWUBY7rLH3zkS/Ml+c4U9cMWOMMakEeiOEQ3YGU5zxplSpcutC0XkEMRaJ
FXDoJAhTn8JZUmT3tWo3G+olebDrHAh5kDOdqkw4VewTOd5qmYjfSVEvWbP+oqNUae6s9oLoEsRf
+99482qwn4oqGt0Fey4UJY0dtIK1gMlzb/pB7FnJ/LMKUSiZMaV+6mE9TeVoskZEMbpGLlh+OHJG
e2iZ4Si74nLeUFHLS4dn86ecP1mRi1b/tNV8qTuJdzr7Tk5VbRsOQdMcsBkGmtnp2xjUXeHlobh1
ruqDz50dyZwq2Cxt6FU26427HGDIoUtw5ETzgDrk43J2naNMoYyntImyEAF92/ojvi0UIphGq1MF
rsPljtierjeQaw+K+/nKMho66n+V1lMJqUnVHNFNamLKRsk9Hs7xSnp5DWOOxXL643AcFkk/QnxA
vOs753P/R+IdmenKVgYaxJ04ViX8m5EW2ABElfAOvf8EEK04ehZRJ8KHBuJpG9WUbC84K425xK2a
K3CEJL49MS1bRP0CgFncuQV6yjNb1aZepjWFdHovaB3tJlA0WCWMucHh2/SLXw8+ECBcSFFq0VCt
cLTE0vL9aaWhA+/o8tKX81lmfU6OWH8c3/qnF+vuTfW+XTLz7wbQmMWNA/Voydlt+UjxrLrUKUtm
r1bJBwPv7Mcc1ZE4syFqNcAQ/0BNumEsUTkMquiP436gn/RnekPZ7vjPNQ7Fv20GoW/iCYCK6suT
qPtkvdbjjwXUTNFq7CxZCNGNkAQ5git7edWvBjUajjiktndlZ+EPQXDVFzGUuO4S3UHfa9JPrM32
ZBzBHFvCYURM/4z0ULe1LDDklhi6qI/OpD4xkP5n7E2otgxb6//LJcTii1z1007e53o6YkNjAUZ1
k2UJkwnFDGcJKg9SjWtDx/G3zj9w+RSRhFoe7U1doIik/AR+oPHiURltn6doI1iD3UdJ/wZ4mjHR
o304ZO0Lc0e49agtvgKuEZRhfi/nH4F/rMAA6zsL0qgJbfPPSbzubnrukti3ddmjQOYwplf+lCEE
s69eRLwXjLrg8SqUMJt3LbTi6c10i/MtjCBm9962EcCmWKQEScAl9ldQ/yj6Y+wVFbNYp1NwqYTR
S8F+0UWxa/UjU4ZfLeIQibzrT0kOkfL8PmkyfFRRE7MWfkJWUeqkfusBcQbFUAyjwzHUR2qoz9Gg
0ktTaK1J5QO9/tzQU7IGuljjQqSo7R24m8ScDUSOQaJy7nYxTYOfqzzEa7CM8pgev9x3n6XigTXb
xGUYEEHcWGTgSDsoR4Qa4ckgUpe/ZRdQLamQzs0t0PwZe9eXMQ+0A9Uc+6oGIVLLrjxqv2uWx4H7
3yu6QKRQ1wpnuTM2d83+GWKWxTzAR0Ch54HT8qA3zOpwIHX4aTEZawbHnUyfIRPr54OO+7TKLJbF
VQU8KTFP+795q/yfyI0p17f63/TFy84lMokce6aQSbcDMiJzOA3kqGA0KLHiSlTFLB8XJnvvqh1V
dZqvCogFh9u2iKnV2pa7vIo6ARFnvfvNlYwLTe/jsfvxzxLpfLwq+GMfJqSOgB3G5WPC4YIxDvZi
tVhSPkIT+SDcYQhfPWHrFX4aMMfO8XyfMh5aTou2ZTeNyoGYCRSNZsecUj0Yp9zTisqzdElRaG33
n3xD8lA30jNfJd9b8dDYgM1afxUkse5dwp3oSVYP13aNvZgD2YwmsgkRcxs9jAz44oQnf8G/sUJX
eX2srbPbwdSupeIflk+JKd0RruTsrgCjyu3FN64sC3/jxW1PxRGTIOFZHDXGG/zW0ycX5ZZrRvqx
CnFg6YWFhmsf7iUwZieN/uyGPYAX8qjxGhEWDu4wr9Cx26yUZ201OMakBKbbLPTO9I5aUXd6bqHQ
ezscQQygRjCm4WZMPrj6dQS0wgnTz+992P4J7hQuXD+Zqt6jwn1ZYKCr2rnwo+G8l954kSlwTVRU
psIPx4YXz4dXOofQADe+lH/mjY//F94JTXBrMr/3EGVaMevFH+BEHy9m6ZUTpSYShq2gZRrGTEXP
K9NXI7z1wzfnIqGTuQFA9Drw/XTgiJf8GZ4gd/siuFDQ4v/nqKkwJzPBjdljTN7fQK4EtPA0YmlG
VuDCUbEO7Zcn9ighGJFnJ46RujkwU9uoeCVB83OBMNwnY9ij9K0MKbjcYB3Sk+DWsFIqalO2wnxI
Ipz2p5c395ZcznTcq7OUrC7WcY7erheYzjFJLDtzsXeL68lhdd/9qt9tGm3wH3qo9PRAK88XZciW
vENlnz94HSqltUH6opDmC5VB3RC4iHYrCtRaZduiQ3Zkr5FuHv6DxeTtrFmiDot+bPJ0XyWctccy
nR/nzhQmZmxoxoFjX2D0LSWPlV1we2lliwRwPfitNJ02nRgQzmaicvJIwVpLrLEaaHCu0spaX9gh
UMkco56CHx7u5tzk/Wb4+mu0DdbvyoiSHkRm7RnsFr647TE42QRoxOKIRPOMp38qHEvwSgjAzt2b
JCR601/Sj1SSfbB5AMx290Y/+JCX1LZ1r/mAGPxlv1jeviUqj441Vp79TjRBJRK/Bwd1ogHzaJQg
Ch58X1o/Xc9a3HMO7q4OwN0il7QPKpHx83G/JQbp5B9ckjNmxEtGKXwUUPCv4wzTgIydLJs3aKoy
fWq3nXn1zmawQWf0Fwue2aleaKOcPq+EtV3cwFOr4S2xUgSuKQggaQdmBAXZSjupTIPHlGyZJRpb
auGpp04vRjlDYzIyp1lEkXEXnN1air4+xFHujfYxMJINmArDDMRj1YcEKicGZmRcS8ty4E5evD6L
NF4J3OQh3TS9jEhEMTh3KlshRbwUaWwwQ3WYOmBoO8hydgRsGCUZXgNb3Ui8aMfWCjj6XkTte3be
MuVf8bCVNk1Z13tjufE2TYj61vYeJ8upjSjtrkgT5saUSBD/PrT28bP9HMmqVGl9whshUsUZ2FlS
yQTeqjQi/KPvFyi0P+FnERFPCJNInsOEnYhOG6xyqN+l/pMTPsjWlhh2aEc7DKBubTP0qmBdXNTS
n9MIkHxgqT+aQvVy0b8XcSh3cz7wIT24l5sQkxrLUxstSsphEGSgj9F/4BH6dPI9/zIsHXAxo2c0
elrZlQ4/VQCR0KOiKmwRAFSNu24Df8rZ2rMHZpDlaBifTttGApFWPyDR9N+Aw2yyczMMI8SVshbn
1JQ94dWwDSUPly0lFMRSSr95HY8JEjvHSg6a2J0wuFmN5C4mVOSx4oLRZIB6qQfNoSYaiwjY9awU
VyEDa21lwjYGtRhdTBqXLmBIBu2APQEy/B/QVh6RD4h2VmSUUFmI/kkV05madCmSdumTXrAvfN58
614LEFAvDS8LI5HeHpoYtSPQ+DTv8TGkGX2ngBBjiHe9uRP9ifoqBrwOXIKYUVjE6XS8l6A7OG7Y
aTXe8CSYZzgfxpL9xmFIew1VBsUqiXSMBLVCvwWnbJTNrlC7yXz1yjvQ2CXZI5kFfAZPjHES6vZR
TFoT2tnG01bFmdwhmGkFK+Kn9uZZLs+I8GhPXvCnDCqkex53jIxrnpxa86xOLUMtRTKxpkQzZQlw
pgLLSiisVI6Uy5GGPtJju7CvF7xGSA5tjUnukwfATu8mWfFSUkdAW5jtOqjMxfircefJZUY7oZSo
cfK071Y5JaU9q/XxoytDUX5vLQKeJnfdjQFafQ1fbSI0+vpNWSt73EOvdtQjxFvpSnlLw67+ol/g
GVomTdiOIXShtw4lUarpyACa3jo9C8pMc2Um+sPcEd0l59ppjV9Aqthnv1Bmtg9H9d7L7D3Q0TbW
Ywu2IxRdLBOVWidmpVIbeJegWLytOLRuvs01YPgo7gRaYblEFMMOJP30oy5a0/6fca1hjiq7z+oM
1KAlt/El0cwtHa8f4glrAlu1vr2HVXcXS1PFYCZDJTuTIe+9xkSkcecaJB8lWwwc8yt5XK2SCgqr
GXMMBgx9zkLZRccYQg+EUg5wDTsQqgGCQ+FVsjcz70hDQ3O3gfOykOOCdKPaiWhjD6qJP9W9hcKh
EvIz2t4mUTPyz5MMFpR/VFHr7r8619WCzEC12+74v+X0mEv4lRpqZXl4/+gL0hOMi0Jk1PAcLxTa
86h4xr4Df2xqVgQxPjcIeXzpy33+HJKvnfeTRLPghEP2E4zhuKOjVcgYnwzzOdmyIqWGFxjqirSV
uNVlbMho7nrAfS+ruSvdaWC/2nn5iZUy1FLTjXGuB2GHhOQkl2YGHQTO8vtwijTe4qfSKKTYXL7O
EOGz2FmxrttJW4qIEiWntd4g6PUfeFZcQkcZZNHT1l/t0Gb9JIKnwoDdu1kZH5WpyqIJiETUa+Z8
J5v+ZvRkuw3qKZZu6KzZTjeO/X85JTA8DjJGYj1uARND9qsCJptFXrnV9dt4aXYh5PHNk2wttOLx
pWSIkEk5i3LNaz2OcHM21MyFp2wR5xWdreJKyw8XlESxp9vp/1t0V8HkqsLhMj5VyiAHr5ySYJXz
zwt/Tlf8M87yDY2FsaAYM4EYkJZSx9QFvEZyWwuQ8iYBHgmWQgSFiqSd5wgCNhGxWSTLu7wTBkW5
/5jopkEnCEF7zHCMyhZfF7RUZZg2cti26Qrqy2y7okK34Rh3XqF53UmpK96MWFCRfKWDHGufadN7
O+2umu60s6iAD2hFQALjmIOVAaSYAnyScBCQQleiIQkD6qyu/LB7P8UB5AwT9Xq/I2pg1pHPEazY
5P2Bk96lAejU6h4ADH5fsP/RmkB8CLe4Jbc1IMbKFwnzgx/D7z4V58IZjxLsDG8NS3AvZDgp2haV
dqkEjFMveiqFwGNBUCqPhBYwuDOSbZtap5Z9R8R8tNhO4ZvoWpG0lBWq9LzrfaqsVmTC6vpEhiQz
oOnyYJbrryKGnOZABRuJGShPonvsz/MY/TWV58UgiS5OrS2ls+rAnGJj7Kacdz/eUZG3SVUqpsCE
fnwm70ILgCBmDF+09l/Bu0F2l70hugYcWINhdr03Zr3ziOVgkPD/x0IvfSAHvLG6/R+ktQakYGCK
rUXwVtUaEbM7DMyct6K3aA40Ea2IIuXMiRRQwITvsQ1fAQ8tYIMuKmwpInknUImjzl/QFrJE/Fhk
KwGXwzoQcXqFPVd4DCEvfHWp3WriK1o0oVgvf5g84BMmWcbXm8gaslo/HJF2WVOj2xU3f0Nxhbv+
qYBxJXSYb3MIlrTFO+Y3elwsFq9kiLJq72ktwUnkTrbJlefT/gdlUvZ+q9s//REOqohBoNuVOnWx
hMnKJGtnx6ld7gBfHBzcWG9Okay6w3i/Ydv1rj/7U/fDiNd2lV0dxLwr56xDFDXR7iTcMTmCeo6+
JGHb0ehPLnkog8/tvDDCD9QRfIEbLJTgmKXG2PBOVvFzAmkB9g+EwJYeYYLBLt6pZwKAaspkOmYm
S1xYCFVtFDMdnfZwo52GWv0tQhp8dDs7O8y67UnUkRC6cvZ1l1Qv1/BTDA3uuYvyPfo6weZpfvUK
XElGBynWdvIF+3hloRkorlrEcYmC13rOkMrrDJLzqH8xO6WPgSyVwKpKsy/1nCg9tmGLty2GWgOs
Ed0eNbOJOPdSRiQuLBPltxcJi4Y2n0EKh8BaIws6YY/t/kUutffEvldH1eVci8NpSQPrgemhhwNA
VIdKmHmWWkSCSVTNp1u1fO3nGaVFwYJk1A0yC7Jatod1Ni4OsOaZMPLdqu3+mQTgKWld0khJX7b1
KHkl/2WI1R9ma1LszQG9wU/Jff9JeQexamsLDT0uYqhy+GPcTV9dljC9fdpWFLK4kT7Ih6K/gNlo
cN2fzSPpepLqwY5al82gmgC7TslNLqCMwNLux8t3JS2AWtlExn0gFjkmNf8y2q32zLDe1eY2i444
kTwoV+dnLEBwKroHr93Z3b1ri9wKpsbJoJqzVk82Dkjw/PoLIAsbv8ejoyk3kQjEFJtlTJKRdvlT
YVvJYPaNBLOsrkrGkweutH3ZXOk4ROyOhcq7PG1O/3JUpIHcznfOh0Pc5Jo69BAUlOJ53dC2dMvE
tgrOVK/cnOijjK35L+l4KxKIIc4Le50UgHgUogKSGrl/nMWg/EDRcSFkXLCCKhxeiR8Ymg7WzZgf
edVbDh1KAPhq/v5Ak3shaXyQJVIpaJzZ/Pvk+auXJuOVF+/ARUShHy9dVitM9p5lfh8uxvm6wlUJ
70WRVi/2mC6E8Pwrqi9nnTfeSYufjQdDxOZpIN9P3qGYUP60dmDs5pQ4pUhab7k/8bp+XP8MmiE3
NKXzLgL849qdVprJd5wj02Iqz/3bDiGL/jBLGS0WRz+FW4lKAfXlZOIfMGXvipUEE757pWXjEwUU
t7jTNm4tBnFSgYdY1eIsu1KTXJ/dPDNyjg0iTQp8pgya68p5fwkY/eFnPlK6KalKaU5+40hBgCQU
PaB04d2RZDDuGbU3ufCQPodLxt0XB5a9qPRfoZq5lxQnR2KuvGuJmRuko1OoioLRWUT1FQa9W4DY
1yhJmvPgiEjVxTKe2ZDU4etff7OLm+I3vu7oevXNg0t9UgU2vmDfWT3XHSA79dscyMcYqGoVVt91
OMM2Sx1EGg28FSCbllBnILvet1fh14OFUUwBucqVcyZRsCxCgoGjJB/ZMn6iGxYWffq34DPr4QMs
tEnJckn5Z7UfKE4K8R6HACkJOT+SPs71BkqnN9CR6beSCFBw7Ya3FT7UUgDTJteWPodxpGUUXhDR
3JF8dGEfpc2IKS/2J+4jG3in68DbKyvF71waahQn7VyRVbxm3Fsfx2DJsXVWn71Moa+N631DrtHt
550Ig6tgKjOvTDfMdmtqYSKq5YcFp1ks4f6HoyiKtjqhYopN62iapZbt9/gaiXghmdLD3HAMt5qR
FCpX8WcM+w1lBaI1OaOodvORt9h1aEUlhFW7Ghr72jhrlzt/0+n1aVpdO3guZJ+6i6Gfakn1oe/p
yeDl8ljR31270gu+/PAlFqKLJ9SU1kami6+YIpJhHaYXOXwmLFKsEdnykOjFO3iewoMJFFLC+uif
E/ENwMcRFGAeVL5h/FFcgAnHIaeqsmLxZLZ4EVJffMhCviIUy4f6zQ18M/grQlMJu+6xhbJihzac
nPwOWa1QFPVRxMEh5MFUCCL2ffxYtlLjGfqpZDzvdSZ6fOQWB6S3914XFFuXARB4Mz9PJ5cZ/U6C
VzKKUrSKGxNXVaxe4TY3446qlzCJuiYTZ/OR8gfxLe58Ww/In5PbyDDGCNuj1Q7++gvfLLvQDySp
u9qN1RQTv+JKP/W1TW8Y0/vyXAYwJY/upUeX+G88+xX1HVZoJ3MQxVo//vFoA9OVbgPFaFomC0gG
vHS/gIKY+uFAdWoEFlOo7r+Avn/dZ2DjVKYPCtYPsDEFZDr/NkfxjWbWCp1+4hEofNctgajSgNjj
BRm3IoZTtQjmPIz5+WaFjx+gk6nnbFYQBF43BwPvBEgGKg2DXvP6WAKMNUK0J6bUvfOHa60TVeya
y5C+w3bJ0jKCKc16GCjlDJnBUoHc3Q1YA/MM+Rs14fJFGOhzXb54bABKtfSEIue3OS5OBtRgdFj+
UGIESRj4zC0xK5+FNzqqe5Q9P30dzk4rKzPiYFf/GM1h6jVG0hGWU7xsuwaHtakikGPgCYeElEHz
cPzTg/QjcoeUtODWoVORPF8xLCNIW/G/HS7UK5hIUNdu0uMR+tYeYORVPagWiHxVbJk2GHdvy+zX
1jVkjGhENApRRrk3Q3U1zC+GuBd9illMaMwy2dGc8QXBk+c+7VqaqvpGeNNczocFBTsdS/CtTOm+
6qrWpo7U97RDJ3pIXaL3qoBzWMZklu8z6pNJUYuHBdCOK5Gmm9fd8df6NAhj6o72ZO0JwbxnRI0x
Phx9itC8ZSD2klRkCqxhrWg7IUw9lKUWtxtqZ/N1ahS6U9K2+zdLzxWlgWnQytC+H8yzP3tLQrTu
xc1x+zVfiYMmjQmNTFYs7DnDRi630m2ig7Mgq5Ke08XgvQwq/foTMjAXM/4c/73+nvpdyjBQhG9m
maHB4XTzqiBEUHiD1rvLyYz1HkqCSzAQk7dK4gaiSsTQuD9uI5vEmTSmgmGqvTPWerhHK01OPqhe
lyV0zu3+Eg8RQfKCdMZ4RpBcb7z1G1cxnslfXrXRLy+nHNdOpawkdU+YEd9luUHIMwY/jKOH4E8Q
lW6S84FsXWmocjWk8JyPaM0r8nnpbl6Yy3u/laykidz3wlDNywg8B03pJjoUl2Nu2ydHPlpvZFX4
IJHPrvcFSkqu9vhSlaNC/SNPMPAWaQAXYhA0mOqG6P7TwSbxMyLNCIyLvw+RWySQfEMezSr+CKL/
BBcg1kYoKIszdNM1OS/M6wHtB7X4zgcfz9pnoIr/On5/SRpD4hxdFYWK7wx4+MaX5rwn7CuK2y3V
b04r91zsYnIJ1nipgTarxA4abkdQJK8q9880x41vLaRLyMJsNISTFmuSfH98PhNaJDXeuzTrT90Y
RWLKZiE4THu1iiMEo80BtCvFsuzR+dt2Q2SVFixLz9vfLm6Z9+uB1JsqWQsYy1lKkrdYUC3jpz5S
Q2dWsjMCn0GXtVjy3nm8GhenLqbrEkOEh9weAlxQTkCsXrE52Sqc/lsZGpF2V1Wr2jaFZKWzksfa
36mJVuJ9/LA1WdXsMP/ZiiCpqmwmksBQaNN+gausGSKjuTrp2Twu9dytm+TA5kjSF7L5ZkzYP3iW
bTQ098O1ZPAuh7WKYrFKLfh7jMY+FnQWv1GasfV72E7BxI4dgLIuITjcZ3LmwiFkF1rwq5jC+AF4
gX3J2QglN10r/+NBo90AqfLocFU32VuU7eAYhm9qAJhQiapwEt8+uf/ckpzN4oAI5rXPxatOvPEk
WAmjB9Iym9/LKzrBZRWS6glHWRnl1pPOINODYcIFiev9fRdo+66erB+xAxwZaQ4ceiPzZQ7yVKvB
GK+QATCtpf55CtTDuoRHACwOI0jnWHuoMQpuagZPSgXH2kU3VfVyX4XTD7nij1BmmPGRcpxVbruV
gBgS6UQZQIuHmETsfz6AjLdz/AqhNpZAYy9MI8UnFsTdC0K9vAmQSpgw7nvvD6v5fgV/yrH4ENYM
thkwcxVDsWI2rPkMVF/AmbIGNbZxz8J99AZtW9TFcrxuLS2vxCKWcTobHy2TuNjUOBXfuiG8wJFc
5d8cf+TO+Z+6RGLjaTJvGALXFy/iqY6IvKB5efo3Zlj5OvMYkG3wTjVkDsLyJcwq6LrxpekJyccC
KP0PomJ+2Sx2Kjpn30bD+TyW8Xirz6N83pseo4lTCihZjD1WCcmyuO3H4RiC7Fh8+TqbXMu5i2wf
BiW+KGrZIIye9imLSPk5/Y4GM7DKuaF4Nw353YB9XgG+TDo6kOxl1DEzx6mxzVmihAB0CEPBhdn3
/Ws7XLMZ7KwQkTI087jybCoNe4cseW/Kw0RJrJVUX/B0ysccfwL9+jW5MtSEU/bZpMmvG5rk+e3l
hkGAYVat6PSMSvM/rEztnNG+v3xfhuAdjAnnB+CwJSrHfxzdH2h19sbDayrXoDHXa4yEEfMW44lS
Kc4r+pyWwHgu8Kd21WUitgqJ4I4TtH8tnuKD2QFsQDKdFueWUQ7pBijjmwGXfSKDEJWOUPaXSG/3
lmqpXjLfge6aqA/RoZk/QR+sr03rMgyNmeexZA/FdJEeR/uPlYeki2Fc2mNeB5ifb7YN3l9m9kpk
RZfZQoL/BUXrrtuOG+Atnu7Hd+r2v4i2VjQJpCJbPtsYp6Zb1oHe8sh1giTMkTaDAz3Sz4Ar6MzC
gXlRMqSpfKpNucOKgCbmts/ZAAp3VmcqdYeJYeDh+Jon+R0Fz+mJewRlU5HPouXIPbdvWwllYZQ7
frCowDnm5VY6lW0dUkBS2/tDXr2LOr5nguCBjZ1yzkxPWJDffxvhbSfiOKq3u7BPcfwNXMlR7Dx4
oztGSaAbuAAZzeecdHuIZ7/40N9IrBoSBwIY5YZbzaFCY6ULf42odhM4HsSrwAFbknoza/tYcmV4
FmIUr+cBsW1uwTjuLRvpnOYfBiLm18JXn60X0shKkXg8VVls2PCwXhlXWXPGK9HvjsFrrYs+XtTw
RPcm1OJuHWG9oUxyHIV845kpnhRioLScGbaZjiD2eyHNpwB+LHW0k0IXu982/NinolGxaHGgV1Ir
tbJ32Ag7ZwW+zM3C9nvwnCrW4OiqNgrMlppcq0tWyadmRF4z1rCvNxpFmjFfmKaPpa4h3POx3L+q
J1UwJfNX6HCmUiASKFy7GFVZkBz7lErY8GjBQJYPQyRyaQGSgfZaOvtbIgaYVMjrFy8gRIv5/3el
6z7K+POKidSmAk+a12ibDQnDHyrrYqm15x2zrv57+aU/hp0VZJF3wz+isJ0vw1H7ZW6wGyYjeScv
SmrKAp2kz0gr4b+naYiiwVERLcZZiC7fkpa4P2bEFHzFLZzHqamZOYXovvy9lxY0v22yNOWPtEkl
UHrUyUH2IlpXX13rNvTTsZt3BFfQMst/8RfiK+CuO4nqY7dWKk+vpmkt2dI1i7vJnDc33E7WLeiI
cHLdHB+a1qM1Zu+ITaMD/GMl+XTLd+PFiZIrvPmyG6x0gV+V2ymkZ74i1wIpf6xHT4SaJSsi+UVC
USlmnq6VhRNLE9dPhuj/YaW6ZaZwhqzpU1DuGX4BJorgXG+MMYeh+Rbdl+fo4mWgXUudqG5tjqU9
Odf5WKrXR2cH/GEnA7PtBRLhjUTNyJeckbaB/Q0p4OHNSvoDQ72GiCetOK2J1pbmwhd0QP3R7x0X
BRpGTqBOVmuM1k0JMFt3/05QDIXGKbNEADYQltW5CXX9kbC90nYK/ILjiKELdHcX908wYGgOVK1u
EAgmMpDfOHQr7GalporZrCY4d6+COb73FD4LqxgdHKc0CsjE9/x30YIF1gX7yJhe1zYrPbT5640W
LGi9+PW8knggnIbnlmdxtkDCeL1LyqRxA2eUdvFVzMXlOpZAD0PSF+JaYOh4hS4/rzD6rN0HIBh+
5OVGTtk4t2MeaWv05cicCX1G+gUr052rNK6lv7ngqAznft+J6r6h/iE3BEB/Yc91q59v8Uu7e7x3
RlsEIEC0EwI3tT9JwVXiNgimy+w6C3GXlEg8g82NvCwTnMBJ5PXfcONz828xkWia4axpAR5hPERH
2uG8Nv+sKUFWC01oVXGlvjc6lMAqKlIhtyRF9k8aejRR8I0ui4KEZhj6aEEvqCUQ6FXC9iQAHjQT
Bm+u0nM8P1khFSqbWQGEY34+QxYQJe/jinvzCBRIhP36Vez9fVdLvmlOfnutI++bMYoJySk4L7Pn
VL+YpTnW+p0XSR6Kow+rDKWUOCAjxbjJLr2Qjy11p/3czRl4PD5LG6t1JzloCoKlQgmDq/n3dZRI
8xMTvvudiz2U/YQDlfpiAg2oggPg3ZOIcpf7/azt26ORr5izYGQw+XxrLF8HZ0qMNnDFpQovm2U+
qaqJAkUqxm+g08n3h9KgdA4O9wolpT9uFZXZojLiflDvOecpvza4neEnddbQF4DdVqFJL8nuM9/5
j42VmB3Vfn4WVukLehabtgPRSrwy56L8rrNK9cjtSqEM12WAfMb0H7soqMSxhmN/Bc5lGbYBpwzI
lp4zSjpGOxc70BfweuGcIQil3QdOGgmLvNdnKMpRwVsFzJzQUAnEjqlYotqRXt5NJw1l/MgvciGl
JGJCkd3a90lM6l/bsTQPh2CPJ1Sle0CyT54Y8G2GzvVNaoKNVEgWZdUpJZwzM/Iy38YOmyLLvbLP
5ZsRClE99hUnCqWq8Q+GnwUK9l7NMBPf9f9VQGlyHYKDDASOFYfleIWg5I3TnrWtckEtS40ML8bk
XqBQqlh1X2iiN3mghX9o+tGkiyjeu36i8iqFzM2hra3XJ6CWaCWFBlIARy848vHrPXDpTgh4IWVW
CkGorhDuaALle04xFyefRY0OPZoDzYoGUanGa0uYAbUPG7YIpV8O5gRD70n4U6gyaP5GaJIVi0gr
cB81okSftot6+flU1+dJez+dl8xGf9urg9jSEQ1HsibPeMsXe5RelaKcEySOYpFyDMyEenCvpy7V
G6MFq6nc0pFmH+EfQ4JKFSlIgyZN8p49U7cRWhXWQKq5aYT3Ru0iaH2BG13qtirP+440lvhlE0O5
S+x1e9++GhwhKLVbAaN7gwv3DL4+JMaAXrqeginH5KQ5T7YJwh++cz1VxRkuzChhEYWlhYc+taR0
t/Aky7gu6JPfOeYhKtulfDX47Ns9mdL5ivwBYS1ET0uHDzPr4FgR4RHKiqEcbkYDWAC/NOTezMVJ
Qc74UfA2T9xlwENd9yoaz4VXDXXW1zTVlc9inxpujfitu5IhGTHpkHPOA4y2YKLvPkjRjRo9OsIP
oiaC75Rv99RhumFwiaH7HW+NUUY6MlDLUcj9KImJH1Jc4JiscpBV6OBjuRMABp/jPeDwcLJSffrL
rOKl/AbRHRXNihljo9PcWOT/wRxsf+hUbPSj3ltrhelXuX0IZq7lLEnJES2oB8F6syDExGezGOVm
jo+BdxDdFRG27nZSOyCOsNtnPou9EGsL+5RXy5rcIBjURzAQs0AzmWMELfg12M839e+vZKsel0if
/YTGNRK8LBrzHzQRUMd71w4g6qcKEw3DvU+bTo7+fYem/1bDW0/cpKoapXZ0FQwFAsS2dyBGUw9/
ks2Ue6yz8MDNiACgJAennkC0O/tutoQNXjBaClqFzQYgucPoLllNv/LQcie0D9GSINc48tJxZE2Q
3ohnlf6T53i5V3mJlHWexMVTGEngKEJizxBg6QS8247Jkk7y6rQXUcaqOwQwNtrvh15WdtS797Pg
fPMzku0TpbxvXCQWRtJJ9rPMZugAbYPW0SeKmJvOt5wEY1HFyFVHnVt70anbslquGRpF7VHskdvp
32p0JGh7Wc2EKBO4H8LWkYolWC2fJ1I0rENSsRmZ2QF5m3UcpOrLYF3B4MDfbV34BqsCwsoCOGAu
o7FcsUmEwxHzUzqDroRNLWHqBrfyNXDXWvWbBEEFAT5ysUNfdFAFOPHPPlxr4ESy5apraucalGUh
p4OBlrqL2d2HGpqZWO+GuibTCdDAWMB6YNS3QVecnyzQYkXi1mlTwTGDUxF+Cz0MVxQdrebzUpBY
k+FM/t0fPC+RXYZSshqKP3vf3siLIeLLldm0haRkgMWILQPqfT/ei3VnuVw9Xdnivu362Yqqfsgi
oavII8Z5h/4XLOAKns0+kDE4vl/Gmf0oIKyVrvOyFTJpBkM/IDsNWZ6PZ2APY6yACWlvEbanvl9X
3zuanVjp9kHDOgCCjOjRxrdERLK6xglMuUMEgkdtN6lPq5+97GoBhShdOge+NrKDV/A7cm6kGt0h
UT7y1vEechLO+Rl6N9S1mCKChPsyCJrrFWGeL9gtsZwg7qmoxwalbCDUI34R8kF6FFZv+6jHg9rW
Q3X9bSnwqv6lQJg0hQ46F7jAGBfrl1Pok6xpLuewymhKsIDItCAFm34BGunFTQoF02Zn90WZ1mTU
23RVbcCz/Z3PeI+9HUZxLZfQdRrufKl9Zxa9wXT+aY1N9nsVJgPXQSB0EQzbfOBvgWKA0EOmTc+H
yqVi18GQSWPlp8KCCLGLSlKV4lWK6Do9xl5O9rEl0+izO+86Qn/6b75Wj120ZFuukIF5fcWCYess
ShXR+6zKFxP51KHdQCNtgiQhVqjP6c+Ni1q9p4tbo881O6a1bqH+JwcGDUC3N1Mll1I3erRbdaVm
qJ7DI/4gftQCFBM+COKEHtANVkfkrhshd6fP8j8FHPH56G+OuseSbshqRo6+dY74UeiwA1JC/LeP
kpQFNLS7lqqOXLoEpSVNih789rv8KBfgGoXt9s2ixZ98QrWSYDNZUS5mVYu0O+Uk20TGoNY0s7ku
oiilKz8CVcvuTvkT4w3Za5ddf0sOvJofpn7GNq28gkxtOlAO6KClHtcGEhcg8eh7QLFSf/Nt/B/Q
fYeE7KRYGA3ucgFkDaLZjUu4yKVDhsbD0C/hrFUAwGfD2ve9eoh4DPAiNA+zhi89JotRFdE2aPh8
wxkFyUqmRwn0LAY/GjAxaq0HFasz4RA9ecWr33HK6GgkWMJKuwRrpxh3kGx4rWNwUrZxI8hCMWOr
KxSDikuoT58qa2YOdW1ISMLislJmyYaDViFb3ZjN6G/Mw+Mf3bxfz2ud+LFZJB5EfSYtIn4Iw95n
JrOOJiWOIDhYen9uFn4u398fTkenIcnFF5l8oYHHBDq4siIfHBr1f/tcE/bmZk+862M530evJf2m
joVsS+LNjNkEadj6tQ4/PeZtT2ENXSzgFEC814aDKeAOSVMlWn9Yo4ViYQ6JNEFTD9n87mnD7WLF
lDo+TNDuWx/qq/yNmF09n30mI9LHZQJ7IYjMxyVB2ux9wKv+BjfBhh8V3ZrSzQDJYvTKLvxUhvsk
fYYhJnkC6MysdHaG9TRmqOUjI7l3UoZPXQVtZMVhIKO+56Qr+zBGbAWHHChNianl1ZfNkj2k561G
7Vw1WtCHxuInbWbvi/KPa4L9vDubM3NXNRXRB06iEhPwrS7M6G76lisY2CQz0r3QPshuZz7v3mo5
kLvDFlUHqykyuPim9gCOi7ScppExHwm4YxgULer9aA8Y0cFuXrdaerQPOOQ9TumgT4cax/X3SjT0
4UZ1r5scUfZARPoy3zeMkvnUxZXrtH0999pvGgd+BhIEhwOgUSKEOZuwlwCsp8GsnkDvg6fVLp9w
zKaq0hfC+rKGjYO4pAtFeA0DINk6M+eAb8KH302fdte7Ut8jyog3gAJcY7bf+jEHcq/Ff5hG7Fsj
mqpXlHid11Wo27667VBZ31QOSMiN50ZIYAxbHPu4HUe5+MO0l0muUtEFGy76hMqvdIPFJkj6J9Zi
4NwQRQ1gr+zwwLkFh6EXKf+gwARFm0XfpamfQMk/jDdwst9vNj1f77PNi2HRvS+cCsn5P6hgK4Mc
uzUsKkaANEKB/cEA9/BnYVN5XB38DLo7dKZCEYBilEXJzl1B4RH7BZiHXRZ/BgUGnxQXqZiyICBX
QVIbNYl20s+R9xdOfIHMGVRkUghQCvi0Dq8alpKltX4oP6kiojwbtK9YsL7AkP811GKYmVoSMPPk
JU3qexlRbwYFRXE5vOeZaRC86bs0svw2z2hutFuNm1hJa93AvN5p/j1UndosyvYojcnrxsPgfA0u
8YQVOyWcLLS6O06roKQGMUES+XPdY/D6GoNr+yemoPoLTCd5zIFvYKils80B7tGeDB7rM9vlGqkm
gAaDnvteiIvsSTKi84slX+eNdywUmvczWCPIKKJGlZiKjGOqulVCiFC5Fl/RTfWYun+Y+qPninmt
jRUqVAnZBAD213Xd94TZLP5AFfw4yv8eTnrYyIzjF9yxekfeiyB8zrozm0Wz/q0rda86NbqN0hOL
azQ4dtpN8d5gtfC+wdCDizjxQ4nf8AyKnz1nI58Cpyrh4kwZIGlirgGVnPH9lXeIVE+EVtgc4gJi
zlsO2Vb/T66oAShpDI8Lf972SwtT4V0KM/Ji7El/eEaPObWV2EQb6Iz5Jqcw5Q+7mMSyiWvfA1kP
Bswp4kSvmwheXPX4KwXWdP2ub3aRQfn1qqpEXPtCyHazTCdLaaY5QSQTPNVns01ujRnTk7VQTQ82
DP/Bh1x+fye4QdztsWZrNWxjBylpO0sRvm+sWTI2b8bSsHPrOFrcFzW3TfgOR6/hPpGGfO0f23Mt
mdEOLRqgnvMiByLegf57ftRGtasTQdFzEm7JiROiP+f77pa3LFMGc++jrVGXU4Z/LcckRRM8FkGl
IvXWhK8ePu35FKWrWv4Y6eANYnD6BPasQofe9KkuRfqySvCv/V8a2J2eAQ2NmL68BZKzAf9gjCDI
g2WhbBLD/V6qnzuN0ogms3I8NngZiL6t3yVoICBu0HUdSFtOor4g5YGnvqZh7m12Lce27sRWqwra
SbuzMmIcYFCw/LKVzm6COrw6v7qgNNUDcC3UR3+FeO/CMHDjMYfw6TvloQVZmZx/EnqcfjY/My5A
zHjkM6WMH4YpH9or90VmRLQJmMjsmAxX3zA7f3yVeakVwo7/k7W+JI6AaL51Q2fqn8JgqUma/9Db
bUIB247TQ5fTSP0a9xxwvaEPNOMJLgY4RJ66JFvfneceFOvZVcgUvZm2bqeb/5VqZxHIuxqBLRFb
hs/Yar/5v0JG2ip4g7+7ha6oGOjUb3fQymyKRc4IDU03NbP7d0OZP4pTKhEXA/tS0etkW2XySHOQ
dKp2ab+M72n43QsBk3oSUJwYdGGB5V82KylZ+o+xxD/Xpw0r+IrRN1lkWbHuUx5YwsikK7A7v5iL
eet33Li7Uz/0jkxKAYxMnNaxNyhUHJpm+wHic/YQye2maToT0n3eEOEhy5IUsQJ3q8pTWYiwxf3Q
cu0KBuuMKDlbo07Vc5tAyl63XWKfylw1B5ZmGhuH/8KVT/FkiHeeSsg8Wk5WoUERrVSj+wJLd/jK
XfKY0voATW31wCUb/+MMwbYcIxIAPejB/BlFNItodK/EOcQBdNhuwQE28pua5htujt9ur3Yb75JA
IqJkD10OVwfTkwK58o2IuRfEcy2pz29qq66k+SiFW1HGQcFdgqEyGNzU5ELeKMb6mRiPUB7f8xb1
p66mpAu0ey4yCs6DfPvVcOIzk8SdLuMDiXUM5p6Zf92nI10wjxKmcI9wZVrFD0BnRo4EEE5Nr5K6
sFmzBnUETkiS8PCeODnFmKRKJzPYSr1pqWaNtwLuuTj8hMuv8I1y4CUDFOwaJqIEuJeqIyUEuC4o
5yU2d+LDJL/3Rj+tFCoGkJfL6RJeUEIFU4Qri17M/FE7Ye+HNXrAlbNFeA3/lOkSGnD5htIaLfVs
THKU8G8iKarEvhP9d0x+YTmpN12yiufFT+pQMpUiFl9XgIvvS6c0NH0G/bwmfjPmpYeLFYTAz6Sj
WHDqWYXNn8lO325X8Bn4aa/0QZTwnKu0wDC00diKEekA05UdJflPVEZN1FDEFQ1qKUfVFvLKogEj
Qs7gyeOfAVfhkwgzwWTQ9VkCP6P2wMOFcAjZ5bf79K2oIsIXTac7ioBUf5hFgcU4CMDC+g39yJRP
H0/OLRzo1DJiKcvaLWwKWT1EH+jhw/U4z/b+2kR1QhM3aG0xRz5Nre415QMNDIJ1pRzG4PxuSQiP
KO7KjcR20wyhs4nO8l2lhGGWpB3HtX8ANX2Si2oM+olM9Y0jXPmUluXHTVEKVTP3B0yU120P8uEy
q+haGl/PQ2WjPRQ2xcrX6pOyNroB8PcTcvrtoiBYtOkBwtGOZJaErhHk3jvr2KJF+7O9r4KgiWNt
4ROrmglHZJ8Z7WGoiFiLfQJNgwcyGg8R0o75gBwt4wmYKGO/Mj7RKEu+Nz61aOFg05iHnLg1NKSx
ZQhqxzvxuYkCOpjTW2r999yRYFdq5etH+H+45VFcPh9CUxtgvnET2VrDQwkRaTBBkt0tQ8FIuLwJ
XyQ++FAlZiSJuFgcKgH528POxSlFlWu8S6hI1djSbA+rmj7V8IogZt9cM2LBr22ynrPNr0aCp0Ek
hMiK4/YoMeAdYLRpEfJWw+df3O9mifctyHLp32ShttK7oeN9xtQumYGpe8UiCt41bH11KU8ZGuDv
9Q1Gfcf6FCnPf/jZZUcA4QWmp2CwP7HWQDXC/aE9b5FaWHzbA1juXD2AudIM9htH5apIuL83AE34
BGghY08iAp00Cgqg8dl9vTf7zDICtdMJxaR07H+gwhgMulWpQnVjr7Su2PrSSqks4WcVGu7CCDw/
QTbb3enUvEHTtwBIj/MC7LdPh68KnfJ27e/vKF0E5CkAjFkTjEou/4HKEd5LVTlJGrloxv3lVF1z
hntzCbQjuVJSHbujTyjg+NLlNARiHgr9cBLJzyPdMUgZIvJdgCC5E7IVDVWrty7mt3sSndWqgjkB
3c+UmUZk+3ZpLC23HxL0/yl6dW+u1w5KYMmpA9B6y+SEqMjD6CP4iPD77n5ak1VIBEHHWv1denlE
w+9ivY18PTfVR2QgNMIfeg/wQli7seLXnUOnMQZCBJJI+VjX+5Oj81p+GJNVzTo5+aK9XQyRjRzr
fP3pvYumUZqOPwzKUFsnDvFZQQDnM/zhGhiukNkj6FTuKvCBK8VNBnsfN4fnY2RdqsAFMUhqd9Ew
NTeuYoBSVISmB9OitGCm71PZuRnXm0rAl07MVwQ1AwBvkFYbS9Gjbfa9HXDi5E2y0J2993Ee6A0K
RN8QEocYKTeo2/xmnmZLp5tyH5rhIApJqofBSYxWTAUGeOLVkj4blbgQSxoWGKv0bUkn71taBdgm
9sVatdQwKNiVbElF274uRfCF4mfR0skkW75sVVQDyX9sBoAGNQZMUIx6Dl4/T8nOxh5Izd1tRecE
sPpvKuZkhc+7rbv++86x2ZzYIeM843KONs4Pv3GnIiLdoMzwiWW7NImwMKwQ4Ue1cpG3GZB6nRkq
FviAAq4g8YkALq/W1DAsBO+iYa3gMTgawcaBtUo/k1Yk22uxAoR6SIenPhKnDELlf/MtFLmonpI7
IAclsGkdau0pMBgbRQwIZTm/EDpbMcjJOQN59m6KZ4JdFzC7eeVpIzpk0bPkBYay5lX2n0hoAp4A
KVI9NcwapGmdrmQz6xttdwXVWVky3EcryNYrDpru7/3VKdo6JUcyUFyzgwNpTRuyDV8FDAzepI5K
kCE3KPHl66IIzUVP+i0m32zGeD2+OI4HoPupky8zebduIdH2RGgGwhNarjhRikx3BXM6pAUpvVAa
j5h1+DvVuXTHCDFWLRZO8jrXl/eJHneT9MMXgJXkKHhQA2Qel0soigPyKQJMsNeBtlL6OEltfpYO
N4LHV9ZqNjoIGIuzIzklJ4RtUXuze5HsSAdvR7fJ+BzM6+ekX09ddCYequRqQxkQDiCmXnMr1Zyj
QPYEhO5fRk8QIfV6uiTlRiKXoJPvvXT0NjRXeqDN3i+OCh/NKtuOPzMdpBpNCH6FUB1g2QLJFM+K
58MBxYL7PixLlcEfU1cp8c3XbE9zspzo8TZ3yicmVCAYtVYUTnAaMU33ElyFx59WUdcOhSf00tvS
V2DukexiilpT7F5TWVyqJTBSHjkQ8KCZjSfnjHCTmqC4C8FCUbckGHKB53nxhaXzf8FO9vTTaU5+
wmC4CBc9TKgmS6TW2RbHqtjipK4MmcDFnJmIxZHmDdEZ+jyxHEV0nUZzwB7R2vvYRIboSs5aIWCb
iu5ERuGoDubBNFy2tN7NsGujULunTBmod/DxcZSk7TfEw6XZF24kSLoi6veQjoaOecCzL5qwSV+s
h9Ess3jKv/1qHLV8cqA9xVwTVzC6AJF5LWxX59cn8TVuib1wCb1wdlG+TI2Cq0AXV4psZAbYW/MY
ih/2hvJVjKNvA+6ttmmYPxxfvkf91XhvYSm+Rrhgu7h5ShxPsC11owXPKB9XTkky+TREN/IMCjam
J3VSX1KPqUhPOFXCDCmIGuSR3BMyzlerp5shzORxrvqHAHVn5xjC6lqN66XzmlluXJlS6YJRimP6
ogBv2arFkYvDcnvrV0GzuVdGb+u2PkRyRrteRhxCyW4i9Wefv2oAoNeQ0xp56+ysNZfCjDUVC8Z+
9qoXVMwp+tHafoyp7ukyZQbUavclDUvZaGUHr9FzhCXGTH1x0mx48a3xVE9SGBy7sYN9lxQTl1Ex
QQWXoKji640PRVv8ztAlCtIcibnCBTW4AXZQFpvvK3F5ILSnRJFLjgGw1JDfs1Pz0nTVmqkrqH8Q
iBIBppqg5Ik1V19MZ3FShs25ijxNn2OuyHFDO0vwRuLdcBujmJrCDHMRpc53cvC05pBq91GxYSCj
SlQbgknXzk2k81qNal4/jVPrA0kCEDTuURLZWYclr7rSlKzzQSAD5wyiECikhPFdUTgugqbm6EUe
BsRPQsOmWa1lbFliRZafZXZNc0dAr9t3i8nIntyx+jpYCtN263ftZnN3MAzPbB/+fwU7MsIQvh7L
sWhp0v+oIWYDURbsSVIWTMeoH0Qz2Z6LVie9RUChD76BnNm5CYS/BuLk0MMqZsUpN67UqZ3Kd5Dc
Kh+BUbccCeSGEoMJkGK90XRNfkNz/JLhiS6mnH506iRpTN+vtJkI/+JT/az03I20M1yEXlLPJUAO
UYtx+tkXUv8+AdAhLiRrH2IlYvPdib41uWatvijqcYyH5qZHrDpDhhw9ubZwfmOgdPwJPIc9BYv9
7OSTdQu/q7AFu+yHJvpYn55omK4euz8l2P30Tb44tgcRjlNfzgFjLnFQwGlPWM5mTl0YonSt4hbV
EiKeBgENhUwA6oOiU/1E7hqC+oinnjujQjPoeA4gSWJciaVD/h5EKEXGMVl17uXNFAYK1vBNdtAl
p1Fkc4WSXIv/R+hRI27NaeNGQbrqb69clRK7AnqG/ZLIczZ7ASHVSfIyLWcDU5Wft4aZuGWkUkWx
+vc2e6aM6NLz7LR9/VOYyvQg1Z3BUVvmkBWxjPbCG2GE1jtupkccA8gEA7dKJJB+V5utzDCOIzLb
KLbZluPIJQ5AujNiDrxRTlt5+oxCGZx3S/dXbq/p9MNG8rw4ZU1eoSehQXn5Gw6Ak2c5LFksxJFM
1+A9C/ItY8IHdNLcZy5kHKtA1hZLxGWuUhV3n42i8W1a66Xl/muffpifhOPJiaSLynIP61TewzHL
4Siae+ZxPV584t+Nor2w9xHil/S6ACU6H9qrX13P2g6F2iQffUmPnNDRooHBrhdPxVq6aCK2rOv6
FRbZ8GM9kYv0oMikrthHwN8ClfKeOCgXnrpuDw5w0BwHuQfJycHVwXaHhmo6dsKMpExjVjwpF5aX
QqE7QDXve2LBrFJJmaZHhWO8DJ9OLkI51Uro2E7gWYuS7P1sulplmwCIJKbAmVpyrqDF4G6da7cv
jFdmzhnFafzXAZZqecoMJDaPkTluvVW3M4rir4HBAvf6vyHczQNZu1aHRovGLzIHtT6evxH4P63m
l3nNBBYp/4WejUlw11KcCfa4bJ9XWQmit/8JMcq86Xj1wayszkM75OuJ2F1p5Gywst3jfWZCsLiS
yjJ7v8lAV7/uppmNa3/oFxYkPEiQ7VTZaaaUBHychgtxHu+pfBJa+d6ONsJQkq7hfTroLQjQlmhv
RSQzLMMmrHG67PMP0cNu8KnRmBNfUKLeSWINUP8wxGbTrTL4WtkM0rRpzx2mg9lyYWDey0hqedT4
3hFZdvCzLPiErqcYmsuI7EJPDt3WV4chQ5KM12wgIwplwxgt+PzlKnQpbGWB1mpoRkAKVlRjOz4N
4Uwgf6WUNeXHqbBdv5L42RWFnPmUEGzqYq0SzaM7N+tuRllZDl/2edsL57gkgbbW5JJN/lmyfjfz
iysmbRPlQY+Oy5GUKfVR07iSBK6A5D/Xrc3SqWxcbeyle52XwKSSYh7kQZDHqQ4T0N2NgnQhZsS6
ux3unvO/H2Im1+wX2Yboz4p9N7veaCfrcXM6ilKwGiw93Xmfuu6HgCWvBnY/Ia75wZHDGp4wbZgK
7dZdPwpqtOVMgMtiUf2X825ShuBRUdb4rd0E6wG2GmbmE9sGET0pdAZd6kgqTKUJTLSTSDJJEQVC
o8S8R2Qlrh3R2/j0MG4jjWAXI7FCELaE5FoqridJ7XnIxlcs/0/Ys9QlrFPR5+BYQhP2lT/C3MZ9
Di97MKxos/A1zCbpgGXF/kxRTOKRwfSOGW/yd2bQFCTq83taczvrFx4VuQWl+YWMzeiSdVShy/9x
8eoWKFsuXIG5ZRy8E3wBrueK8gCebYOQexFwZVl4L8n+IBDLt3tqy1Ud2gQAbUmzlpLdr2Y0z3RA
rrohBZ5UmzMNPVCUAooOoSPDhUjj6dDI5656HPY0s7fBqmJSVKi6AighlMM+33XLmMD9SIA8dria
y4C/+9ns6X2rboH7rvfNDxA5UdPvuXIj26NxbsN1ofi+zbvDgSdM0WY2IarQieNaVnb41zI5F36y
kaisMeT6+qMK9jNEdfVFxs4iAMxPMRqwOX5LJNXaP6/jhT7Wh3+AbnTA3qdfDo7bRmTXGU5P0SPB
cguQY5ztyQDRvXhDnChlV5b8z8+xCafkq2sguM/Gu+OqRcS74iG2KFxD9ek7PPN9TKIVLytI0Khx
Xy5INHhffbVsjh6K8vyFZSGjEhfcx4Qo21Vzp15F1B6b1qBR84zIMF52n/Ndd2yK11bLFlMC2xSd
8MIAxc7fMLyyIvYYgN8jFCAXoFV3Um4qu+lLOPXfd8UFbzkTrsm6LBXtOGU50Nu313P//JOi+Wkp
8reTRA62LykkRXFomtjSSmLOXQ87/TL4o05sivd0BqiZfVH40ePSYoLDrcYPU/IuKh4WmG/f/skq
AKdMK4MX4DvvDb/fssfDvLLf/qPWH+0kschHok3ziEQTvNOX7yIqPckVEQkE/HOXb70HGOr1Db+w
yW4E80vIFr/waEhYF3+7APmO586xk+cawJ1GV2cMuHOs6Lq0w3EmxR4U/CMqiAHN2DwyYdNems1A
Gp5Iq3bkaulFNMG5iMFQ9ChwRqMDdd74I/cch1w2iEUzE1dpbfV0r2/cN16stYem/C4Ot5sJLHjp
k7hwVFmW6gpdA/6SbreHvHky1OiRUXtwufzrHdWP71ThZntc57022asRR1//Q00/jfFUTw5BSDgs
pOr8/AZCsW7VS2pVrKoOfq8hANk7cDLqfk7r8wqcHkqDUVDiaDr7x/qQ1xTPdn4wMrXzN88NCkvR
wmYs85gjjl/688jgyFWwHMPH5F3Z5iin0IYocQcj7VYagYpP8koWs4kbHPlqQaVQLeRQz0gMPU7o
nJdS/eqPiIkDaolMev/ELv0ji09J/wadB29Xx67S0/LxDgBU8BRFfDZpD2TSUc3+yqajVl9N1mhF
lQjkAnWXoYSFfX2bhJj8BHXDwomAnGL7znHyyTEcEjji0t/W2FDOw0V33hsLQULuaCC7jtViGm4v
fN9SD4/cUT4NKMj4jpd6rai0b0B5BwUsy+gBuDe+mCwzdco9Xf7/yOBpdd8M+/SfxY+zY8PtY2a5
7tziHw8cHZZ4hMj5Os9VDTMSu0G8ceiw7i7lG9xnMOJ2Hoh5fZDw4e1NoLgZIYpisD9CubK/2bCr
o4xamk7aEL9b6ad2iGkfKrn7dqzD5r2d/E6LQniPnYdiaSeKPvY6Y750VAHksamDiDk6L+DIQZUf
GfP+/XOfoo+2zla6iS3e88CW/BJ5tRgU5TW+bo5yrhoAnhogGGiVNSBVM1mQRA4IxYHfuxz8Tg8Y
aq9UdmKQ4u+wVyMMxdvkI6idlu0DOulAJHe6BMbWSdJ62LrOrxXJ0QoT9DnM8EIWQK0sqvBYICvm
pgn2o0O0nM0fR4sHGWmt0Q7uup6/2mRku1sFLMnjifet3axbasM3jmNaosH15HhPh/WjgyQl/rH+
PlQ7bqEgG4f+/ZQDYx7Ro4UjNDgDucWE/PKN3u97DBa6MarGU/dVpq+3ikpSveCaBGjz3VmmZbyw
m+FeMQaoGlGN4Ujbzl+kifKcrXIBzbV41yClEv4gnEBruDAmb+ZfCCsbNIGguug/biHktQYQB9Eb
f5aXSks7lP0QVfP9ZJ1vI6/4JJ/s11CnXR7yN2BebcOh47E3nmuzNlcAU6Xt9pdSho1g+3/vVXYT
/zbpwI1pam7rDk7hFkMpYdRPwE+sOvXzI8E3tRsRj9+9TuuPlZH79mhkow7AZCNY19nrwXfXsRrN
lYTOhc2YiThkdBG5/mu+ngzdqo9OgTlU0U3U9gCBt4KWhlE0t40K/3XbBD5n5/Bsdq6oFzuggY6C
v4T16GSOEvUJtnk0MfHKZQShDFW3Q4VbHvgx/sZkTszD/7SbY7IgyxLusHKywrCPJuLTFzYv3r15
XADbsSGZ2IIbVUj2nGscVSYmmsyooM25PTNQCsGT6wnJTZ9wMT3/MJ9U95PdSq2ClnBn9ZLg4WtX
9XcFTlBA9SD7201EJACAFsW+MZwSDMKlInU98c9Tfw4Akhth8ye+mV2+7Ic79vCAzBVDIBcgznKG
b4+qBWm/uy+3zxsfCFtHqZZPanJKAgdkhzaa2ThGG7em6ntUUDWWIKlENyJrdijntVSthHr7oZiJ
ym7RJHFh/ebFxni7+W8Mrr+6EJvBywUXlhe/j1Pgz4rqzLTaVU2WWgDLBwM8pmo7JqJHacBuiWlw
wEJvKEyaU8foImMzQyukJXqke+Hswu0qdanSsiCF8unrbVkomccHEY3ZJWfFUqnTFGKJyPZiWnXm
v/CjTaY+lUfUpTBmvW/RJpI5bVWyTmhPomLQOGd9FxzDZhRm/2VlAu5Vf2ni5DTuS3GIja64MJD2
S6awZkJDz4LzdHyjW+Eir6mK4JzQQX53CkaO/Odc1vutY9k6mLCo32/859sbBiCsV1t1/eaKpWJR
m25tudgkYAVC3u/LBCPcGxsn0JrqJuOVVXbq7p7nltbyAhq9xEANQUPreIEr5ByK13o908A+imTo
iwlp8uZRlvPC8H3I6fQrz96EP0YZHb9Fr265uDFTJrUoTslampB+7OpflGJ65L+tX8/zu3xxVDEB
2i2Pk17hDlnICTMqltU1N12f9kD+SdnBW+ol7JnpMGC6uW+Dw5AdOckpZk5Co+06PIuWDU2lyuS/
eEsoJNncsxNfA2GdoyPV4zsx79yjrfh/OXHQv5CAyPRL5kS4pMulGcb56ms1o5TZuVSpB9CtDJIT
/xMZXTzeBtnL88eg1eIqrCHBqlN1RNZO3SXJcNrvXbC913eCcQgv2RasEvGW6ICCEY6Hx/zRAK2U
bYLNuK+IAtAcmlgwtrJ70Lc5sWzcfxMLOR99Kjh9N+s6FUWblB4nW7IQ/7P+t/Do+23S7bilGl5J
UvzrWZgg3OkbkgRzJFZdXMTTXbyZiESFpfiXYwwDvscSz2ZaS1Ub9l2GouPpy5KUCTgjc7w+Sxcw
S8tlq3fP/XGWpXN2UUk+XaxAnIn1jhgn3EUWjutoO4G300wYNZlZo+8K9USaNAHSDpvsMT74GNoW
iIo/0XV2wXybbeNTFofTndpxbKy/PFcbntIq/xESx2xdrNqYFCPuN40ypC6RYb9WsvMWSENeclZb
ZO516DEf0LK19ckdHKyZD0vg7hSLGRxrbzr99o4/3sh5ICOkEggcY+i6DbNkWfblMJDBow1IWeY+
aOF3NaXIhQ+4fIZdTpK2JJs/fmxidM4degRIunn9Bo+/kspbZnaYmcm/FQ4uMjoDq6ocb6ISBjnc
paBahHf9Vm28Pj1GbFIWf/J4FRdVRtF1tz8Eull0vGI1hwC0Okj3do6YTSZTF1URB+5OXz4+LpDM
kS/DKjIeVQwp93NQKF1I3KHQkfz/K9TEVWoYjf+sPdQFCNjpJyevoTckhbYQPDogDhWkTztlgyjl
Uba+yOZ4ZR/R1odt1CbftjlZTe+B0UG6IkH/+X7o5K5ut3zse9LNtqzCaw17EJ6ki0OtAF1T9JI4
FDWEx1Lbwd9hGJpSEXjPNfHqHbAqwADLrOvuSSzGaq5WQg7SNlRr5H8nPAiapgxLbtmW+NT8ybY+
eLsOSDyWM3ClTxB1zao94YI9pqhrSUV03aDqyKT/iBXB8OJ7A5vxvzICGl6UT1O+QvX2iz+hjOom
eze4/Clye+FoY+6WOib6qxUTJ2LPKzILYm2ppkxvGT1Es4tVHonQt/dJSd3VSB5TaSM50Pr3Su2C
cMml4BKqD3SN/Wd95rV/YRiynZbEyivqs7zdKbHcahE2mtXEAom3AOnBd5uqvJ1tOfAtmliMO4Ol
vv7fcJCraQMwqEuc3lOQoduJenDoGmyWgpKMvaNBiOk+iakgn3ikH2MnsR80QIdp5uRb81OMes7u
fDk0SbX90U1Z2JZmm4/TQqFo7M+q/IGQkyInZpe9MHR/fcaccTAucBbuHSGrO77MXzJbYspPj3Xd
QjAb1Zgd45NvhCieCzFLx8z3rQybkT5nAIJFo5jTOEe3XtLlQK5LlWsnlzQX14J1FE0L1A6p8pFY
D0AL7rKjwd782OtxbUa7dGJf0nMQ3GtAenUA1yYndUz5immgEd5VNSDh1CXFzpZXlNpyh66xnqau
muT/LlYxfohd/xx4hNlB6iDCiZksiC+LeBFK56MBFf+zqNjZpsZGdCK2sV7/iEXsZSm28hznrkrE
7XXvCSEyFEm9dxvJbDi2v7aqH1+wuj12SUdkOSm0Y7kd1A5PfmIsfeZoNrEjY037bb3QuOMWlO/D
DrWi3/6mWbFOKPh01iB7gvc26g8W1TT5cSWgEKfckodbgizdRXI7GIUE2YIngUU8KGgrX+qN5POj
JSh46DFQdzjAwjezoBeBKDjlDvofIyAieIwsYpRbGhxNlv0ajNWTMI9jAxf7+Pch7l5YXaTnWjUY
22wRZtEzR8hbRqq6x9qZzKAbqwyqZoz7ZazEaKy2Qd/hCxNIGW7SVYlWlXDJdZqb8MBPxbd+hKlA
kUxvYbtz96rA5SonDP97FdcNTF9GB3iyAbOwPYj3j/kFbri2z5uMJzNrl8iMEQcHAEk00epmvnwl
OG4Fj013k/6DCy0YBBQoWYg6+7yBXs5bfl0UaMOyap0K4DJu/XwXo1x6HMV/aNZI9ZBpD0Hbs541
TJHPLqFvZFy7i4KPBr/kSynny0pclc0TujK55Hu8nsRETKQR+3z9oZcyZZ1OWPsLBQg46JKP0Cq3
nmQBvWRg4dEqCSoMN0kIVbVQMQVD9STs8J2hDhhWNw6z35oRkBYdf/agMwl9A6C4wUXX1qlpFscF
BRYBf8N/EwrK2qfpwNHnwQZtuOeEFuketuXA325pf/rzzY60tVNo9m+qhBSRHPCpb4n3GQx+rq58
d4M/BiUQIKqKSRIsMxd+MH/AmQ+7OpPZor6hJrxs8f3+J2g31FcX79+05JrRnR2ET4znhmDuBZma
+oj8bLuxGiW8EwGccFEDvCpkirSZykyzsX6h6oYCYC1IvQCAVNpdWGdxczfiaaIgXri/Qb1WJH/f
JJQNAGed1YH55T8H6+ieevFNjb2qZ83+K7lUP90d5ruQwUf9wkKV0gq2xVU/+hP+hfOEojVFiMcO
g/uCrVwjP4QGev+l6JNvqEJdxVfWgK7nDeEu89IqgyeAi/MNK9ABo+mdSH83fIYfchIN7HxdQDuJ
gtaUK1c/FwmKMJWOAfZ0QCPyd6Pb1ktXMTFiJ4wzQTl6t9Tsdg/oHXZdlHeIgj/34OFAXpWLewgW
IvkaSJHj9p4Sm1NAvgfqC/RKOtzOMmzjtTQfajFDiqDr6Obx3VZ+2LCNVJZIPdewcXvWJdq65yu3
f9nC6Iuhwnba/U9o2RkL3zQwh8QQtxSAKgw+/15oWf5xqhEF8OyW5LwTMjxkaJUiGCs0S6j+mPnY
+7513YELMKyJydr+2VuNeZz/bngH6skMtQ3u5DFvPg2EOVY61aesafsNYzC6yycsU0KvosKybW+V
s/O5p2y7dSO9rur19W+XgX0w5zyScuV2B/c0ejB0XcsOpXu605ETv6GN8hAoGgh4oiE0kMB1wp/Z
tPtEQO7s/6VSPXZQpNSUleRRkz5lV3U4mR0j1wxftGe8jrdAHSgbb9RkoDbUA9JHkOHMu0GGPFiO
kzueZaSROL43cXqnSYSHXJ3YpnW8KUnHJKhnxijtquJfAHdXrBIT4ud85Dlbcgls0iwn38k3pOlT
Wi0wJ3RG/cbwjV2Y5r/6l2gPjU+bHPeM4MerfUe0sSjCpPJQ0xb1p7t+qCmZ145rhLCeKus5OpMz
Cz5TTPUQt6aVmk+/3EiY3JScAI88MJCuxHe/peYSshCxtThlVLx9PGC60xACDwxpxuIYIJDXJrL2
2Zalt5/bWD7ad8tX0tcJKUBsCv3NJzUST5/UXDVBai92KxJRe+u3djfL+fjdLUYsluXE4p02ddwK
3TCi4XvGSjUCw/XRQWkNB7bBOr+Apnl37FyCj5wWAAI5l6rznd8OUB8mjnouJhQd5N4VlKkv3wRl
LW+++9EQ7Taeok2XzdrIU6S+tsEEySL0zT3o+W4wiJlq7yM6WRFPtqsoThILFkYAQ7h9S5fuDoBT
VKk7mf7skHZmQjFsU296MFI2kmokBVCWyXrB89IDUy4T4PpONOx9zOYkHU+fm+n8kkS2IXZKI0m9
xZZe4X7nyjWKzIYI6n+PHPEvT6mXZP6YmTrdj9B01F9QAUMyAHU/nW+Ue6AP5fEa7Zz/U1QZW36U
0AcPqsu7dS+bLPwnCTeptL3+1iNlfIBzfLt0vIAAHnMoPielUGFi2UyoySUnTL7W8IaW5qZELHPV
EOgW76t4YzlxgW4nVENWrgOYulWyrSFz4we7ilEogf0hMYodNH7ZHdCJBEKQ39d5FtAxbkI/FY/v
yWs4gZVHPsw08pgUnV0/aCGfuff6a5o/reVwkfL15jXuvwWVSta154SWJzUG/Bb9bU5TAw9OTp9J
aCQqZn5RQROoAZwin5VziLDZM/HcJLWLXdbSpfylBpR4qs6HNYyddeRiKbQ36FU2dTp1zG+qMN/u
PNEAH0XP43NkZFJuiRcx50V6XC4GroFZ2NsYTFFZpfV04Q9gCBL6gihYBxgitzeuZLNEuA+SA1xH
mwdsUta24fPWNagjduh3We3Qvxjvzg7u0C2D19LctBhPZHSzhV+ixB32qPKpwsC3zkCX9hdY/T9t
K4fL6obbpFsVvYN+1mKUZEjM6CS/FutnrCdh7D9LnRNGK9AfSKpAoCFxjEUDgdEuW7IqU6DlV28l
K5lvLisj0e0BMgRgXDSiAaiejP/7yqr2ZSlS5KKjRjrW6HjD5SXERlHYsxPliT+p1uia78Ikt4JW
wb2AT+dMoC+Y5PLnZIKL90XQqm24hHWsNcntsuDLjPQ8Vp5TlimgCoWGjY6LX6nVfWlXs9zQMuH+
VNw3urRACnI5HaUa277H3crIFHCKmwxQt9AElDy2MS0IEA7bt/pf0yj9zx360LJJQleYJsV3U17O
XVG5xEegkNH8muYjI3Sx89tG2wdpPLQprt+STn2k1WK22oW4nTj2vItSgVIjhMm7on5mDOgb3hA9
vq48anFK+kcguNN40sEP3gf9UFKyBXwsKYvpDb4BSdij4/q/oi79RK8KHeCJ1L7M/i369ippmaVc
hT4CCqWTFDmK2HeovmSOcksstx7A4PF++DbtkqGSmb6MDikytQL6ZsuK6oCMv/A8Or87jEAu6sw3
59Kc7+EhnoabjhuhQ+f8kVf0K5GxCOG0X2st++YPXw5jBwXfJGbO4BGnByuLwkCEdN2qvTWYbDPc
tNouA2GgTKt0/D2kA2416N+3OKtdCK9OWjtf4wLCUwbWsK8Xm0NwSkKhd4/hR43nuyAhT5bLqqih
xFovRYc5SniifNZxU0a4V3Towz6TwWmPgVEvYAgv+oiJvcExUTVO333OqcX+8WGLgcxduHCCzRJC
YwA65WGl/RlgYoEeSi6QvQoSi9X4uCEbOYqtZhnBZ3+TKTlxvmxgOLG2S4heF9Rw6/aFekj8DoR5
h1h7hOCY3Zz3Iq5iNSXmkpWINAd4JEigJTtpQz2U/w8kzTBXbbbnPQGy+jHi9kbR3XqwJxD4jfMx
xmBHtpYiJTMiNXt8U7/uVH+JQ++cBmacG1GU6cUD+kaAt131q/vSld0doKGBOwrsDEV8Y8DfkErT
ni3M0OceVpfRPuCpXx71NynPj8gRsJoyrQCxHJewulgoJNxk9JD3k8ZwZ93B6l+OlLI4NQkbTk2m
udctvyW4NoQttE+qnsUOERKyWrZ7Dkkg0SdHr2Bd+9Mqm07Orj9F+7jAiaPjCxLdfCDEBambIDvv
jO/uQPxzKLL2JXjQdE0HBUsTCMCB6dhTqjPUb4SVTFiV5FMn/z2IJDtRI/I4lzrRrcaURZAb5Z0X
oupDn9TWJsA/dIR8TSowqwOXRwossEXHuEyLZuoGTMb7xRsWpcjqWhyRCm32Nf4H3YxBBbjXcV0J
+5kTxNWmK5VIkF9D8Y4hdw1fyLitpBHPb91d0ay5r8DC4JW8QcoN7j9SlTGXJ7xNk1uw+sVEByGz
UlwJqlmDrRSt6KCRCnZh6P15IIumoPdYRX0bhOdIwBBKsZY1GGF2dE6c5gbaV9BP6YxAr5DER7a7
cbGEodUNzZl3RBSYO5n3EZcLVlnkHOMWudjmUu01xOjpN/VHBXk4aaicO9kCzbtiTmsjyyNnRdiu
2GfCqxMNxWY46NeO+r2YvyLiX0fuDS77vyUXSqfamGVMf8eaVC0pmeFS07EJGDer7W0tktJ5IGZN
A7KewJ1pN0gNg2TzoK8XijsHWiv7We1+G33VMAuxN3dDkhg55w/PhGJIFTpG6wd9WQB0AWkX6FQZ
7RZi114whUrzlu5XbR6IfkcL5bIaPQ29TmKzSMypUIBCt7HkojXVSALLmjAMMGlUHQdpHu07GTmv
MLeJZvgtbkAhHWIQEdFPNqoDI122XRfdeZvM/6HSeoOk/hJb764TtqXaPd9+tdz+crprmboYjxBF
nMcydcc1sXJOtAig+unRXEtU+mzxmh6L9Wf7fHuklCCBN5m+g5m4ubvVjssxCkGohWBiI0LxHC2t
SgTQAtgn+vuxbXz85cvv65kewrsr9qQsgLgc5ZKfpUK3zZ+8HQvU6VOv76rqD/ozTG54hhKpXy4d
dy99qcStNey2522xaW5HwHDaccRB7h/JruDQ78QwVCsCVRBG3iIwexrtCNejcu29QTjfyLZBG/uc
iOx6crh6hlzRp/a4YFpk0cNoUq6hlmiZxQ1+JYYG1K40F6j/UsQplDqZMAZ94kpv5nSZFqKenAg3
nq6W4Lw8FKTq73hYpYQJl3vEq1BcvEGGxpPbeiO9HAK1kEQ+uxO2wGEDelpU8rRjwUoyMF0s6jbq
rZjWppvdywv+wZJpkAdXpp61IAYLxalJpdILMwV8skhPJCq6ae7dISowiyj0Lg0ZnPLHw2FFk89r
/ORzAcAnzzsB5+pLd07kb2d7SNmKZOzFEpyZhF9TpElMmTYr9u3/ZVqHsxdymHqIOUSV8OZxfAn3
xFF4w16fYaD1r6cXQKaTEz0H9WQBJ97luVA9BWbB1SV8iotNqS+qjHG25SRh09/VNdCOSUgV35jx
MufO5bY9G2b1qE5ETj1DyryhD3KQC8KCHasvsjcI6zclj/SM1jZHUgipCEHvOgrYtCIIeBhK5KHU
4Nq3io7/ihp0AX5uBoPy2h0bYaOdf0xGPAlH6q6mMNpyCkqeD7hJ3Mpry33OCqbRVu9AaYEFKAdb
PEh+NHjDClN9Dgx3BRlKlMYvh9Y33eROE9silP8ygFuK1cHxBkQH5WVS3RFocXib7EQUNwMk6cv+
3anQv0s2Cd2yrrYGtpWnIuYKAhgwc6O3v+umFmuuSlvyOhub6SCtbm71CWSq9Vkgoo7ggOBTE3K1
PvW3oqKfqh0PqDond3OKN05KdBkh16ppJWzAhL8Q3nQvLmmRwCxnEUoZwNzsusxosqslKuyVDmjm
TwOYBy1JPnQNy08bjmNLw7T9JvEY2ibS1YSvj78mtbjJl5NXn40CKayetARjCmJaS8PHP8PcfGgu
HGNPE7gYHw+8J4RubL+PvOhwnTVLE73NHXZdpbXOXOUvJrUpd8LP7nleX1KmolQzihAkfEMNBePY
giL2BeoCK5bs81HcLhGtv0bfCq1xS7DRPLNA696huBZ9Lt7Xy6t5Jbqo50mUDoDMAE80ugiOciNT
NiUea2MD+XM1gkba8uI0MqH6el7fNxufzBmeFu2uOt+FqL8MT9tgaBRNRnDyZKzz8Jogqh/SPAni
cUneYnaVP6+h6zwPVykdIgBT1vQ0Tkpw/4BZWNHYzW392VHhXK9vILUdl6eVghjmV7eNUS3u6d2Q
rkYfkjeb0WkggEEjJdAOAYGLXVSXzsK70qqALbdzT2qu3EUKl25eWdUCGBqmwj26ILxIiZUFLcnA
qlXfipxcx2s2a0mf6g93AYbZO1eh02USEa46cQ19rfJNmVQOYAMPqjIt9yqCP88zIorOpNWdgCtU
m03LkJkrWgyjQTWohdu5Mkz0rXtgHAULjKPXaemyysBAuWdXGV8K2Z966HJRVWLByz02+CxQEHAY
wLoeqNjmYyQrOVLVkhkEZ/Un750VkNMhRmvt3AoOXZqs38hxmA3z/HgJgsWsV60zM++0+UJat1bA
3VT0tXOcEDe7O+XxFfeeKhIPTfZ0PgB1BG6IPWZ2GdQ3ochL5ph6u+ZZLXhserrP4VPJE8SDjYQ6
y2zWAsUUtCnMlNB1/ZYYFRGZvIzCle6Qxvw7IX2MQh3q36JfTnaF6CfCXlTV4SFOcPRHuFQ0NXaT
t4Zu0x+p9f/vWbAky99Yo4KaCZqsYFINV/Lezvm/0bCu6zadXdKcRM06p6SSy5bsEOgx65Q7liiT
GbaNJtbuw2m0FLfUSTcSiN3WrPFv/zAyBsFcX/IRLmAcp2Au6O05irYkmQDlan2vTB+hES16xDMr
zpawLzcpiLUaFEyRd54TYLxedpJ/dnlYuQjoguJSnbA4owA/BjHwZgfwvzEZ3SVMNxsWiuAEKIpA
hpn7WLgrxav/ZLOyFwfZCCsU0GaJuMcjddQHO1OVrLoyDYYg8UeI4GVCosMn5DVeU2xCdZ0TxqmE
yWHxLVhQf4HfKcJfKFbBpTMi1Vpw/SJy5WJ/VZTJLUHI9VkgyrclxgNY0jEevq0DbkHh62E2HQRv
RDTkhRCzZXKfm8FSY3MvTRX3PX5Q4HWUpisJ+CaHx5q3sVpzaYrneTmCmPQFUlC4A8wGTdUMEd8f
pEGuoPnR/zVQP9vIYmruWRA/bdYdwYS0a8WtRu3JNnTUtGy0fVaN3Ps03411mrZgXpMU649Z7kJT
dJ/RghT6qzdDbyFbiZqhMwDJUdUqc8prTN/1TEmhuHFRvQ8HsXKLuAm9ZGaX2ICi4uu5tTZ3pFB6
M67LPohvAJMB74yxITXTTvd/a6CV0kveMLx7oD8J9I7oul0mh8jCVuFyV12SnxMxUV39fUopvS1a
gpy+TFjSBIr+PJRzNtjkD3XUoyYGrU7yaFLcnFHm+SC4WHkCvEqFw4ssWnn4oBANeKGarX1X5hza
pXSNkMdra2UUJpN/2SxMRsxRGn5pQPrvyoGy2Stot8COnCr5AmyxgypLwVmzpCG+lN+BkogWtF8E
K6wIoqdRsZe3qUUhEmyz7OJpr92f9+EB6tIXk1Brrwe/FHBn2Dx6peZ31P3XFpTrd04VGvfMq6qs
rjiw5wIa1OOjuAVhYebh36ICiu6LY9k4u99ZUdlP0ML49iw6rDbhShgtcnj8JrVduT9L1WOt6Toy
Wxa+i4qgyuNvcibcUdoWKDtps30yqwE7ga5/gj/cWakb+CpwyEH7AnbULBNIB5obx36VRNfsBS0T
bYdGaS5lWFe5DDzjoCPy9Irg7d72tXKq1CiTFzb2JNmvS3OBr7f11NuZPD2oHwPdJGzCrTsu4Mar
HUH/Pd5E5pbfrjKsD5bfK+e81upw7lLqYznDXYsT7cEx7PpcEa9IwdO3d/7+O217x6QQvPUeOpkV
z0IC4lZamwyQVMgNi85WhMH2n7fQ2SAB0Y4KouyAI0VHqP7/omYYtg2TF/IBqUIMes52YZDfHZKJ
j6fqf8XthRRyTWMFnbwYZ/Qips34RqWWMFWlE7p25Iy1Gdh+1erkvYJOFDz+wTLhLuvHl1MNLfoK
nXmbRSGPDwQS1nmp+za22yeBvB4lDXhvIcw8rZZzqNHMhOdOU4xJzUaVGlEruW4ntAglvaCVwiSH
QPPXlgPirecjlMDY4+dg0j1PIMwrqT4U3OD2dL06Yxf8/15v0xM7c4ruecILiLmMAP0Zjl9cXTeR
MsK17lBKNhLzzgllxUI9kSVn8AV8d0jUfDXgX94KKweuw1Vm7O5qEi8CK4JNUXcujjNJDIX1l8g8
15e3N8nPSzWpHc8Q/wxHSgrU1ARuFkjcydKEpFf0PGU6nWHZGw4ohFjSgATICLzs733VQkt4G1Pf
m/SyKZJAzhKowgdUuuuLyL3ElDAKkE+LdGz2uBAKgFlwDtsCUmASr0Y3Yuqgok0eZL54J1wjrHFe
BhlZ2nN9vAh+XGlBYXom/ifoMhTE/nYpbuDtQb8ujZHUciYjHqcxKVWji9/Fojla3BilxyktSTwq
PTiZCD5b3FOupctBjUK8dgmdrudo4h3tH//+ESuE0CCGCRv94GMsH/jZBpKehO0AAyz7NthikdIs
PLjqgkr6d7bhFd/f4CTTkBBGh71T7FWW/yQmmXmNkH47s4ClzBu19TG209xBGI9AxnQR7himR6nR
jA6vwqrSV41zk14QTAMV9zSGCoDOeLEdnzQwSTsKpSYrNOOe4zEY8r+gNmdHLzdwpBizFOUkgFmt
sMspXOJDBxbJ7lZK9MWasmL/NORsHNhpt/VC0Io8r/0kb0eWqQjz5BI7QJY/kdj+Fdp8eu+C0cI3
x2OdZ9dql+9qGu10YUXv9SX8o291qmj1JhAoWp5W2HrpK3GfSMdWgu1w/XR8pflNGIWWDfE8SiBD
dg7G4cZ5Rud2Px7IWzTyce8h3IesuQ9MuzJ6TgdWqwSLqAFZjNqQgiMO6GSOuSTB3hU0yPOGGb3Q
4GAGgm9TnGA7vzN6aPPGLbVFCNKAm6y/ZjCSFJpP2D7TGAPu8nYdsWAlev8X9XGxlfLNilQfHhDr
MegaZswKyxymNuI17syTv5ggOcEFBY5/A8Ym5NE5bEa4xV8YPDFffMCfRCGMwnHqsmUykX9o5EqG
C6X6vbpXWRdyvsdNnpZd6LZIY2dUEflzM6PHfXyxzbdqcC1qJss7bznXbdZeKk0xmWrpAom9UmWX
JGssuwCf8dbse3mEjlqPuTIgxIa3fROv7+3Pdq8DIre4WYHsge5lz/2yy/w8nqm3B1T7gsym0kQM
abgpxy/7A7r5CWZ/Me5yrVb60AC37dLdXXvWQ8klolcqO4lUlETKFlxhQBrRwGDh22VBMv4GupG0
/+JK8zgJ4p4uaNhhO/sci/n1uKIn9YJOGR5iTb0g6jvLucg/2Qglw0nY5FAUEKr2uTEopyBPRU5e
Fpx4k1ipdyj+S+5OpdqHHI4dJoVGuQfz8WsA0869MPfGcvp1hnldfz/QJ1cBFYtQsMRzvnDGlOx2
mgRHoab73wNC8W8eiWLGS5Y0RCLwJFnX36/nxqBanpFcGWw7OxeNDbSZGE7/3y6gM3nDcT20DCss
QRxnd1e7mypQF2L1Srl41HV/Li8hkUzDLZPfMWvR/rLnyc8hYv4UpFz60Cb6h1KLmyW4e4lrG40O
NVOe39K4oz4sxolWeaQPkIVnHfpHA3RQGZprxGf7VA98TM+/crg30RXc3cAMYEMJOtBqGmFScvtg
Rv/PAldLwpdgF0y+OJKMIIHv2NsaN8ePIaYuHArl5DBzzQ/qFU39i9nWBMgFgRuNYbvjf0zUIZ26
4ri5x9ICvL3WDXQ7cJwER3JhiWwKYULm4cEOuLI6ERCYE/PSWmsvOV82NZ+gSy0dpvh9XW7uj73r
ESfdvU63b37mctqFLrOCn1CmIorM7efiGf7ED8CPuaY6MCaDPTVJGIOx939WopMqQzpn8/TMmJ4E
8LDpO5QY0J/BUqPn7rlMoWmPNBEBq3db4+W0Eg13cj4mqQF1NmxMhOY856cPxyOchazcUuKpWcwU
mgk0OhNap7ZkJRRR6XV+RjuYo014Mt49sqiVDDTQJT6CSnpcf2PLw1qi3jXVm2C2Iwv8IHSlff4K
ExPyptyKeP6Dl+mYaHtjpdAz/AY+Qk2diR1xCfktX4xBWZQARiR6W7tPQaZMm/smBoGPgjgF4diT
FIG3X2Gcp0YwSjP4mXkX3ofM4J+2fpsKH8YSiJ+6xZyXr6Vu48lN3t3xI2YH0QAXt/JXVezLp6eu
iGWzPaVQSFySWbO5FXHjioZU//gaPIZDcWeaRG0e2YccsUt5k0e8Tyu6+jPV57n7H6XX5PbcBNtZ
DDpW2uoj3eZCxpycUB79qAWaGEk0L+H9sRfun9yRRp4vYhQw14wj310/GULrKHD5XIIsiDer0OH5
wuvRpvjiHpVykLEAnvDuDHxPnOcD3Ahwm/Ic087mkHftsCHfPrO3VQSNYlV9T7Zdmnlj+/18Cge/
bwHcQA/JbERZJgCOPNpEJ+rw21OiB5Tn6GQXY/UgxopEPviOK83OY1WRZkPCJ8gff6iq7+4ejcSX
6/iJ2RuYIMQd6FM0ONIE1CQ92MxyDriNQlcQZmLnWpWNbjiyujCpjIPFLvjHGODRc4fj+ZO+VFh6
IgkeVr3geCcP4KyvLVklW2oX59y9u6K9lVNIFaQ2DMmnl3Jk461iCzTSntlUTQaN2Gf9GsBIqR8E
t7iZTrQUbdHMkoYKuNAPvq39pnl8MPQ8M2WhAYl3UUmHkdZ12QogWZWMpXyKvNKlro2Vbqmg0+he
Lr/3RkHSmG7IKPlmCJHWtuyyioPJDislFEWPd3n/2PKempZxnAROAhBIEo4MPK1UVVMjQVAU3831
7AaJZgpcYRdqAHxhQDUmJfnJ4Xt7psoeZLbReVOx+z5d21eVOpXKZTg0Z9mIqW96RwZhbHj7X7gU
RuJbvB5yv+/aE4RLp75AdihfgTnrDeG40dl17Sha7zB959YkON3+LQim71hQWS5r71EUmj0otW8Z
bVadHVMg6ut2ILxPHA16aHUuevXOKi3jsHFPcGNvIyfR/TfAuoVWGer2MgFgWy/UmAHVfn8XVLLz
u/rrrjIUeoIPwTRle5aPcvFF69ikW/PYk0bVGd9QDrdOwz688OYX/cKv7seHAddPMAHinfCTInFX
3mBXo+dsGMxdpyG1FGqJ9KbGgV2JiVBYub6/aZ0SYMIEJ9F1UB9OX3KQdodr+WhUndY1DYejKlac
AT4Kuukckp4pN4M76kwE9+EBIprLBs3L3dP0nFQew8owMKyhUmyQ6e1ynBmmTpzvrGQVVxLmxbTE
9HBu+pVI3a7iVhInLscl6UCExPTDivYa0Zkrcl12PR18xXx6HP/apOuKgEzCpNKVZ9tq0nYdZVkj
5GYucgozpvzNy02CKqTQ4LNniQSS/rYC9ycWH3mDWiHYCe8Jwm/mAqKvHd7Rvkjuu7rn7vtcbiEf
XcwHnwMv85SA1LpZjkOegA2CNXyFV7PerWpO2UhnoJUHkvSHnYhuRumfFTw3vzhNF4ltbPuYuBuo
R+g5GN7TdTibVL1OccCSwDEA6cS72lKfxq2suEi+t5sApw83XX2HjUS1w5/3vaBdiDZznMwffYUb
D5qEamjD+wTyOUfoLXltpegf9NFp87BkS8h8p4SIwnQciYqunUOs/HeEuE8gD+iIbtZjvawWUHsY
g2UMHYjrwtLIZ9WNCcU02AVB56I0y8Vr7ZVNtocaUt/UsYkvJzQAKfFOrcAavYu3BnV3lJEK+dr/
hQ4lHmHTpPU676wq+F28h8ojyA+AbxhWNq6mxEECI8GU8qt9UfoWOWsmGD5W9fE3A4s5PfIq+dcU
Dc+Qjhu4JUwZSgPssiZvgZmWPk5FQZ80T+qcyaRgNzpm45T740BmrLCBmoBzWVrJwaxRDMMvCt03
RNwvKQNIdpJO7rIll0Qo7n3GEiXqTBUS92LffBrxaBDLslf5GG5nlIjlQodZ/LXuplI4z7H5TehM
vYHyLsa6mgnd/+vz8AO/ZuCRTINKUv6F3o84aXEdZWma2VyV64mAc+M1/OQtq1g9NZiNpaReFR9K
bkKLSTZsghvqyBCeQMzyraC8IEHcAmzWvjSBU6aI6nGnumt2PeFijbSwv5sBQdfd50Q0FLDRRmqM
r1/q6z77tIm9X4ZYPs/eNya75LxiuEjL9/OthdSP8a530ZJmz4QsugDWhoIBbsQXvYnjPIPVOzNC
fGmo4MmsyMM4osFASZIg1zhH4YuXNejw0Uzu8rXqwWSXaouKvsr1vHuitUjW1rqRw3bJsE9UeyyJ
4emXFZbY049JZUCbzRx/DW1gazN/WVeeDPKglk6ZqfTBuFF6c2E6f2tsJXqeccpkXIp28/7Zn+kD
o3SBVZUnpoZT0R3LXa0EWytYkGNEFU7TP79yJmy4kknnbOcF1IgkN6OIyj9VEdXXw5k7fK0XKoZ0
1nVnIfrnZjiAqw9GS0hJe4G6vetPHP7MlY61hP/lWRTZuCCUNjGHX4ihS4eKQx3wkgMs0moKqUa0
KibFmDWzCBKQwfx+6k7ZPJoilE60JTZCtl6UHRiMt+UNQmDzwURrHO3VtGzGmG7Vn0t4rkQIyhIp
zpBy2HUoNhFUtobs8SRtQUhyvFvPc5AsNV3YRCLGDxfLwnb76hy6JzDH7a0mKT2X745l0SUR7dKV
OR5Id2GHQEn6UJfpjZ7rd08Dpy5jMDbG78tTqOFFBu0g7m6jKLksuHi0JZpLG2eHyBOmZl4qwrNR
yx8R/EpxxEOwDQx2aQeDiq7UvY6PyQIOHXynKG81dzW2IidYgHj8FrDXES+4ycsRftUaWMAEb7lT
C8mreLrBGc7BDQycMbWZi4o8llFLmYS8INkWCWacutXTqbYGoO4ROv8hF19A+UuKuBsnfYFW6bZS
1/nbCVGlI8zZwYpwh2HE37SLlEE8N1Rv55sDzEHirCN87P3RqYG5c5D3E5KatnrvhM1nPsRwRsj9
Rtpl6TfqujI9sukI/IPrkXNSXAWXCsVGW0lPNU5pd+s/OHzZhyuicKnSiJx5kN1KFafT8a15Clnt
Dlsa2FHN1rzhI3cmK7Qm7bfUNhfaa8SwG/gPsKOShVTWeFnCev2JCTHD4TC2FHlSE16xYveXg9yI
tipmsZVPW8hZtjYYyTUjM0/y7xVnAUAyikwInbmsIJ8ljpfg7BRVXrKtJmNFc8J4+161jjVB4kXy
pLOzXb0oCQEsfdTzVkP/eKObvxlKVKBGhi6JuZHwfartA62DfXI/f42K4FzJXqZuuqjrLWFv2a36
kVqjRuqonsPyUvIEvP1/13zYfzzAXd3GNUL4PNqj7YWM2pdssL0hSYCUUCvnOrAKOmtJpuUwcj3p
PLlbzXfCgngnAb4ygA+HG/UjsfHO4CG+fxc/KxIle1RFnNK7DhfTn+L7W6VL3lkEAMa4SjeYdANo
GY2G4RrCHtgO5JZSbvHvL56rJ2SlOrTvQbq/t/5U+WJQ1NOONYyTXd/YiYDMQGjLBE4L2Ow/PnmM
/MKJPAkg4em1z351HXWy2bwKndxGnLS+nQ/HUkhS9uuSUhCQP9+/F1Zv4KzGJGm+woT5vwfhO7NS
ZPYs0VAAtbrFknAXkMdeN+5byaeaIsZ/PryMU83M/WDgJjFg05tdwNMHEk8VucnXjYKl84zgX9hJ
0jNMfzXBBGlkrNZW/oNjwdLpBXsHShXyjntZQOJQtugZABxvO3wiw4rtiP4iQeDn08mYB0zrjdj8
u9Q1PE3DTQpQLvfl/m2MaMuqWwdpayvD2TdxzQQb9beOScIsraNjKB/rchCdGPjU/p3lL9NVoce1
BxERhx1AQAjSb0TrpMLjeXjItF/cj1koZB1dNqA/bnIHOH3Q/IcoKTVP7zXi99CvbhdgsKe36XJl
YXBFW8bS6xhYMyHtcKlVw8riocFoo3enLiJJ1NLPY8pvPHwc/sqfBEPs/C6oSm8k9rZ5zxj3l5eV
Vdzem+ChNkRkoOsoJvfMEvfFmOcAYxYYpR8BF4UJINACANd9gcxVtKnwcFthiL4NYL6wXfiVbgJ5
QsxmX9ZYPcv/6tx1ZuMveRUk2AOK9Ux/IdCuN6LtCUh8L+9cVJDi0HBGI1EO1xrxTmb+7X68lKF/
jsNx+Ny1VZdOJHGuZsBUq4Ah1yM0I9v0PEApbdwAcSsCUTd+4RsdD1MFWWGi3acqaK4t8Bc1f/xP
PG7SH8s/XA+9LVGPBPnE/zM02qFBXc7N8WuINMtm4BRTZZoE+O/ktHWeqQQ8IDdkpzCgbanEJNHd
4m1jV2+1qJU3sIgpcT9xDxxTT/dwXkap3nAOa8jMq5pp+xdu9Il5GKdLi9tCe5XLIvLlKpvICumM
aG65dzLrDrdkQiQsd950q+jNT6v451/dSjFK+XVcx5jmABus2Sl+dYGMFMWwjKMoz/48Zb4XZMqO
PT3SxyXwy+MknULTPAmyPaSP9O/hsNst0ofUnCu89fQ1X/vXm8rkwZpsWssItC/i3VxJc4+ztJI/
8+OXvO5GMBPni5Ysv68nPkD+3W76LEc4uR0gG66GYgC2QVfwTN8ApeJhiCJPWu9A0MfUHiQyrC7J
3/HREEuwseU9iE0L42LSy/5UeKYRklcLbmgXu1qsZUUJs2tqrRW/I5oyDo+mwkMMStg9BFfTloqq
EdAmD17Ume8H27UWUu1BX1xXlfigul5K35BYe0VswKFft+w7YayV136Ud1EhqnjYip6UljRuKVji
+ilUNFqww8k6pp1ty9ZTohQyIdSGvap1djqMy74hDeHLc5wzZfFisejW1tLTb2/IESixVPEOaC8a
sJzrkS/l47III9qhcjIoctKUSG+dGSGNRWKpkLf2NvT17VcnaFh9yfPNnOfS8KwJUId4pKfPgiS7
Tj+TMobMcTBqbmKTV5R635lAOHUHcQ+HiLsreXoph9T5WlCBo6nskZy05oa1eJ+H0KmlYn1ZSMYq
YHkVo5+DrmIlLKo1wdno9Wxg8JONzmgfKAHyW2QQxZSug8frglIgQoDgwFfbbbl9bjP4MY9wq0h6
+lNviOeRz9YMlm5ujyu538O+vc2DrL6QMFuTHDPv2b9E7p/qiifwjsLQGlEXEr65JgL9Y9KuINUE
1M+PjGRaIDi4g6bGfXScFnpULMBONc6Vi36c8PlgL3klT5mJ8Zn1A8ErS3TPwikaZ+yJFEtet/UG
2dWyjGOtDAqlCDGSUKYtvjW2sdmWrcTor+9AvqN2TuLEDcFmGhqa4OJNMXWyd5IKfrvJQgRFN8u+
SkZTD+qof7AeMVRsQ5WyjyLkUMFGyBzdu6NhcH7FJsUyvTfqRR24U2Kmq8xy2okC0/92oR+Uc9wz
KOX7/ZaMvcirv/cXoiWS+iHgpoDxDNdoyo4HSzf6Nx3bojWE2X/RgOvHK1LStJUK4y9eWk7mvtP9
9TkD/vchHexYS0CSpxlwinMfbsSBXRQ4KSs6KE0uwOjgOhidB/4NkmtxG21tTfDLLxvIIkrARLA6
A+/CtsLDcSo0HmQbynKdZEzp3YmSRcg+zISXU/T7aT1fb20lUKbKqzw107upTf3nmjcSCvnY+YuS
BjnSIMGUfJ6WzdOmLOdjP4hDtoeO/qEhf1fkFP/z+1/qtYR5hGGztRDBwpYoZVkn3q9BasPcQqmu
lwbZsngVr2YgYTSFK6SE4P9cpvVpSEruSh0UM3H3CaRmkZTjePwS187rmCnTGzuo9FPJtLKsnPCC
tIa3YCbNRa9l49+ozNhwcSStci9iXzRD/TGGVmMuv96vhUSuhvzS2z6H0GYorIh3IYAEPQr+COdI
fTPlWdg5ajrFeHELfAIzocZWNkoiPwiF4SxvfeshYyU6UxxYXcqpSzS5VH2FRYW49Ssgics8YQCR
LqXTCxbrWreDmyU/AbALGq/DFCgQ7mPahkZaiu8mvtLAzLtVXysGb5+9qg80tMi709gqvW/WKV/k
y44MGjYNFqXCo1vGrgrw65ioNuNBZV/h1coiQsdZ6Oewv6ydPcSoUEGfTa2nPw5+MPTZRuP8tHMa
DhNVPTgFWNHA9/ENj+oO4rAIUvycqu8/oHD7ppw9NMwAxm+bUv2EBNKln3+DPhIdtEGDBBuLRXz0
Km6c9YChqPw2sbUasC2sQNNyLn3sFAroFRxdCVAcDx1mZLg/4laOxUkSsCOBonJbhZWxnWh1rHru
apSwYiDSfp97RGkc6tHnDnVBNnrITxRLLGSEyPs0cj30MuqxsBeIqp/mWj3v43xp6+rjaL3u8CgC
i7baVKjU7L7+ubH/+fzk/MiddXYO1kZ00h/k3htQcS2di13SVoPVOoB3IVMMFRZRLkcnZ+miXSdS
/5E9ajTEsyb6UPPh0xIKDu5YkDRL6Y5Avl3h3qIHetrFRduQaobG82iAmrn5ogfDwQKZJCSpbnE8
PItq1wD7Elkwd6bT9QC1To86i6AyysI0sBFr2OWWmbPT3MFVdLNxUrQjyaH0DQbJedgSvj0kttEz
q57+r4VJoV4h/7VBxbXbu1e9uilDI4/h5A8Gqzmgp8AtYuZnQ5XgkXK7D5in7kFi/VkmXnY6Sna1
AReqGLL9P2+EN1AhHvx+Zuqe33TooL4Fw3YJrWWuXKSbLCW7pG7NxdbYbL/VbDqGMdYWaCq+egmZ
uU7wIfjNguWpCjJoFlEx3vSZmQyPofhk7tPDDg44NUME4wBJUjglRidMpg9nGdOCuTR0NFUhM4q1
K8q3/Xi96+SP3TG/yI7GDS7cbr2s11cP1CqWJO3cL3DD75UElXglko0uYTpl4GGUXXWdv+VfNk1S
cpyMkFPcAQNPc6hkTNGNy/YAnEh0T4oB7yBIXsWHLYaVNIyYyJ3T5Ir94lrHpVtEtsn23mPd4VAe
56M589qdv9UqhJT03XmLivUayM33LlToef0iif+4FuKpnGNRQH320aV/X93v4Ww3VfCCIuU0/2au
fsKhUtLhW4+OzYLlWn04bNiMw1PnysT9ekp1tGYppIe+T2Zxa49gXT28SUhI7CxcT+uNnc9/EYPe
oxdxp9Ozqhq/YLPp9yYj2rhRvdC20I+TD6jIF96hN4y/yDo/wyvrdOzinmk5YcWjlU6XeQ2Ff5Kt
Dm4FaMq1gH6YfUHJdGgjR3DGb8SIgzfL1K5Aya0llveTtcTDJtIaQIk+QUKieLk3nnt2GTNjrKXM
fxPz0JWJlBeM48ZTD6fLKByJIF3EJPkAXsOrVuoaVHiZE24HegFL1Dk0R59hN6ohVRpQLwK3+5gk
u8xGV9EKbocudpJ0M5O6iJZ/zIyJt7j5JnUoNjnqpgyWceaRBxWBWKb5vEA7ClxVAW5Bu3PKtoZ4
JEK4gnhRu2mGLeeZZtH1R3Cqj33p6CneYKWhdY1JWl2Vs4Zqmw78ygCdaL+JisX90QxEgplYtJWI
vn4x4Zi8uVeoeQkU6uwqeq+jPOUr6myAlKdFbhUoBUh3w3ITRnKKq7vwnY7nAUBRLnCbUjqr400P
McdPZqaZzx39x45lBKgcyBR2BbkNyqqohLK/+kA5UauteemG0H+vTlmO2sBwUCEG42q02wCLuuWh
GArLJJTiDN9TLiZqrxTTnDg9T6Go5C6DIhNr2MHyDPKr8BIppH36VMExjsLyndM+Ata16tsNrUmV
5OsnGmkJ+hUzhIuSuwbtbN6VUC+tXZlXUDH/7BNdJE9tp//JblufBEEDsYeimv/NushcqokjdOZ6
Qww8EvhPe7AKGEDAtJXRSYIGa5XaeNJGvFplOrvlMAiyvW0mP4ByD5Wdnew9kzA4cxNmcgntIrQH
ySOc5w8Qttb9LG2MZDtBGRqzcNtWDSLawuPBP30DjGm87Ykc3Zfw1G1rI2GW5ovgNw//mUyuCEDN
zxZCpwPiW7lQO0SRgmq97SRzLrnKh8yCklYMgpYwbYaxhSnlO2FC7e+AHJkpYBiBTQsOAUtslh7m
ZvrNBajvmjmX3h8XseqxXQgdEfkx0uazyRAka1YKi7mwSbroT0SffSgJNmcWL/+ahy1ZCv485QiG
xBLoLoNwmVIwNS3NbwP1+OPxJ8J6xxww7LNF1IjWuDGKKQ88WVcQ8Fk6cG8+Bi+GgRGfQPuL/WFI
33c7Cw+I+Mc6rTYsC8y5QDWntwJ6zH6PZywGV/cs7jBgrhmK8n6HVrfRCYcfv+BD4wpDADzffljq
6ch5fDFpOixNl9VtjaZhl/mMIy9Zu095Lr8jV3OFb66pHb+8pYVdF1oasOBSJEflcIMWD2SgV/LF
0dDPNc0LQEPI10itvgz2+mLrSpKmLE38sGXGyra+jUyfX22+jEq/RyhCEAvG9LudoMFH1/vX4GBQ
znMFZIRN/uHzZYfZ0U1Xiupfl0+kWxlaDeLGnju9TpbSGnaucNTbQNbd5l1/Vu/j3p/p/e/8nbIi
d5TVwOw1Z0rJD7ysphjUCA5gf+Sv03kiV4W2E3U9vNtZFoyhCZRVIJt9xsm41dF44yQt/7fv2n4k
DsGau4MUObU1rzhqgEgSz2SIEFWXWQO1fev+8/vBo4iivmWEJBGuzj2p8yt9otHPXIOqO3XogLjz
A8NVshItdknfyHSiRGMmvQoJBz16Bw8UTzfMwmzCVLt0b/Rd1TyeMs02pwrextxgmXxcsa3Cp28U
Fejj8GNPvHcuCJUxV0ty2eRBIddxRcQ+WZ1BKU09oeVW1elWHB7g3KgSbhZ0afRJ/zzfaYBZkQt+
5UkJGcyehCLC2LPrMXuSmP4x/bXPOqnCJUO4uyTTbYRYkA0h0bMbTprg6a/zAZrtnyXB2+pHT/gV
iSRjMAzq1rHANMihHxIDvS0bzv1Nnwjl+R3c9LrKEVF5MMkucFEBlXwK77s433yE0UnqwoW+RD6S
87FTjiioCr+1c9t3rYd7Q8qOviJghHXAAWPHbr2UNLFNXQOp7NF+i4Grl2POd04Sost5Tm1lHMcg
rSGWUskQYTxM5xtAFbIv5WaI6g2ZeIeYuWfZPq5CpOtcLeUsQsqjpRd5ac+aRxa7OhgvWPScY0zb
ZKt6GzmiU8FXVu9FLoE8BRlvULtbZjkSRp4poggZL5f5QGOY7lp2Av36b3BFqeLrwH2Lvz84l/MJ
w9ZqO45dh6tUImi8YiYSurvR37mQ93es6ziUFprLQIANwme8T/HlCNUn7Y9r4GKm3zZFuEvakIgf
RKZYnIApIFnpCnMvtx2JRVb8Uy+5cXNXOxJwNJCZ8R0K6BR3M66mZJZs5qxvkcC5BkM3CrmDSw3q
feRCKHbRi1/8VIZ2moPSMxBCdgHwza+e5GSSv8d4AiW84WH6creXvlPMee7sDSm0cusxNiWG95s4
gKD5KrW/2Y7i0ZGI95cQYcqzZm3uEu9Xs0wmTnwHcDSip2FUt+cahjYw1LzTk2sIybCz13BZG/kr
E4cqMe7GVSw8qhDAETa8XSB6HCpJv7s7iBELEBy9Lrsu7bqNyHRudN9ZLYntyYx3CzTe9RLePPns
nZH9UZnAiDq3rq5FzXdh2lKsiR03ZEGYMJzBIhe3nLtW8gt/wgYCT1ZTOVKnKXoNMYD9N6TR+A8h
5v/PwptwNNM8B849grPMIOlgcMI7X0Y6lJCz+Ug7EmksdDAMYRzkjtjOC6+G+pbj+78kqAHnO9uj
9xZyevEt8ioHNJi6cjU3UaLHoekMWyxqTgVhOtdfRQ4UY+ZzhBBU3p8X8ZAxrEY3W4RKshq0qJt3
vMkE+VSlbLuObJLANK8WnjHCb0W+fmw+iMSnAvUTv1wuBu96n+gKUsyWuIbUawmxLYdeROJmZc02
lYHp5GxaYi9eH45iwpt80wKZOA7QYpJReGDM95IGmsEmXkhdWoWE6rBsnbSu9iGC6uKjo+V1U12Q
1jgUxkd92FKPOtwDj3YJU+Vbdbc3eS4zU9Gf+qOrSXxvud61UQIy0rdXuNCUOYNnOUet6v9dKUtA
Tbwp2IrLDt50Udz+LmHu7HCGD6S7lTL5i5ED7w6MyU6u3yoqZxNvdJGLMsTBx0TnoY9LZZ/jW/Qi
UCF1p7mudx09lqCeehWYzR5BzDE/RWkaJ7bcID7DrbmFuR4l8ON3AWAe0WXBDG9Mp8XJOZ+T+90f
qlxh/4okH/PcIbwHfJmyIAybIcQlBkRQfayw/OlsYzsrMpK9UMszW+eq9QgLYWvY2N8fBImaZZX/
axJ52+f+XXWIIohPYUsBfvTjYD7OawHEVWeCUvBsB9IavPFAXBieVJjQ4iO6XEx2XeYpGN8vxDB5
wFVXXnFOb6B4ghBpsTj1gvOz4iA4uCfmCxm5/bZKD7ZNBwLEkqa4NpqMB00PnCULYrpVKjHYI30v
8yRHTEuBR65SZKDu0jzinfIB2byrvPoW/rJ43P4dxF53SKdQlEbYDWKWYomfZtKnOb+vfFlmIPu+
x/d8ivhE5Ep3UAQlR8A8aLBWUTEial0B9M0yxPoQdxjAvDL0CSZJe78/Gd/9VihbU35fAPtONR4n
mqt/6itY7srDpl4ncktxDR96QcCh83m/LDBiPBXpV54xMw0bctXPwkDNK0S3qFJ75rpeUlzB5ba3
kYs8I1P015yumFsiWjjmLpwFQJ10Q1ROePgNDqpa7mJrnUOSUP6ZmmEtgSSIvRMxY42l2Gn9iCd9
OeW7mtFMqBIkaf3wpnfK8MDd4QCFGl+0yOL99tDKKPXNiL05GHFISoTlySPuTceZpoINE1hDoXHh
NOjFIY69Z4+tgxXZtXl0CLEgvFE0ya5Yv97ZUXY6PzBDTqBK+qZBDvyYdGHGU+Jxorm0Ckouyxun
lz6T21iot0m+dmnglBsJQMzc3a7rZ08CGhZ8zkrgB2mPEjr1d+oqGPqYo5i76vUDwcTh+QJEaM6B
Zud6siLkYAUQcft4O/W54wNoooRUonXT7j406nBDhdnYiheXBa/u98n4mNUnsOGKNkyOe5LC+wvf
3zGe33uVuptHtWmX8Vt7ePoHksIPiAF5PJ+1DzCOQ+u3sOMY+81oIVF7xQacKo2i7WC6hwbJFybC
GpjKWtIChfVR1qgJqEQ8TPOUVhfBM43Q2uffYMP+LU0a0NGq7btK9DtIsQDV4xyfWnvx/kWl0Tn0
bg+fMq4YtCidKmAUScUsNxpsYE5LqloAJBRfJVuxnQPYjvEQX0u3wzkZMwzOYcPjojDvmsFhUzWk
aDRuGAUAr+f5LU+6uu5XMoxtaPPO9jw0ZbvqHlPLw97oIUJplyKbmMlChf7eD8A44byx8/1o0PgU
xbEaqYvzfoDNjajqWTzt2D7VH29vCSIh3MxTEAG85EzBJepDQKh7RW9Oj/9ep6Swyj2CvZdiTmOf
Jj9tvHx/R30meyKP7RyzE57Kn8by/pS1Ll6vqH3u7+e/m+9VdYAlSi+hksd16M2pa5zYp9gaGDMR
zio8zxFx5mns2yvkxMt2+2EpNsLgEnt1JHtftgZyegxp3kXbHYZSX6v6j8+nePBOxV1OnqpCSGLF
BbnX7GtqMRJRRtoOLrMZuMwqfAvGp+/uKCFFBgmZX1AYweywFdy/wwGrfd3dlNuILMoCoCSOuHEI
BOOp2t6zX/xE/zdXXRSDutH6RuaZ17ep5lKBg8TK0gJdfnDBj76MqyueehzBi6wqqOtmFHp1c0Z8
f+Y2e3CfkQGw2Ez/itIj5eVgHP1VCV3vkuYyiammOeA29ewpbBWTiG7pg1Z1ThByrdEUb78ORUwO
YMTZglx0kEDXkKUVgdVot0K0OZ5qaX8Gq1LvSvygiygWapipt8E5IH1wc9cFvWcEMMCXZHlxCzzq
KviVg3pKxSiFf+pKZlNdy4bMystCUfv/P/856UGE9T1TtF0sKHO3kOnJHGOXQuEpWy/TWeyZ603l
4m9QJiPZUlJyAlJ8guYybmRTsdHez6FIPL7wODStsmRk9NLTdhbXL7nocats2ELH35QZjZLFublL
cEc/VaDir6ldekUakVudSLCq7CavXSvseBwshda8qQFkv95I7Tlq1XJ43H/zKnb/WByyXaiELR0h
VpAoL+eEkwKl7M1B0WD1OQBBDqnNUT3YoEw8ifVLzXNbD71bBpsiOqTuXFyxQAgnT1cNidRF5PDo
a7KGZK+6d6uqsF2IOG9D6Ov+fJJWbUvTMRRGoI6uhOLjpih+VMbyl+yRlrUKxdsSMS4bnll/WRwn
9HPabA1oMoFl+SFkWhBTyEH53gUcQHZvdv/K9CdX6hqwAKrS8vzF4LRYBTIdNiAMl7cPUnYSJe9Q
ctrp7IUdm3XrSdIPZwBg4RJcgsIFMm/SN6Xrvx6PLR1a68sCT0hAebwxpXzevVWB8uGo1MfBcAt8
OBQAEQOPHAWDhkCrwmR60flEe+WK2fiZbN+vu4czJvvrLemT3/VocQpveeCKvsm5R7QHvw6tytn3
zz8lwAf58Bd7PLOyYtH17AnZ3s1sQwUqiweqwqlVYPda8JvEWlXrunJtzzq97qsVCx/TZur5MbV1
OFLglzfOEOo01VhR68AKpM4BuzXHKheuCuXM0myCWlx4OhpvbG9QS03nKlJjiXwiPE16O1SSXjhB
J+N5YTlgOeCCIwvsQX6e9ZM4xKYv42asZ5ZJ5kYpMQC0cpBBbZ+nzFI8lWnHjMAs0CjgDgnfwJ6x
OZJn+IOBeYtZaOo0jeNMnY7gP5N/pE+jUQPS5aX7vFdtGbzPV3h+IE1rrLf6et+z52fMZ+jttvM9
mTkRDDnuFd1geZI2j0DtqvSkZ9gnlFRBKrJBfa7b5vj0NRnv7ofUkbDd0KNNmcAy7Q3T5XBHwgOH
CShcWcEIodi39L1P64Fg0SlKMbAsI7HjLwZwIQvax3enMB2WjokWZV23ggNmiEZHo4KGuQQuh+aY
NizJYfzi/KKnfsOWDjbiom3DkExRiCfbYbQv6HSuIr2S2PtJdkI0v5vTkX0PWRPvgyIQDRbHuEwP
W/PlmwYsrapusvTSizWE9rKV44vGjL3iFIyWpjGfycpmg1TzWiGjeLhlMignKpjHOpTMZnk5ZxCU
vNA9BTnoWQlNoRE/NB0WGdzcwsckwLRmmdXHIk8tLFOVclcpZriOZmHFjJ6m4+7YTDCOsj3uraBg
veOLVzrK8UcAM9HmYRc9tDqf3GtdRLODG8PKBaBoVvszq5LjXotItyAzkMK+oMHfqKOW6JIhOJj7
iR1+JTAGEOFnxL+QDajeZEPtcRaMdbkFeaXKU8SIhcGmUQbV5ip5eMzlsnivr2KoXakoZZWcaH/K
ZL9XUkp6olCDAQNvmKOHIFvYp+CxPw/jA4zplyy0Gp1QWT5xNB2b+rH7bLNN/iVLVhbCfc3dKPl+
znux1RR4Sj4NYCsm6RlICtZB0mKJkMUUJ9aNE24l87uMAq65Be4Ewe96p52qYBasqIQri6yj/0vS
O04TlM0BlDJnT9nHI6vfDqIY3iHOwtGtyJju/4z6s7MD9vxLd2ZbnvTIBh4g90S2K+uQ4iW5t7nu
6lxI/6IqGtpJVd0RzhixO0mbYGuicrWgszlQC2VD85ySrjAkouT3DjFdL5OipLeHBnLESab/HSxN
CnsNlS6B2hXijs43pN6ewyQ0j1/De4ADyhiBTo0H73Nnv5pmk0f2UqTusBozTcBFDKiACfiaq2g3
9/cfIXcCrB5rwSJRB6KchQYUbsG3DF1uuGs5TK1x/dSaOb951JBihOvKKLyh02k0Qlfv0+VlZYIr
StewnXH12k0KPa2zvccL+oUmcLa6L1gLwFZtdW1pRBEnHMLCqCDxq1WdD60o63/wuK2tEuIRcG66
+b3hF72duxaXpB9NiHtwOhJJ3/l7bq28tJseaCiAaQO6xhAP7yjN+h0JXrjQYGEc5RTymNLzCszG
HB5//qqbywiXeNf/ObQ1R8hyoii72y77JvSJBiO7uLLl0VcwTQTiHSCk9qba5kTkon9SwqocscLX
1h39lg9EmQKwtKmZD14QiIzjiEmhM3PyRaYN/uM+4jW0D/5FvpzAEzbqjJ9B4Psmb+pXxpQqJl7x
bUmY2GngbB9xCJ2R1fLkNfDIvFteLQlVWLm2hg0PhUjrdiBpRdqO+AeHys2xt2Rn2uGZczgiGV/Z
nf9nUkUzxDa5sgUyjntNKM34FiLJkmBQ1/MOL3nuXG49FOeAf9TuF8aUQm5FhDkLh3VQDgxFQBk9
x6LbOBN49+c8vbtSOtsRxWbMt5B+6LwL2N5HX6CDmUl5I/IttCWsjNYNZ00Yb2Y5UfIbJa7y5ABj
cvrwcFXyQwZzqQrFTBbWl75y3uCj/Y7OD21pqOThiXKusMd5OXlSx0yIdyMgqeRXRd76v2TgqtxO
H1GSlc6oEVy/KI5GdkoFMCVgGQVOQ3jSXhU8Tcpcji10/112R/MSgji/bh67eLuFkwci/uMX4Fty
u2VDlul+q5chKxJZJn8pTJPlKduOHCMlDdqRfTDurG5WrYAF5ocul2+uA6yKh9gdODQAk/jm7qcG
HTePld5g9HcnmWvwOm0QV2pJBVQfgYHAKKRat422gEsX4lx7ESdtLe6aWmGMjJeGMVYsI53vDeZ/
Oh5LslF4Q+934IwJuURK/dCSq7+t1QwzQbnJ18aNB4MBbOtQ45aEaemVHYHcjMk8TfAsM17DvT4g
+saki673Xg1oxTTj4EKrYzs1APzYD3+5Qah3KYGeAKBYwrsEaMCNVDiO4aM8L9WNGrAlEhHgp+6P
yO7RPma6EY5Mdn2qeAl2l1+B/pvWCT1KA9lg3M4uZh+taob+yfiLXFmdv4tmojD39WuFqbFfmbbi
8IR97IPPxP37sfaLgFAOLRGJKNLYORCFMM4NzEvRVir0idr4yxRNRpdNOOaZSut+BFhI4gcEFMPr
2Fp8Qd0RTZgPAD7w+EAHSQJ+A1VDL+vlUS4RWm/Gz3jbwfs+/P8ORfpt5IFSHOK2J1H4m82v9Hbz
oMq4/zgXniBjehG5za8gEC8pcxC8qRKbYQ4G8S5a21oNAiUQSoSx6RSoy+ENV8LLJNpIczQa792i
0FbUEaeKYTvBoKXIeXWKxzxO2Gj2V+LQwwIj66+wG68BTuXBStn2KH0ZQyCSuYjyilsXMYQ/89mL
909O6/+kTdV4f4LH+CjX70GcSEeVHIOJc0CY7QrhhW7kZhDdXmtmb6Te2L01AN3eltD01nyQU8Kj
rzaQSSxzt++ZRAMkJhe4dm/HOAeIJ/ee97iE+JELNngbrN0KaNErpvGmhoAmxRolUAxjgDzjWdUL
Pkgwi34yru9I1/rF2Z08u2kc8XaRkmKMMilCr7lS5bvSWQ6SbwWZ84FAqSomVN8VT2JL04d3V0Nd
Kt/uD2IvWwuy2svdrwsHGmkYwF/tst2TQsOhkL+oMj3AD4MtIc6TxG4qo3C8Q16zl8Ap0UkguUm9
RCepddFzy/qCfJZx59doK12bGPeu5Azh/lufv9K7brvICS8s3JvxGRKe5dgTr0FGCxiw2oRzOxng
SGcPYzPT71HYMRLtvkivlVMoMrsLUYbIODWXxw6cqK8WduCTdfPX1XVMY3lYet7rqe4SpMJtT2pU
gf6tk7s6IX3kV7xkLD3zOn4jmQnBiwg+6+8iyQbzudXW/KwgpOrenp7x3HfcJxmDNWLpioKNh3ip
VIVXWAcWfvbtpeoGHeyj5MLTE8nO7EH70udKk5y6PCz5DeraOJHiJx8XgYOobqCGtuNZEoEFpvgz
s7ftp+6wKKMdpLWpsURa3dn7Y1yAVF/rrpXLWoIkMX4ynj9PKcRmIoPHxwpEtHG8u9vS/bgOjSGi
yjEz8/9haGM89zzPbBfodLnXMZ31QQ9fYAyDGg/d0MG1Op1RT93R6tFNIsaUpeR3G+WXcilqdoO2
wjgW4GkVP0ndOG8fJq3kYbTshs52GJmsnYYWa2y786MjzChLQsz6vkb3XPtS989jj7jkvPU8d49F
MKvKRDq7xnYxj4aSqtDFVvHR3kweEkKVmJzreWdWWGcU98EHMDLFYLTQOgexUph9oNks6RH+jDd+
dvLRWRSIcVjMQe+EXPBOphz+y+yCL89ry+LGnnLswcSz8rvlTiwf50F+qgxsmhYYEiaFQJOf/V8W
TMdfNdNhFP+OrK3p6i6CeAf0CeAFLPR04rkpjWeMkFlyCy98RxN+sJD7lDpaXfDyun8N1Y+18I+Y
0MxvbXFEb22gqI6V7bWQISPO+Pn4pcgDMHIHefi54ZdzswdX+FUtGqY0Ic/6uYj68gIa4P/bAzmI
E9r/kF9tuNJ1opfm290PvYdhloGY6OC+vRBG6NRkvBxzDub77tnbHNqLIh853eKt88/yiujfo/qt
haydXZqJ73mq9t3F+DOjBxgUz69FCQ1zkANgojhLJZKd7SCeVK2d1dolOoHxQhm0vCQ7YSS8Ud5Q
FA4uMN5xk81tzEyRuckcAYtra4r4mJ18myD9IF/UwV0HvINQN8lXNY+Kzcnjao2eLpfB64xKNgqX
IfzJTITl8s43SMrA5zT2GTvUBBQMTiphbgxnKm93mJ++1SI5Gtf4I4ld4DaXdDz4fN3juLkhT3Qf
mqqFY3wDEVsNKMyPhJU8nSdrjbDenBfpKPRMY6ihCpZoshTJHihb8hcCITUKEiwXAS69mRriOWtE
FuWb1A+YPxhBwivSHL1LxpCjUF1xxNQfFbot/Ku7EUM3UdfI2hSxtbDo2UYg/T11yisY7T82Q8yl
fK10yYw0zhJuhJsNRapdNjUGD7ekllA6ofaIjoSqnI1FxWSLLNwIcCyOO8/0bVHvacUzY+UGTs8w
xJPjkeAB4fPZc/zl1z/htQo/SJFR879e28sIIlUYt7iMpn34sgmNoKzHkV4BBZZ2t3XYpldlcS9G
N1/8qNfwvx/SSU+yH+CPnqxgCstqQTJtfNDmdg4kcf9vTnptigUQB/9fTboA+EWS7BxIwoio1YK8
uzI0QzXJ0KE7MVtXZbb5xC8Ljb+sl0ANd2IS+AQPQ91neLCeQNcuff/O378RZdP2OskKY08DGfNp
bkCjHZLl8Eebiyd6ugVyvR6V8Jwj5c2w9eK8ZEabOGJ1FgOmVHZBTIURmisgGQy47X48/JzYJMWy
Hppcjv5LKWyiaSDNOizJfMZJ0vG+XiYXKzmmTd3U7N5bvkBF2iFLx9k+z1nwmw1Q0EnjATaiE+b/
Iksk9pZ2473z4yjjrsloj5FviUdmKwiXiJaX14Gm88nx2Tt++50KgxSoBxRchYxVZWP5IZnDryG3
EalFdiG4EcnMHAqpg4iNHy7L/YHxOFtFu2+qVfVfD3cJpxVXpVV5TOMGgPhIl5UkN9TdyH433E2U
T8yj/N1YIrMw8q5FWQTft64Jr3+oRH+u6+OmW8g/RofhisXxCd/gflxxMtG6nllMufK9TeNYpGYY
YsKMn4chz1GOHzINnGeBKm3d46TS+d982pu56bOmYoNnsiyzCuDZr2m0+0RNw1S5HJMX3I6v3KsI
OU95isQoiKDkmaFnEs9kAODfWITkVZQlMnP1wGPJZ4v3pU49P+F+vquqO/akc0VSdCgWpyDMovia
obyHk1PsoPK2Q7v6Fn2cOkJNeDcvJ97kiN2KdynSGqKucItSUNBlZ30x+/JGDi2eYcYlTKyjdecM
7VHO8W2RDneqO2fgq6szqoxLWeo6vVvn5bSnAE5kp+yQjJ407jBo6U3kLMDBWYEVxa2Nc5TIGzsH
0dTmgwsIfoMsArmEjNEu+K0uHVeI62ulJ/drsSKlf5rICd6sAMlHrZFiK/PU3qis+aKETtbwJ8P6
0pTqJujsVneuwS38MJtFJJdyPT+YmBxzX6h7w+CHPX2b1Hyv55BzDOZo3x3JGOB0BwKBNAwxitlE
22Xee1qg3M0Bz19znHiUQj7KgwccRkDA0gC0y0c6++caumh+iEW1fswcZY1bUrWeZBB4H8XRiygL
dE0dp0LtaSZjYJbK4vSa2pCmH7HqyHKt9VNJ8hkfbJGIgAt6DBzxGaYn2STCA5IxIM51X/ZGcTg5
BiwqX2pPUFQKShDRyYUBO1AOxzzPg0YRxzm/hjA6J2HjDyO2K/vgnXs53xtMy48nPuORj06g2rgl
Zl24k0MkvNwW2fY/y5WpJW28Zp62SrsVaJSKeTM3ltRrumRLRYxAQK52S0eF5tylqqEzTjfcBm32
vulqnSK6DfWIeTejOIZk1Q4nLG6S+MyUsTiXo6RuaQZtR2YyXekPmcxjXDYs5jGB7QQhyfM9DuUT
KM4tM5xPm41fS6OmJ8Azv4+obeleEsyDh9PAKnb8m0Kx7JmJTqXVfAIXWwTIzid8DlDVzvoSw7wM
BwWIlTG1MvhHAmuK8ot7XMzcFw7sYI7iQoChMiMTrE42/lZLTq5lg+h2ljBb8YNXbGHyTZkijS1g
osa78gmbGpWq1ky5qMWTDh9WBUBiZQrFKkEbLxz+pAx1qYs9oAj4789tORlfQ5pV0gkKnd6c15qD
qvLmzByAEa3fAAmi+7ctX4SMczhApnDTlhOnWK9EgeA8ciC9jhNrHtmjaP9+h213jVvZx49CnWoe
SAf72hiTiF+MP9Ks/apeu8YlzidBm0z/6wziwEZfPNxlu8dD8yWcNW35esY7moqfaVny5WPTOdaX
wECE6GT41B4PEQSCuZH5vH1pLf881tNwN9G7V7Oq++3H4SQ6uFFFKFC6yupZU+RLArdzJjOzPZMo
Mo89J3MKn2kZGc58kTJOeJ6YdhCjcubw1P0WZ5JSppMrObnervwYLl23VS2gwSzw6RP8eR11piRb
/9OOYBrPMVjPWRskkPaNZzqV8Nwy824qC3xUDJkabZWHs5pIABcADonGr3EB5x5CdIpPnH7S2jV1
bhuw12co97yMpT43w8WRXAmCXeuZ85qhToPbMLMi4yLJuaoNrqnxYTRB/4gedIB8turoM++6VwDq
F9MSadSg1+6DX5nqyIy5wdv0veJLPWAu+NHHrYGWNqa3xL/gs6u/t4+OplRW6C8Q1owwpG5e/wTy
ZeYTfbK/SPleSIfnwWIFQxTt2xl59UlepQYwHnF4wo8uctz19FHfAb6D62GG+im+gF5lL8VI+r35
2Kk5GTK8VB3U/M7xhmzNqikUeah5wlSlj1n/1oZU2974xOlRrHdQENU5iIRa6hM/xaJp71FMioRu
nYLrmlDuqSgmvmtekUfbpaVohx/MkzZw+3eoDr02AGJaSkNc6HclLlm5S/AN4pSWqy+Ctmm1B+Ko
aADNkJowc3xZfBTjFi0QbTxl8nbfIi2GVNcA48S5eSUsS+z43/6DQdmRf7NNLrk6/NjbdpCyxke9
4wUGLnDr8ioFg31ssYOtNQrNwIL4YwmoBo7U1VYQVD32vAwz23ZR58Dho010s+3N6QL25FRUsoTG
CFDygsN5WyweMmuSQduXlzNNGlCxJwMMdTiksIIZIIf4ZRIeHj0/dZUb4+1BkcDaUd8Oj8mPJBbH
Y9PgxFpIqOk1/SPKJYKjD0qMdbWzrPS79OS2O6Sl5+tBEYbNZsMayPQzWXZ+Aa/UOaGd51vVJ2/H
DGDxMRreF0CjbLcAjj9PdZMWuNB4dib0f7sYGpPyz7WCy7XJHXbHpcI47Y7mp1BDhXPzxBPeIXLF
8ZELlvQXAHIHQ8nIU/YMARfqMaCNCkTzVpPEnAFuXY6X8Xq0ZQBTk63j1uMBGAXX1he40tQLD693
RbPuQDSH5jELomnmMMx8ICbtBry8GTZlmbdQThMoXFwD/meZtJFAnGkUOhxZ+sr9GrYxhoIrUtkj
GiuIlRbbM6upjfsAQH1vg6hMRjd5gSwZnpF8UR9+oMaiIj45F7jv59W2j2mx8+krsFNYQ/Q/D9G4
HSB9oGdXfh250Rp4vckCnhJLOz8m3b7K7GLhoj9q5YBPIWTJ1TEZ3bTQIOaaTSN3v91SupJogvsA
a4HgT0/M2ftTEV7z2DoaxL6YDjK3ifwi5RAn/QAidcrdVm0FMXM+uAZcDHea2stP2uXbhmzxCcZ7
FIuATVe0V2cGNRURYguc1E04QIxT53z2TxuoQRl/tGwEDfUA2Ss0J7x2mG/flWkTqyGz76hoJa3h
iagvfNIcJPCb3SZ5X8+PxvkCtD9SBVHVKbFcwAOB1sp1+E6gCH9B7JTrsfs1yjrUdJp/XUQMPge9
TCMygaVVgHuoZE0pcZoZSxZSef2jxA7KPllYAuG7T7TMjJFZoWHrurv8v0C7i4ERNYmxcd51MMXo
48IpNXCvFMhR5hnTp5FQAbt3qHJkecd8vCWfr01d8UbZkj0jsFeVDJlfagOAOU/sV01pJ/ssugpL
q2nzg8pMY/PzmaRHAJ1+o527wyMrceFPaAZacvUL4MUfBJlN6FwV6+U1IWepQJlz+twh87W5TEv1
SBf+fZ4cmqG6utFIRpv9+gtEJaZYwM28pNWGSWb6Rwl0M7gAz9FYPuu1MpkjKW9gRitv/NWNz4X1
g4UxefiEjtcP/uJclySVfqh8KSm9ulnbQtM7HkFTovwpk5v/iHnuW2EVZTWxRESyxzwi+9ExLzGd
kW/ebDNsPaNqTcXO35v7Kv8oLD1tagQHnk7/0BeVUci0X+LyJ4GpDqYmehoVvBOa2siqEAMojQlB
hJzz9wiVjOBFsTW77HKLzvdiPjAwGYt4/nFfw87/cdd/B6SEY9rRXhZe4fkz4bek219dxnZa0Oth
6nwHXNNO8RSvDGfy/vGOaa2DJbG43PGJCRNvsJRksr5pGaWrZEniLlCdTPwtxvUoTmoGHiLBO24J
9v67EbN+mjcZIBxWyRCj3xTFx8+405CNIvxZIkxdWGDgx9c8sWHrrNI4ybbjTBNsOB+TLzD6osod
VY4DfhCH9ZOTiEkaL1Ddj2NizlXpRCYNAAc/ou3xqNG68kiGYoDYOdd9Onp7wWsLxhpUiQ5vk/Ib
xy3YyzAkqZ2YwEGJIDHqSCTlbzSkOnoNnU9FwXBmm0AG+CQjo/masLxo5qY46JuP2Gu4uEaHQmDT
RJA9kDcNeXZtSt/jp/mnLzr15hegzjPswcUrMXWRWmLyTOd/yLWYWnh5GNNzIvGb3Icw9UV9zI+7
f7RgYmFHLjBnFq+Xm/5/PKuWQV3XIr0SadqK9RPnxQ3WgxBsVGKz86OLIgctKZfvAaIhW+VdMAMB
oH3OzLDNqMNYmj6ITqzcS8JL/fW0MKZbD6e4Ud8n5jPL0ULekaKt2uasIf8XJ70JZLmTT3Ox2BZn
ESnf5hl5JdEQm0zeiS1QpmBy1txH7rrExcW35k1lT5o+6EUfGpGySDNce8gJD7KT+FlACvf2Gq5j
Z1wk35P3RCSs08ay1urQNozUsmErLEU0mgEcSKUnSNH8aCz58rEbHI3fyOvnPpp9eBzwc8G3gL7f
3R5vHEFXnFaTLow69yDRqWqZQ59t5zPO3Lqhtsc1udMRRKiJsx6mRceVD/PHVX9SruTBArmjiaXW
BG8JMWMhrXiRf+7N1XvRIk2V0T06p8GWAunudcqjiUcvZ6wfyJWnZKNHAb423sh/J6uXZ+srSGpN
+0mj5jvz26uX2kJFSJtQyPtalhDdZ1qtRnBA/Y/V/KsVxmQXyxMLNylzwWsQ1Y7i5nP2Px1yoyPP
KaHhUGntDJn82jDDzLxRhu4qWIYDYJWgX5yg8jnLzBKvXSME4RUssVjqIIvGI1GE03kVWrqKmZIx
ZBUEsYUliSFmrt99UOGOwOi3OqdrX+pPnjII0iog+Cc6AP1UXTZfaafWXJXbyCqpJ754dCklMC8c
i3QfH7Kh1Pk93fHGiSHgkWyHWQtVsHzyZkb7FgTxv5cBLEwKwyYyEVPfRqIbN7i2I6HSAVRgLU3Z
JB4Cs95ooCsECZh2fpGnM/GEaWbMzPM22FjkMB/u8jrg2relo/uggZDK2PfjPiPS52jKiTLSNDbZ
JNoG/HFqmlVvfwKyVr7bsbCV3zP8JFxPaB5aa0PvhnJXp7YS4jFJkHzeR8PxAMzQsXmXyTI8GME1
v6VBbYDqJNTFj7t+cHWfdnzzmf/DXs43MsbeGQPyNjnEXlXKApGA44Pf4rLPV0dJR8wHoKOWrT70
m3/mKuBYJVcJNuiFxKxT91LncUGUPY9Dre/lzvBJEyY2VlG/dho9nlqY7ky4Sbni9EMFma1DRcbf
YtEqTcIKbZlNFTAKpZdxkFI+BWsOWDmQDHPc/hNOk0Ij08uVUWqAQqnpJZ1n2atg7OcNPrcPZ7v2
U+8V+mDgVi9uI5IWqGMHF9phAruLxhev6nT8lWgqicEaC6oRe6SJeLOeGCsu6gbGoUSE91upScg9
0JMHArVOnnOAop1OK82U2RDhfE0r/KeGWXLXKwDVdVBrmOv2zHTJj/Mm5fbfWojxFDGR0b3iBNDd
UuMn7HlweBiBZYsRLALyaCiNMtiMDjnccIy/XWy0hZq3+i3jh5XcbQ8IJVgn0uqvrEgGdbO2kSem
8OqxXxMGPZL6UfWymSFH4scAkHK0YvCmMktbx+6/2riC/97Dj78O5IeRFPBL5giMOxZUVFYrHXR+
VgkKPLPUlTaKgUFNuEjkkJbi+Sn9X3yDSwVCI8196bg3roTIt8NiOaYlmaZ1piUGu3ZJu76un8yw
ynCYdIIZd1Q929ATASAeArk7xl0iI0QYs2K2ByU82MK2WLUr+M6l1uwF6k9MGi5CCm60Z9WubGxk
oa1lXbevlnxcJa1TDxOkpt4RCPJwigcaC1kCiHl9NkygDc8Igku5axK+9BoCagL3YhjhoO7l3WaP
GCQa3dO3qJdhTuwF3w2BmqZMlTasOsy+U+7BWV74i7uB/o+qV+AWIz/ChKVyMaqgNj4Xf1kQMU8o
7V1yRfzJevcXOSs/UdQlQRA66uJUO3ZspsuJ/9CZ0UwEgGY0bf1J4ZVciwUx2ox/5UXPz809DTNZ
EMTyMu/6fWWrO+tfdOtyQUwcD9ZrCy/IDbWPvyvX1yjAGsQi3PfomWUpyHf1cNn3aubh9FfHRxzH
9qb3zvoaoUZzQxdZEW+ijA6fhU1P0j4NA2zm1hAB18tTZ32q8q+o9A8E6rsALc+YSN06HYaJHlo1
NxY8MOC0H0gLdqHdLfsZ9X7xTTzrJKpBSJESORe8pL/RciQx0a3Kb9AIyLzUDTTz5LAaoTwWQsMW
WNxmwqJpTnTWtCY2g8TbP8Ye9YyLslSjBAznz61EpBARyab1XqyC7vOkARslG27tYb6SPN1bdeWz
pvSFM1t1qk0fUaw8eHSCtPQD8lmvV9AnMaO2s7TSONN9Yy15MYddg3zUa+4SrKynLDUB4+84nQOs
cVLZ4f52bJS2b+mSTV7PMwGLLv3+XobSkdStHvud2gmPcdfMi9NYP7TE02iDZmU+SxxbXNijxxrm
Fe30UF+aVr00HHeQFxtuCRmqLenbhT46KtvqfStXS73lXCulCMQuu/9D/GiO+LX7KPYj+6dr/lHI
EzPuJU5fYXNjVGQhM5XEjL7eAvXbGdcbKdRffk9mcKgqX9+Y+LoBFAKBvTaXNx5ySONAH9xX7vKR
ZlF2442wNRMCMatdj8KXqtOXSRA2EF9jeIpvjPH+TNhd5kvq5mmKZcflvKg6PtUoU6q2+uXCgjUU
MSywnPSpwwj54vK1UcCeBEz6qaL6HGo3U1QYsNc3ZqRq60dOk0StbHXe9s4u2O/FEbzyLG+VKVX+
OVu7aUetoTNeX6h3O2MF7C+Csz8Brf+rHPt/R4x2WExKcRDVTN6nNaqFM6BCz3wYYtfN/31792ow
PzMjV84wQ9KDwl+UIWuToz8tfvqN2j15Few98caGPuLICEdhzZX4veVAlBX6hjrlZ7vba5gZr+ES
orIqs1NKSHHg/FxqyEnpdWGzF6Q7E4PcPY4XL6fy1Rv5oks3nL+XqgNC5+NTTKou8+NCgOTyKvru
BZGLa7oiZqD/wFT5c0TU2kAzreTNtLaQDjzjK52ln7txjvkGhVEN6QsIrz4PDBVoTnKpFJ/Jhk2Y
4W/xn2Z/tGDNxR3u3Ps/YeMMhlHzyGdwBbb7Gq9Fq7jivhGCffNQsneYBI82j+3d4+1mDESP92/j
tpytqGq91DMXFtwAqcfgqoFKBxJosE9lsQDNJxR+c5lUGAIqsa9eCEG9x7cMn+JYxM7+edIaEclK
GknlM+dBZ4Y2s3YAaDN3CbtXQqcZU1RzzsCqNlOkwbr840WY7/FORbTM83rj8d/J5S8ANNA2FQY4
zpnhNIYVg1tHyuwLN3zgSqAGP6mvwdzr+ogeym6I0wYJt2fJA6Xba2DG5a0JlRcTa7zWkIpFLdfq
9kfiQm1JiotGGI8+NNTPTdiRCvlY80gLOTrfevuqszS6cKLzk4lTYpVx5vp9z5cCBM+wsFzQNziH
CeFuHe+TTMz6fd5mm6Zzujv0um7GlK+niBqBTyY0Xln/zB4eE7O5g+tBe7jcGGhQa0QEDoEaMsB3
d0ycdvJ2VGlTkFv7nqc29Mrz8e3WLxUS4oDqgDy/Ceuo0Yc3mVF8IhzE3J/YZOMoTNWm6pvHJdTS
dTxT57WdGqgcA0Cd/2zmofVvbCAsZP4+4pLtGwrWpzUw6Z0uYyjfxHSlZv/IAOPtOFLHGqDdqdO5
oslpjiPJwSu2J71kT+N1Le1kcire76fNWUW1biqvOztT49rA7hGozTPlsR5RjA96E6iYr+GJPlYA
CALa22KX+pMeMn2UtBSuDD8ggFXafv/8KJg+BnFGVgqQBKOOaOQVP08MQmTDvlXat4jadS37tXYr
51VcWSg6aka08yU0x5j/iXTvm/6LNuSckzXCtKRIQMEqW4oZanFbpXDOuZgAySarhF+HeIRz9A4s
qGfOgBhL0VPfOQXgXp5soGu7AspVOYgYr2adX6VnPx2zKagbbxVH02h4spRejEjGgqdWP8eojrYi
8joWwb9DPOs1Zl7xj3dyDwseZ2ggzovrhfEqddBZ3H/1G1emRqqjBfOynIO+dHC59wHICYoH+T7Q
DyKi69PKigz9MqO2DBOB7rhpKUBWDrF8Q9FCsoDeJk03DsO0PW3lX14y9TE7FXds5jIOxQRWeIrx
tcRCOYHReHS7lbExn4qahveNVD/aQIBsCLkp8zYEXznPfTHRN3XMrAWd16o1PL2rupfEi9r/752U
OJsAnTiMFTtWuc8q324l18p9gT+/Bpyaahq09v70KmC5+jLKUHkj769DEq537mzze0NUjpLR3S//
06AY/uDDO33HWWYayEU45O3esfLdGdRbEwu4eZzBErUFo6LL8vddeId++h/q/sg5+gHTyLhjsvbk
m8xgPlZCqnlvPtw9H+BsXH8kL1jHEqnvtiibo5ME6ILghCIwTWRsnFBlekS/Fuh25Gq5drzJvuM5
W+jeUR3hsKm78hyaWJ5UBwGb1avDPVgT9GrACiT/84WbVQNc9bq6L8B5ruHNWvpEHft+akITcp6x
s5eiavfFJKSxm5o6JVQeeKSirmkijoiOVNV71S5lKR48QxfvdSaf8rxuv6SLKq3x5AMcuBGi0lKX
ynsSrShzJU8W9FZTCPvmUIFpOd8B8a5BcqV5hq43arVE0XJXcx/5u5lMSnoKc53WaFOBtiKE/q30
WOOTcFFhZA9l9kcb6uotdQ7OMOwAcOrtsTD9PzJcK8+U0dkEh8hBLPClzcX3OBHnC0Sf0PFdYXXF
5WxE8SoLkJXv0pamlI0iqGltUzPwQCgZ/8sNoKPZSnkR7RIPWA14cMQbfk+DRlL7ru9FPh8MIj4f
i3XMYcmYwelsDzMMqnPMmo88dhOW5Z4X+wPcit20zUvHpDQGjCrqTWYWjw3HFwSJwA2BBDvDEZjf
QiFp+SQTQgny3Y+44JIbNhslJ964rxr6as2tU0s/Aenx9huu0nLRAQzEhnRxp9Ems3lEjmbzTh4l
c3hubnx5O1KQ3Yj9PcxRoncHgreLR4d3jxGfQ8c8TEA60pNqvQRVnO1Vsjr+5H+hV+HskJGvF37B
1tAdCd5PRF8Sipg7ykiL8QbPHIIEcLEIjoK+c8RnnmK4u/tSdqoFBKXjRrRDRQIl5pnlC5yXWkO9
f1qLCXzDrou/AKdFTBj/oRoAJVcMsJD5KbKkPxH6SY1oDM++L2UrdEXD47GKWp9MgS2Vt/EHkcQv
7tjKnNP/+WlUWx2r+o3ygGH/y2AKpMafEzPgPUyPLCC/7W5O0sVXFDZFCgqB2upBEqw9H0hbP89D
sg3+YAVZQ+K0C+5y9WSSJdI9N+1gbEMgrA8MW71Zus46BB+E8RIb6u7ecP0Q//zO+zrjI2xSEQpY
aaJbontx1Qzg4vGU/gnrwz5DXZcmrZSc3CwzWzIL74gWtMrw4ZXvL8g3+iJqvXazcmlqZ3RDg2xt
ZZgwMOut2dYuYDuQ0cz9ckJv4wtouLLmFmC7tZhcNbIT/nFY4DPEYmKASJrIWf+4nXttnG65GRyQ
tgz97Z1szLyuA4UGJ+e2++rh6/ZlQ7DrbaWwgHW89Kv52TAtqyUPDJWjAJZ1/rGmH07UPkfca39y
y2V9n9yqRIMhdxrJpkPj2PmZLvCvi4mcPgz2wVVwyj8APzRERLwJI3tDCIObQsfKsdmbGvp1QpGN
IGTFPrWqlwm/MnXHDPytsCSNj8XjHzZk4TtyjkWWJl3RPnzxU1mKHg/77MQ0jIsrpEBrG7aRFJJx
uxnQH7DX+4J906/8F3qdZMk98hEjHF41jpKlshr/qIKwiuRTZ7Ax/M5rZ4OPUjPoIaMsBfUgfvH2
TeMf5ln7Cr6XPWH4cFQ5utvMN5Ore61vpxFUsuwSjQyAcp1zPpp3bFA5coQEBtdwpEeR9YlPxbCi
Ekh1WVltxtcVdNk+Pnxnjs/jhlufq0J4Oi4xMnOp4wf9dKgzo41b50faDRZ0xGMsMGXF5AbT8DJa
TQx5ltE3u05+5TYIaonjd0WAGOv4+9JoVuifR/M7F3JKvwvyhEA/kei/AQhdQVvKRUItuWTgo5N7
PMHZI4DIgvDwxv+/bIaOU+BB+cwRcbJ/TbDnls4VCYg6DTkN61v2oS6C3PmbS2y5g+iMfQQJ49q0
TyuUoPEI8SF/aD1Q9B5mCdiT6eT/WeeF8BDZbl6vZMLolzyVsNPfGxBjpkj1GCn4hdKbrhN5UN6R
frhZXYmSI8IR7MC972De7Mcu9PuOFRvhwiMjtUMScroG1VWj6yTKrobHaSKkOVYeQiogBilvh3jD
Rb9GaaV+OH0EOVrKfcQnHOmKLtFlD7Uw8e0QQmWLuFmOcUZ7Yv4IwQXE3KoZ1cb9sLbYgaAJ/RYz
rff0Qr3Z9r2aBsEs2CJr7OvrxyaQ9XIOUeJ2qWcf3sYnXEIsUWFmxETpUyzt6cJeT56QzLghXcJi
xRqs+zEpSDiJnP1DDw2hR5X50Yh6J+O6KAazBhYPnr7sK97i+Olda3y4qCWzmxIzUeeOjyerkJ4+
MxtQvkIIDYhhzlQSLE0rDU3mBApAEYf9jVLwT0cPjH1tWQqopTBDR+6pjXfJcZkhbcbaICURSs1F
h/lNPEXsajuKdxyW2jxLeU3zSgBRMDbJbhrphEYPJlv0Wb+SbUVhbIiY8W5vegPgTLgTNaT65hgw
/lQcfck1ZNOXAn7CSbvauzKkrvWdTzDJ8zGFn7W+LLWosNWAz+kWe+Cp6REWIgi/cPmSLPSVek4i
k9ZyvreQm82VWs7mW+IFcFFlFPjCC27DjZ3hR1E2xRTdxwpcRjC9SEOt4JyFnI6gZD8Dt4yh87zL
8A2g7Mdiu99AOzFWEZbm4Mqt6s4rP7+Ta7hvTU232o3WROmLRaOZyhfn2S+dYyn0cvMly6qArnvg
XhLvGfhE/KbE72Qq/E2tLMK21/sOIMLJ7+hRrGiMZKaKOQJFENlLxZNV/geSudssnfZX8JbTKwXS
L/p/rCh4cZuiki/aqnoY3vGPa2H7Ei0FIHLWf23qmwtk9LuADo6+rFfvx7dLeZP5HRjhOMKkzv/C
TlV6NbIemafN7CDSTPVcRFL8aKzHs8UT9JcHgyTKamfLWmgBq6rf5UtbCdl6J6uraWOcZ19JvFMj
GXv4RbnKryq+lsTtMdT8P940bD15qUGzBZ/pesWNJeGf3jJykvLt8AacilqnmURWup3IzuPTOvQH
RuYGhD68p9iZOWvXS0224apgPM5G25VZMBqvlIkKh79uSYATqAwBdKAvRd45xs/mge71oUBlbzOR
Pp5UdwreTEWLOHoCgvz/AXFxtTha8+QjjgimZsXevGuQN8MjwrZ3HkgQLdAISYhs1yPbUu4JSCjK
AbRj/7iqP+BMSPGjcTQFLqbhlIxk+cnzXOKimfI2ld/zYPfw8QpcvgYlUTpNSBDlml6e2w5DdZtY
JkHzVSMnCDCFsjAHmZI14nLCjG0mSUbYQ3jKctYMH3Oojt6miiK/gn55roigxNgW92B1qxmWWay1
eoHmlbwlWmkopkFhynG7aq5pZ3dYrDb6UqwTagQ2yFl3r2e0B7a57uP1v6CThKaPRT1aYWVgAF5o
KD1U9bAkBRS5Omz/6xUlL7OnbIne14Q5mRDnw7Am35xJt3eCGykLc2L5EKyhtDCWuK/hOvnSF4VH
pO4zMxVnA9nSsRSlgFYS7IlEaqhulLoGl6d9SQbLoTo0rCFxICkpwSLfjpqvLaEZ0NoOwjVNbxt7
/xQh11dxUlFihK5CMD7LyNJQjRqEIkvqlFs8QEYS6SUW35pe2O1YQGMFiAGfjtbLHrb9eWyq99jn
MAfgXUDZkl3IMR8kcZtDm7uVEnV4shzr0LWNQnCYfGNCFM8KIZcuXAvNwzTXgM9tjlfg+godbRPY
tvXJy+AZI+WhRO+DZAXDzg3EOarjIPDASgbATV/j9dSTLPG8rrVK79ZYQgq34fAd8+livZbzEQUE
X4Im4j0trW2LWgA1q4phy7aC/ogjBxHEGSbmXeP4BPRfcJ/cIZReJaTN1LnhppA4UxCH/vPFBj49
tmolrIwGvPW5NUNCsTDcL25BY7nUpDoBtjEPyT8kVAarvi7rsgeMW2KNvj9DyL3SG1INDc3mZfmg
XvGb31h4jAflF9td24NNhh2anaZ0l+m7sQt1NS+ZsmmacNnfln6Z0eh0qkRKsN6DGAZglmMfN8Ui
OruTvvNdOmapvaq/+k7Sd73fWEX7Ytd5IVkmMeA8f7MvO5oSlE3VH0vCOJBC050DEMXJnpI6JgF5
zIHw+dTjIZpRbvarchJjmLAAwCQSzER84/ZxxdpxoKElqN9DvVc9v3Xm2Qn6hbeYt+ZMyA4i08G5
bZlMDHgDtqIcJ/EQ6cignr4kTXcTkTTCOBNpRilkwcJWDwpMdJE457YmShmaWbwkFAnvOOgrHLPD
PIwYLLWMyJw4W+T5Xo4ZA9C6h5w/ZqzrywzhMxJJ3+I+QBStW5dIeTtZr40d1q7EenO3GdZ506tT
FLCzNAKe9DBdNvuM7NKd3vl/AA1BwIK1vbacp1EGUK0pp5Rg5MJfj5GpWsoqeqkGlkFhruUMxBpv
Cl1sFY+3clR4N39DqQd1YAvEPU8fOOs0vErmxQqvlnrjKZ+RhHDcK95HEVguHLBxJ3ZeM2EiJcqA
RAHJ1BUg9+iHjGQVLKXwlMm8OG4w04y1OC6OlI1++TBozKO6LbNPB89PxE3CWhQiQEPlQopP/1UV
pToOmH9sJfE8oaOoQjtxJaiKOAKfpLYNQMdz0bAmdbVNh5DOOXlGZGLCmnV6FGqTaW55EQCwe3tc
zFbwieFjTJvCO2XRxUTndgqyMr7m/V+fQAJu9ygnFUoG9x27d6rPWNwdJgIK6gKuFYiyvyNReKpO
fAXH+OnIjeIKx7nDj/etC3+e1RUeaykKbUW8f/Jrj+7booLjyk2T17Z1N4W4BTQmTjA0o1PME6L2
rUEKpyV9EZU/esInCEo+pdmkbhZ5NLiMQWfzPmZouEGZEz7xXT5PlzCpRVzJaU0clBT1+a5YE1zM
HHXhBci/h8RYMPVrANfG5Zl8iw2UXcrusS/JSCS5p3XsZ4KHTosmbCxMNpYm/aYyQUGV//r75rtG
3OPtWmsyS8e99jglrDjDhav/PliZI8v4Au6PP0ubRRipSyCRgu6TjWbxbfo1SYNgWxObQOi/xgqv
ltzG2XwPFb0KP7rIZ4hx5T+C4oT1z7HmgOQ86kIy+cyD/tGCVYxLswPug5exRiXFwLh1Y2k/NtaW
UHfAEIrIBhtIhI92w1bBEMf2kNzK+D3BlUTuqCYFrRPwI2O6HXErEQ30kEbWBAahc1zBzx5bDIwA
lqfqxsAS4dcI/4KKupdFDGqVEP5Dh5FQBLKzJvR5x9OrwXuwe3xR8Y/fkwLIqYk0XOKZGzpMtfEe
mg/LJWeD22C6+spDiY8hGauF2h4b0IM1g/WggzxAYfamvYOdGbPFp3TaxOPLqvdpPj4je8ZcvFhu
+TJHh7rsWNA982QfqW50buZ6XMlWbE4ojDD+tyqI322//WoHiKAWt3FuR8JTvjr2N7w6BopjPn8g
6K/eeqQ5xi+ibnnU1QbY6am/oj28hd+0Iwut5MwQz3kwDSXVMQa3sI4REZRLjQFdnep90JhXMH4u
Ewubie7NsEqrtS7Msrq9Tjntnb+Xk+8Zk2f2S6EXyi+0vJzZrww6XB7xJdchgwXK2b20zvE0VXxy
BDXhiboCMPJCubQFwx5s7I9gWFoXiUlImkukwmf8UCyIqR2mkEX9DwIK39zfB5okgVGzoWEgPmMm
klIHR97M5xSd2jMaGDcONGE+TvBzxmQI+rPbcq2rVs8QPhSDEc1YuEEszen7bl5uELhPS3hC16Bp
I39WGjs15tXRS4GbUFpoj6aYdVKv9BZ5viSDGP/7iiM2z2Q8lxw5343k9M8CCqV01eNoyePue8tU
qHwKPOpnmagHTDjk7Ih4s99TeWdb4c981r0SK/RC1Ph/lExI5rc6EW6TSOOq7+K6r41rcw+5laNj
r2eyHcR6Q99Zz5WvgB/Mt/bQLVBPN92zYIJjeDK8K/Ziw1ROAM0L+8kGScAD4M5FbpBXYDstGxwp
N1V9Q8QKzBHOfTM/0bH8DQKGckVxnU1Mex49aczWrlDlCp3WllxBtk+Wg33uIQIT4VZHD4sqq/+7
23uj3+/Nw+uR58ldCxJrbiXCJAB13ra0evHPFje5GV+DwlQSykNabE2UlzhWtWpgrE7fy0LyigJn
moZ3L9EgkBjS0WUTERvkMBRmxRc6SnDpLu4v9mPZN2xybo7j43wn5gv1KpDwG1iNmo8S3b6+iBLc
8S42Jz1tMOY2lS7lghCzXMMxISUidn1QsRobJ3XsaQ70mkXDPMug7ygL1LVsKkuXN81yDgqX0gQs
Sud7op6UdtRzZUZZqkKVJ3T0I0nBpiJa5dWvPM5/9KAt+sYzsB/HdLahtr3Ho3Oj/f1ErDqLJaGc
bF7OWoi7hj3RTyP5tdI54oChO/Udw+WiwrVwYZ4yjoD+X1DqlJLhh077HR/2G3DfL4OhqaDdN38F
4eT419UOGEFwprljioLdBGfJ3wZc8qTYAnsX3XFG2TYjCYD46bE3EKVMeyStX+PPaeqJqZddtJKc
VP5ABZxJK/sKPz+7a7uGVtJBr9h8grk/yXXHZ1K/H9730qRr0MB+s4kFynWDO+mV0toTlzNpEcEE
lj63LHZVepPOsC8lhwHDqo37R/4FUk270tD6lykKXQ6gbIEU/dJ6TJTqsNmo+mQ/IDInz0bHSErx
Oqx8tXHniIp2UtvFnRAQdChh28bRj0miyjAT9TWTp4a41sAIiwvj5Om2mRtGQYv7ZcBfPZcwOyw+
tBl/vH49BeWtdqSDxnPR7aJg+fkhHdbIqHRMXLEnFkcKCoiTxCa3bHRLav0OoD2BwlGiuuvpbPXf
ZuQca0be/jhegqSH9yMvTbpddup2DfB8iLnsmpNc88mJwVjgwvsasoBP+V53Yzu61mXmWnpAXBMF
jqradJdO9viz+NSMGqf/D7Mkk6F4mF19ah2FEwJCejBfVkGx6DzhfTHl7+xk9RBiKKK4Y4lGDBDz
fT4VtSkm7DOUL+dCW2oCPuEde/nu9RKUI5UvCKIHrSftxqOBBSPGwdk+uEdVLuS9usKZ90WuG2D/
jsZmqqLAQ/p4myYgrJGdtajUsggaWBePFsx6YsDK7xS/KRZGcV+P2tIOhjUBFahzQrkQneYFYmvG
TRJ0rSzkHltrbJr6ZOoL+J3eZQPPak5BE1TKmxfaPy46VA7ewAcK63dFibiBbLGRb++bEFIaDlRn
R7JwXGs0wOVcwzBRrY3PTOzJRmBBYZLqdlzzNe10P1xkRMYCVKLtbfp87BvIlrql93HHiid5W8Wy
BxsbjQHdyOmwCy2p/iCCqVwBWifozW6LV9Y6k+Uu4iFaLqNRsQRuknt2c16d0jr98ZdUG6VdYexO
xhPsJzmxr8I9H8ftBE3CtgiomF/ewCncje6WVfan+/ZaFuErS6bb3sVuoHNolJrF/K1HbTyCl7Gv
y5PbU0I7xNRTYDRPENmKgtBO24Wgb7NjiFGg5rdny+Ig0i/rRmOj0bOK/ItKAph7R6YgMLfwwnSk
/kLoHHKeTwEZNvdEkDvOktBCcjRY0wge3gzEt9KchgadmdHGXc0VsjRq73SWFk+ULVxlB7thILH+
l3XVxdf56Rb9LTUwXNiM+CoaYVurcoK7PXUxHdamDWuo82P9aBRynvvJk5jX37vnSLQZQjlKIylp
9oM54anYX9TR3WQpU3FgrdIW0l3XniGWa7K9eirUKG8qrYx1bFz2MTOgqs28mnYepqw2GUWJdEJ5
qZ1f7DNP11bCGtgv3aJuXBIgGpz04knXZnLy6/7EEdQC3cZjPqWYSzYzawzj0MKkCiHCAUfhRDE8
F+F1SZ2S7KEZ/9+tZFePMOIFgFY0IAz0wOMHuK9DpnzhMo+HMJsOl7PkQj+I5evoWKGVUZqsjoZS
wfWwCgjb/pQH0uxMWNS/SsCCVJV9j7KLVX88M076trMOPQ21DB4DkraGu3ByKK2oY+CB3OdDQCUC
cMa43XfKIaoMJNa9b3lvybbW4tFTYzORMxN9DKFbCfylj0tchlsFIzi8p1qO/myAhxs1OrsK0BDh
jr5h59+l11G3lBqSjIyCBcWLHH49HMCU2r4dFliwquYuSLAXtp/tky+KElJelLaU+ZY7klg5bXQH
cqxEePIJYAljX+q6CF3SIa5pZ7+jDAmoV4+L/ECVL/xKh6dqNnJPL48gpnDy4ksdyQH4ytKS6ZmT
jEj2rpyVI2QjAk4SYgBr9FR9CuC/2caEE1V9FZAcEiY+l/hJMoz9FmH5AvsEvdOeFi1hF+sC9bfB
IoKGaVRwnoMA+/FxTCukRKg6pzjytpvKXqv3YhvvCjExXSpK9o3ljiqBoq4SXUPTOaisd3Swe6/L
LpOxP++yDxxCwxXnX9dVt1JzOvLbTWiuHz3ogIejCaWksEFZB9AWDMnIrVQ0zmNYvOrZYfIcGFeR
tNQ526V0Ozq2jnIRNsUigRIqphbwBwjJ1OpBGQm8xUXXBC3sguzT310tikk/NqZEbN9eLB0vg66+
8j/0s4mTRFrr4PobaBPGc7aOie1FvVoRIQvXFGLexZQ3ZSWsWyFUhA8Mf8SxEbxrrjdQyWQ53ciC
H0DRG07kCJ15419hLcF6MwZQGd+tHIYuKuGoaBLIrYINIp/k0J1VAKQkZqRUk8p4D03q6AQTBuhK
VLVC98PpPQJFfLtC+kbsAcCOJTLFVoHqRFAfAVRC/BeRTssvO3lsRN7Jw6jYjYysW3VkuIRquMJ1
MzYIcSt3NfZZ4wIMj2kypsJzO5X2+NtXySl9MRXiQJySiF7TnLGBk9FmV53Sl1/ltnUoJ4HRvxmj
0nLuIxTEl5vZNJdrN5CamX3c91EAj6emm3AJlQouMHce/8rrdrk98PbNv1Si4Xvu6M3j1CZF3oH/
jA0+Z2y/cSdcz5YKXoDKNJKDk+EIKcFOExhscvNnDYGL5EdioGeaFRJWqCln0IJUphhXmPq9J0du
O5bjcPYmvk8AbDET+OEcbm542VBIHq2zNOX10gqNbKl1ZrnQ7Q84sh5FNikinCfqEoMM/bEemFdh
jNiwxAb6j4cWMUVe+dnirQ7oHLemk5TPHAYn71fnaunFxzkPPnQzVFS7/e6xF0ftJYPkJzLpH7Mb
eR9TqW9cjNfCQ5wLImwAPrngDqOzJK4OfpRNb0nGkO7croppg9bhR798IJ46fbkdvhNIV+yAnxIu
avgevQoN/wCWdVJ6FqW9t2Nl3ywAMUs3P0PblhvzhfOQU1IJ2VKwL4hChuMPlBUBooPtcsSy523N
uFJC14fjSYkCbmgjIzK48hTQBTpm51yLAPp0QsIVwBEhuXSq1iCXph6anmnhJZig2tvdCFQpsfir
9GOVwJmqmHtvhIBUlh99IqbYolED7IDWv6IK/onOx7BhZ9OLKHeO1tSeYPajB9GlUNo2r1tEXcJl
GCoItMNyHMZGew9hVloZmMUsuwdBQs0wiDs3+NEVpCYnzJuV4peDUTRGm52M3S7cAkPublMKjV7X
EaSRZ/InJwp8R71YbqYo/La8++Yn39GDPeCqpAFq76UamVycpGCLToVvbOAejPGtSB4gf7dae+RS
hV2NUxoaQHjXjx+Vtfz11fjNvIatQrTGxlRL73UJU34l78F/fVEYa6cM+uN342HT/ujPQTtSRfV4
fzkOhwX+2+2ZFLulp1Udim3G/YdQyE/usfQp519dDBcYkC7K47bheol21LnZoGsKgE7qB8MVTuxw
OETFUpZmWeO04c05G2kL88aEpyoGGx+dvAQkWIguHm4R0pxvC+HRfjI7bF0woH4Nt0f4asQkdHov
UYpX8cdOJGpTPPC7FbHElGYkiR0ZMHOICHrntwyi/XMjAfwraHgvibWKMgqd0ngF6Pnr9uSk54u9
bum7PGFUlb4ag/Kc/TD6DAKhq6xKIcY9+dqsSyKbgVcMQGYk7E9mwhb+Kc77V/cxvTkSuDHQ07Xg
Zsv6PUcZpTW+ebZm2NAAGbi4nTcHmtiVSBcZ7ESw2seDLjRdD/IhQC6CvoNyIRNGP03wYyEij1Gb
aw2yEmFtGQSEkHJhGKdYFUTthYS116IfA95JbRrfv5OfaHH7Y23EN8dcwJHwYmkoiG+6sZcaS2aA
q4QD4HkRqkIor4Gjk8s/m8feiRPM8nTuRV2qcuPRvfpefi7kp7lfrfy44Anew0y3Mvq09KSM4DFy
5JoCQTayM3jIlsNKhRnlu2d3Jbv7unYvmnOP2PzA3hwBJgeTU1BA5yNipLneyOfzOjcPbu1XUinp
/mICa/5WA/QxhIvotxC21njKoo/RguJ4yNDeqzAMv2BejWBHvvo4ssXlgwXg0ZOkLl1PsJJ4HEar
ib7V7V/W/ZVuILvD5Qn8/b/gg8an7aLBAvVBTyNxDfhRoQylyoMd9yj+NeSd4zYVyTlacaoRMok5
1RH6ZTBDv+WizgExeKLxlNVctSSedMwV5uIJb3QwN8+7/+w9JVP4LUC0MYYvUI2ZEkKJfH452sU4
Tf341iRXwrCof412BurvTkU1DdgMMMflgzdWq9ccd63mq+e6MOZDjsn6vkcZ/bPzVE9uvozsMJdT
K8EIzSJWUyEkdFjuNdlyZUNY9BIlHzJXUcspfdrgMqrLUH2r1oV+aunLZYFJMBOamROzfs8vLnpo
mCwv4Dyqxb2bab+gVwytuaBioeb8MO3d3CyinVFYVzavju+qIum6zZFuZmbdqvb8rfDUl+w8/mJx
lGGbtR8Eep73o8Jo2i5cyi9Iq5psOUk2bnrImqY+HXDztDwGJ0/6MoLZUpvSeOWD+z1cyj8o0GTU
dHMTUcNxYKvieKfJybUddWtrpiYkkyf2NdftVdQyBiBd4taEWeiY+ZVcaRwNvdIR/0ahnTat/5N5
ikHpE5S4KDdv0DDwPCVljZXesjyiYKpkZF7OQQbFOwVKEXXtQZjsmrk8FIcsILXNO8c59nSBAwDm
KlPh/Jn13G1JGVfiZPxyE3lz3REGNiMIIEEyXIpyMaXvr/qyFilxKYpXFncVwpzayYba5qVeKHfm
/RnIjGXuPm0UyAOx+hylDMMS6kwmguA78brE/EWSi8EevpWZ1I4Le1UbXuQbFOWZbahtEcP3QXxO
SHzlV83bsojMadRv/dRy0t7r9E9AT86veDbJp4EUMKaItMMt9bwpg9FKUhGDymQStFOXjhPmFBVd
JnwLjDpWzEEWv49lV4Q/mTIROAIYINcKtaizICDyozleHEI6FpvobgxlkRj8UqSkSIAQX85usmGZ
yBEK24TPyn6V4ZD/AVwWvwlCoAK3M6J14wfZj8NnHFdQ3IFzdrRQl4Ny9vYH9Y+Jn23o0NPpdfOG
RAmSv30yWRcj+KG3/DNfbkq3+AEckjGTpZa2f4renQrxjl7/QknhipH3q4bS31Ao3NO+nBMeww1B
1xclI1kgg5+aYa8BJ+sun2hxrGOOqpGMYDWY7LeUr3mg/Cd/mRpLiCStJWTjR/gM6v0xT5HHLK0m
D/aHQvHpilwYPD4Zuh1cvoLxXBcn842DbbFd9oryrb6N7hJyrAwx6dR33QaPkUZx8okLZkBk53D6
q6Aod/qypZLd2feAo0hhOx8MMONqQdmuKhy1t98zoF4CAncb6+LRH+HLQvA0BpNEylwWiCvKY4ws
Ntybu/qRXhSey736GxYmPqR9u/Xew/W8zQh4ySuajAm4AX6KCfyo7tlReoReOi26uwpgWYfi+M0t
Bc6f7p8x01CHlI5fhxUsfNpweJulrr1m5CR5CAD5rBOMxRr11R+9NwRI17DV6lPQZwR+wxVLqSMu
sekBNwtXt6IrGTPSFSdbWpnRa5zmfVwpwsCrszgO2Id8gcITfen+NugPAFOFPSrkEavtqq7yQJPG
mZVIRwWdar8wwtW12ZuxUWYrNDY6MuC+hDwGIHVi5UGTtlbVx+nXRCKAWXuKoxEL8feQNz52zZhp
+YtzzooDldMNF+Syng0CrQEqwwHTFp0irvVgl4YMqSSBHKhVbItu34mzZ5o6AQctGSmV2/ScCeiY
/MERwsltpYKn3yUKUYFY3BP9g6nh/0NEMRta9FRJPwRJ6VKpcaqldJJynLIRyt6yMF6pRdp/ykZC
866XeVam73dTUEn9LO3A5sEVNLcjCu/XCuAet1kOPvgL8WpJJ31K1FzY6VJuWLzJwU/G8/VNpBL8
99Ch64qJShLkRAzuFbB7K/nGZ4OzyKRNoD1vrSDxc4FJZ0BwYOBGXhK9VFdu80PkrrMO1atQ8WWm
VVuajfSr8cpXqN0YLuybTkmgq4mOqKmh/ozj14kyo7NK6GthXi3yENDXgX6ff5opDFYbLy5SEhyh
FWGTJgM/lyIii6SyrDaCwO1m0G8bxkVn4d/jfX4d8FZFDK3JU0t9coGtLVwSJgZh+R90cah62OiE
w8bNsfWMIfidfcYiAUXgG4TJda/Cq0Td5pnhv63HooWbp+BVnxQu4huYdfo6VS7hRSyecLG+HsYH
qc+6jrWjngHDchQI1KaHp2iexOgAHU6EwmAcQDYVfBnfIjFBxrVMHXAknnoYAxYWxVngEuHxBg00
Lu/SJS121TOJ6lBVe7Cg2Vy/LFn4H9cU1KjPxuGx3OhnUHtlp8qWEDcqntR+w8t3t7ipMQpugecf
ms7xewfs79+pCtbZqXxzsQStrtq/V9NamOOV9RGiCf5HdmIyHoTX5wXM/TfFAoXLEJsTUeH0ixru
1uoJ6tom5J242rjm0WhSi1NPX2WDVJq2+AOZZ4VMKlKBmTqxPoWQbD/XZ/ib2lVwLMg1gG2WC+1p
PBqCClE1aIzuP/xauMeErSHiUFn9lYWUVDdb5Exu2/DfJR5mHW/67N0NPEYwDpmwRBhumlV9JWVG
RDP3mGKIjpfS4FRZlg/Djkn802kW8Cg/Xta/2W+0XPiil4LXp/RhkAHBo9aXScZf5ioaOXhs/CUJ
MwtWzw1eYoGSaDCAvLHMxnaDXOSSEXPBOM8mO76CIKtDIC7b7waCsERC1R30kQWrjcjQBezZi55C
vF8u9mHqwAkl4SZqmFuattRWOx2FBanlDsuHYc7it2yXlvrTjSVr0dJwazA3NaS8gFmLcXgnIicU
lUT/U8//gpN/sS6tSgPIo88lD8ze6DjnUuMa5HPBsZ9mwaDSqSQgW8FvaAPbxaKQRzFYcRotEJ8N
EiPS3FqBpImc1Faa5sB9WDN5H+WXEpOJraW6mhhZfP3ukTXXOiJWwoc1NnJrLz+nqhafAkQxlfyp
FWYd/zRPV16iRn0vLkyg2yqPl2ri4aKFobEB412L5oEiECH36PiiJVrRxSRjERJBhVP+s4E3/DPl
wGTAF3dmWBo5woEKHoum8I3dTJv1bINoysAxpKlCQsLjnK5MGqA3WOhpljLm9rVae657GQ7n9b+i
PZTuFPfXthvBtOGBpvbK+sa2xmnluydjfXhAGClM95oHvXZil86To0TKd+JLfDsY9WF5DQnF5dF4
Wwll70hEMoqD46RrucJOWH55VTxEFU+QiT+6HYXj0ZUwx2kashKELPiDtruLIt5asEnC/G/xwRfV
f0GoeNpOBDsoW4yqsKpnc4dVelxwr5Mglbw4RIhN1+X4R0BwOyYpCN1YtZ18ptGmU1TOxzpBGLsk
szZUhZnLr+VBxtN1ghKA0YeSTfndRN6fMF9cuIcpMaVCDPzBqdxVCi8ZQcJeXkKhxnqeO4A8SS/Q
1tP39g+b3bELQEQc2GcQ2SO+Ij2bp/gCqYmY29KDF7rpVznns6NTP48cc2Cc9lYWSBJ8GMq/LxwU
bHljikxb5oclqVn9rrDgzYALGQ1ZDd1TCmeW1FPYbomz0wsC1uExSrnZfYcEQF3kjETatHZwILKG
oFHrApt2FUOfU3FXnLGUOdGmunj6C6dje1amNx8DXcvQWD2x4AUPKGxqqvdyrHvMWbqcSV4AgwoY
kwUfC+HDAhuF8AZWI70WXDHBLEZPkCuwijph+OrNbgLRBKAeCRSb+KMYo/hvkJBFH66J1DNuzBJ3
SW7PaWEW557qsakNkUfqbKZfiXOBsJukrGz+piiskw46i91EayeMxh6a8x3XireJlVfqoQzoHUoM
hGOTJ4Q8is9dZInVU+x0TFx5ImMOkwGFikPHhv0PdWaaCH1ecyM6iykvXhkfmK3TDSVpHm0i4aqC
4BuD4nGmR/igngoMk6DNmXGEzM5Au99r0PMvzci2kcBMGByAegXnjZ7uxVqLMo4ySkHXyqJ6hGk/
8zKOWFm7kVF4SjJ4xyfRpQPzxVuilaQ/aN+hk0LuxIxzOKGOmjl6dG07umitSFqf2PS2nyUS7iGK
9dH6i78SQ2JKSivfklpj7lw/S6TpJczCMp5rY+ODhJ9TZo9YRuAH/RLECcik0VjLvscxYIosTiPH
OVp+ifA9cgR27MDvYlaF4OZOt296QUhsEvJx7F6+AItKjTHZx2I9EyLK+5J9vWBB/kAwXTk298IQ
HgdBSrG1LhMMmoXmiBAdFMbQpuWtnY2K0TttVgmv5H0NplxzWic4uoc0P5MnD4/JuD8TNABaQ+Uq
tF44V+lzk/Yve1ticsnMzGd+6Wm7PJOuHngpbZAFhEbzpUOT2mIePUDA/V4K4x5b16y5G09pDgsP
keewMjDVp4XmEmOSAsTpLojtV8tBkbo/F+En93FZVdJ8A1HRIIlJMYFfwFCnzjN4Vuk/cX77bCgD
tmR2CGr5zY0TKfVfIuiuUY8k+OIV0Ojg0qztNMNjBxGxSZp5mwPJ9Kb5JSqyK0yzPns/O8MMGKyP
UJrozw05WXIaHlHOlTiV+P3cEHLLNMBhnrZTWFtgwe+hYjkz0xb7syo/er/LA+5MumNk0f7gTKg0
TNVoWbHcudFIi8QJ17y41/MTTn7+7c8YMURVUV7DyjjeIpnGA6Tqz5nsW/fSFpwoPezGmDVzs9ql
BShojG03G6ACULkknRx4PwzHmLzO0Qf4e6f5ugn898usRZe7PRCFvsbfIp07faZvI/O0smmdeBPM
XCIgm4CgAtbQJXHmRFyd7eHcFYu14oQsEVrWiPH4nBkkbCzZjL6wng94Z7zP3kYrLHz5FLpNtO7B
+GF43dM0bDiW9a7JOB1EONwPRA1qc7r9e+QWSPaNh+sdJ9MEPzY7KBKLVfUpsXYohhFmJYGg7sZK
+3C8cHzWzim0CCUt6G9nVq6SVx8/j4kaAgxnY6o+9nnnXwhTUNTz+yYasKnAWLmBCU5402cXxZ0I
VWlwsSuBAkFK4IUvmbUFrtuqDFILvqAs3cDi4R0Mwwlb0S/tBQkpC/1NcoDIhV8wC/Xa2PWfu0GR
Z6veTBUGsG+D/kYJVEfnmB2+rz2C1ZgRZtZGiBV+95yO1fhtDs6gMoBQmOoVxsJ0c896JtXYa7gV
bUf9+LC2Xmkd13vJrD7/oHg992sMlQ7L1TUdWHnXoGc+Qj5E2G/M5luj8JJ7u3bkJLtKYugcAQbz
o2D+8UId7hz3WN0EtoI+f13lwGGOlxk03+cSZ9pgyP43iFAiFgrhxgYNXpRt/w6R/V3IsXJ/95Fs
D7x3VHCmySAvdmKswukmU29svlClrq4GaKYpCNuLn9Ubi0cEetNZX3GbGmuSckQA1szt1f2hPI+A
n5T4dNNnrfxAZfxQ8WOkbUBMh6Ogbu9XvJIKkvteKreUfbk7jrUbciIez2rVnjIZH/sAwAPL5iDS
6el8VAx0pUirJjiINmceQnZMA5Yw18rzf5elwAa4BQeyolBgwveCtmvZy7M4VSW6aDJwSqarZtyn
qFwZnZo2bUZGSMqwI8qIck1r4Y3xQ4EJ2+nFpGDOi+R8rvWn1HUWG4zCm48alxQqfw05f5eHjcp7
0iWKnwaEKoO17a/wVC5XgB7mRII7hrvyfbeKE4V6e8JQdihbLZYLkgNJtMoc5j8OBhD1klMEzQez
4ScPrrw4pTdG1BbFWxbpWgN+fHILYt+QrHdtIq5J/rx78QZJd9AMUXLWbT/8kQu7jmwXPIVPZ9gW
Ks7kp1uJppzoZS9HzogPa05tMb7qek6F1abgj/+wcnJ6T14bOq2TK7MXhXHp+n0ZIY3l7aVkS+e1
ZG5sosZP6qK3Au91/Bcg+4zPXWB/Dmqi2BcgOzM98cH37c2yiz56oOVfsw3WFMY0USaEe/FPYizn
nP70rqtF1ch9laBD299TyUv4BCi31sEpyT5Y1HHi10YmS0g2kOE3lBd351wlB0yqeBmHXVxfnagw
6sen/3bqHAnqqiXZ4akzuBBMOn1Z8xTfrMd0yvVZS5lSVMdD2Qf1t//fdO4SmCdxTOvPCKQ93KJ8
iPzD2d8Egzyoil6MvMZxPU3XZ2gZDbip4njb/myRrWCBmUmgH9IGt7c2860kyd54Z76feyQkXlFo
jjCAdoB56XYVT2JUjVHtb0DlgOY0uWCHUcgI5e7XSWqF2YTjV7eDHCJOA550m6mVmWi1ejQcA3z0
UvlA//auvsGyu02YhdhoE53fvyoevGqBh0VaEz4DR8LyY+AQH2E/yivYyHTaPjs+QWOieTRH2gnf
+iIOtwlisz9A/FsxzQ4h29kAqgKNuKs9NqBeZoyZEYHl5Ivg0Zp8qukA1hZXCj6z8+YSWavVLvjK
q0PCUYbAEI/uhU6h5AuIhsoNlqhQLf8OZDJLSj0q6T8PLVIDbq2W1ZHehUXU/7MePQYo1gjothb5
TIRZ2Lhb6rV28317WJ7Mpzg369lcdFufkLvDZcvZtT3KkecPw5fQIiNn+Q7+luUPWyehXPXdjJ2W
JRSYuadhx8WrZ4Mbt6y7nfl5dY0NgwLXF4ihv9JYuBiDN+1SxalKatjzdrxvL4QDPiKkonRdOiDo
5XNCVf6aUhLq0Y10K4w/wkacJeiE3yw3w7fs+tLg8lvHhgBBZhn2hvyng0jYw7b45NzGULrsEn/+
3awV+bnnGiXBrEiBx1lAqPTv0+nepSc3AOYJ0h3g+uOgLJfMPtTmoIT+lxoibyq777fJak106EQ6
2aiQYc8p225N1ETzOEk2rgn89e1wcRkf0w4aQzGJQsd1+8XpJI2lLCezFzApUxzSBC/M76I0YIhR
SIA9kcSG2OJgHeEx1WgNHvGVvlcOVMmGANtVQAUwZo7Rk0mCwXV+ZzRkV1IQkSXcMnYaiUVb6DmC
nfWX8lmBhNek/oBIvDxmll4bUEKt6NxRsnzL6G/QdZxz2A7Ctv0tshuhRGoNQukMLVWlJa0CuArW
PvhbY1Njod1jqji1cHqViUPfeLv3+Wxx1frsakUJG+/rx51sEa2V3FfBUzKmKer1sKtUBIHyFRnd
KgmUVBtEsC5G+fC253HIiH52PNo84Tgbvtoj5jipoiCNk/z6AUcsbI0gnECw5OSUZrOzFzRWLvRZ
JMGE4cTSO32NJmgVT9xYCzR4uemm4M/swvuGrg04a3X/79NDmqLlxXWXj20BOu/qg+AEtLdNvBhn
ALnKynxmAu2cju/9pjpBLU3RE9aaH27Hpm16wgM0rMIvx/h2Vsa+k/W/X1kvq2SP73+gAij3QqZJ
zmbNqTm3+6eJ24MbesJBv/3VXJfCQJhrpPKdWhXFaXaSOngU1wJnBVx8pqUqTLNOWZWDO9YuGcgA
7JYGOmRrMeLrmDRB9UYk8kNoPEtawujV/f8P/gCPgxoxhhVfsz/SO4Y7LgXXG9kKJg7abgp/vDxG
TES8vH093LFc9T6IFc8x3b3PaM+/E5ZwPfs/6uZ5riCllYORQNgQHvkLMUjbhfryd7knd5ozXAxH
rZV2e/uo+Zp4rgkwvK16PGEMBnqO+BR8b0J2zas37wJgcIyeEQI4uEnTCNq8EBYf4RdjJjNr5qn9
kgun08K37tl+Gt+w6J1qHqR/Zf7wgcPRD+owLe4Ghgg0+P7Gq9n4c8OujH77DnGJxg+un0uWPxDD
uRHGjkjaRIYfQS+bhjZZZsw5MHQ8rT+rmHa83Gv3Nxn1V+Haq94ax8GqjAFMAtzNTB78QNN/OT1w
A8OjQFrJGBgP2sN9apfkRTEnwZz58vmKfJWss5IvKuxD4UeYMnMR9AsMAwhv5SVHN5f45SU++tPx
6c3lVdGDw6QtI32G4k68uykzbKk+3nY0K0lnDjxkaI/6MBKU0loJa8ey0fyQnPk5HEzpZZ73TT8j
33dGox2UKUrVIIdwlkVRyAVykdGRje3GUgw3UywRkA+J7UD5W/XgVzJSPVDbWM62Bd17fMeBMP+o
BTmGoZxCAzZh7NWz5veoKN4NWP3jeiuX74rdzooBG2nYK2MgVE6ZPFJ3OXVxikyq/Gm6cKdSxrD0
YEh1y9BHlZ36oXexjQRC3BLziz9im6LhmWJgHHqrAGgAq4lKSVbqxLpiaDu9P89XUQydJ23ZNpQD
TsLiB1BoVR+ScBWF/xe2fj36iPKsenX/KAhWEtCS+mf22CtFzRcUDFDtnUlQyiN7ySv9ytauxWEs
4HIN+6g+6zBDwEXh5NRibHdm8l3eKnFIE/djhBQoeXVgxKX7JJ0shwsDAqA7d40J4/oGh8CfMbtA
xfLdl+E+oNVRApPTAcOd+S8byRhfgf/WbweZqa5K0HZrNIYoHQrsHYAf0aovsENyCj9ctwwH1LAG
SokxD7vlE26O+Fs1b9usZbHmYGvZ7yNext80np5CqItmCnsrvUpQJl/z6FZmNG05et/EM2AI/yUu
wYsfl82FCtzDyLOSzT4rgei76OAEf6BruLlcZJONGqEpVzzlRH6odxoy+TOl9NucfDezJ8DyXX8D
SLWYugczUrEqxnuUDJWH/LiBI2ITpq6xTN9s+TOBX648PzONlt/tmqNkjTSNbntEnLj4aPIP82IX
GrpsFloLtoEIYkSuN+P3dZWtVrKGsACRhJ5k7VynBWB7gPFVW1E5J+mxghX0NuCuqWSMRRvkzlXN
9v7ut8v+qgUMba24CucOpZkTeakjg5shlYU/rlqBc69oc3/5Tk4kbp3Z+uyWMA2sx78P/4Cnw31T
gjtJ2mOQHg4LTDFI25iSE4LZaGZ44/EROFoNulu3DVCdH7rIsii1J+yA1lf1ZgiHY+zI6nymYpZI
URcO8iWjuZDq8MxjcWIVf8pyTh5urBA6bvUjw7ui80oURJ43SHhgofOSRz6nJ4S2LcbUNoucdw17
aRAovyKHwtCJmjSCkqfUHN9YxIsSdWGcfKsez0RBpGCe/SyKXBbiXzrIyf2e4SZ2GqgBwIS9a/32
YqfhQLDMcPRiCmjeTUdA7/QKsQ5mnwMYs7KeqN7JIrRrX+FeH3HPdbvo3KN6M+eG/iATj4l0pkQS
YwlPb/NMNaZUGkHTBoudQGgIqF8kHbwyq+A/SVk+jI0EYMI6tcTPLJKqhEvvqAJW750C7nN/tVqS
9ff/J7gAu94vdQ566vQgvsSrVQ6OY0HXWUR/yEG5LmFlN/nZY5A3xZLVXMKLq0Ym8dodHRYIyxWD
nzwetQNS/FdKcV/L3MU64dSFAUAHPiNYnWeAXukVssaeP/6M02Ux9iHsVvBlx0t4Kg7WEYcCCREe
XWkgGw6eiLI/QEk/Kzr3foytKRhJcbRWdewt0vlq61JIe0xBoB+LF58CF2yXrYOj9Vm2B6UUmgym
xik+g70cSQiMjhMMRBulP77z3MIDVCtCiFNWdB01wW5A5hzI90Tr+np3+f8wVE3NplMyaILmVp6n
FPFd6VvGNT2r1ZwzLIikYkoZPS5UfMidVtzdEeknSqI/Erjolvv6pPcuFAx2Bti1lJSntTKqi9vt
w5mSEAvlYWpUFGDd9hmlVMdcMLg/ooFL7cXBhBY3AXDFZlRJlhRPYqedPWv8WYBkFc4Y37VaT21p
VIE5+m6t8gOe+Ns0U6lLBaIVo2ZjLCiMENhp/gYbk+1TI69wjjapww9uT4hBwS84VeTs74egQABU
wYL2+Zul/f1dMxmAP0b9JzsKtJ9IQJlKIgfnhnnE3HG4wh+gsyX9kLE623xRRlLjQnjysAMKRlwa
5SIxlqRVJ/yMQNCgth7J1qfLneURHOa2pBXWqQBF9Xck5qsyW4cmskXlCBQqOcAiAiLOJeqFA5ce
IJF+q5WuTOOhbYSEs3mieqluBKjbQj+/fZ5uFI0wBlv9E4yJhegzNjZMqWzyQPjmoimnhh5Eeiku
PXRrXWBWVQg+j1JBdxZWi82ODKC27AEgu6tnUblxDwfV6OIfM+WvQMa0VrcD3AVQ5gLBsggs2wXc
eyDqnAtzZVS9PArujK7M0ZNvemNi+cXkV153qwv4+gU9+GkqSmW8uU74WDW7hA2zhRYtImfB7pe3
elMlKFX1v2GesA1IMbJloZK48J7pxGS24pBX4b743hjOFzZlAp3XCy9AdD8j3Fxw0mBq4EnCZNnj
j/SHj5ZrxBXaAJqIJBD2Uv7BDbleK5FJz/f+5jL3elOihewrFet4RkdW+k5I2CPfUmQvkMV9nBM0
Z6AdaiOoSN9290/K07Cvr7GDFW+wx5LKe0Y7xk5FYczkFgJTczGG0Qqe1JBJMJ+X7hgqhEYB0nGE
007wkHLH1G6uQvmtbBuOLEUkvucLuZAtEpSUxJBM4Mx5sW6ilyrut6XS9HZ6l8qEYiFzM/0UEt13
lv6XfT3rq27FT0yGl09nHjrqbHRflNqaEYfWcutjmXVWwlB3dJCxr8zBRPtC2gHyIMNc2N5td1mi
fZPadPol1ToKk3O+2Sco504G9BsUIveVY141wyx2ZveeNO+OaYDAI9u/sgWVul7bpfkdez65lgGq
WoJm5/7oEqTngPXOSICGPlVQYer8k01BwWTo00NLy3Ilqcco3nvbLU65JkiKCul3aTgwKCerFePv
Qslde7Dw8/28BA3CtOjCQpKWJ/irMlum/1o+M0n14KcrxSO+pIEREV4rhsyIvj8+0cgZwLvxbiqK
mIV6HSrkfbsW3Y1eEgn+FtZM8/PB9VsaeLI1gySeMaRke7Hkq9WF/83yYz4S+bbpRe7EA8bW1PEX
ZfZRtZ9zBmxF1uKJp/fikYFa5mVs4KkmVzUejaleaYOQ1nmqX5IoxGRW7pQeLRpwJuFoejEqOiNY
tIe2zv5AJjHF9mkVefNCfdl9Nz6fS1rVECAo9PCa73YMezyonSHrNN8gOhfbekOILjCul0homRV3
o4FtXe6N/66JICWrjm9JNF0fzw40mEAWeKFOZMRa2SRJZXtKsd2PbT/RLhJqOsJtLCwzs9gQGCyB
TIMqfcJ1XB2unvHSGZotrfQstE3hDcLBj0KkSi0sYVXV9Qo7uerFmiI7xxuPZgOKEW379Wqjs21J
BcX2v4EexwyS3LJ9KhsAVMQYeKNSfK9Q8zqs/aMVXtIiTWck5CjC1dlysI9CNOn1IPmdm/jBFwB1
CzweumPmARLRHg92KpOG9MogNhDaHzS/R6zhqTs4AL1+tqqezyvww9u/KRgZmbSEDPPojOErMA12
9Mlzj4GYpuqvW0ZhgBac6xKTPiSPxuQsrtw+01SO7dg6EdQ7eRLmgS5uE7Vq70b9ZnPDaNPrFAcw
aGm//qE0Tj5VNUohzvXeaLT4NPzZG7C+c6mF8ivBIKag7tolGTG+RX2Ux9iRpZk3QRCWmR3XMK8u
DuWVjbCg2Mz+Tvj1ZeMsV3nmE/pAtWMvQhcbPwdoCTrBcE/3pvi564amAMgddZvKxtqJIxlBuhGK
+tqaM9Xmz8qYk9rlg+ZmyIWaEj/zStS1NPUFTH2yvHRMP8vxXtR2Hp2+ag6YC9RVyMrkd1zXxbst
sbgOvh0iVDY1HwkGCh6IFXa1gMmPJMW3MKL34HRSUWbOUtxHuPp6LA2V8IrcS0XzMduBHo/AEgaU
1ax3AUqLoe5EolPB/4ZLBLu/z6FMAQzPDoBzYhnErviTxfNPglKhLJD+1vfffOlOIpXHCigo7OcH
H2Guxte5kbTzNpV28GdFoB9gJFxXFEmfHtcFesydHyezCqJP1c/YtO0ChPyUErl6C4i4hGqwRkB2
/hsiSSfCYQGZPWZs3ISVOQixR6D98kdMyJbQ3k36F+FXIpRLqJipEf0ZDpRG0dGciB1NGxJAXvMf
jpS+8T4HkRJv+NGlsqK2cOJTz66O52jvXA35yVFGOaC93gAXxNoAeBQ67ha80GkxRRtL5qb2E6At
Fl0in17o6G2TKddS2fCR/U5nfnVnvYh+/kPqByZgJF7p2QJm8eKiRjc0kQCTGut/tZ8WG33eKuh1
162I+ugcn9p0RS5OMkXXlgjD2C61SU3Ht0aCf6owXyj0sLqbkF82el2vRLMYFNmd+6Hz9Qj+BWNN
RTMsu2us3vbJ2d6TEdBC1xp46fo5Guru/90AqUT/OG4we/r6DRM+7SFKN5F4Wwb7d32QDwgXCkTv
zhHVOjoxgThHe0EkVrPkgA9K8G8uu4Px/TLQVYH1e1869nEHHtri63LT2+rFE/Yo5sq1G9dueDIF
K6GBh4s73G8VNb1b2VQsMKodwJEHMdz3mpdUOEIv+qf+0V1W3j/cHEJpa2/e4h8Ea9AcjXraIgmN
9wampfpMDcbtnpr2tIwnZrwSuTU9+5x9IUpEPKbty81dtI/duFIubbK4IJOnQMaI3HACDe23KkWE
aP4jwcfyMXuOvFyU1NeQgCdxTFKElHIqB5L9LsL1Dlv12YkEE5vHkXr/B1xygxuyMp9b5l8Xk/8B
1kJzAIcGRo7Uc24chZ6wGulSC6IRRU+uQN3ulgxDIBVCx+RR6i35xhW5U/BXzcTuZZz2xQFve0ag
vO+PobKIFRDvdy//4l/jTbdoWWsnY/fVhOXb4/pQmHKL+3sL1ugKmlBNNqY9OLw+cJfziDBLa681
pF5joEB6bvzOBKQtD14SKNT8J11CuJ0sYQHzjUTxDiD5bYk/L10AryeQl59/6hRn1V1Xk0k0JWDe
WWRXu0JbBh1cVqf7YKInubjX7+KEq2NgZE+9Jpqcd0X8OnKG4yhlVwFQEHrqoP6hyy4TDGHVGw+q
vMdS7s0V1IIfGSbRklq5l8WfVlHfDdgBqaiWvlInpwrdkGyYJ/L7RXVwO6TyEltrI8XoP8tAfmm/
odLSFAOLqRaxRgu9WvjPtf4Wk2uJnDQpk19BXuyR5fIPGyjmSzMpMAmZ7KgFeWEroT5Ia+CKbXD3
bVXcJO27BrzRUXKBoZJOmLMpqUf8rHRKtbitNIk607VsJUzH2Fais794HPl4hneKCCfdbJhphoEH
AxFiHDIHU9lOnerF21EMaBIBynQSm2y8qfZ+TfBRn+AbE1Q1DOqNAE+H4/Pds0XsRGFXADVTe/X/
v/+3Yw6V7OFVIupooVGDkrG5x1EbmyrZqO4RTk8Mu8XXpt2REC4V28Qyt5l0NApaTYfIkAjxPr3K
4xkeKC3mGuF8FPdG8O9zYJesPNnMRi1Zg6TKmcnurGSf/BbXL9XnbmmZCejoMSErqSJsX3vtfKFm
utZPGPyEbDpU1FeKAJIYABfPM0Y2ZzjVoafSdz9FpAWt3NIzVDuokQeQ8aPTO57vixg7g0I/4bP3
myoKe/F79uCtZK4btDWU+FnqVAUuUIJj3AGfASTiTDZrKXBEjsN/CudXC2G93CMuflRuglc0rS+F
CW7Mzm030RGw90ngkeImvP/EY990EhrdGbkxk7C9Wu8R7GxBPSgTXOKjA+bomsb3FRXOu5BRHZ1W
gLoywGxVK+orEA9dF5sFaTlCMIlWa13tXmjg33xR8w2HEUV58WvYwetLrmFvozB5go+jhWEoj80p
BPf0KUgnYQPKKRMteVU/OzLtERxbgqCDUy71RK1xd3cz0HwMnsbdK16uwflmHs0VDQQpht9L6g5g
1NKIZsdTpLSNYYDnmNOD+/vGxOBAupS3kg5YksoLj1YjVAua707Sgd4Nuct6YvQyfnZ/pAn50ISu
xl/X6XLumnTq+7LTv6N01XGh3pUn2du7tZtvo52z8MLJY71aZbD4J33+QUXeiVfPonLNvBF/yLii
3dOegz60WxtJi0OREG6L/pQuKCjXEBrInd64unrzJk5FQS7G39FGWU+JILCLfjM2VVLFQPvkD3Sl
EVM1Mha3GWVFiuV5V4O17SwA3ZWzuslLGwNhqNLoHcYIs2wz8zYC6L4E/U64tXC8ug+NghP4DvW0
I6+p4/dn6p4zPA7yu/UP0A+j0ru1t9V8vRBeI+yqj/1qtmv4UNZjI4ixbbivuqfjF53fSbW4MWU0
o/GUEi1TPeFuYB7BW8fdyD+hGv+pk9889BjTQjVjYchBbbJbzmKhVo7vEWcoItyzP4yKJoaSWd9b
1Lb9k2J4jlpXctR2cS8o5DKgkFtUrhk5S72NGWB+JevEEnnYZIGvKtlxVOGWPoJqCxyh9wmOE+9k
/PF12GnVsEwxgCqumNQDHW/+x6jNsxU2pyy+FD+1O3ITqHfxDgvFOLBzPtVHRoyHAbEOwCCil3m+
iwEbemnJbRZjMokujP/OyIQ2z4UOhsDppu1fqxvUGTcU5zLniq7b5nTRPqRgnLFu++1h8K61LxjL
Yss4ckAMEUFQxZW9CI8iB4/NrTIIvB07PPtNJdMei0cRXm8396DAbG5tkG1UfvIboy5ExxlnSTv9
dSDn7pV5e0UBj0dv/tKHG0QeqNQZfjKRh2n/8MgYoA8oshDodQOxD/D4Tj/f4N+HGRpmNFXquqnu
lhyjmwMWJHi6UeAeZqOagJs0r7ArqQi4q8+Yfmi9xyg43zhJHaBw9u7V0n2lMn1T3ug66lJeeNpb
fDLsoBkEQbo8DRNvSOK+gRDN1eKDx8b5o3QRkf3aHKX1NbXZzUOQdOSYKgflPS5+vfORyNZArzLN
WPaeQocazcgsk5DUXiUKrUVg9T+vUb7U0MEyHb4HuqPPIKiBXQAVe/BY07YGKo5iPV3svrKkovK/
WLNgxLkPqzfnibb3yiE2AeiPRdNcQBMaa3uf+8lQTMNhkD63j84ZvjC/FaprI9sI84jPdZDMQkxF
KbkmsvdKhR9qBkIeZgePiBT5vNIkNua479YyKuaBqK81Ez6MzN8PASqPXZcXW8lmFeybRghiMRVj
uV9S10VZJzQTOnatNbkdaP5QOLLnb255cbtcarEmWaoak7dwzCwDpjc02+cLKtwkmxSrGxn9ExRK
k0CZRLO4hJnxpN7Cl0Hl1++ec26AFWiavq8RRJx/6dZ+rIKzW0UEPOf7BdPne2JSBxgCWor0ZklO
JugWqs2D42ZCknNU3Dx+hCpDzH4A+4ZJbhKbYFI0NvrWfZLe3WgEmaD3Y4FlfKsPpzQRwjeMBgql
zgMxy0LJOvrEculmVdQ1QMTAICwKeco5q1INwbkbNl4pWwB6HpXKqmfigTrrbQSOLnDuEuiQYb6V
Y9R7IYMqvrbrWUu4sZcF0s/DwgdI2qO6sq1pIccqXLivFhS0oYrWUdP1P2pVGZc2x/OWRI4GVhrE
IsxTvYU8BKAG870W5Ka2c8xyJssYLLBPfxFYDXkIH9dMRooHM3RkIbEA3WMoYu2QN8pfegPAlbkS
oLGLy0RKeWff+J/pc0uf1eDfVySMO7c4WH37xFH4CrNAIxGzqPEyS3Im9oLS04whq97pp/Qz1xlu
CU5WHK1bCn2KgC2kidnpkv7PoLiRHwCe1GzcOvOvmEjy3+6IXq6aAQshJZ7ynZZmEeUSmZhP+8m6
pWemrsPPxa+DwNhGL3S2VZqZV0czhmvlk6rZzikkc04axz2So0TmYwUqM/xUk2/TiAgA2lxnXc4x
MAwWOPf5aWuameZQPH0J0j8mnPaTZCMc+XnuGWCOrTsVv67YPRsrVHrYjXbz3D4gbbBOIt73l2bI
oMTUJYyeLx8SnhisLQHDqdHKsvupz7wgzhRtIPeDV5HQy2TQa3bLUuTpnh05mm8v4vwFJavx2Mqb
N3GW567Iv5/K/Nkh3VxxtgKi+sWxUCcybthOyVkRA3Mfp26rKNXZAfPl8z1UfkhrVQdm1E6GYFy0
1DsDUWarIllCXubL9xdabBFCjLObOcNkfbLS7LESRMr/kF0v+yH22bMR4w5xrpx2P4F2YCJectCK
ViunTtXUi22gMSJJlh+0T9un1a+/DqyLMrBsrGB1vuDiEyn58L1rTFqreuw147iYUpoiKcYwdUv1
QXSrQyTCMAOON6AL7Bn1yKpbLht+xcEHM9IiSy0YdU/uiwJ++MdT4vNRrxVzGrqnWctPAskEIAUh
uF0S375R//eMkGT0IhEc3fXBfmcbqUJayGwxJ87YetMeNoNpV5gmiFkh+QBENbaDPUhDOmgurVr0
4o51Lywl9CattQB6bFi7NvtJR45WKvmuRuxhnTn2f/z9BMZQPWNgwhmo4V7P74Dic7FmXpE5U6Td
B+8QFmK3iAG+WUMJjhDYjBjBncL3LJlkWfAZqBfemB1oLZTfigGDj/dUDFuSzwNBKVPGw+4RPlKq
i/IRtnLCmrb9w2oFj1sHw5mr3q6iCl2TID+7z3cJjg+lJ1HKowzu0y4cJve5fh3a7rG3olWkLKv8
4btgVZJc0sZUyMEN1NdbDoa2ubdPagrGhZv4bBJzCoYF6vk/IUDLOZe6MNlYD+1G8dYBBVW5Oa64
PDGiNhQBKME5cnkH7bdiglclZAEX/KDJ63BmrC7bqDyK5Bcmvl6QZAlUtyFFLrOwUSIZElKWXMKs
Ht6dsh9byD9QfiZ0Xm3DqBvr830Cg4CyOk30ynoUdn+NExQMWxk6iyb7uhFltZkVmydchEV1qCWg
jJBOia/FY5I8WmqMoVmcC08pfblYJCmY+aBfH8Xdl/hc5/0eMCsEyvXJTje+pzOgOFhtkh3xUiWQ
zb5Ev2n933nAdUphdaFuwEhmkGS6VGpSVKWQ1SpWoTMJXF8T2cROwJXW05W6BUmG9c+1lgla3uAJ
/Tw29Mt+XfuJm2ORa+/jwqkYAGC1y1RsQ26RDak+JXNCVQ9s26aZrb7gzXkcSBOLQGmnksA30FUN
z3KggJ5sRraZAeick+/WVSFbf+WXbxkvkcdiSWqxOgYI7g+C8N16FumJQTda03byCMTrLXnSxiYl
4DC4DuDqj1nXzwU09RXHFQiqR8uikEiaNvE/N604J8gPU4r+RWNP2xdz96p9HJOZKh2iP+5RMgQz
44UX5AqSkpJ1uffIYYRFVDf1FrXjh5wcnJCnrE6TZvDSDjh8NhkO6KF9hQXC8j+4vD1AcbNtSlH0
K33WinTY1pLN6uwiPjyUN30YRAvlMMX7Mvl/GawABzu4adM631am0hFFlHqO0ygEcsWogx3Ircxn
xSF6zOfRvHDhh+5m9jdn2zL7LLrLl2MlOjjpyvvQgS6OXBPQVE9bQqY5L3tnwCD2iQXJK3GEYvPV
S/6E609eHvNmEs2Q5OL6U6F9fVvbnNlNvEwaq/AwE8FsPXyY3r1EEbUS4oTmRUCZNPgeWwpjaUuj
TDqVs/c0nGoj7OBL1h3a+jCLCKOViRzF4oXTOacRCMGUNmOkIdBsqyjnv7F2P0TJoz1qYrSKnTmn
6+1eY8nAFMmDfMjNopD9dB8pbR5xmjknJZ5QCN9qX6LULwwfRqqQ3m1dwcjvUuYsVSMOiZNVOn2q
ZjrU7olBdhRzHXmcDBlV5ZaVqx5AH4sKgZkRLI/+nAWviIYfYD/6A886W2zEQq1vQ5AbXIDIsYXp
1KxUoFSj9efUC5HMalNezb49JNemSj3SE1Y0wYr8rKN9IVIKF1gCY6f04bjTHcB2Oi1uTp0xdeZR
mWRjzGaLOCGjs+lq4GSL+gELNBs72CgVzgtIKWxCFuhQO/ciNyz04VPI+UIAr/Kpcs5iPn0dGePi
+p0z9LzvkVC+jkWAkrn1Q87DlYjBHbhVwgc2mGBXdenkqVuF/Ep4Eke5OPISGNCddFEoLwXe9gmb
+Rew1/kJOUVTEX8kyx6U4eVtqKrF+laAEDqm/EDixzdo5nL/pipBwJPd/vtXVQq6IdF5yqzKHzcd
koItDMLRc1UOf52B/d82+T02IMT33JyYL2qsCuyWwAR4LKiLzb2Sf8E+8HyCvT6xNa7bDHCrJmFH
51xIffn9ykhn6u3Oly45HgVLufpCgedhCl7hRNdWRC5YkgluP0wfDn+pYCPjAnOtCnurAQbDI1/9
vx3SXPduWDcW3szKMN2F2ceLY5H9L/LlPeTTAtO7AJQuFJkzHBSbjGEVEcbE/pbn1TIw2pXdv0Ac
oKx4eIh+MaZsQW3qTPSegbDUNgoKGJaiL2AC7WC1pwlSs1dX6m2i0HbJBqXE8mEVICb/BawQxSIr
1fRBWWhBDV/LeiT3NAXSrU5+v+2IFG8lH0TGX5gkMKbAU8Jq15E0do3+1CJgN/O8SaihwbzqoE0h
sOJdD83d592UABRQXbgTake4d57FqVo+SkLqra222JBvOdBjbHOhlK0ynFYk02n3KzM1MZZo6jBU
ToROAXSXbqvolQKGDrsvZqoj/dcvhwBtJalgSAP54kfQ2h5+Mnxy709EQnGwOziXuqgLW7c35Ma8
jhm4mEnPIZjJSyM+p6k6pq1lxXuoE8x7yYxTVO538yyWxo2h3hFrKyL4bG9dRV4UPS4Pk34EKsWK
q9h5n3e2q66Uxlabhu6TFsLO87pnL0D4qWWG9II66Z9CCTQDOJQkIuf2jZs8DA2DgkSY0dyKVGjJ
C4XOIMunxSrlYwPAnPll59LpqzZNNVgszxe3PZhLRR73u0NnLQ25wFtLIojIGXZQtkDOuMGRp6R3
FCpjuK4MxXRovKO+8y3mnv+LTAOMIiZft/PyEyqc/3s69QmLk6Kig5q68RmkT3Bla9KsXi3pN0uO
yn9dvUZIMrkiUmf5LuVDB2nlohnlElZavLsHT9xmns+Psa8xN3narbhfZE3wI2wvu0NFT9F5LKXL
ven6kvjCrw6fIDoM13P6TpLvYLbh2OO5MJsQyNDavKuSla9o9F5iTI7+aXZehwXP9Vc6ruDHyaxh
emphlJAqHs366SLFkHp6jv85rKgO/VxWAcuBM6DenYH1K3cpHJ4+2KOy/iQod38Lc3Md+WfifDQy
A/6xtRRqU6ZPiwDVvmhB3dPkMuVRTdt8rSMRGlvZFB0axk1hBVTJSFXmCk2o3mrzCjdqUjsw3XLx
A62Amx8taUSOTJi82e3AgHGKk7fFYzNSvL6KYHapJ8aJKPa3uGmbe4QApE/AIuQV3MjKpp2uXn6Y
MVps/ImRT6OFEFpUzTklPiccfT5PfCxAijEOm7Xrx5brfi0l5bMZiUmaN5/Q7BPTK8TqGDgZFpsU
e/DhQSloDNRVepsLBZ3ogdtK3QYa4SarB+gf7YMkLcOxYnlOTvbeztPi+8iywMntoFdL3iobwZob
C4JAZ7aWVnDXL9AZ1ZLkO8oXVwGRZH4bL9u/pk9UT7Sa2bXveL1ZxfngGKKvLSK2u6uwr5wNib4r
zKzXtLK39oGeAMqnk0kJI/BCa2gtdi3BP7oEIyCnROciwTAi902QPn0qrtogX6cyy/CADuwjWpfS
e7SczEx8tyGheqo6L3a2wKzTQflWSd3K47bGIr/p1oVMCR3DY85XFEhEHZf36HlaQC6PCRqlm0v6
U3OlibKPLNusSzX3PpcljuL7iaDJ2MQkz68C6QBdRr1bI8hyxj+Zm1yr2di1+Hy5M9oczlitneca
JfUH9VExnb9UO6aAutWKes7hD+RSH8Rht3fpiO8A5Lb9pm5WkDJc/0ZrZfJOhaMw54jdyIkILqkr
a/5JU11aYLtWlFFGmgibq2K3yseaHENvTLmVCw8YkFskdAQDHaGjhm+/0QgYOLl0kAOUV97S4b9R
fJ62ndhwJolAPhBb4F1SR1jXBe0z2d4MD1t8ufWeSJvXzWdQZoe7Si3bviCGvQMNoMaWVI29eDRA
41mpFIZ+2oKT0Q3p5dUWFyTJNSS1ot2tL1C+h/4gLlUsfj1kDt6UlB2NeQcT54iqU1KVA0e/dA/Q
J9Lgpi9NbB78KfXJtuKuCQ/bNwIq9vhf+h+M051wQ41cKaBFD+y0a5Pmva22Erii1DbSTsrbdhXJ
Wx+UX3dM1w/Q2rZ1zc01ZoLr22I7J4xwbVF/gFu0X/LhHdjEB9uL8PcQ0/JTI+6RKDfoHlzcMsU6
X+PtXvGYfC6RrNtSJZCzNKBT/AQ8LFGyfQIHBNziw0IIG9CPp3qEpMB8TgvTHl4tNRt5iRTd/f1G
ZK9+I8tM8374Xx5by3yrYECBRNoi13N9+v7NQSwQvutXBKT3i35IG5d0a96tnTRH+rN2p8d4ouom
8g1YnmRxMDioSu0ShEUNhFx9ZUoOoL9QVFUIFEiYYkd400ZwjiZdmbLs9pKyuc0qWslvF4wL0+CO
dvhODBKhzvkw62nsdjuNqyGj/QzU0W5VlnDkyB7sDK6tDLYC7/K05Ae8h6WkDxEDwTYkfnNekTkO
LdOR3Fic/EmI7VpPkdLU1YqjaLVyoltB/s/BiyBRPBRB9hxDfOOmik/el7L3SIfA3092s0WgxNKh
UP9N9L1p85qKr6TrIYJ/THa/YGcD04Uc6aKM25/vlT1oKC6ESK1vjLhPy59Tqci+8S8CuhFgqZpL
liMpl8XzxdL5snS8SRIJ2uMQvnuDsic5H/VjgL+l1GeWXM9QIFoBYi1mE4MICigtS4/fa1Lh3My8
czsGcie1PfLHzCSFWcpg37QpnVmwkkjE5cOrLXT19CwK9jtn8Bb4d1zJJ3hj7Y+OsiG1lBzO45rJ
M+Ih2T285kDJka82rek3sUGuyIddXYxi8jYY4V30+qkVEVSK9xJgRG+dCUC70mzjN0E2vYrEZql9
3j/KMp437xQ82GpHXK8OlazmH8bRZQba1Cv2kJzkGc+nXkB1ebb1Ptzoc4RVNxQQp0xmzW2UC4mc
wWcAqlrQSZFL0Sb3e1Mv64OakF8SOeV3lNV0noY/5aCg52oPKQnNdvjLwy2R5mp99RKh7kbnMKKF
GtqwtPqSS8NjCOwf9t5UOfm2BftgSomR/igXttddaWAry1NLS2svb5dZaanDc784d2MAMZ5Nn1L8
OgmrbXGX7+8PQB6OLdFgg30wINN8UxdHSs2eZ4tCqV4nV9hmxFE4OKHK7RtFt/h6voKuLx2ohoTr
9PK2L/t0SYDdFtfMLXcusBdOeM1dKBnKz+MD9DcM/QwYFYhS2mLZQwBndhHjE9ObhEMkSe4o5t9G
Bh6DnI1mzxoP6Bk9G80u28GcE0pkniqvs8xrQLHKV8FcKGDjhTVlZRzTm++SYCfAmhkG4Ghze8YP
kfyO2Cubr57QhjTgSYSN5mcriDoA4kxyl/1/bUsd+d903SitNwzoaSZxn2oz14vU36jVKcgHV9Zb
/OvuykIc0NvVhEkecP1dEU8ww1uu/aeGbIV7K5ZytH2tqxZoLTA9NOK2hvIjRq6nw01nx9bJ/wfH
VPX4D5eq9vQPIW4ob2zUqO+xptzsvl62/VWcvDxUy0kPCCEcYkNHWvpMJuEpMAGi8Fetxxh2ea7x
vzilOFLuNNSV7xNSJtEJYr/YzCYPxGnPDR6mq6rzR9gAYwW4DWAw2wN1wKcalnUJh0Rmst4P2/W+
UkSHBpoozeGUPx4vKMkKT8Tto3lS5h/c0A3o6ok6SUifr9z3HiHqnmP9zJzl4QBEFjLDh8e5wX0E
wg0vU7Yn20mNDyZj3kuVrvctmf1M1q4EKdpNh3EnuT6zTpIXQ3jswnx3oywLq4Z2btY2wVIzooPI
cBAG+oovor7c15P/lps0Gd5ENJE51xMtIrbsKwYjIds4C1fZIV3Mw5HFJxvpp/v+rX75qRUMz/42
ZPC/7l7ukIyz0uCK3O4Tr2AEsw6e96Pcd4IsxvIgzXXoBLah7JQWWcIP/SMJeyPenGp1sNYt+QFS
5xDfuSNaF8bQoZNS27YKHsv4wbp+az2bnwKEpQMmWo+nLJwX4OSuyJ7xParGJpbBXlRX0IP+dkws
iSDprhU7x2/C9/g0JvcUiwAXzB77SxDwxLiI8w3ZzCrQODkigBxKSuTlwW1CiPCIESiV9X4XmBYv
yZs3aHJoFWG2pjhKSWfpfequumI6SpVNsttUtZ+CsL23sbgQ3KwmGAV6jNBdjfRVI6+r4Mo1oTV1
JRFbIgpZLADz4aTSYoRRIlmkFmuPvBojurRpSAMCQSyv3cy6u+XBqzFkcLh7OCFm+3l9vA2JH7JX
Z00RDs/YrWLrRd+TZZuPKvUIWLdSJ8WxJlK8N1BPTmhU7sO1xWtcGWjnDoNX0XwlS5GS1a7rIsyI
4NMY0ecPOmxHJeIlR+VF1GtqGb2jbH0O1+cgDOky6ajKcrr8ve5oLuQBu7KRmlyF54eEdsM+5L7Q
HpUrSgld9Gj6N/2mEEC9y2gHjy9+hFJ6kb/uCO9OeT9/OKqUM7ZEf+3B5Vx7m2+iL6s9Fc1WB+dK
tv9dw2we6H58iwCLtEtXdicIwvS49Fb+JWTBy+NGTL4wRhvK2XU+qYvoNnVTVFzk6F/g+4t0KMNB
aH1tBCX5m0jsK0HoBTVeg9YYw5jKxHATBceKjvbtCoCoX6WQxp2HjVAwRWFg4t0IqQd/tSr1+Cvr
uYfvDr4KNX2A/xZuLEx7p/c0AJvMVlaZG6FiGx+LWS/WSt6Pe3Fr2XxYB0Kqf7uoPLe/WpbRnJlt
R0omvPB0wFQ7zQmwDMjfZsEQzBhVOpn3Bx9FcCk3UTTxbkwohqPoqSXnmJh+htuzgsEf3E1L8miN
+pWkKnaQzedMXF32to6cIneK2+ykwQml6AalNGR9rVpyc8SRSQMHoLqVj8CQ0HktQnnpPi7cQI2V
H1LmuFK+3Zk7/h0vCQ88tsQSMnYBleH8YwxZkuGfBJMykUMyOG5iKzNje91nQDWGn1Lurd/EGJ/N
wCvpuE+754906KJujTeTLK4AjGuvW6XS+DscyvMw7h4rYshX5wMsxfCI3+hbQPqwh7NBI2YqQlMB
LTkbdurVLDTlidwjSYdLg3A8r4P/nkW0uKM8B/tHHEdyxhyRAOwsdBedJYWsdnZ1GTsCzlSLOeJN
SjSKKzkXSYl/qj2I4AYRseKvas3Q8jkC3YTiCsI2t4KWyGCaT5RikQd+X/ABYrfU58kM//MgKaRo
r8EXxqPd1W0ghuD8Gd6f43sJPNfHsFKFnD0o7gwIQjfRwIcn6q3hjDUpGiZ+CKf5Is1t63MscoC5
GWdsZDsgJB72iZLSlcKwxLqki7fg31eyrHI1BYYS9OY+bkfONpQnKbqY3gmUos2sPstPHBbnCfGe
1l6nasWNtnW8fzrzSqMvyTStEtJ+jfHy2FaG8QsuC2MKtdQkg8LR0j5Tyl/YqUgqIErDMTzJnNd6
DSkRz1hC7vRPxY/d9gtg39ki9F/Dp210XLhQp/2gK1mlhjrRRy1bcFXOs3HmS8b+Xt58lzq5gUcc
XDI5bdZMCW1LerXVGs4YsMbNpqoTwsev0KWHsiqCnskUjqZXxjZZmMiimXlC808jCO54Jc13Q2Ny
JGhbGk1CPMsPptT3J23htJrRiKOwu3mc8RbOBRUbK8dM8CapQ8CGQYEUpiALrJfSzksp0QLL0r2K
U2p+72Flx6UYhMfKYu+qcB+R1IV/DtZFIEt3dlhOP2/h9JyMcYtM3NewMmbPBsYOadey1LBFFb9j
ku9buETA8MgwlAx4bSULK2dY1LWgqLMq6gkhrE8BSXWlPhurOszJF2vMMEJxa8xxtZ1E5nXyck36
4lncDybJOTvMPDq3UBkhLjY5kNxYcc5Tf4Hwfoo/qeApP/Ous5oOmrXErIrnCHqEjmwJ44AcNdOU
g37rSEzx+D5CesFPkP+ZnJq+v26GslNZ+KlDurwYP6YaK4dH1JZbK0YEx5OYKVTAjTA2hXl6fqmN
nX5ioJ1yDPEORuiDG/z69HloqO8J1QcTjgHwHOJqebqB31EyCnLISlfdwqnUlDRJGKLAuTT1bs0M
OtTmz8ENOmj2u000Zyr3JayZRdgxAQy2tSTk9NUi/1J9rNvjrMP2JRti5G04zGmKUJqquKqt7gPk
WzUzFN/FTe+3A9U3gb81oRi1vIfqiVcy4Xg5YZDPwR9fBJQHwIUuSopjkRwjJWC6Pa9bsFirjoZe
0KnwI5+e7c3dB4IjSVOSk8sptykUOhjo84VRAxT64VoRB1D+KTqL2+F2zT+2t/sIMyTDV9FrdBjn
f0C2FQ4lkOD0Jfn1iTxuyhk16zdUMx2KfnQsCFhPPxI7CFmfV5dI/suk9pVTeFwDhHLPZ9B9Uq6O
97MIpYD8IZdooCR3aEgHqgcfAJIgl80627ftC0NyKABaAcNqMr5UlP7vR7gbKOSvbbR3vFSPLLMO
MQ/E5PKV2jF0fXgUoHCYRTcQVhQkN3bl7T2B2HyhgwSDAoC9n46+GIV18QF09tqXIUy37mS5K6EP
Wapny0cmheglGC9Z/7Ied5pi+HsGOOQTjD/KHME+odQ8704Ld0+qhYAmAd1z/C0PmF21XSt8qpsM
0SQZUjlFcNKd4MQgYU+zDePeUXVqjLnP9Kdmb6PpwbkQqoVy9Xw4pNlew0ai/1A9BisRgKd5Masz
8pNYts+uA3z6U/MFE4/GYraUbk8F3Rgen+6Qpl4nO3IPo68qs/DNJPFDrO46GLT/hMTZg4apjLLh
q/CvBRtCCyTjHVRgn/0lGYVJ5875xEkvLpZ7hS1JurWNHBGZ+vmJ2kRC03fM5/17ymTCUB//i9NB
T4yVWoR8fvYYLPtQ2FGCVzl/J5aQxZW8f1N+sCbT6o/0hHlfznUWxjRYJ7EWXxH4P9GIyDwMTnOT
2uP/kDOOLiQZR29cTVSUJFfv7sW8kQ+qlkGzIyPJ4eqCsMCj3MMgby1FRsMRnOSR4uvG6j/bVP4v
jiEzh8CcHBjk4NzvX8wcxQ5hv1HXsJRV5PwNIcmopKnKT4PWdT9wnQDgrTaboqZVaj7xMvXxHOT6
Js81tVqEzLPJ4oeg70Uzjj6wmnKpBmiPgrzZMl9HXA6XHafqsVIxbc5iTwgDH5yJ8/ritCTZNja5
w2ymGPwfpaJCHbmwpgwaer1+RCtb4cXu7K12YFDh7fzch9LE9x+Dj5PCZ6o9em81FdL3i82cfiFq
+ZRbjk3Bhroq8swCZDTqMuKIOGqDc0kvzAjH9xT0vQCyoU5uSpBoPOTlzvb+74LqmB9GcmGJO5iC
yD4AS0PeAOT6gIDGasa7Sy+m3wRgRj24YtXTepyn91YQ0tnd9XeUZ9NoFxXfFuuMWEAAb3ZeN+5q
XJiHXk7+Sg3AeYaS9Rd5aBjV8+RVgHyY8knN6tHQO/pvzrO/FR0FwnX0p3eePE8VBd/UF5fTXgI+
22Hg9RDdsPGZKx+djF2cQZggTjPvtizLd9qvnGiSmGU1yWvpZ4/H7jzm5G7CYDYwuBCc73R3wm7o
hFRiRzXg/zVTzXPOf/CC3beLUGpzF1tvn/a1KDHC2MwS0+To1l/HZWE5RsklViPfjUYMZOPh9IER
vUm0PftPEUuejGQCUYog2SRisAxs/IdjnRF9IvdsvLhWmzmM7bXgao97nQ7Wi3hnUVSRUvIGiVhd
kHHSm3ODCkEdjIfZGa5z9pM/Q77GsvWDD3Tl4B9L536vYvATtJO2t7vBBGHjz8j0JyHWRIHczUEv
OFSH52iePNMxib0G37tBB/ly+ki8k6adcqfLNbrCrWokrmBB/fQVCD8KGtkLfGOWfwP7ZeMl8Ft9
Bcqrk3bTmqI7C0zXtHs7dvB+RLE5Yx/sszcKEWMD7rBQJEH2hJwoWg8+m5gDYNTWrTcoVwd21JYk
bWELPz+m/o+KeLm78gNdEVtfYNMKeevVdn3sirFnnNQHrR6IHuP8J/W/G9wHQYV+7wzE47il4HUt
tJ012lCudNDh+9zvhTJ8/Rg7wh20r5ealOjVTVDCiDvEGgBEF6kg6rMyoUT9Hodhn1c0h/0FHAKf
D/PHY3+X5P+q0AyhX8OX1u5t1kgQmnf28FEu4A3J18Dm6Bo0KOYenA6/wgU7nYdwbFvZJ7LtOu94
gh8y3VYj74rXkoxVc8lOX9Oqfsf1MPhzi+rXoUPSRBPDwyvRVYB3hWbB4U+ir+opuNxX6qiXb/tM
h03J6JWOOxLjp7P1DtDhkBYoQqqp97pAYiQptC8cApy+HL1puWfFjiy4ua4vyWD4juyWfNMrs4ao
5u22NynMSpd4QJ3h6nhrD1TdIwEbHdBQPAkPVizhgtfiF6nOc2Ynwth3BpyfxoJs4KV1ZwHHa/dt
JWFyjSXqy1aOTRRwJotAXYzoHdOzPbV9SXo0ITZI2u185fFVq0InWKd9/LR7/UGT/YG0IFx/MKjA
FZrLDv0WoCpBBB0D+KE3qjDbjjDVb1EUc6QaRb1YninEjaOZLNy8F/09Zcl/8ff25XtfzRrv0EMm
Tb2poltLe3NVevmjwti2q1b9y6OPFzYXSKTJvsLZBCoW6e7U8c1AxVOcpv1gaLwik9zT2fqJ9HaI
s4jxPpYW5XwHrwF346nX62ly8QRpFCxr94CQfG8YGyWyoVMIGh12M47cMUVxQJwFNBwtvxoKOqly
StNT8OV1K01B0mbjYJIkGo8bKT1aQ1DevHUemFQiiYL9kHVKuAcQOn90416yUdJOMx7fyyCOCO4s
EjhlbhTfpFkwbIRUb539ArP9mz//LsZ7T8q4vmBTpByW3WjkT+6R4mN2HEeR0Avg2q/pM8pZuyS0
5+y5zHkXZhfrxoh1lr446YqaW6HKcICJoNCQChQHgwzrZ4U2mSNEPT9VV8AmJJ3mvg2hHutgv33o
H/wcaEkT3Xy1h9+zpHOw2ngkYrk7+dxK6N8S6EnMoFC0n0JO1pRV+g84UmrryEnzdDoR5o5QmnXM
DvDoeEqC0EmrTp+zjKulftnAM9oDbBfNFKeEqSnpjEkW1MYK1joQa3M0KwxOWLsbkz5x5f7QU7Uz
4TvS3DgIoU5RBMWyS2NeAA8UItdcCslwCRi4TsS8xgowzDIFj0UaUYeS0d4LkDmzYv/HkSoygGJ8
MPlaRakKtJnWPK8/kTTE8xSsHw3PMt9H03T1E7Ch8BobQVMUzUfV0z7rtHoMRXI06EDT1z6bey0l
YgDpiBgivao3sHPJZfOySDVTI3EM/xZiRhmitWJbLm/sdaug1MZ7Ax39tdMvm1XZxhEWobmiqKyD
daPeLVtpDc49liwtta/m4gZIB0nuwBUB8z1tYOE5rpelddZcx6vBCTZ5BlN2PVF3Mb8AZcHGyQF+
OspBh89A+1Vyh2yFX7IAJcaDx6BOsbfBGEAiFe5iMLNENgRwmNw1hRIq0kcWxC/wFdVwv3Zj9q4n
vx7jhRe8sispxy6RiFqDGAZnYEvjBvHwjQnLpumCz/ltX9B5MGGnqZ05n64DaefMudUDvIisMRgt
PF+Zpuz2ARXtxD/rCUJ1MT7Y7G8eg9Cug8NNodgqQ1ma4W0lcuuvTlXHYzkaJy+qfu1PadvMHIro
gwOVNcxU2ZWQ/2mfbAC4Tel/xn6Y3MGSsH1nQqK8PIQgWFV4FeQn31KUJfELibPLjdf5MltIVEzj
++NJwtNpJJr3c9Hk+x8by9B++13t2iOXBrdKTmIqo0s/5QfEmR8K0QqaEMOxl4veYNAjzyw27/mL
V7+vV5HwU1cMq3k/SY3k6fJ3hIPt3aGejPFtMhy7ITTUti1Won93xvSOizXdO6HkUP1kJQj9Uv5V
HVcpzWHUacNp+OriR8jS5lH8uy2KMyFkBPElsp9o4A/qDmjK2Z3Q316yUUMDykwLyp3zmDIAVkDB
thbh9i3ZDQlalE/JwLvsbwJDmRTNB2nHbIRNmXtw5HXMM9p1Lr1sDZxu4G8zn7cvPi6uKQ81yrQa
K4OT3S3hrKhQ6I3IV+Y6SMTUAw3sAbLYBh5e01iTakxlPPhv6Uzx6Sr0lTsQmeOZJaAhKYKyO66s
oEhmVm+kAcsBVrNDsQYlXoedDEuNJ9XfUj8yjZfIp7aW5BZ3NG/dY2Ooial0niW1m4/PQuJhNGXh
SXV6hK87hYp19cFCrMhDgRsziNj7qmKzcHrlVXkbkWdFg8qFuoOvUA+YGJgQOe41prB9t9sPjr3T
6cIakzLP+dri9DE/UHG12lP7n59lSO++cZl6LAVD2exMYI0CZPb9pk5hS+CglKLQu9Kb0F7qti2u
CvYa4LkYHEDT0okMtwuj48zqMA9xpVijDpnNGh9Cip/0QnGCMyFt0n/9JklOZlDnM9tKwdLOOfd7
7OIKfm3LO0v87Yrb2m9XD0oQU0jCMKRYGM2IFI/VneZnC6IstGsUyMNelzrqBsTIvPpvlAzKTGjA
E/QjpmAN91XEc7M0YqypMQeZVGHGmPKm7UEp0OKS4pVvHn/gtx48iKPOW1re6hzdhX9xYjxjBfbd
JpuEu8Rb34RLyywwMvEVRTMUxcjEut/Dm5mLU0/QcOV5TUGLQekf1Pkv7MTBAWGazL78TWfEMUfJ
I/Lj4ilsNM4o/SUhbSgZkp5nwekcA9y6sviDFs2bTK3qvpn/NLr6k/VpVotOh0mzVyCvbytTOeLv
XGFi6b8v/06nWnnPTes5D5vZFT6mm0zDeSeRc0KdWcNw01zx6gBBlZn6rhhehIm7FhIu6vNiOtNm
nv4srz7DboSld3o1a1NzHznTASKcnjjNB4UUpwSgicqDgmUvACLBCrRfi20vAvylpLi8ViwSM+vN
WoC9tlUyyRjJ5VH6iLqK1qm0pxe/dAmSJnTJnd1j9i/21mpul1J0IJ5wKKeWbgsowO+aRwwX/s71
OoQvQtYiAmfI0JE+5/56MDQLttyLmBvaiwGZycjfKcvy9AayytlzERnfE6/7s4rJftM7xzvRyXaD
pnkSumuhCNvAv510O/C1b7vLn73mQU3XxUaA/MTKfBwjPPFMSZ0uXU8jcyIKazVE6QB4svRieqVv
TVLZf+sgKfg4e+z8Copb/7SHlMJlFQe1uKrv3vcxPWFyBZ+5j2daBA+NcWq+DmXO39g+lVE5x17d
YgYRwm9KG3Err8Qoendn+Ype911XzgGwFdzSGFrDTZpIwMfib67esAdi7/ttochwnlEkJNDZytoi
VXO76BOVlmCplLE+CGYRJ1HUdmOcz5d4r6cclHI8145d7xwkDJW2qyx5A5dFYjHIGc79M2LUGz8D
zWH1vBfNgeW2Sa1M392YXuK3mTHF6VpnRZT0FwKHcV1/KtTYahTMygK5foeX0iTPzPv7x9pol2Qa
VnxDHs4ZGcjWAFLyPpETMD9kv2yYqOWACnw19TKAykyV5YESovShOLC8ob8tQzTT+xPLMosR0/ZX
7pTSMvnMdbSefpn1kOKiEO+0oz+d02UNM/SlMKmFnFu2DxZRyZgI1JaI8PYKAn2mlWXIQTz1HJZM
/r4do/Gkuk9AeIzomEQ+EVpY3h7JulR4XeV/tpVldeiimh4QlJsgfaeLpmWr/OVMfPDJJqmGFf78
CFBjlM8L0kHULK1n2FLSjjpsKtPqpwk/D7V15ffQEN28wq0kiBeGrvY4DlyrDjdCIdd2CR/Y6hKF
0jrU4WkLEYIMmLPVrRhgj7il2d6/Wf7Q++UfVZbSJYcbpviedaQkzXATCRw3wxWPGMqJk8gZ2oCu
1QsnbSFylwpXhWC+ngDuyD0WAVo52bhJkF4+LvxyMeqxblUPZAr+KIYA7zJsWVFA46a5cai5xDdV
pZWytq2X0wdU0XaJneai/EcYVgRN+fR677dMRD8aoVEEd0J0RZ4jq1xFic79QmbVemP5p9SibZa5
4nmD3p1fLpQ8c0eeWq08CPl2is6d/RfO6/4tEKFm/OIqVcAPBTrGZmrg2e3iI6G/NY0CQsoMeYZR
MO8j0YkFjlSd6Wu13lt6M89McO/uNDdKvR5hJTSxx+JqqtD7qGDMkVthw4o410Laszygn4ugDlRD
XGsSD3D9AroYPI7QlxDOwPFya0maC5UyzoCiQn3skq0sku+8QQxo8OV/3u2NVCXtia9lIQCEP5Df
swIeW7iKpvwnDN8CrEpzNZitRmLu8BAHCfHD6R6JnCLqb5/i47hNvCHtmpmwCLAvw4eVkGiDyv5s
JRMnsLGJ3a7T4a7Cs1EyMRMpebdzET8cfzwrG2NsoV4dh5z+pPEdFT05JGsCW51nBm2iHciBbAZi
CPq7llud0J0+DacZp8V1AktbM2zKZi+V1aRrei3YTx7iqc1bD83STcRiqBxcEHjJvn358EHw20cU
AKTMW4l+gjZPoNsp2lxYAljfGTL0wJLEzq9op5T58wkIKss425XlH+TKOszZL3lEp3eNoNz84Tqk
SeCAWozVZx54PL+7rF7YR96jq2+bnBvlAk2IXKkhtn5BnfywcAh8GWjUhnseatGg3IFEA3bOBNAW
r7Sl4w3d44N2wtuFJ5+JAcE+hTviG7jLrHJjNQu31QLTQvyn+B6RFhqm+ksXgJvqb5xUvN4y+5UD
d1GAYY6Lcr+V3dhpnuewyfbNJeuNIsCXVIU8qpdhiHf2a5g/LNxCt6j0fAti2zAWlIRSqNdojZzk
iUpdGg0S9mVFyORFjF3UQSsiXA82sWpLTuXZG6HO44aC/dYdmN1iqtPw/z/r7joV0IfUVFISni5N
CrjYZ2YuUF7ZiglxAffwD/2l0m635SgWFdJVltSLxtOJyncGxcjYn9o/4YoHHNN8ye4fREx4TnH1
OqocDx050DMfPNePbRH6s1QtLsFQCQBNSl7Uowpuwovj+hFu4jdVFJggd3Bsteg3eI1kjHRGQo41
tW+YPHfINGCMh8D6hjESLUQVMvSZzAY/5JoXK4kwggz9+pkVTnnil+MVF2QjIvRU5wtKZy5611dt
cftOOXlGOG7Arbrdm/ALMJXCShtxhcaJjnlI1h/0TPyPhRIaGfkxnVDxQKsxe1l1UMgbbVtz+shN
KOY9oHIbVnt1BTV8R0De0jwRht/Fop4/cNSvIg9HYF1t0QG//uojPVqOLjPc45p2bjQJJnyDto0N
ag/IkWfKvaTeGdTHwphzK5bh1PHnIDSyzdzg5LqAK1V+TaDTstBefAfTa+F3N2qqeYjrOyeajNsa
kXTzOPoP9trP80zIzSGGzFjw+AIAL7RjMJZYvHjQXwWddd61fyogFNodeubzcJBX26ZGaBWj6/Hf
jQ/wI6GMtHyuMrKZvvOrjNWgWOVuSmRAi8StRiqxlh3uDlTUcTs/MkbN4WWTyaEquQDp/tsk7IHW
vJnngCS24wvjpPMT+wPxu5G5f7mg1F+OKyehTNrI2rCm5T63JZYVPuEva+jGJjVYjSRMJvnEBCqz
h572b2vbO9pDpJn5c+pKut4th5sFTitLRFe6NkMset2IpLP2mst5znJvaIs029a8xQYEFMHK+udL
B85HqS2avP7vjaDDYqpWUkwKrz7BosU0J85Ghhgcq9jq0zTM//V/relXBHA7iV3rC2xthOPKdnGN
kAbS/qej7p6RBEiukx/8TsoTRaRzeSVXqFw2FWz6P5Q02kP74q2QAKvna68xF8pznjTXdICUXYA8
TKB8Mg4N1ERXHDFCMZQT0JqqAtln2aOQxMxPAHZgpk+W5q0gdzKDSUKflwIIm8yxbYRH5pQxXvDT
f73w7k0LaeEnECj1BkcKiHTCRGkSlUWu6mql3nl67bYkcYrfOrCeyE+StWAHOR44cmdDWzJYHx47
sVtm7yv97401aWAlpn1AEvIDk5qGGymW+0EnflXhFYVMWPrqxvvehrOUzQyrSUDPR+PoMOlNU0ap
k2YaEuXT+5X/XeUfR5KqMbwQzsd+/sUoia/ZCsArMVYeGz6RNnuA1VR6Dlk4XhRZrpkozifh16gQ
tQVEBBl+VHyU9OxH0jK0gpTC4ng/4+QPOyHtuIIe4CabDBKrR6VdAFYNWK5aaRUPdP2QFZgV+qi0
HL46tYYkuueKI3U5JuOz45VtKQAYL+cLqcF2oLQU+OwRbW7VPYO0BS3LO0enNkzQMfT3RTIFxkjX
/LnYgRW/XfIjWOXlM3S9Wo5W8HQjD53v38KmAH/ZxGVr0tslrZSIqNIxFDFMuv90EuuxI0ZHqATO
/0IMSaS+mOh66xPjWW7Xql1CRC3jtKtFB4kUtNDkhxZmB9AxV7l2wHNRSZzbUprfUHYoMLzvfmhT
JJ/TKPEq77/7biB6sweeLHH8C0Hgv5ePQKeYSOMB7E4rNzHvXREHNRLBXWjSIf49jxkNq8oNKyvj
p49qehrd7jVakElaoVRFSbMr14vR8je/KX4GBd729jUQtf9k7g7bUNyhJvt5modn1x/a4oeWsQ9K
SPJBowzbkBP2coDpLaoDMWvmQL2deXlZv5sXS1u1opWwGBP3JFbwtXUncu1fSC+aCZZOBteeVNor
yWxhuGev1rYsv6hjgPx+SQe8nJ80FGWPr5eWCOwXXLNZRmf7vrJfGv8XoLCdR9LbWEpdiH/6fXz0
QTG7eU8q+3N6Mjmay34vKDPN10s58LvQBJFdB5Y3tPV6vVNwdLXwocyKOp03MiaJsRy0prVdtpF0
07fSYgxQjfUo4Kd8n6GTjyS+qSNQHerGcykhP+JwED0lVxfBU4EEHbWwTIgq4B1UIL5Q+vDaKyfl
UNpAe0bJ9ZvwK7QaloJUwaHuzmVXlxJK9rRWaszutly7DwI+FwiuwvxPqpYHDe8ZCy6tfjk7zIkw
plf3odXNnjaOfvRt9Xs3BjpX/lK4WZyk0ZzWUAFMggA9QToBPqkqOl9hMD4865lcO0PPBAGsYjAV
tic73meU++HC/TesCvWbvlLj7czMlS1eej7oKa/9Brw72Ve3DbzYIh7mVJODHVM898vm3AnLFBpA
6wt79nVONbv58rs4rDUMn1wV0R+wnK/pEikN7uPCC4dw/ToeyXJv79QDwzjZ+r3BsPoMREwwi26s
6PPPCd9N9KCqBzKh8YoYus9Hr5n3uoShwFeFS7rPfY0dlgL1FwJ0nHD7Gi4qCZdBKw1u/ZZon9Pg
uNF54qJB3dO+QqGsmdQ5n1v6GMX3Rvnm0QJNC3FBYolSc91fNKSHAMZbNrgMxCAk2FsTnAOqTrjy
3r2KR6e2unRpE2viZi4bsWSkURU0GVx4WHdpGqu4e2X0Pc9xI+moaC5Y/wu3AyGe6HujB+sXGbZE
Zs3w5La/sE7WAlqLUahOLpWeam+UCLnYWwLcwyFz0ZUmSCSw8KjtK7RuvfF55Lb04FCp9tn1WMw2
wWd4R76z51AIgUcm7Bb1HFnw/07UUwUCzFjEsH1cBBDDvG8HNO4taLfK9Hj9AsIk56gyQ+kO7e2+
a4McPCwK2QNhwtLp02bCpofLuqmSZGwYKpqovvB7P/3iW6BbpjEv/bTeFM9AFWZDIUMuTPdBMVxl
NRkTuj9+E/91eUWqa21xJVO1QQLmPFEEK52kjCXbsJ6PGDd31NLQlU8kuVbVFxHu1smTtIuX29Us
mxBihJkF1hvjf67OeDtGgB0wEZBvFNnNYP/ONxScc9pAVba8MUM7ZozlXUPuOM3IFIYgSPEWsPzp
VvEG5qiKQV5C6BbBN+lz46ubvElj4bzhgs4OMWh5SgX8TQjQOZPvnTWQzZNuqaoCgM17bkP5oepT
nJS1SllyOKFcyitkv/3Ut8x4pzfyrb1JXX8i/cDWRYeBSyRR82YOm0+Mx5jfR2X/szWdkCgmJxIT
45gU4/TUxMTToUFZLS5P27sUpUCp0XkOh0N1ZgfVxn65NAEddDz+1/5EmH3T8rP78QNro0XaenzJ
BjzW97n1LlxvTJqtcH1D2ZHALdEr9o9p5UZp8ma+zhj2BuILZegnVDAm2hKNRfcERBsc9+Z6WXUT
Nt37O0wVkyly4yAp7SAoNZqwSI1DXvek54g8LAEPdvee3oV1hGwwa2k/66HfqgqF+qtUlD/EbFMR
zev3LwhREs0Ez2AUDZPflHfcg7pM+kOsH0HxA/0ilfIVocgNdLZdGE6aAZ4AWq0IYRshqZ/08YjS
XV2TTpeFCWNYXweKSg+puO9UM/ogDF3p25uQ+r2+I2OhwmNgnLdHG3meWeFH1ia0ilIkOpGzgT/b
3RP9ndSgk8D3WPQeMYm5AGziZggCMPwyF9/ymJfemBjICNzfXCi2oERndPD4kqvAMklh8p7hCi/7
5SVXkpOHvbqWYhWTE06PYoId+LAMdY9ualRA9TCrWRGK0W8IIlVMXxV5Y3hxJSe14XszLtuSndOv
A1PECStXcElSjhcSGRpseJkSTY/0cGepPu2Ex8q0ZXfMz6IOlxYt1klqUjOUXCnzCnSqGNDA2jXn
ONHVu5bmwZCh1W25e6C/Bez5taCsOdjkRoXMS0Tw789XVFMMpDqdVyNDKiUE77HOTMvV9Xy0wYuf
AKwuabuKO00aXoUD1Oi2TctGuI0UMCFSW2mmts1BhRa/VuWTMwLyFxZAw8StI6APdSmk6rTO+A/F
GGAb7OW0r/rZNCJWn/EuBDTvczUgZSHNA+CqalmLcRMzvQgMzo2XE15XOajTZn75KWTF+U2LRm2q
/bmk9/n6YoPGFT5+vUtKKy7iR6KqYuvZkxEITxIq57GQ1iBmkN8uLqu3LzTa59lTJccT9FAR502s
PDXvTd4/xsoDRDDk60AQN6FEhTuT0YT5KtXYy82IJ8aCMDHYWM9HGWRRFf4CtHJaodke4GDs7KMG
9KFaRaDu7RV6XUU7DBmHQKmm/OuTABYFmzzVK8CdLBaRTvZdSZUnC8C3CZvtA0pBZk08e1tNcAWi
fmoKlBHgq6aABRQMNihgo3lc3VN1HfgvS/gKEvj9gXUKUiSBBXmtXAKSRn78Cfan3UXnWw2l56Dj
QCgNcBJxzJRzx23Wjw2toNa8zK87XT3U2sxGEI8k0R7GAk935XMZfNWq1U5iYjLAA1vMoQcOpBH4
SRzBGDFTfXKY9F4szktAZeSaoXLZFhYzc4A0vHKbJZQZZMmfo0oD/vvQpkjTajDdOfzBGgGlbcWM
vE2Tp7Avk5+6T8mHAM5W74RkorkMfNNnpweme1JiYz1L4c8V1BFZ3CAsD034WWKGvfIwsDon5Auf
BySuHV3YEJsuhAv7odB6PBAEs7bq+VqLTQl29dGdikATkz5GsHCVO/4WkgiexOCKE79yl6TlOKLO
/hU4+QtPBeZdxxcONyZ0fyzFUeyc/occ5y/iWmr8ZyclwbbhZFLIMbAfKW4Ai5pR+JdQ5RXbq6Ap
3iNG/QT7pOorqUQoED0LABVXZp8FcO/nSEbsRZdnvgd7KNd90kL8RvG9tcwA5alDoHBIimN082OD
1Vd+fgLVBfHoAnDeNhdMoJNeESQpF7YsjRR07Kk8DQWh1nxasQ6ePR/GdPdwUBMP5BlmkzPoezHE
SUaLSRY4VXevyv196ezXEmP6y6kY9uimpJ+YPImHWfUPmll3Dt3dDhkwIUV1t3Uy6945ndYBFSIo
oq01jvk8+PuGSDJIX+Nnr5P1PRV54nXPfpCLhFZVY6K3rpzldeHfeo+7ME26E/pKdzOQXl1bjsjx
EZjMRgealnXE+PIbnbqgA5CXrI00mSheyPmFBWuQk4jyeQbKe7947qRqmKd6C9p4/+b58haXJZGi
K6Ki9T/+3euJEzCKOnT5fsg7ebJwCMOVtMubAdXPjRK5Ril1MS0+jE3UA3D/fvLOaqK8M7IyHJH2
PKi76VqnGCQQYXpqfDEOevBWraRezGRGUwTfxeMehX+OXNedf68E19aq2050RRKCywxtPVFvN2bz
H6YWG59Or4eomBW4t+YDA9eLHI5JeKb667db6zIIEoBRrXo/A0M1GHwlISjrh7bAbP3rY2Bi37+P
Io7Mna075B2jxntHwzlj/a5k++OX7jZIQJ+VLsm4X+L/tOKq4fkbL1QIwRufsc2SPLwbPHJEfj/r
avqoMIuKdtdZabL4uU3SXZW0dvlimnYvxDJQh5ZbNaB3xe1Q+KwpkL3OkNzlq6nnrmqVaG0IBYL/
H8Gdxu+AOiLqqLRkSUfq+ytazSCt1MsyZsqFE3UlxmfYlEehnsWT8ttOL7BWolMknNkA1TMHdyYK
0kaVjm+5NUC3TNLmbuwgZtMr0rLAWSflnHfjF69CuWNeYPdTADhAq8hMVXnc87UduRz3tPHjpOm5
kkB3dySz8wBtOp8qKHnPn8k+QpqchNjvOIt8ebtnCJH8Qe+vQMO+mE8MnWpeI5siUgT31w5+N4at
Ug4ku0S2SkOZOhk9HCS23nHX/vkWu+iL60py3PbQXpsTRKxtEX1y7UPNuvTUZsJ5ZMlc9bt7iHTZ
uo3aqxfFC5t3W5koTrj/zuyaXcnqo1BrKp33FogrM9xrdbi8jYINifM4ismtNNasUiMBaEjDAiOE
xEu8IZVe81sFiFzpyTsS3lHDY9nCHAO3A9PnCq+qU3Ns9Bxv1YzFTU2Yd6DPx1VtPH7alsV1C26N
Gkdaee9Uf/pWqQ1fnHaQu+a/iWMHpTQ651viUbUjy7bT67JhU7rSKH0f48T/ny0Q+bq+EQrkDZUW
bH+02qdue+r4SSjALVSzdKl6a4NSuaOm3D2mBtC2Hlb5ig32A6OV5bRtNuxMGUbRERmCxpbN3PIJ
5f5m5pf3TV5ugoklMqF7k84mSqWsB6jEmO73trmhpOqY9l323XVuoMILee192pBnVbM3ya63Qw6I
y3/RVNtz4q2Ku2ho5jenoywGh5VI2ySIIuXMzR8F1i+yYslyvBBmW+kwcrP3wEOV2A17l1V+lhr7
rthDpRKwLOnyE1U0rVb8yLfdc/65zeuTMrq5oKrqngYC3Wj1mdjDTDG4AuPEk4a9aV9ZsmLXF/g0
RkiOEevh/FjCzXFzU7YMk0GzoEsDcDCdJIFzVcBfzH0FVrAGhmLTMndIHdDQHkwci8h4VCLhzLVv
ZsKKyuoqsTT8lk7NPGNeCw5qm4/87nZ6FRB+Cz6DnvQt5JsvRndGddUvCoXp3XKzTSFdedGZK44F
rbUWIS2WVItFYYd5YiHTab5tosYuNgBBmF3ZJEBSrvLnNaCgrUFv3IuUDPixjbO7yRFLUyF03DGn
SKKyYBYBH7+NQ17TEO/5fyDsjfQqElQhhYc2hd0pQKYmQ/bNsOmr+sXL+LQeQpKTQY/7IGX5Oq3e
CRTVZkhQknbad0qBQedDahcnJUOhOSo9AUVirZovO4GSzepYvxKDEZtUFWIeTCyUgd+UJ1b4qpr4
aZwy4NURt4M/+WO6b7d3Fdkdept0i6bGmG55iQlpbhdQvjiKZhPDxbpl8uxd/U9Qv7+mVux2Diwh
kh3OJfTBoiXhMDMNKMGgQpxbjVZgXLni0NbwguX7/xZy31j2C8n1tYitPxBiXZT7Uq1IXo2Vvw3p
HVO/V5gu5XA//MVHWu5FBwHnGLzIfHNFDMgMD9jc32uURYKClWQsqo60kZAd6XFueSpYSZPbxceu
bFnX+yCIXGCuNYky0ppdF3oU7PpZqgI9VDbFmuAGwc9pb+5nLU02Z9ymp4BuLCipqMcI2+T0Kaha
9Dd2d7TRpYzWo0HWa7KwDYbQtNeJO1BRMO23bWN6m/C2+pumEVVliEKTZ88E3uRVjDHtOJd7wFrX
trSqmQPv8u0D/jm7Qg8xk4S6r1z7taUEAXnjHMqFDpYKBuvmz37WRYjJgUXfKYxJQhDVTrFlk2Ke
b9ZDqOE9RW3KHUtutRPjj1bRFYS8KqLeOtickmYqe+pliy5YZY2hdfwb8widfAqBOd03hlD9EXi3
B0LceLjI+h6szZzvn+bG2NL7REGwam+RdL7q6Ag9alehngs16ke6uQ8lV1iPi++6cc1XKo5Y8qUc
bQvjaz3GKZADDSvZppE6UHLS03+1VImDPWed+XcGymm5TZDGxqUVaKPsDhsXizvLgaInLozgZLE2
LBV2ry6A7YKuYRdstKqRdFFRb8TKxkoeSgwQI15vJyZsM3NUApxkU++9VjUBhV59pZiskFe0tTlg
fpK5JoreM0PaPzoFuIyQZD+p/llCun6kIEGh60linXkyvmIu/VjRRqNxwWmJg9CRGjCyYfXrd8sm
JlU8bo5GQkDmQXwXu50vZn0/PKXznxa73wrGSAuiqP66XUpUSk4xqlHHidD7N8ya57iLo0LhWo3F
fAXIrGaqAksijWavP+y0GvWwh9xK9uiE6cjx+hvI2ii1bZlaRF8mtrKInaV00vYweBnkxRrOuAO3
mAR/TMqR57qS5GUQKq/VnQgvD8MXJR/G8jNa9cJCX7fdSrSry0XEQ5LYD03QZ9/Ph2IppDb8gRqM
4OPKhMefZ+tZISwlDyuR1jYkZUM2lkcfDbnipNOvYBoTmV+jU077XjDgdwAKtzSLYw5WHDRZscJH
0f14lTEZ1dqDY2geQm6EvIbi3rxRvzGG4Tg4/UfqiEAimLaep3lXLJzh5Ian9+Kyib13XwlwBCgZ
+tGZtfo3wdUpWMNfEKwO7fIaZKeTWEDVVfJA80mHM1OD5ptvV43m6VFqEVrg+fmy/ZTGhKTiY9IW
c+A9+9yuZxbkpK7hihtfQBccmEKQF1XUXk+4P/1LbQnc4088lCAQCEBytqfON94QuPT6yXwWWJ5y
GAMzSWL1uObPbdMz2d2Wrq49AwFFjyVL2nN0nG02LjdTpYZIOnLf9yms2irTdKNeIfdIq54TKsZE
zrJUVWCdKhBtABcd2pEASI9Dztj0b+thpCuXt+Qe0A3R30+ypJueJWjCJlZjbdsmVoXAZzj16SZZ
/Q3sc+MSoAVWZvNvfJE7msT9zUd2glBcdGs1fLXpOMqxUPw8xvOb8Grfvo+V5jx5vgKlxaDYuLhd
axwx0ZlvQetmb+yX7mUl4u9FKuxfn5aUPdADypupnZEiWjlLB37g+j/inBqL7t5SJyP1LW/RDnt1
0j6TftE2XDlUX4dC68hlfHR2hwBqhmy1LfCxnhvbnDdmrZWCwj8ekrjK5MXxJ/9ZAWfgw5e/UlM/
qoQKVcuY+G4tJb/7uEFDlCVigMoDPO2GYu/UPG/9sO0496yU8J+0IKiW7JwtcBQmUUz3xj5F7CJu
qvCSU/NOmbzj0GnL53A7HYcBK7kYP5/orw/QqxZSgGhbS8S2GK410WgEvxDP3lymAf/xLrNTHpvu
YSnkkanz+KaJ1pcShT2ulFV/CEX7YDuqJvUQmpJsoF081j+wBkHLsctjTXkQMJHzYHh8KWfGu1/P
o8FuIGvC+fU1O2hKFcCM5mCd5qKgqcB2XSE+IyXXuK3UFKQQyI7JvqWl3ynRbO4jEneEGPr6Jgrv
GG9y/302T2+oS16oHE9eKk4h0KXSoC2w92xlKzRw/DOqODe3S2oGcH45P/miNmPOMTk0gIdLUJvj
cq5gmVoNtgBni5TgOzmt48QDbb013WWMmeVcuuos8NJi4pTu9S/jDLC/nAMNLIZVUG7BbkGBsLnv
NNVJm2xXcHWtmnNN/R5fsFgtIupfV4s5trG4sUDwKdYEeU7qZD9MINf/YBPIzrTHXbw8bhMvJsUh
pKhi88pKed+yPnYc7gn9m0cR8GW8zH3gQegIPQAprCU+eOGvZRMfHNc3p2nkpjOLHHeUQFm6A7oR
i4n/e6ir/IKtq5d92b65n3Fv23LrdsglwhZvWMwHaUfzMGvnv7XTTf0UrC4x2pbp5YqSQG8cWZLJ
J54vHEoruoz0izQwNwmFHvu7rfUgzXJCvLizm0u1DBxha52AHuYHDG+Q4R9l3dZaNwofqyOQfHID
9R+qCZ8z/8IqYMblVbYzEDkH2yiTfDB8aWxB89JPR48C3rg2ajHZs90QzhfNocuIwQ/ZMtaYqR5s
aQ7m8HATBPVYe+Sk+6vR/+1Uhd97c8VsC/6jlTu/O6wlDmR+dTXlGvdbioxLLsjob1LQHu0AZi+t
iuscD74SF0UUP8qqOUO6gdRjs0e73g/TJzCu490RfDZyAGUPZlCVBfmO5d4wsyHPUA1JZB5kwkOn
D2Ffzy2x4+WKoDxL8NBPJzABlcdTTF98oV9ZhjRvrTWVM+hTRR8mvnK6cdGp7nGFTRY6voVOqwbK
rnuD8Ts3lq5CQyMjlCmlalO72fFhb2RlQV4e7xBX/t2Ln7zvDFOD9bqmZlu2HTEiw9SsUmisPucL
kwWJTDcfpOsbShvaiDo4fJqswg9LlzCui4aSWXI9WS6U6YCnkdDApH4otPRWOjFSC4jsujjR4V0r
K81XY4Zwc7+WT/tF0J6Maut/Vkq+oSfSqdbOgNcygauOl515xpU1k5CQvy76PORenyqZ1oieUkgk
7trhWzMV5uZKAAkDoK0UE3HFJJQCgxfWu16aMnsCx39G9AGhX+qGuaHN0QoH8f/jXK4SBUMetxTs
dLcooX1KkVsdLV6QJfxpaV0TaJKA9HaDCo7/6CZjZbH9UUElZbVukUK090Ta4w9EpEayOLGCp6U1
tGn5UkyuAqOmHQilxTICmUjAaWoGhVg9feaBpjVl8dHC0gW30gYOxx/8RFJBILNIdfwK5GVpFbAi
UCot8Kb3fmG66ybcl6ZiqKcjqvLGsTnHaqDlQkrS6ngekMiMemekKMf9ulSezOlhIdCB1I1WAKNq
FfAsvsyv6cQAnv0NYfW2pnlPgEGiIEldYRNDZBFuI9IUGi2tkSKGQaUGi6AJzFZGu3haecZ21OaS
1rOhA2fXREsa3eMczAW0cv1IYLkuaKdOsRJIkorj3k5jhww7FofWgpVw8CgB6acLY5t4FpA0bsBK
i/O/9WLwwk3WYwduxiGAlaRUGxpCSVl7NJ3VCODYifTuyevcxI2jTH9Hl3ndvcpPruGNHvc4KSPP
h1dmsgjAY7fBMGBnlYCo9298L1EYv2kx8eR6GpARjSo8lxWMINhzM2xtaZArILLygQnkDnpvZAlv
oCroi/uSrhc5ddpZVbznEJBWaA0zmbV8dOorcmFcqdyO7i5iNAyQlQUzCD4vO1sDKDIAE8AbDejI
UAV4DqppUNwW3br2V8Us1Wy1wF81fmiFR/M9JvsFVkYjijtWgs67N4ahH8RgAgj11n2f6li6QN3f
jp+cyKzosb4ltgqoQlSTQjSQE+2YrKTJXsjsBZ/C+WGMSuzqwt+ka0hKssEvG95uBOJssVA6rOyz
h6VizcnUvZQ34pQzn8RU8BNwZtBvojjW72B2aFUMkNTBbvoIIAH6tE7RYmFfI9l/IFRhwp6QgrGp
0/DM/tLqjwrzPi3xVNhKUZPI+Edaq6tIs1NNUqnChuoImNDj0iJ4cjNG1veZNwQfY92RWSv04Xaw
nUvkWUGzsad7VilwEcFdGK6A2du7LVWiZ/rhoW1//E+704hYaYAM0A72pXR2EB02aBWIAohFXgTk
D/z9k4mY4UG/fHhIUZcLKdg63fyawI+VVnyKkd+o3myTZVAyu0plz8wWa6M7A2arpP6izsS+8W7K
PYosZIzPwoCWAU9FG7Fs8UDfVGyaJeEbOsi65ezKRoFtKzN+0/+qkaQ3G00GJfbbl2t94d9rF6zA
aabhEjzEGYC9zy0HA5zEBgMqmF4UjLrEqRQZo6aHQQuL89SiSR8EapSip4nLm9OP6kZCKuVd5ihE
Whqo0u8DSLDoEBsqptkq19zFJ+wjuywGIwOjHmXF1o/l0OV6U7mr+D576XQIHS1wtJVqWfIvJhMT
/4BgYkCT8EDfYKScTZTaGJWHoslrV4e/I/Atxj+LzuQUCxkc2s9Soji4oRqCu6V+N1dnwTWsKUF4
JxpgCmm9Yt/n4tq4NlyhAi8T8xB/lxZRsVL+G2ruQ5Ne87u0NEdeJwPjMZvXr/6ZKEHfTkn18RK8
A+rs9FJ/pKrMGhTMdxvoF5YGmXORmMa3+4CyZ4mvb6diMFPcobCHQUwThpD5FHrByj/WaCH5A29g
yQC2LxFCCGWSrQ39vz+HvNz0WaCkM4HypXel4qgpE8jJqOEr52iQAb731qpCk3dJYXxJMtU+io8x
7iEDRLWE8injeX+cs3ZnoV+VLUrdT2Zc3xYZNrRX1bY+aWSniilo31/DOk0Y4gz0Pxj82AN8QQII
yxMnLNDxFBJ3SRHLkLSyc1G4et70I3rRdc5hbzHYv/UY34ZfZiwZJmcWhUDetiIpVCz3CyqGGHC6
iwfC40PETVJmD1Pc6iL1U9bVzXsIt13KkJSZ2clxcwyBRornmx2/4lRdwIEEsvQxPDnBxR8jauBP
gUsi+swpjXV7tX5WfZgSRH/TMScJnqTwBPGUgB6wtcXWsErcREXDH1OxHZ+s9wwgzWjhOIoeg5Yn
H7nF6tt0r4UcGUZehWbYukgJATp2LmcBMqOcSqNdv7+qJygwZqnvZNh4umNtfOdql5K0RPW2M01Z
pXviV7E0/lt0iAULNjS1o+iPip1CshZR7Gu/Wzs9VWkbMz2l+/gD1Q5yVuzA0DSKHgJn8oa43M9j
37OEY8LA5+lb1PSo/1DnM88pHCdOoqUyYHL5x06Lth5GunM+A3iIoUHZyDWOCyr5m+R8XRQ9RLcV
Rc1iCcPpPXv6d9A6TnF/5XaKyVFxP0k+rJvJBNnDRj6nmtt4KRcoiLJPetMLCRyqi0x3kqWBe3nH
jJcMI5dnSwqGA0+tuzNkfXwV+MFJexorghUkgnaxkHZkbmVzZUkIvLujQY9SJjLdbMMVaYtHKdmo
h/gW9W90CwheMYXtk2eIMRqEpD6Ij2280dsiqo+ogEqzn+n71e0VKtxjGSyS0bCti3/RDCStoWw+
XA7GX6iPg8KDFirOyCazplATedyWbYNLXdYjdEDTqxLznhaKhhzEKD7EcrGdaLu8E5RWHCYdDVHT
IlIOCUg3OrTnBseBBbd4oTsaicoZ2JIyiCbrQvjlapNurlUnUwxz907jYcxynC+YhmVI/Pi5y681
/eKr0FsATJ8LYi8cWPD5fJvOusosk1axOvS8s5g3DBs8f2ZWtFUOrLnN1wwlmgeoCE5MLDVVZLgg
9+V7lQtPLmZFwW7Y4kHFKWe0PhdpKj/kI6Y5z/+si6gMOCJOzOh54jJLddFpjUo6dmcClzvdvhp+
J2XEhGb0NcoINQ1TAYpLFW6AQ7KqeHUYOhbdRBzUd7asd7r9ggLooGc4YyAdxbPYLPq/QDOJfJpe
T+AGov4CxLOp+iVvc0Z+BQfbymBHcQ6nbY+XUUBKOcTYFHvf2KKB97h5Yj6TR/9mNUwhrABLcob3
mBFV4Su+rqtoLFT4F9RWD6vUnOywYEpu6mNQV6Q8tnDhu2j498vEd/wPAS2DlLTzGhnZZNX65Vis
iYi8TyMFfQEwIjiwBM4vdsAzUjmKWdokJTclbw3IdPBN/1VKnbal2JiWehsMmnt7JdI4AKfxJUW2
9k6K+AfSxJIfpKp1/bECunzSlT/38kBslVY9sTKQJCI1XJ2tchGRQkqwEXN9rhatGHvfeUmU6i+y
HEckv/Jz7ekw7mE78f/VOY2+7FkUZ75EDQ2tLZH6sJXIwzDX9j4sNwKbf5/Ecv2BMquHAy4UnLZp
LE+KbgEudBvKJatnQJIErzJoAa1FDgDIbIvkSh5N2MngIi0lfBwU65gOrOVfjmEJ9VwGKbVnD0rb
wnwcM+vETQOrE7/wTqsp8ZoIYEvtNzml17/WMBoHVSoEFxXHjzSBuowxVl9WeLH4ILK/6n5LpoQx
ZrWhg5tU7khuPAbaFVAdDNa5bhTpyTgvd600Re+huWBIO7rXHeou2q1k0OI2ZtncA0uOGiEZ/+At
GWUee4PuPdnwRrA+9ewMjrl8R1JPg4wD+dTStCshW+WyGWRXk1fKYIAL6kJUjkXc/p8wLRxIDpD7
z+kitEKi0zxbBcWm7klo4w+XdOWJeQBlsCMXf62x1qTeFl7D8/S5dGqy6DYJmB89iybDRM9xZ6VH
9qS44r9SGA5smHjOw/OwXGt53T9t9tgAJ/jnY2r9OBYjhrMIluvHq4PObMaBGjuic6vXET5EgI7H
yglAqtGYUHaJfF+TAYr5KmcfBqsOmAzjf0om9ZDJFkbN+T7ZGBSfAXrOf5ROxyldWIVAHbKZkJom
EDzGdcqpGQ1JRCoZyLSaPKuFuyRZEHLwkA+yFo1gSyGbpAhp20WSzYbkSS4IXj+rAVgZyZp/16By
Xk4IkOhggaJrj9aTbRkUsm7i/Xnk+DSkmNpzC2rh05bQSkVVKRvAbbSYrM+M1GsgzGDDq7ni86eg
Q3o7pzYEDAe2PwzIANGFSaGgj1P/MsWJN2J8SvvLfcyQYZscew3+OiLktQp+HcCIKNuRBFYcco2W
mgPBLKlJWBymr+CqOQZBTAWpOOYHAXL8cvveIEgp9/GEwoVco0wG+AMXf3qOsycr7nTFkiY58bmt
oYSomNAE0KO8PidBsgjb0NG9fF9hTrPzu178xm0eRxFpVBSLOoguWdcOIPYFcedqD66rHr319lyH
Bctcrrfehoi+Jc7v0BfGeGo4GI7GHjVMsaMqjAmT20V088IwwNi8BTp9FRcr25X5KAbaQefTiFM9
vyrDGbPMigR9jMql/LkGNV84fnB80yKCDvhvXQKZmLwU4Tgy+dmH6FanL5j444aHwrf2rSlYsSiG
ID6SqZad/1B5PytW05DBEJ76lS9lAjEV1ShQXRx3UFlS7944A5faC/HpyCgD3NQXljZSU2K6Aw/0
kx0U9XrjjWwNQPl9CJICLn4oxak9643iTJUJEgn6lbnPZN7x7FspgmhkhN/Kr+afkU+YfAT0YQ3e
RpMYeq1Fcpa4/Zu81u4cwbfVd4CvQOMGL8GJWFtFJglDCF0B+UvKyK3S9qJuCUa11/O+6TXZeHTe
7vs7D+deNqXx6a0A9QM9XDsR2tbcBWuH+Q0d+h6QPIFKjGUv/3FuhbuP3bdXjIR1gew2wKCfkpNY
VuMo7bet/AApeu2Zn46ofCGlSHkIfsYaQEwJNFaCGAAg04uQz6se2UkArPEU7h+hjTb/S6sZejcM
hn8AU0gI3ewqOV60WotG/0/QI8cEJrwe4sE8zNpmUvsAn28CXCw9Zme7S5f/AIuZhs1SA6CuUbgL
Fe73o6QHItroyRk/zmwT7ToUb9kZRmVQ0BsxE1agGEB7NQjLg8mg/tEyylyqeT281MlzC6SYXief
wG9qgsnd4ss1WIyI5/mLyElz7x4jt/Q74orQqGIKjcktmoDZvHj74LI5jIO/eBf+oK59l63bIY/8
14x1Fa8JDonjWyR4ESmU3bt5drf3Jp/L43iozrFe5xwEAvz++CP51NMO/KI7wOLHM1C8TQ1AGY6y
IbB6Vhs7r8s6y3JA39WKjmldjaS/mbHxbD3tOxs0TnHrAsTOo6NsNGVtNwyJUY6MyLMLFlpUXSdA
RNoIhPv+T1kWUKzGlliG2P+qZDFJBuaMQbkowdPZfNO1YE8QNaGmXgpHA+kCQ/D0mu/1tge1VIzq
VW9R6By14ExfwDX0GC0GS2h/6IisoMIyqyAr7FPKS8IUQ0ZWb9I4EooAgHipxUTnDdi4pGXAt+Pv
GdAbE2ZMcRxzSiFdB66R/7djM1R8ayC9SEvnRq1mBQ6CsvOWa/foISbiT8y8kHjUb9y0e533McCr
pacy/JIw+1pb4VQFMbK/wA/llrDxK6Qqre8fwaygragFXrEQAZVVqJn7DEbl40OhEXcO2BZ0slsx
GovvKgionHYSnL06FyPPOsKDnjC3hiKbPIOGQwX4hVUUwptIkDk8al9cjCF/o88mhzff/4md2Chy
Jh9yOpij4O/IDEdZ+vaEPK1Ei6+BE4s/+VWPfI9gb5wfVGd/ZtODWg4gPSgbT22X8xaM8dL2Ow0g
XDlVqiHu9I5Wk9HXSIOgzsiggSjAeqg5a52DOkaMErK4NR/58f3IlAQAwHOJzeGbDmmdFjPe5Yal
yKPmRepH83/FxrbBUcFT7MYXetbcJT5xdxS/JP4L/cMf50b/5nGtb3ygF1pRZpHImodfxhuzlA/R
/47PLAKykrEFrIPFFCLWmxIMUK2k5lh/Jky9Vfo+t+v8IjfZNqyd75LAR1aah+8vk43z5VzGh+xo
2ApTCJ38CJky/vB6jUpfI96jLL1fZRe5gWq/FiNHxk6/xSwIBS0tf+9L8lKA5aoIzxIKzLypRpyL
b7Vm5hoqiwbd5Vs/shI7F8Xw3KD9WmjTBpT1MgwJgDaiXKgCxqMIMSJSGmODQXbrCYV7cDHItVmy
LBRb9xnKUS3ddClX6YOIDwoObSFznA2CBZOXiMP2PV4Ll8p7mXj+ppTgvxFubfbHZteEd3VGUsRg
NPzXEIg/i2II3ytHZYXln671V1K/R+ipaiwLJ0SLVsoPqrlKyUhXyKVkFKkEG1honB2fe5rnDtoN
G2doQwRmDbOcJcNMmiQS5fmqgbu/VchDS1+Lza27PQpQ86B+RKnODJYSo1Se6/CvpS77/DKRGC4u
qDqlRmuEX4E2hm9Y6OgZGrsVC2hUwRQCpIelR6d0F+oYonr9bA4GncPBF5ndSWfDwIg9T6wbkg8g
lN0BVGv4OsEpE+02aUcxD+xaULCEIrW71nXvAyb1iCgIezH0TYzvg/qADM/mjaFaDxhj6T28oD9c
zoh17fwl6KFUsOnorhbp1is6X0Y8cS1AwOqMny6MWYgkFaIvRSc26ZMTQQ4z+Pr1kPljd2hfMuz5
sQY3ny8Durc39Foj2CwWb3rgC4RWzaVxlQWTPWZaIV6qG/2iI/H8gs2Tj/EtMU7+B90YRkAWsP3D
ipEi56WumyRVMqS06RgzNXNF/9hf4adc5PwoinTIVP7ryzaF2yE2gbG3+OtobgkdwDEsF/cwj0Lm
P/74Dd9+YUV1m7uDypciwMMFuCFxjfVeASVwT+xhvIKcowMlVqHz6AkP38rgqzMLKDlx0H3JPwMo
WF8yeEV6wdaq+FfowXyZRmUQlcQ669QEOTMRqGigwY7aBgB1Xhm544BoYL7V2DlJlsB/3o8XCWFS
GGwBardW4y0yg/PwFds3uxwULzTmChCypKhIB8ExJRHL6f9PnN+OECt02VStXUY98shMqsI4sw3F
l2hWhQ3gws6fdtXmWNPXiVN1mBRKyAOYBJcJMmWRm/TQSVlQasNZpiQgHonRN8Ha298EmVu4dlZg
dlq6cRzzfpTJXGUg2xOK8aKLSVzWi1oF2dULQzxwTQSOZsO5OUA0WbcPqKHy2ow6oOeO4Gjwca9D
SSoxVptlmujX25eIEStpITPeMkmm18+Z/1cUOOZSSMnTAUVIFXcSvds6/VaTvKWYqzWFAV6Y2O19
j2Q6EA8MQrgJafZws1e42l/m6auvJpYMj7WiE+G22xTlUoZn+SDs03w18NjauYX3YqGdsNuiDM8j
wupBf6TvsaiVIHc8kEiasqj9M+6HMBbzq8Km7Hs2kTXPml96wnzrGnADZn5YaCOPIy2tVV5r7P2g
AjjX1LQy5AUK4+bv4lGlQi0hgVl4ZWrliTIQRMKWsarEbMi6vY3GFwKV2fvDvizuvFRNtNq5ul51
Kepdm9FeR/Cupu3NKBk2Ks/9FNLDdlr487OBwP0xVwejujaG6/AXD3p89jJ/bzSI9ytT5OJ+J7D5
+f+Cf+E0iAMIIhISB7hkjRpTHb0P7aHYya/IgtYCbnuLw5J4KNvmU0IQ1TAECN8eLSVgKOGEOLsg
RWVYkRAZnlOXC4P8XHx5wTJfrjkky+Sa+qtytLF3JfAYO3SBiJ/1ecg+/0ua7Yn2yZtX8v0I9GUI
rxeWWoWcOOKcp9UYatjUThExudURd/1dT4Ck93wI+Cizja5qYGTL2RTPbAduiwbjZoiFQOU7RtBT
aXSv6NwPUQbvTLyQmdruXCengtW6g3d6V7TQzflGnR9CGMOaxcmvQFjC8V5Ua9iW9qAIhI8yqG6v
6WETyF6j9LgjTS2jyE2fMch9BDB2d+9QqyzqZBF9aM0GqNF5Wre0GgaZwdWFIEnuJ62FmOI2sCUh
b9kdSc41IFh1sK9d0A7uId5UCpWMh8vhyZhSAU2s7Mnw1OxGYG+BzD4b3B35ov1G/odjiUmhWVUj
871imCPDj4m+tkaAF5NMVkcPINIMVXAHtX6ZWPHcE9AAWnGRfPcZmI/DqoH6H1U32eidJiCYCLSA
wmbzfeWJNs6KEj6xS+dxB4jeyCL4raBsYb4JmvtjxjVeXkWWXi4XWY51k1iwaex2gmAyxGYLjRt3
6tX0WuZyaWyiGQghvFl1iBkpWjRFI3bd6LpJjYNgcHF0ojzY+Uvcbfwwrq/4habqm0wYsgpQOg7K
8lcMeTsNBpHSNsSxg/E83IYaApXd6XTGVu4AbFE8erUvtKSenKu72eKHyw8f31mXO/USvL9m3jXk
afBKF536/KSK4vgoLTPhlDb7q2SdY8W8XytyX4NNWfR3cSGDpF00OdnE9Gc02f2ncdfLBG7/jVjD
dNjNTNWdV5qd/OhcF0m6bnK+rpmBfaiJcRNpB5O448Evmh9cran3vphr9bSlpvoy8n8f2VBG11vl
pjXlhAwPPEyX/NnQWmR+0Pehslb1Diy8NbApipVJLmw0FyBHgFSkTSHqM7H0DRHuhau+kzO/uEZK
MBs7kJLhbdSvI7nbX7V9T4ypNOQr+0eJMC8ugmOJZgVF1Tqdo5ZshzKkZZHNNDnJ5XPpLS5FN4O+
BDWycI9RziHcBiHcopsDqekaM8Q5qD630K0/xEepvyFe+C/K4uJC251IqhudFzqYNsbKlKmlSovQ
3DzD7c4sT8iU6hlQw1kMC7SC/63Ri9z9srWiAVaeICtt+BO0o9H+Br1uRM4q90T+cO+l1SKIJR4a
HV8R/zwtTt7KhUh5Op/Ne8XVqFSbARW5mWVRGsqTJfXyNe0BTHsGKX1u49+0CajxpnJTHDPF9I16
oK9O0yQCEITjxjfVIjJ0/P27ycBhXzaJjOEFv8raYiATdTdwOrvxN4mPvGOtxz8YNLOBFpcL2lr6
F2aXmN5bnmiAPe9ZgMaxxw+MBwNMTkVHKwU/mFBE4tWzrcMxwYGnLj+Z3wYvPHlJ/V1bchZuPspr
WeFum8hAryAuA2tPPTPi/ZKp0DgIBRIyAOKNDBlywajy7AU/YawROE4nZLwRFBsRn8rjnXctlD+K
tNYbaJwiz0OviAeemCRo7goO6g+gCdB1KuKNlFrQGmWLRjKoWKTwCYACRVF4R6MXLFqrSMQQD6Fe
1oYe6/sK0TiyQtigWnP9LDJTJ6GC+2BojOMF0ABVsAJlHJop4qI14SAfAu/5bd/2kDYF0QjT78hN
JoTt3gMUm+aAkkIMyCitPPCzf6zP86ympqGrIJH80AM1zYD1l6IpeoXeK8pCqu5/yBvwlKmkVqSl
IxXmLFTGqYijdWFK3oky32xyhAS5Duj6MiZ/XBDrdlqufxxi2PIcUTFb0wvAIXg9PSwtwpPHCiYM
9184EQqfk6y93670y/LpaaSxsjyD5uG+89nQU13eav2K89C7L560cUdiODI5Ol2qw2L1Y1JyPgID
2EebpxyaCrqUCJqi2RsfW1DhX07/G/PLYlga6h1dPWbM1ihdh4Cp/dG7YctY7CPmdRdwgaQwJ+be
FVH4ZooST7UGa0xablp8KBuw9t16jHsaMVWpkq7Jh6H+eNS+B0g/Uo5ErxGJgqew8h7I+69rjoxE
7SvW4yCwszrM+Vdnq9JRHboWSbSJ2FBKl8yG401WJIfNaaIVgTZVzRO756Gl3ZAv4IGTbI+bMlUG
LLfiLhaUqqRyl7mllk8XFLJS1aRuNqpsrXxvuRpVPvYUq8pWyXxjd7YxzYlPaWMeFkhcXIyj7I+o
72RZbTHg2bzCRIhTB8MVCW3DYQpk+pdFm4VISUhl4e2fFEdSwS15GfogpNLn8ZUOPnXvsD/GOUZa
L1pVtgi4QjwR8ey8+WaweYIzpABu1jAoOrd52ia0s6R9X5OFjhHuCcJhW6c54k9aGNNP7XlIvFcZ
OxA27Cvq9VDRnDRMOBzu6gXL08rKoC3Jv53aLBWG7Y6VhNP9q2z57dp65jAFUEd4CSahaQuAuyqO
wew0u7xlzlgoGXx9CRZFkR8b4YF/rRwhAvp5ywOJxm7OYba+cTgWch3lII9ouyaF6DpVxmXqCTO4
H8mYl2H9uao1RmoZOBvSp+mzTvUkGzaZA5oy99zKcu+F6QqEAdFiDSMsaw7RZafpu6vvZm75v5Be
gL/4MFbICq8wBfw2LHPb8tOjTszNcfloCp13KfP236Dd50KklO6/0dialhkib5omnu+WwkBcjxTW
WPqrc8kKRcbe8F/F2QbT8/hVhwjwhthH+6qu/3Ks5RP5zrO+dyT0wT3dIPk/+knsmGBeGvVSE8Bg
wuVWbOAuvMZVAV+3/FEp/PAzuG5eznvAIMMh/S1YrYtMBGspI3I2E5T+Mbukzx8RAI851B9i5g0G
TRtUaYJL78e2toUHIyYIxK9BYU0iu2YDM3fzXzHcDv/6IckCuggpinxB68R3y4In5WwkUhu4wOEr
OT9bZyGNeHW+MxmuHUdIcdVyEa5dlUyr3+wffxs6uO/D7+TLR6LCIafuFMTMYmEOxvXIJOMqJ2xC
KsOoF+2J2mFoKP1urr9elV5GIOJw8/f1QJJK3Rk0qGb4FYgaJdplRvGpvBJ1A0qkfNdUkqU2YHKw
n3EOz1ap+C5psAT7XF9SSBDXL1phPxFpyoynUCOqQjVh5PSQF+doHFWw1bDXfUnl3NV1h1b1KY0k
7irNIoTRSUd7/+qeqq1L4npi4pVcYOB3bmcK5l4lIaOZ3XaamFacfEhFyPCKLR2DGxudhyInlYZN
iU5G81koDkYZUE3I1yUtyiRYdeMoyK3cxiNSEXvtmhLDSES4KowHNhbai0xRqZR8WW+CXyxHc4QR
YBwuZGdatV3VQOlpgzpgOkHjdb2VVleXNZmjTG80ZSKAoiNYGINqmH3BJU+WZVuHoo3DFyIc4Am2
53Vt4HdnaCODAbRUQK0qd4qnD0RmnNcXTw2uSiCnWN2CzisGYkYkr9KuRu/HQgXn/5rWndPpVdrd
p2gKt9yueoPMlsI5Ul6Ca5dHHeYDx71JGFiyL+QOi6g+BgHFqqwJcNxnwuYB6HDB0ZEAd44DwMYi
9wtTOZKlhqsnry9Uka1cV3QZ3H80UbJ2wjmgVTzJfhvkJJlnXM3A1GeKawCGx4U5UE/phzsOtJH3
+4f9Ly04xd2DFFUVv2z2AUK0b3zlR2hg8vXKuZ1WcfFL3h1rxurt5DDZWZSeypSbVeweDywiYTdI
irfTKqiBqsrKl/fsYDOA4kZIv4zEOIDxDTGv9IY7i6PnU+u6BvO4TN8s8Od7BdOSSUJ0YBClmzJz
CydLIBpessEel8S6DbKXD3dK0GY47NyYf37guEnUvyuYi+jXwCqkV8ZknsFP/1ejPKCwzi0t09QU
xGDMV6Fe7PpHndoprFJ7l3T60vzHqQeyly7NM4vM39NPvtXFQEzCVKk5uiWjERL3RsVck9wdo4UW
WJh3PA51hsdfRIUIoi3+nsKmMlEK+HKrshaOoATwRYPXi7gHuHWf20bPZx0vekwXI3ModfDezBr2
ma+nGxKEKwh+t09Qx4ztzK3B7xkXYTL8pJCmk8EOW6DIB8yR6FxifL7KSx0S867tNMdPrLrIs73o
6o3s0Y3eOnC1wRg/yMjZiE9hejwAXE4zEWG2pq/FgHL3eATzpznKdc+Fx+N6V5W1aPSPmk9Ztodd
cEboTfAbQwjS91EKRrvUQ2sxhHNIZfeDIgMTSYOVLV7fcGdjh0TNak7x0pMpymAhF9Uiht69fXjw
gN+MfimK5LZLHWJmMpC9Rd1TEtgcXb6c0ShcWfbDg1heMhm4TVZK4SXkMExeOfKu78MCXv8G48H+
ezFjwvxVETNCrsLd/xdL0WZso85YzmfYMCL1YYKXlgmQfkWGHRw/X5cOj47q1/nLI1l2KwqeoELn
P8E4BErGgG+FpefoN9pY+zKCX1AZIJsNCYQJ9tZcvFbEpluwR7x5qN8vrgZ3CReYH/zetdoMZqdI
SPNv2eL2pOkqe6MqZ0ivkFV/oMVrcArCBQ+0sJGVaCINBGWc3nNL5/5OY0Cmx7rZrAphrdOLgrMg
WiOZ5cZ9yah5vK4Na4g3wyEIgAUOvnPcuVg87IVX+8lwuEcAUuHmIAS79lGw//C6tdZjIDpY19m6
94ouGy8Hr1aZM3TqLdQP4GOunSeOlqrXWHIOD/XKn9ZUl33RXlK6/WKLbmG2G5O8S1HaSit928rx
uzX4kB/LHYiczrW7WVBsddlvoAcvRI4VKHqs9t0NTda1N05UQcLn868nF3QXpYXQmFCuaQDlk6sp
DZsMJa6kiEXRH+RC7K0rinzpAPmpQlhIJaKsF3jiPU+K6Mfz3by7L0Ih5l5UFQmqb8dWLj0q8LDB
zDJyusOXr8ixQlB9UqqqrH8iKJxeEyIpRLKpwnxRHm5les4sMNgX6pw0MsNTIIvRcN3SgDidSMdh
yD/JIhwHPn+izB7WOuc00wyUFxqNiVI/FcD5XtAtfRoMVDCrjb+7AmwILIAGJhZ4XS52VH3xp2K3
qaSJ6e+/QZx4pffbLUbnTjVnVcm+VYFtJHAQmJQkPLRqaRsfqmNxCdmPHyrrR7zztSpzXESr/LSg
vN82thF5NwTj/Q9U8ZJvy+vLf7cKmUR6rujPqHRwQaRFIvkmSxcHCV9b09d2TCrtXLQkary/T4A4
QxD55fcwShxhZ5Nor6pjsTuyU1Q0c6PRC6xk27157P19k/HQA3kDyeksVnYzh2SawiNXIObpmSm0
C6qJNhN9Gs9iA1dpxHqa+/hlfgOt1iK2/7X77eRkZr8Gkgu7X5c7xYo2Qs/IhVKpWN+keXa3Icdk
DYe31TKZ/1HzuQKccHHIORkkrQvp+GWwHzYBSSuW1ZocFYTWJ0zoxii6QzYZU9mKI3uCHjXSmoGy
LGXhE6gzeRVSRUWfqPcqeX2UZSlrJKrKjBBOEI7qKyuN+lKpz5g7fwiX5B5q7NeywRhcSC5xcJc0
G94wToKPUhjI9WgNh1JlTfF4rZnwuXlwLlumDojIjD3FQ4BozA3PAgCvt85zEmet7SjR4CrQFgqo
dnfB0o7+RFvwSxXHgSa5+yZ2P1P+UOh7rcz51e/Z0mJ2flClHkmZ8I4hIwZ3waJO9TuD52cjteK8
4wIW+RdPKjPkl7/tnJTxAexFi7UeYsEOcbA7DV8JrGJTc4yjBn6PSMJle3MxTygNJK2mZIGFgct2
ph7NwFHAVCoYUi4OfUMugRTVZhY9ypRg8Mb5hIiZIetE/vciPGUCUnHFPli5zReH0Kqr9sh5XMy5
mGSG3cjJo4639xVWR7ns/G9HCUzSjMeIXaoJhJ9TC5OUj+jjJdxhuBlXltbIwx0e74kjRT0NYGZS
xrF3G9k0FjES96u4eb/2Q7rmkwm75GawXmn+tnkKobmPDOS8Br/Meavk8Tf00iTCaDptFpNxWMLw
YwZDyxqRZg3NVi0sdGyMg176nZM47VM9pJ9nIeiohjACir06u/m+S52HsCCvvM6Z0xeSoiRcfOvU
wcs4VlZcvFh5mXfcfOyupyMnXJiKmDLQzuPyz3xjQAseJYeuNWbAUnd3UWvfvMXQIZsfq3Te7Jug
FELJWnouORfuwD2Kvlw+oC+H8cA2n0qoge5MmdJOxiJ0AMB5J0HQXsC5i5vDFJZouUEk7QdO42RT
aZ9L3hF5T1zdsmmVBP++iVnJFwi1tzji1PfeD90L4rgtKli2KugiN/RayarOH3wKakbXCA3MJomn
yoEYrNvN1sbTT0M1p2yOKnRRDxNSUuQk3sp/rTucb8gol7bDde/s2bewwQ8HFqTnRS9Kht+42XI6
R0PI/pGUCHuXklkbWP6kIP3XfoFkjiGA4YmEWdNI3/87Q8FSzmWCEP7kBhestERUPbeXcJInjGQm
RzA2bNiqmFE8mPGzt9PBJjlYoX/8fUwFv+JoF2BEhkQ4YGLX3APBQ7E143KvED2G4oxl2atGsMRK
7wPCsQBoeJdqVcQjrdj3nTL47kk5VXrCUTdpEtm6FfA6kSMqYjLNIBijZaIP8jPyLUh43nWJJe5h
JH0vJvuq5Ce2LP+iV7zir/y+hxYvmdq/2L7S0KjOOpXciZBeAbw5B8znUvSxYIbmW4hlz2J8va/s
7sYE38+qsUE7cvYl5FHkdbH12AnkxOpONIx7Z/SqYYrGnEgQDGiTvBY5wn3rt59Cgumu2FpaC1gI
vkwArMtytppVZ+YkV4NgBy/gN8kBDsd9qwiiDljX3M4dBWUyJwjtRqDOFY1efYBlb6Za23LVsje7
yin/btPudj/kCA5jqFu/XScian+5cfc3949Qw2ph8/4VIq6F0BvKB53sscwPFI7J64rU833jSJp6
OnKGtaBQvd52433qvNEAks5zET2hVFSM+weLftJ+GCGP3Yl7KbvTQgexxKG6QYEFXXoc8qCaEbGl
mSlNF3RPXGctBr2SsPX9exY/E3YqkL5G8C3Vyw+PboX5KMSKIpx3mHHFqvJj5OOis22CF4k8Zxv3
85U4gsj/kyQIg39QLWAwT0GnwESuv7FPpzTozmXQM/Cwj4x7C7eb0cpsnVsa68SDih0jpPHxcnWE
UR/eKHPpgVl7hGtCZ6NKADea69mGv12tN2MJ3+Nu/uoP0/2ktcSHiCYk5MwMiFl0KHT9d3Tz4U27
XU+LPqWHsojH0Px5d5zlGUoCTQ0JQOjiU2nybZys2025aK8n+Wj1RuO/Vkj90Sxf49JB4ojzgsqQ
RiMl6QK/haaNyhDCA7/PwC/4ls3EatQIPjFHeeAaYUxGuS+p2TOrbWyQF6D5UOTU4HpQIz48mR2Q
Y4d2jxW58fMSWtVcd2m8xGMUIupXE+OULQcUU+WCO3D/sxjcPPYZZK+PrX9OI/l5WAJS5h/BcSzh
5FnHkGFHyN/cpGZHjApLlF6TJ/7LnV4MapWxdehpjV4gmpwD+0gjbOzKknBt4gm+YpZeE3V5ROZW
P1zub77+8WyAWFosM/fFP9poiC6130LjgVufOYJo38arQANaMjsc4lL1wHenszu59Arn+db4BulO
gPPl5a+D8GoXb0/dC/vwruzeL9/0hqKNa3PmCB0QsHgG9s2UzfSBTvCYVJlmU8/Nytsn919MCC3K
NEG0MFPulI77zguk1prc9BpBnXTaeTvQQsW3ZWVFj5WvWDinFTf7kDcCrL/aYKgATXxlWVtYKGjI
N7fgCvnWhWcQNmRLTbdH0EzsUi/cTiyvWA5ChSRUN3Fzt++xOY0H5xsNVm0dc9iSO+5URxGHXVyH
8byNKk4B79itvUarOE56FviOvr5wgaBeA4ZBAp/0RUpXq3YXVcnUciySt72pc8Sg3LbSYxZ6viiW
QacrUWyMEE1pRA3MadCpk+r++9X9oMAhFzoUmTBJXCReJOEHdVX/tr9xYW6v2Os0Lu/E9qDCZaLj
7y6jFsxbV2/onqHw8rtSXKrRsgk5NH7jD4XkQVNqd6sI+pgkRLj5pyItg5y/H3s9gVOqkvdtqhY9
on/Kas77oswDNHuR8/GkbjYT/agJwJRrrAx0dG5Kc2ocklHvbszApYbR+G/9YLNR6AUOL3izUWap
GIfS4CXGEB5lCFTBpiuGfG80W7q36IvTkGV9EYGcO7YZ7aGbf01LX4HuFRw79Q0OJMcjo2vpwugS
3wBp01POP+fdja5/ijPbykJrXrToLMckoIcfK62u+o+umK4dAVm9gLXKGUtp4tHye7bEWkk9ArMO
ZFJgeSkKzccqz7yEVl2swluT9vxQJHjhwUJXYUtJ2AdcGsulglQ4RUxp31Amgu/DpqZ8QDss0xqF
6QxGbxGuhLX0qoGiuhiojj4uAHfEgg0XD30MoW7CRpkPlI1o71iiHXXbxTYptJscTmQjzyZADOMp
TjFWzdodQarbxJEh7pbYECJUx23NVYvs/yf2ykTUi5AyLYmBrhLjseuC5zqiSGBi1lL0Q3d1sJ38
D04bU49OykUl9BRfNuS/IvchNWxLNCIcHsCqu+GxtDGHD9s4rArC5a3L7/r/co40CcLjErJO6NUl
4aGmB9PEh1mTUnUXFb5RLGSuNjI8FmAZsRz6qGZU8LPhlVXHiuz7jJtN5CAksee+260Xk/IAw/h7
joJDh462UiLPzOV1fzTNPBJKzhnaVi+ircvgChzPOKxp5DvI8MFfAXscm2vRF2ALpBhUWpiKGT8g
ilhkUXN5Nqb6liU8L57l2d6L0yaZKltyfpIlfnSuX7QjSozefNifqKb1UkO46VHaG/47IKr5gaoW
TYUulzQcVzEeLgzTD55tf6eq5jRpk763SvdN8ZbKXD8KucawY2+iSPWJuVZj2q2+eccxn2R+8OA4
om7H11GgUDWrCDu9rPiMeinbyylbxq+fjE66L6ZeQbslIiETPn/ewSSZ7t8JdxzYSkRhtTYP/23j
wKUwmt7NvcZGFF6DNEvfosyPUCi9FW08yICK4Mheyy6HnbjZu94fQhcnQXE6YIqQGegMtJKJksc3
2d48XXWssg0Ebt9PX5+3ddiMy37MnYOjqE1gm59VxtnRoTxhtbaacmHDaF1Yy5lznvPc7Z0VOjST
uNbHMwwU3QiFanfkFdmfHhBbwUl5R/f/hC85TmQylfDWEA9S4IQurh+Zuu7v1Egaotf6j5wtDesR
ncF9dC2zmqrFO0AcjQCiPMKX2TE/G3YMsofOBcHE1GvGk/qXcwdcb5Eu7lIcNLS4Wa3lKne5+M0y
pr0r64oCB2KiTQs7xAz/5JbtNTjVpBPCAF7o562nEJYUjTub1n96X/dEThp2zbzZLFGBz11iMCSW
eX7BUD0i8+nbQDBpUNV0784DR2QHIcErft1cpZkuC9sAJz8jdcrjJRzMUAcg1qgKBGexmWXmNt6B
M5HuCo720qlSO6tic8ImbaabBRMqywicuqIyRvbsKuRyKxC0wivcIz7lZcqzKvGzjCUtrcrkyhGw
GcOeXhwN/dcL/72yqG4hclRfWp+i5sRpKuLR/NRyfAJO26mwI1PMdqfa8TfbLNQ3DGjfUcQfKVRv
HOSo2xu6Jc0i8OsP9N+w6WxNPpRjYuEiXm/zCuaIENJUWxP2Kdtz7j1Yvjw4o8DsH12EAv2NsJ/V
lvV2KkmipMZi1sMtWksKwb8L3xcYwOedBHovh5zKv6aN10Bom0lwHOYvhjFuxVWc2LKNbJwP1Qdz
Ae285TRFijI6yKMcN0O2Sm/ptdxh9hqsEbQEuHq01i8Um4q2uH3B12RNbNiitGjOg5nV1P5TkqaA
o8lx6p/al+A8DCcKtZ86itD8voKgCIhBsLEACsK3P7rKHFBcUZ5SerHifZ3YTVekQEjoJyl4E8BE
bHKF29ktMDoKtrWYJdrFr7SGJeKloRwrIC5c7C6/FY8f3nOr0RDX1ePu3AMnuV4ObgxC6JSMI1I/
HLizdFqfEcMvfCcgCgUbpLrKZ5PwX7CYmOe095h0yp8ho0oLdB1XBx4wW+i0wj3ZVQIqFY/o3zZB
ji/yQYXpChIHzYeSeh3tM+SvBAbMyS/a1ka7y/sODPWmLk++GlIwrCjVc7b8CYU1uqX62pYzmqX/
z3v4+acq21Iq+hw+9/FRB67IzAPhLBpCPscg2xMx6PG5bYNljK1shBIv3HNL5nmnWh6CHUC53T2u
QL7fuTNqIUjiHrt+X7YNYls3c8Qd4759KPh5bOLYFszn87BimYbBE5pfu3H0/r5M2QbygKWNqQPD
JmPO+6r3fr4jJxXfH2LGbISUfcLlzhgQ/OllYNTHXOMC+Rfg8ZSO3Ytfg7SRRix7tSrZ3rRv/ase
wdVWtqvhlsBhV0XzCUuKjwx4vom5yk8hLMV8CcbZsY5wP1Yhdi8FXEQ7HOdVlJb8y6Tj6xaMhs0u
A0tAo+nWqs8Dg7UMw7LvFwMGrpOYBSB4ZxWChw+2Kslegij/Xkh8ciQFgigXElLqTpmSV99dxxkA
B2URTCuCy/VhIIz/+4jhkWBHDhu92YmNyqI8CD6CsaJnKTo/sAtFAfOOu2Ca8bojMa5qYEEvGLBj
9NkaPUWZDHbGAus5ONgmIjWnRzgfaN8oBWCtSVdk0qcKvA0v9zd3zDgVmP2mEzFQStmKLZOR9Hm7
9PSe9eBTtbi9iECDAos8tVchzKBT89OfStPVWyY1cVcUBRf/11+UXdrl6kVmTZkPLeSQNTVJma4m
5n4gGtAusTPkHgn2QqdSl4iR0S9fsKkJeO3QnFqFRicHTfh94AlKtEQtDxJ4t+IhVKAiWbdq58Wg
gwenwXT7uRASFeEgBIuW9xqCKVdPMr1FaLTWd91mtKWHwvi9KsFAK+jl44LklNRlEgGEX+XCKUob
bkLtXSN5usa41q8CHFMuwTdfPFA6VdjmbSAu69Kfv8ayNk+aITBzjxvR1SJ9YaKqry+t31FVF92g
GjhEeaYIc2P7fsFQgTo3zT/EeVatp0G0310gzQI3Ne2jOIMI1RmDBfNgwqmi7PPs+Kj/PFsegSzs
hMPvwKoQIlqvkd9L+7M9yFQHxAgsg8FZYNCmjHuZN+ILydrRkeAMtPhGsFEi5zy/695iwfwjHKYK
NZwJFkZSMrP7Oxu+EKZzWVtbbQwHGGaIelvqrFJdbqCFsS3Xc9spzl8/zco+5QU7ZIisJMlekAEk
BJZpS29WLsQW+Yv2bi0cYAb+1Rn+bfsGj9KElR8RYWhiAMNJ92fUS6q8rQMEcaSsN92cgf8yBtnp
W5DA8gVtJV4nB2yD77b5oyhugZTjfPOY+2+VUnnDeeOqBDBUXq6pPMZBW/G38GexsccMawyuabaS
5wylmpMGQvjhRcXojjD8WwTqBY0tGE4NBHiAsDD8s/uhPGovbOpbCOOwmvtMME3xUNSVrltkohVz
TLMEF3962NkC4CnXOxdR9OBcc4ryXggz2m0cK/Vd4Jspq9WGKGAMjIFVMA0P3qKMA0jBjU6f0ujt
6k//eeJOAUML2qFTJULGTaYo5dsg8G2a9/OyL3/w84za3kpt5/Mfg8mH69l/wT0mxLs3Qr1TlNpA
UMPNsa2wJCZmjw88TWEtxpUYM2lWe/xyPbMJrO59HpGw2IPB7Tzv5FpFduh0/ezWGbaxW4wLqoX2
l3UXc/uLtOlg7yU99fPq10WzYaqwFSs8cg9m39Jt4umQcpgK83msrYt7twYt54OTAdsCWdmhTfVC
vn4s7SonYrQ0Tegsye6/tKpGhCYIe46JMrdjF2ctA0Jyv7tMlO8j6/qScwut4L0bQejQE4D9QRtk
QqDtkW9vWEXF7tZ6PPGn1i0WBq3b8Efe6ydqkOIfJJDIA5Ze4RY9vydGJl+mOnPJijRUSqbfms0n
rzr5SrT4DBy4a+xidUfcB9MGrjlKheEu5SCvt+eyIQ/g0rMUjGfx2POn62hmI96E2tB9JUDjw9sE
N22KOKV1u0ELQdlXMqvhwX8eswrhIOI6ka3wasl+Vv5wUg04WD3fKIENzP5ko8IvPnW6DaC5gVcY
3/ZL0bhWw3mI2Jkao8ZUFAEAOiIjUOyea4AG/wy6DrEUzc6EL5sQqcXsdzsvsWr0mCKw8fsN227d
j30uDPv+BcW5C0xU690pqvyUYtE6YLX4pAihlUUKoS/Z5NEagQI+/W6nK+oTztPjHwp1PibGzkzb
toAERbItNLAfKpEf4cQ+nc1NTu1tqwSTJHVdV2PeSFYVK457sAkpPllvSQiR1KxEGSdTuqDh5uAO
6v8B0Vwll0ZvllzUVHz7VaHuoFAUmEtFBL7BpHYVv/K9frgdiYcgz+n/wLwWJKNmgxGqN6RIGRW3
wtZuGSM/ITPWbDosDtPAn9S9jRiPKty5z9LOA/Zq10he3uPh4BlpIWygTrsiYXCf8d5A4PA73Jy4
3QzAW/Z9r7IzwHGONb3uxEgOj+qcTCrYZuBKbcvAxMcpEXEe0zgH1SeHWR7sbX7GtUsXyB9yeYAz
UtzpTfmXgkS1+JGLqTUht+vXZ3qdIt833d52SBoZ2CotG8I0gkEldY1Xgl74j+gvHj7ML+XnzXl3
KgSAzyvItKhIobqfg8wwRWmc7glquvzNigNaD/G7PZmnI1OD4gG9BKi81opsmVYYNaK296qNSi/w
jjWkBNqfwkFc/qh6NO6cEtArl1rG+PfjxttWifA6WqRTJIg7lS2R/kUMTJcGJJA44LWf2W1MzIS6
MZmGOvg0UJpfeOYMrmG//JMxCWwCLrjQm3r5WOBLboVH0U0Pj2EVUS0WO2hhphM9yhmWE6Mzw90y
cTw+kkjGLzfzi/JopDgW8+vgzT7XMTlkE6CCB95CYPk4s/2pleWNL+p+Wws1x4djeAMvuw649uyz
Naskyn2T1gz/+Ega18JgiPBrcC5tZL9AEmXkhB7fvFUmjws7rKLaHQrWIwaTey5lPlHKdWbVG7G+
1w/HN3N+VPkqQMAsnLOM0d31zMLLId+b6wQOyHDIZkKJeAHR7mcoN9z//Jpfqp3a2Ylx1qOzFLcc
TYgYfYGIt5ATzZ7gbtxSGTMY+z0S6YT6eUVXoqKQG6wNKGVRhZjZ3Gw8KtU4y2Cy6+3Czc+Wv6Lr
lfISETP5fcik/Dd5F+frKwNwQ53hXJ47O07uUJ64HPil9/i0Jbyn+Zmpbuh562xYs+O23o5xXA04
kuryCJd9Ueh8e2SpYltLCKj80vTYIJSlMgYq89bs0mCBfuXcyCY5BmbxUK3KOohfKv7a+7huLNqK
XO0r/CLplEs/0ngUzJiEuy/HnubyDPK/a0OBMo/wAEO3mQ6CfrkW3F3DEP4iKlXdZKWav6/Z0EMY
wLh83Obcc5csh9O2kttMi1RWWaBouAVgJ2uAlUZM0D4CQJkeovYLgGOQHn8RuIXQAmlF9z/nwyUd
ZMc0Sd40YZF0ym/bL6UejllBgBBP4qug3fCOjq1Rp2DYYB9ftV4rB7aK4NC8/n7FZWma80FefkzJ
/N17xIviqnX1eyDBfR7NABO7uauarka3upygLoZ2mpcCn+pDbIeErctMfU3kD77LowwYjJ73wkMn
jQfri6+2dfh6M/w+kNxDWU/EnSrl57jU545jpJh5e6T00G7U7oDohcsAlgmP5pzZ8zYjNInIED3Y
uwFq3eHE+ARJWYXTOpiVwfIuUnMitCni7EknKT9vv1znBfHGP0qCm6z15msU6LtnPIdgnOWa4iMq
M3dCd4/oVkBN0HFUwt5vQYCrKFrZk291lrCm20Ui69jedQhRVUz47ae+TyfAl3XsKY0HJA1JK/9H
/zpOV0L7Ttbsr3/9fZksmchOGeYV8CJRzJKUas4TgvHJGtQvB/lWI8qYAyU7Z4EmxtZKmN6/ixCt
j277Lti8LGeeQusd03av93DeOUQHu64zEFGTpHiaEfU2XwINQGxzddLHYblYzkncyqbZpxCPGBvY
Sxzx+wUYyGFnxSvHKSwegZ2QMeHqNdKRz/y7mb9OG3TWuKrctulPtla6J1QU3sRmcuRBSHoTJBYc
FgkUJQezB8IgF1k6O7m6G6p7715YVgZtCzu2qVxvhlRMgH/Y04Ms75CbJhU3MKDb5Mg6qcfOkwQc
2RKZNeeI6pEvGBJ4XRS2AO5Sni2h52N2mBx2vUzsL+feV5uZyJwFJI6qXVBDwg/XW+Gny0X5YG6z
jJSUfPUJ/VgNz/RPjE9xoaPvTwJdkgjHK1UVybBjbkTSQtiVF4ftHrEhuxXE74mGWsRC6oqHv0E+
eVsmd4FISvnuBLEmrrOaa9p3brfIIfA85vw7ApLUx0aODJNny62OhC8J1iEi5BTYQb31ldQpn5HF
lvGYJaJDwbdDwd1xMsn5u0P0jUfv1znrz8Siwg95lXzXvCOZ/CCWEjuByWwu+b/JlC55PHx//r8A
JCG/aXYZXBnmd1R+60jZ8Nc+WSWPMU54GXRK7ISbnY7jXG5b4Utblyk8cTwaTuvgyE9WRw7ZD1Bs
S9BVBIDtJNCNrv6x9jmtaUZpv09qNqVqHjA/ijwzZ4Z1pg7X/4rdSMRBF7F1rCv9yNhoJhdwc+xo
FR17zYWLoHwlBBsb6ok518u0LSVFfBxd74ewAtDOwjz0bcRvgIF6Ip4sEqc8NUGLcnwEi9g9A1N6
QchJ1nP72MgQtb9ZqOs0grapghPwYLWZb11Gk586iSbj8IJ1Fu+soKYZX/0/tLqoMjmj6YfRmuzK
KXTFKVyAmSB8Xmy5gKHZdaY734MZk+khKAjanH/9h6SiUhfNNV90Zj4FdgEQlnkSKyqIS/v6vu6+
w2XurIW6KlvgsfjHgmhUiWUizZIkTKTKE69YfES4QT4YPz1oD3hlctnr3qx61kffo1w7CP8koMf4
8KqgoQkQ+/SX++yqEy9YGdRL4l8iqTTGPbnNKDNSKGNyYE1KTXolxTqYH8pMWzvSHfVEdU3MgaCJ
mOkJip6iqHiiY5Zjl8rgHaCkjJoJnt52/bMg+bbooiMj1pVLJDtrc1+IV0FUyK/C3WJzRT/NjGHd
uEPpl76pp0x0i3AEEoy/nm31UE3BndX9XJKHHQ2WmyoMoWIubTsdqbZ1btDhSk1+i2z3eqavNpJ/
C6pCQ4nv/YLAIbS4N2hevIliDwTM7ylmOqn1aBFmvnoTpal7XesUxeWUHkmZGUKwQ8HhaLFFi8//
UhvHq4vjixdNS9y641ABRb8wIHLS5/Rb7+y0pnuTg4qoQFgKVlvErG6tygQCkgM8WkeA8BSX9pHi
2YDp2aE/M0nm82LudSo+4eSAw1651BeYPK78zX9taS6wxGfesw/lpmPTWJ2bB0yz6sMhXbBu5SD7
mKUX1bvMqrBUUGCKds5O7OaRcpgI2/YiXKtH2WxpQVMTbd1ME98b9ppIHPMJ/7vqG05l77kr6Qas
7r6BEQ6PYp117Jev1SunAPEwiKwjdgVb8BPEwLCXL5GRJr6n72JtpybecCZiXAG2GuvJT/mGXqcZ
ddwWG3aKsleP+zvgfi46xfll+4NfSInbZcJWmymY3BhB4by0xb+9rn4AePlbaCM1kN9ueUi9WzvA
U83DE3apX5kbFqEhmhtbv2LFDbmMZQ3t4/nMy+O7TpxG3LLh9EuqjMUykSE3v3eRcUHA99XgDE9b
EFGwV53IPIDJcNliJuhEgAr4btTWnjij/5cLLQUvotTXWw+yDeIe2iSxoeIxmMExn6nF7ipf4B5J
KZL52yf8Z/DMtRqhNmk9oVL5/uqykh5ySjgkXV/LqfvaRJiku8EJ6XGjAbk4Y0r0AbwJcxzvnNyC
HQRSXzthUrmRndvZ/yWVgrVHO4OZMVFURUJ1Y40Fww/Tl0nt4GWhGuxhA0GIGvl6z725WjJy6Nuz
MhmbijhgpW1Mj0kQWfCHpVkyncx5SLJNwwidrEuLBiG9mXJjAzj8h1MggUnUM91AWXjawJ5io83j
8+zA5P1ojpLdaOtmcLATwgL8KePcpbFdBzRwNLsbln1EE91Scr4CqNAekGRKx1NR/7EdKU5DhytN
Zj62sCaHCyHVPY+n4RhiW8uhfuZodonRLT8ozLu+DfNS4RdRxUCF2CRkN2Pc9XaRdALI56teVpIx
njf+9aQi6dzjhvKFhXJwzLF5FIEynXZaznoUzKId+0UHjaem7VhqSSu1dGVaofXuG5bWBBOqzfdI
nuP3sgpQ4yfyqfmRX3sEH23iERz6PT+Jk7Cwf8nURbKy5TCF3EvxGBlelgcW0lnaK0PuSHJEZAbG
XYG7LmrEtDUdrECcY5rmsBXiVLoe1U2+GKTvhsMh28H22lgZPM//urpE7lROhXfnkDJIH4qg0Bkl
MpOB+6d0Y7pY5TTKnOGcvotwvmWTd4ywOOJFtfjtmkOVTPi2way5xzB6xiJMJ1W8pAS7m8yKQBFT
OMC5Qtw8MSwJy7/kDTwKBYRHrw012KuH0VJPlFRNBw8oFkM9Ess9ACvppFwnqz2B0zgb5yleyOF3
V+vAZzjQ4FOWzmyYsrxzzGdvcpTKYRcAez95sLCqWaatDJWd4JE0olROAjr5JFauKMisoVbgHWIJ
4Ol1vFtdyTxW0nGNV5tkz2Arb/DvhnAPz3pSmy5rkC1k1fC+duIbkhcXNeL7JeMN7ZhvItAnsvcZ
sBzXfNOH3moQWhGD6iJJdgENinWOE46U4DtfSiPkhOHKiglwQgaQvnT6dS38qqZq95EzO/iuHiIs
IeUjcJgtImdSRgOFfkaJpsSPtuxmNSPnlytL91OQTpmHYA2GSd4NaYcSpndvq89mmdeV0jeJtmto
c4Ci6JX0dTW47bfNW8DM3HzjFzYKKKlekNoAzxzx4ZrgxIajpDGGO3l3+wfUUvu9N8DKQ9roMouu
T75uh1pxd+pggacprDusKCS+Cb/J2eawFN1Bxe7y+zvpMZCulEP5tmTbTwifjdSMXUhfuwzbj4i0
fWszLSt1fhYpb3LR8YIhMRk9Hrk8hSfd54hGo7R97KNwbSp9CekbLsBCxBYZNlChajpCoEZWiDi/
2A5F+ztqodWKWbhBL2dsxMb7wAvh5AFwoXdAFwEf8uNxqnfQYIO6ngaBfRViUVC5n9O2AuvzC7Qa
+VHlQlqNAWC5HElmi42+q95N1SDIAdwUwx1ufBXfdycsPPzHAIclHrStKCXxmWsBItDna1da/HiN
I1+hhmAT88ThdKprMEZAKwDGiB9dzi19feex8hqk12kFQG+1jTfXAflp4eMrhg7FCNV010a6MM2e
e8AWVEgkyUqoIrQoqdx2VZQmWYlrmO+7/RoghqiR+M467BAMU34ITAWZ3mt5YFvU6Vxx/bugJSGA
vleFzB8YUMJJg3AoV/MoY7x1tRkDsCkx/vu/0HcXF4pQvefvAaXGc81rDNP8LnZxVzTltHWOfI/R
X7zu7KEVQg9Ogk5d6tKe9xM6L5GQACoHtXWwQ3nZMhP6bvVEy3D5NTw50p6u3zvqN/aFIM+NA9sa
Wa8f8zDlWJvgmRFnogmFUKmWV5ZhG8lsb+926IzrqIDgBXfmwUvn09qBX6jekDM1uf14XrFjfORC
eSYiRAS8e452rWvCEfbs1rtPGySse7yAhcRqFPFI/3lmNOaOAqwfdDM1bWIPcHErBC7hVbbjSCC0
NhTVtHu3pSjbZ7IFxj6qZZmgCMEmIP6CeWdJkI/PARHghO8s/L6/EepN3Cz0VF5wTJKBhJT9Np1I
cnpgeyS9tL5jwK0L9ug/CxB1kQsT+qYBzBP4QV1REunmgbK79l79/eVG9OA0APZiR9G9i6+xuqEF
6aboG9ZuA+yed8374t0yy2GTYQHNrTF3J/QxcbnRZFn/NRA7gLF1utF0cSHQyubRDQoJa7pLNNLL
QbZ15xQc0BREBVhGhy25wlT3zX/z3PavI/f4bbPRZV2gStNzSoM2DVNi9hgsn9Tm+EN4fTWv1zCN
9V5xjWqv3dsg+n87nPSPcPhUcuRr/3myN/siySdFrVFJRgmpaA0raNSbI+m7xq4G5krEnA839ygE
nd1hyFWvHzu1m1/R7pQ/B4T8l/SaADKU8RTOBID0K8GPMxf3KeEOacYMqF5/H/KIFD/GE3ND0bji
aLai9Hfl7M9EeHvgt68YO0A99jhFEO3UsrwlEYfzpzZSMyET6fJpoOYkQFV1e2fwAEUcbU+qKKZ3
sk9y5cPggYekhn2wuEl1qKcTIqED1wLUiJghpBnGVRxOIjo+9ZiXmOx7Nj5TrpKphdLoSHTtGo84
vW5zg4972O/sWTHNEbcJtb9uASAwoOcWWT4BhyFT01P2fFV4ZGJ106Z4Uxi8VauNHAZhZ1xJLwt0
op37eHwI8NJyVL76MCTeUl/ElDQY6j3KJxarcWd1gAbCM5HRwyupykJcf2EWLTCV2c+OPGm0DSA0
fvIvCQuZYQA9p6XR1n+vQ69r4AtsW89GXp1eTYaoXHv+FN/e8NISiAKBwWF7C6/IvnZ/5os2EHQv
yYpUiJlHBV+DdkQBcWSSiYyYg40S2YrJUGhFABpJowtrBTMCt3s1BHAFz1Q3GXnMMnGF06c6WhBc
5i+JZhls7WghvEGGUnm27YB8+5OIFkOcvKUmMeraztbVP3e8EI9GPTyHOoFibx2IIecHrRfpXVKY
pIoJu4whKhEqLD1ksdTu8GyumZDvtf0JPiuDFzUDZO4dX/KKHur/8dZFqftBuUwT5I/UeEcrtRu3
Y+JAlahaX3qFie/8N4hSe0IoihaxvKjEq/aX/RjIBngPJV/xUcRwpSCEaq2tu2xZhqLAgViji/tU
HnTRvdr4onpALZbukdNwxgjmkFD3jx1lMUYUm4W1AjVJRLyNiWwANpkxajg3M5zSc7yNgs86AzJc
joDWoX85ZF7h94Sz5NDPrU9mD9LcyX2SWw2r/uQl7e4agE2Nj+EzpxU0Z9SFqDGQaJcfE9Ur96v9
O57/X++aGPs5xnSHqXvp3g9zBqmxSP0Ar4QcvsWgrvP81w9NO8XLRZSi7ThpTa7B82YmQQwFRbUU
BuGaHpO8KsDjyXYURzPP40Q/Vea+nsT0oC3tmmsVDEz7Xrxtz3btJ1f+bjQfEy7Y7xc9y3Fngmq3
EcbNRMJfOQoQBWngK1Vt3/jW3m16c6mDX4yXI8lIIaoCdiD73p5YzhHmw9Z+cF4zcZa1pI0CbqaI
ZgbHK6Nh0liLo+NuBJugC1G/Co08B7fI3WDnOGzL08fRta9g0EKHPmFQ0DpqI27rlHi1qs93XFWL
MB9+GCv7oNQILQe3qd8z2vje1ra53LANA2NAx9TuxVifRtASZlnF5V0VSzjBI3K1ARPQMPqQrikr
OGJpf2MhEmBEpPR4WZU8JxskoD0cvZBb05F7MGX24xdtHQQav5iasNoiqMlT7YfAi4/50yAcb2fC
tIE61b8PnoDqt6RRhPNXSelTKE2eO9hEQP+NHmH5h1oNhKTywi2EZy14Aloh5wfJ6DuuIfLz/OS9
DQ9zjGpkn7D7TyVg7tYyKj9Th0gzlHZwYtt3OSWMEWaucezxwZReNTawwLAnAcx/HgZakyrMpfea
xcjKEOSC/jVCDgAfcOzLf+AHB6jABB2hMBcBP3TrmOC+5kGg7H/Qc9Il7fCfzmIZ3n30fmO4XzV1
XeEpaV37o/Qh2XQPHiYDdBrK0i9Ki9AiEtez6ec5v+DpTKicYqFanayh7IAuFPxS+a7dZuOU/YXB
xiXxywnU+vNx9Zso5BlcAe3wF3n61UsmHl50mt8cQfmWoRD12lZIaCoMqPl4Pk6XehtwPwPOQCos
7FQb2+QtZVP3raAofFeO7xmsNYB8oYZEBZ1/+k9MqTKSjc4TmS3wp9XjXb27/fysvf6TAOcu3/ia
uNbw03O6bz2IqIOh1bRqLZp3+7XB2/qT3G+SpOjyDVZDAFJphJtZxHl2sahPsMZkaA8QsWbfVlk6
CBt4+HG03KG4ryKYvlh0M36T3xqKhJqwBMZ9cVqXy66TgeIiBwrvVlVdmU18S9wnPLqQMBIysAQt
i5k9qN8HlkrzKlSNikHzR9auErXafVp4qCI/xFIr+K7gmjaqBWIL5rRHiOTBMAzqFUXjYtZ1T6Ca
m4IyPUyR0NVuHR1oBT+YDsWBbj9SZmUMlLI9py82SNM7K+a37oF94dIYK1aHSLqNxxGdz7cGhPW7
4Iy8GsnuEjg2mFYC/BBA+8qTerJYaiVOsUjZqjso41BYCr2ICzueHX/q+MYsO0s7l5zmALm+5wOA
bWPgH4kEe1ZaGIo5gI1Gwonhd1blJn7UXFzP/IpTS0fui3SEn5aMNmplKGk6+2jkX/ANfEHQ4MTK
g/d2EPgE0UwllJflab0IKQTngEnSDpXMxkt3e8R2yYqwCODTB54EUeD2gqoH2CNCu2hqvgNRnvBx
mfA9dmFGY6UV++6mE/NV4YPTTqfPxpqR1t2sdlshGL4yP3HKPtGjEQnh1tVmGBeIo9H2UK8ihDyS
FrOQUcYsP/sB5iCDM5wL3wjNEe86uAObGpCAaWZQ7YpuVQYETR7rhZpuMX19xk9lsyv1LiKYRTcY
PmYc7e6tFI4yuZ5g0fxYehYjXzUt0fGMXOk065BpFJGfp1EX08SkJpRI784qcVUwQy3fmK0LElN8
dMV9JTsf9oKWiGyjDIUMn9v89WfAZftmDi0KBiJoKIhVWSIscfF5bAu6lS9yPO+zkl9Xq6GGYqOW
ROCvl9UuILuqCwy9Z8hsuKslez2gEpcz06kft2rilFFi0nDvHwoMtDEaV4/bEXF7VjhfIcNhVNHm
wvVfIocCtgkhQhakV09IFoGDHMZ1BLjrFTIEvxH5xQg4VgOP8igc/LAbQT1u27Vnt+3lO8pNNw2M
zKX6u4JQDX0IDigRUt0RWT75wcdK2ZY7dNX0ZL3Rj4j+ioOtOqBWJCRn8RO6RZJCvmrCuE5GACUf
lQjiqHTw24y+RNotQZdFsAwohKBotS1Z21TqBUhfaJ3lMYbn5RMP2JjdygxhOPRFCA9bySsBF5Z/
KwbB09JPhuOLYA21cF76+JMsebcyJmJpvH6rEuBjdt1fjT0dtgYcAil4EzOj4K/HI0ds4ngjJdOw
XFKfnwHo6JOeNUoS5oPjQTzri5cMNfqsm+opDWrEIT1UBzJs2lIToEU3sNAqxbMtN4My/MpwZrDn
Cqa5CvxXW4vEUUv0h+FZ1VlFKgSBqGGL5alreiXWFjBPSANvtkt4ewPQIUl2X6p3ZFiFUUFfZ6gv
TK0PO9j+3WG54fbHeCByuOFPthohkW07GwRElTOc1pODM6JyT8UadUalTOBslRA6WsxWcy+4ev3H
1DPTCaUVq5hr8rysSkQgIjwJR8aFCCxaN7DET575YNKXuaQP7nVY6vqyGSVicUSc2lYIgw5mpz8U
XxGDh/0ZLTQbwGxufRWuZho62Ey6YrtBd8hdnFTEraTcbVSTaNNHB9vKUML0dM2K5VJdIGn2I12G
5apwbN6faLw/02xzLeaUpIm1NuJ2y1+B9AKfTHhFyYfP5icAPR+k/l0x0MenqVMmdrsYiVcaEhXd
KedoWFmcG9aKkSramelQFrVkN9kTMmqpWXUr+CCtDAWZL79Ga0QP+PgVGC1pAzaK2YH/gmPq6OMs
bfKNjpUlRcwLHR/KawyACLGE+R6UIvhl09RO0LN93BKEOi7v4NK7c7d9mHtjLeP5GWzCneXW1E/D
ywUyOT5veIMV6fb9m+gKA2Ab6P7cr4PtNc2Ix/a4DBB0sd1xdcVXFwCz4MUUT4qxeilwSLOHcOW/
rFXe7aGIoB9BjNTmEc+xPNsis6GHYoR6AvXXwve/G8X5qtgB7KegEA4OrF8YORLjGejtJu7cRosY
Tab+mhv1dcEBf6kUV/5TUwnhwOf8rmAfjfk9l0Wkko4hsxGdvzxX22aor++JrKPnAA5+YhpFHLti
Lo/84NEn+wXaVp84SWrznmo3rEHxg51kq8eBveXBgelc+V47jAQzfF86RqZbzOD/LtgeMzoFdLnW
uOBsDKas9iECfXUiOp/3qWgpKMbD09o7BVVdhAnLovMh94KphhSzUyFJgvjXr9EkdkddbgehQ6z0
fzW0+0NQ6abh+hZ4TOQdTGfAyrKekTar18qqMFE3xwd/IrenZVpCrFGDcza5/8yXa9ex2fuZIOSq
u4TrmqNWmGZDKTrpDaUyas5PDCnRDqXpcg15do+XNFlxPdH+yTF2s02jHkEvzxsAgPkBw8LKSnSO
C/ntyDTLPygm0WwdSXB2MMEHbNWOtehHiM1HosrzYreMS7wIEuYsXTN/03S0dB0rY4q4vnIFnJvy
YH3PmBljMSpVmqfTzm5MgcFVQ26V5Ox01KgeBJWXce27C8QKTZWutmQq2776cDSABV5/2gwxz1b8
RHo+u3CtbeFFeUH0N7Jp5wt+oBqRujwpVLS5Sr523mWU+QePHthgHnb59NlAbspZcHct6Hh/UVru
t3zXAES+L2hTc65Q7xk4+k+UIhSqmspMdBM+eeTxDi3jfOAKkvyQEg3l2jLKIebJsNdwA4v+g+iH
ZJFFQECTszOYGPHDuHjeN4y+XUM9Z/3s6AYG9rGbRIAg1dDG6bDkpelbm/6tS++SCmDjRgMABGv0
WuUoXXBA9axcMjP9N+oyKOBypmj59b9EWHTihC4L6BQO1G/lcivKGuSn8DVrKzldN6N2KRGK90Mp
uPou9D6Pm+NsXp490t3uI0FQQ+C0qF+J6G9pHaIItB4LbspTPPtYzlykRbpHfooa9CANoGhRqmE4
arobErCaknYouBmYlgq+6LKPT2UhlHvMJkiEcWZ4JZoVyT8mru7r1SJEm91Gi6xfRxwvf05lW/CW
8Ge4mxneaVPFwv6c502INSYXGBkiWleQd1SEVIVqif3iDto8HbT3pKBiyaM7+wL7lbhhcZuZK83s
l15o7b/io8/ZUlG7K/GY9VMIJRPhsCIO24pheQgQmEU7+mnx1rImtK6t9O3A+Peiob00Q+pxhkIS
wZYkwj4/YLDy75mvFBjYwDs0k7eEg67psrjGD//CSOAnJYjxVMNelIXMyL2vVD73f7BosI3lQy0n
d7o36zNy/sbrx9ub/3wG955ktW7QTNrfWxZ1HsQeq24XEwyF0NFAJkHgjgnBwgD73v58XcndbYFt
rFHSE2xD0hUIsInkT4go6dO1+WWjetuJHrA4S2Wd5MXFMn3xl+GTZ4YUCJtVEwl8HEd6+uDM5gv5
YWlW2qCQSX+mizMnMYVZPjBFIYOdVzE7Pnf/VHEZLvOJZHepK8eMMdFJ7W9+9wDHlKzULWNF3U0z
H1WHjOkqo/LHAQsYjZKZpHpb6+zzu9fk3iQlFI0AC1bqhzwlTMt8fVKvG/yjhJlc4uO+Y0yreOG7
EylhlZ75FNHJP4no4/g5dC3nWDI0PaT/DTo6hCjHtGbE/XuHQuUmYiHfaeiDTxqoZAOL7JjJX0m1
iuENZM32BE+GLnqYLsdT9dUDLsj/5kG+6Ek5sShNNCO4ojRui3EmwokPSnitehkk1qYY7kI2PxjO
1ITKc4bM8TwhKc67aBVqEL539Ep0Zjv+G9DGoO9qWxpZCzxmI8EXnSoJc9cxTFSK+wxIfObXuxGc
0g22e6JnVatPytlVJOQnnD5jTgvdxJsmbNASZ8HxPrjovdJEVwTJv5MhyQr4SusF3lAU2kXzXDhS
DFaHHoPm8DsQ3afpl8pjykCLu++3vb2EEBkr5cwxsiRc6Q+93QFFzEde8mAQtTxxa871AjiJjuJw
6ykqe1WxkTosZdIzodHxj6S27nvUFP8EoXvTGTfbjy6gv7nYZ6SZBpLoXwqAEwyD5hahKEeUCVrC
fOhp/xEMNfe76hgPWLr3m70j8TIAtvHH2CvciorvCt8gq6d1nghNNQYOnVYxM2HQ1B80MJUeOl3Y
4wbicwJxbzfdEqOsJJBUM4a1c8je8N1E5eAVEEpMLj08lkL4vlJykoHCzb68UAr1OwYXZMI0/Sxy
/28pR9ZK1/8AyhTOId73TKkvZnTyaV8r616Gy4XQx6ABmRK9MqLpHYMe/JZBsJqaeRzDKtCnMugZ
1kIgBbVIy6fMRgvM7N3pQJtNVJSoZyWUrEUFOac+bkdlDS4JJyOIGR7GUp7YWt2Tpc/C6hBjPWDe
RRfM9zQmpTznhNKzOkqAXCLB0Y5KWgywVkOkXkECne6h3XGsfr6+J3isW0S3xzZUTjhAeYQd9EPH
zLLvyu/zFiffWiYUg369/dY0tWV50Ghfhh6XpG9iVe3tHgXeOJaQeAI7vwmq4sc8AdJjeYHhqZC6
AE0T0I8m09MlZCOFvrSsnvSDLY3wZOSqYQzOLgS207FONK7KqnynLY4sRNKPPWmqpQLuCF5yKZi/
kVqzOcDYbxvBstcZDgc7wDHhagEv650rPe0Teyb+hnPegXSK9YDYLWCyZgY1t/dtFoWxhT6QJlr8
eYxw4J7uQfUUsrEzT1LYH0EIGsk7VKtChbuM18XV4dUIq3F+48nJ3F1qc185ANJeI1IZIemvqAsF
zGdKgKg1FVJ2I9DFkleP/kdS68Xeumq6+W7o8cLJoK3JlhjdfFeabI2qtBPZ+61Gzbt1dygopXjx
tPbDfg/wCiBvHNsEp7uvYFwP7VYp+JWzL123yg/vjMTKgDI8ebpdkYW/0P11huIIufRtZpMUjpAE
JHXKxFZ5p7tkIc0voGvPjs30JvqPJuoIWbrGkEUXjCbgYOfUa5tsDxo12tscE7wK31Aflu6GFQi2
9EzXpxQ9m0KAFxbYOCuPjMStGcaBz9f17qFO6BcxHuqxYlARpKbW9HjS5aySSH7WOpxaPmoyyZC0
dbSwsmyAdWzdgbz0WCPtQyLD0EoYifOyIXXH+FOPmrGHc4IbG1ioEY/Zaeviz97fM60ttgTGVMn8
X0UhONK4PIyEfqLAoQPg4LeX4WdpDZsF7Xp2TSPBoDuB9xd1xo7xPyVoTxHmKT4P2DIIFqIj2mrf
Bl1u1Ddoq7e6q/5lHHr/drrzv+rZrpQhK1NkQnHaPAxW2AZsfGEcHIqcFfuS184pkvCuYB7vrTPl
OoYQ4FqjGdmoWo0e9JYgwGsXxwIKRXM6sxx2Wy8Iup31WsMjFvLczuHth2375jUT9M/uhkRckbrB
iH5/ySKLzQI6uTCPD9KfDUYJj4jwss2uc3PxM6Jm1esFES9D1CC6tSMCaeGDCfeJrxXSm1QHu/4z
CPkFEcO8JyhJUe6bnPmZiZxDJUy786oYFshO+m8KTQ/DmBEX595o2SM9URX2JDbQL623cIWqWmwK
KZFPavrCFBWHt6YVALoma+7VMX97qOQ2bDt0yupEUJqUsCXojhkmeGByqWhz2UpGvR5SAC8armtz
iycqCoMLSAcLY/+J/09qvg8we7nnKSdSCH1EYk0zf1l1jWuOcAXJCqOeWBhSqRLOi5jdHFRCacuF
8dbfr5MmI/nT/Eo1dZAoGjAjj04F5ZerDzBKIhfHu+qF1U8GlHrMFAskpvaKxodO5MJ00prgbYz3
UDe/JgpQ4lkS1Xl91pce3HfcDydHHckjF4D8lB3nxFDNR63ViXGiu7/kXlKBOaHH/asAvSjF4zqO
uw3UVnnxEHs2FtqEPbhRCn7WmNgI99t/hdG+udYKWgXvshZZrTOroGsV1xqhHDxHo8tBggh1VYRz
9clhfrskiEGwfJAQPqS+tZxwjXuHVu8CffxyodjC9bweejNT2N4f74qphTAEMzvYkqLXglDifKpD
GUuogQiOvK5UMwLtPhYCOwqLdY8ow5qGSDp6N2CjTdahgdR+6jnOIMI9RxP2RgACRNw3/+fTrz1B
H8WmJlxoS2lmt7iD3RB7KNai6pQiIqPmoPOK2AdqNiazJ/pl38NDZeraVTBp6VHKFT1oQIwGd6Sk
yugoe38A8CYbchJNdA14QFsT3N00BuhAmEW8+WnPZL2exqnH1Jq97X6QW2ENfgmRQ5UhwCCnWvfw
4XzbgGV6pEejAcbQspeLlvIoGs7b/nqUjY0NM48fsPYxqxfnXXzQUODswrAmvBDwQvZKXlivmopo
MpZMVsc1c6oh0zTuHhqAmhlr7e/QTgSEVITajfd3z1LNCPfkjv4RUSah15CrHqJ5BBYwOISQua28
IIOqiu1DtxPs/dgPU3yjW/Om5NaGY1Fj6XZiWR7gyfonPbxFMi6KCnQ7eyW+DZk8I7H4FowmUiSZ
bvcWHX2CPznLRWiwyPTUtc0JxpEf+4PN0ZWcL9YaA3pKU5LOnL8FH842iC8VDzCNLddxjRAL74UO
VYOf2PfnD5T44znpS52x2NyckmIs/y2Zrf7P0a+4SNz4lQwVBc8Gsq6cRYvMzsSEciuJtQ5DBA/M
sQ0gbfpoM6Qbo0rq5iIrLftHTus42uW2Fs0+IL5xhHCntki6z4Lam4x6M0QWCMLoeSVmOgJmUdRT
dBesFG2qVAUOvCknvwURWfC4snKeoeq0v/mL5RrpzRwwSc54fiRrtPHUTvjIVlmfzIqfv40N32NN
cEKBN8zd6aLTPhD214pHZqhzH1kDjAUtb37SnFuEH6OJnAsSjv0flapeYo33JfzdXXf8F0ksIJr1
XYY7ii1pva/62q3BdlqUYC57i3FXHG77NU2avtgzrFJtvSHS9Iogkl7sSHMuPe6gEfViIGr/f18A
l2/dRAOa0vLuQ5VYAFMXm1+vjtDIKOnT9LQIFyMIoUQ3/+00eGw8gAz1aTbh0JftLrAxYpbFNV2p
YpZBBAptdgrQjvB+3SH/tmn3Jz9rD+nVzx2al3Lv0tU5tTmu08/z84dkYV+aKiOmvECi1jARCzzx
gNjR60JYu18DHsPr2hrUtpAVZ/9qtn0uz7qgsWQ2gaUbsvVrT7UMcNLMFgMpEawYzzq3Wso6uoS9
JisIZTvWLeYk6valgYTRGWR58oxM9qJBhWoUpkHua0oyrD14AcvOCtB7Lhr7DwbRfq+sznIrM429
3uNtjlhHEnYOUcqROkhWUDChAflmkObSczKav+A6G41BUSbhmLhEaMcHf7lBueNAKFP3uoQ0MjzS
PXu9oNd8HiUjlGpfeJXqO4d1iR3ZPh9OnlGwyZfYWrcZxrmL906OgFDtKppRp0UEFXuz758+kID2
4oZt8vPJhZ/nfJLSyJkLJ92koISxdFMF8gGXgKVOgQhmalgjuz9G/FhWeJuZSti4ES2rc9+qPrJz
rhUaB7vMaNhNhd2QzWkBqAoOL/DSMRRAb3H2OIHbXDpx3E4K24UgBHmICfbwBhIxDvkJ1KObAr3u
TjXRUG4U+utj9NEOxNgCb6o/OFdTgGkl0L12Ej9sSu8h9rTjMQuXXE1URR6R7OAc6jAvdQSWe0TY
j2SL37ii/ck5t6v4K7Xfbfp18bbG22rvHKWIRbkY/mSR9MdLAegW2whEv/K0vJqQPejLnOxwuYni
lb5f9erT/C6+CE05xbt+iyPxRmYDZlbfqoWzPO5CWzSlvzWSOAOS0sBtw//K8WeCvXkWtNNOJ/Pj
17kyMcjNAzXQcWEbRMMDap5Ggl4hBdBsCwbLRNgSkdHKp/j7/cyKtZ11D0qSapDG+eHgirxUwohB
UOZ4wxq5/Xz206NmjEHmp5jseiNSsApbmVP35jQXR2AkmTdrWI0UXDjKfkrmb2Sf2zNljBjDmJKi
+eUgliXfxjRSbOqHkd1SoxJhUkspyaqLVSmNZpCf7dpwuHNeiDpPCX0Y9vs7KmdBELsK4MKmI+TH
5wVf8hSBnbgxYp8Mwv2i4RwnPm7B2YIFk4ApegZ1NG8Mi8X25p3sXhelJGK8Rb5fZy0ttrDZgpJ2
mJguT5pVwtQjHZPt/irZ/qIAujvNoXggbfGTiiBR7JEY0piAyQ/1Ddf6H0J1/kqpciBW4CR7Ky76
MLcHp+qMckakcvP00bB8TahPbmjvUpLFADYUHuwNlm5+V03QCzGZkJBKbEIGHoh1ib14cIGeow3X
ak7Sz2lCn+twL2h/kZJfXP6zaWoqro1rKyOugW99H1OOwbtKL9ThLzybwTs+Y5KjoewPtaPrhLvq
aoMRjLnn6prZr6FPpEeQZIiEkXoCFEx2G83j5B7XOa/FwPDIiXC+hIJ9/eP0GQMV0AX6OsX+Bxzz
DeqfLTxj0uYE/OCvGgZH6ynDIruG3VmNy7s7faxhRsqsUrPLCVr+2VZUcG2b+JCpMHfAX7jwpaYR
jO+/Jddyb7lyVybISydo495f4mltZgEs4/p2n7H7kC6gqIAPSp0o5ZgSgdzfjjLTF1wHpo3Bawrw
MUOb/ytOl1LTI/8DUBw17h0VxST3v1UKb6IwYQOdVwmi2bm9Ukh8I0XJi0g68SAp3I+T9JHAHGOW
uZfbWhxuGzjSYDuzi2IsT+GAtZD34oHxEzhCEg1oU4KUlXOJFkk8bcJ8ZhycTL9XpbJQF2zYNSBy
iOuqRzFon7TihbuUL8xzxPcubizr9nQLpUFO4RyA5S64eXNvn3y6qz8ll+FjDFuQ47BUq5fCODdg
YjJ43in3JYSdvk/XRFROTIYhzMc+dMuO4opU5xyMruxWcDQW6diWNRHtuqKSOhd7g7Y6/jEMPt8C
aKtIJA/S+ceCO/z6Bjn1cwChFXTiKOmBUo6vyKCyEb274cbT6aFq0t5es3MekexHaInIZqZij8jm
EoMASu1yzNY5nmJ6W5d1OHG5eSFqcFSpNDnrai3JRdhQpeXVsngQ7iruK+GKO7HIm78IE2/T0EjE
flIek9zt6tnYMJxdpH7/WPJ70aKo+OFAidHX0cYBHPeY3nQDMWILQgrAcM1h5bIu7WfubKffKk0T
ZhkqfzUdRh2dRHAeIX5kcmIjU68sM/lTqN8U0sqbEr6JU6UYtUIIXsCcBoKYUWtVoktFbao/Nv06
1dRBBOMwNHaz3GvBM1Ne1MAdHatSPChQywtboHJWwPIEBslBwbekqVrhmcmq1eUKe85GCV6A5sJC
P8CkPsM6hbcscTk/gKHnd6foLArO/DXYRk1kkk1n8/Zw/LQTHj2INUgKqdibp1oXyKGYvWW4zVIJ
bigq1Bne8lLiq0vWZ8izZ6Tn2hLYS9V3Vv0UZjUkYr/m2JljgQ4rgA8PvzZSIHcOn26NksqHJje1
ndx2Y0lWOXZU22PryBWSO8jxo0U+2/aEwnihGirACy+ixPZOzP/7Ci0pmVpmGUX1pkzkKKHfCpYJ
p0YasULEVpVQPpD+VHGcbMVtzSxhTtoCzIXlgQYo4qVe8pBciKVInAiYdpA1cuiHCLZwLTACB0Ei
v0t6UKshv1IiXaGDSP2rWdjSUaN2q31ZFLicnWHpcDAYvP6jiC5Ul9R2AhQdrMV4SuQmZ9pzIkoW
pXqQdIjdB06Wy/iXFYxw8Yul4cYdQJZ9m7Le9K3tXvHukJfr2tRKlmxpnX8UPTRnwR4V7jjImtBV
XWMkw3Ssz4/PMAZsDqAeXNJ+GHHaMhbYXyyUp4umLT+XaU70qDeEjIYLVTea5dS1LVdIL4llHg/N
+C4uIC7qydlw+x6UdiOZhDroyUxPodWLUTjXjZnZ3z4BhM64Y2SCB7SJ3SE205k1Dwr+RGDr/O0u
89lnlPBFqh7xycpPjRqf8LE5amiKGnsO8aFdAalA0D6RXKNVlP+myZp0XPlNv25LT8852vFp15zD
WspHsn4aDQv7lHRUD+tUh0tGkv7FkvHzWOCpPjt4/Nco4JjuOKPRyezQIvHjIwpnKtoJCbWCIBYf
Gdk+U9VSkWwLZwHFg9MOypyvmMGAaBIaOF843+aTgdP/Sk6PujXp38wPVyzMRCm+H8UAZBouXQ76
QdUf58QI0w3R/3HjMhVmR4M3fQQpy8zYgc+2tQ3P4MaRj9x5SiM+7lGrIMNKTkzwhqaP9uOTcdyQ
SiimX0eYbbnpdMqS9Iyiza9ni4hdAr0MM8zHntBiDsqhtdQdyFAw2LnMuIYDtUYo/NqVSIIZHSE7
OoGeYecNBbBF95zVRUJdm6g6F6sWH7wayK3mTyPBo9LS0Kngb2QHE75qFUmjp7Q47Pgms7comtbU
Lw3C10+BJRqlSLGZGKkOu1G7Ls19H+mi06uQkNU360CmvkzQNip9kzXPzw/5aegpJie+Ipfq807T
umpR/QzrrdfN0tLpyJl9O2JT28yemlLiET5Bkoop9NgGImw5Q6QZNPWcDlAdaZQjUYdTxFnCb0fT
vBTVceCOCBj8JXEb6ZaF7qWEAgm8i8+y22GBR7Ij4trSeoUXDmXbaaxkIM4tenHQhV8rKQYulC9B
TildXAw3U8SDQXpHKSUCh3VrdldBoovYqR3RMtQtFHbHkeKwHAjOW4meKvIc0xJuSfS2SyqTb+0b
TlenHKUOhHpmTu0zu+PUltb5rGP/5MvLTE/g2AkPgkuN+6U/QsQAW+86clrTPwaw7r4muF+lMMLC
CTNb0sv40aHIGo7HytJyGOI0bLiVXBtAVBMWtwNoGm6QdWCbVbAuaUGNQEGvHCvO4rGy4lY3MiKp
JaP17viAnlqtZv8e+BhtB4b2LP1T7x6Q/VeNM+ncMKeznHZjWh7+4LopEKTELGAGS7z+YQ1JhYse
tBG7p/bYZo3eVpXYd1P0OrXK20sgC/QHZbSdtc4XNeop0lcjb5TODYLJ2xuKwLZzFHL2jPAqNoMj
uHXWLg3IKqoK62etmxniLfJ7bgQxgxE1KmGs5gWZi3JI+1DbgtqjfNNmAFpRvL0dnwiz/TNH1eFF
x5zcfBGLEcSQtvZtZnHp7COWZKn73tffpUCUlXuxeUPpYgE16MAiJzRgjvpGx6C5/iw1GbfmNPZk
S35GKadq8lP/7QjCMPvSQYxPfREr1o5lOdRmPQAh2SoB9D7JwuxYUd7nu0CgdF4eAS7BkoEQ/bZV
4EGMXJnKhfBzZ7vwC3Ap4jIIvd4T30yRnJk+axFjOkBr7xGWPTdR62Bl2bsjd1hFx2CTvcZxl0Wg
f/Eno4w75XMd16lJSxs7GlNg4/x5fv0SCw4UYnEo5udMA4LYYRAwBx0w0QmOIzJxN5HZc63Tb/Rl
cKXEsIeoqv9Wfbe7kURbSMh9QOBA0Ru3Z87TygDWa3mFqVSlPPV2H9V5pzNNOjtYarRfZ7ZQE3wL
LRqlrbtD6AH9KlCLUsoST9P680JZc8GoxxmCLmgGU0gCF4NnBvaVNI7q7KpYms2AcPeEgLt91lJh
MGenNA1YqV6E+luJ24t7xtdRwKaeSHzmLQ6oM1oN16gpn80pJo8PnKmthTpwFYdSEHmzPSk9LaQv
sjqS6Ic8tvf+w31apmn10a0iRi+V4mfwDagj6PHqrNxKP/bDkefY2+ra8l5q6x+MgTVIdqSFVF4I
JgBH6NYwJzCaWcli3vVvGFHe7Ru0P7m1JPeUeuksfNk5R/0sD5uYXa7mY29bkOJULObtYaZ8RM+f
0qzHrPxDIoIFPzo+45Z3c1OI3iI1AOwlMBkBOrnuO2zLLX5BU1B5pTpNexNsFEKB/b4WydJljxAG
k/DbI8SIyGXdS288JMZ9cqpqlQYPTVAkyY7L9qfYcMCKi/P6Z9mSupZ/+uMXakdSdJrFx4zajuNa
PnyFY4dtBU7+8qeJGQuEDgfyomsn3t4fZ94IzqdEbxFG8IT4HMLN/fFna+cxjJ8cSsYZ253PnYP0
azbp5EZyvbMrL9tmodcCiFeDjXD0PqkmfED8ynUCGxOEwnAb5ms8HR0ucxZISQ5T5/tUTVYxQIc3
unElTdzYT6WJBZ2gkv5b8U+K0JMJlLaUVivSO39HQrrjwYjWZ+V1vjSskNHcEeUnZA0R1qo14LNu
NlfKv8GHcW2W6dCc8qc8LuN+B+BJWGQ4m8la+tRYTJYNItxB+VNxMkt976U8ZO2VxtXqgdFrJLgt
IP+ZdG6GbV6NmaVKLrotQpEt+sf0eODGuVjqSmWhizJxGr+gfMu6z6cqvfAU0N6TgcGgTFl14fM8
5Qq6GWe0AdrUmnJvM3AqCQ6+zZIAn6OUmoEZaVdw2zQqqBSt9iNodL49BAKpqK4N04hlxz2c6cIN
F8hD9PXw7ybUHSeEBx4vp31x/nw9sxhKN2tpNWcLeabPir0zpdaNwAiCaNX9O9gInxixba/XXiDj
GO+qaBb9LZ3umxCVIkTlEmKDIvqskUeCtzwYj1DagT8i/1J8QdYlgZNV/m3k4YN/YbwS6h/9nKMP
9EyD0EyFaFUxgbE9NHrsMIPAgHbSbk24ybHFlM+f+rzrm+YhDmoGrk1GLtc0BXTrOzwcN1krmoiU
nsLw7iD6gLqqJfbywW6knXWPnZvpmiuugyXmEd6gYUZxZPEhPM3FuCZuv1seWmqKgEezjYt5LJ9O
pt3nenLzUCBVUkF8PhL77RZJudil+23BAdCyvoCgpjswO92L7+EwLb8bOfnjmFRBoUNA9aD++3UA
O9E2M9LjZwHW9pwNY8ym+ri3q8+HzMXOiYQkrnoBVySVWo3dVEnzU1CGxa4S6YGOOXCziCub8xBO
s5oYC2GFRAiR8r64RwLUGixdV+/XFYreyuDfqnkNrn4bwcTPDJNY0VJScPPxhtAAK9oVOpDEWfMo
es0uQgYX5qnP88HItklkOo/ZlMfEhoTDsLXqI4+GMU53kIF2SYgle8p2qRGcPRtNPnj85cPPW83f
ykDZUZAmZYdOCt6B4Ew7iq2PKhFEBwe0fJws1JsB8IXklB4XXCr5TcC2ZsKvZxl+z5JrhqPnxc12
I91yrvbN1fEeHSHABX4h/0BBNv0qHWv8GdLZOi2zSCopZj1R1CH/ACZ1ShwKtN440yXMOO58rRME
IQIsbqPfCq/kD0i2olq11Wtqmp6AQqRD4Zsui9mqDf5KeL8W02mJZ0EmBkHq0vrZFdTbdQe9zIvF
vcBcaOWRQmaeQ5Mi598EAymlgeQwhwfY7rG10aeeNFj9vU0e/ngIWOvP46o6iZhhFp/aKtfW/ge+
IS1EQyvBdL+iVMGcEIHmYcVr67v3D3EqB/T1a/AYekowmtrJWCcuntaA8wM5Qe3vO01Uduuw2VmU
9cMR7RBYNl/cBJjugvOF8gXTfM//ePuI4v2mUGR9YBDhFPeni4bqZseDx8tSQbzRual4+bEUAz9q
mB4AXXG10MifdbOqGTRNWNIkgQ2Ri7aWjLZLUSBz1iCLBkyGppqJTZFg2r1pxoClKthdXh19/oyv
BiRpBtJufD8jcg51SZ6KYv7cgHR4RjfZb3/IBdeU0UarbRKiUzjbcHNcLTtP9QPPA0pEyfVLYKug
d2vOKJu6LyzwGcfqNy7lfZ+2wJy/AEqcNDer/AKwo7quwweSO8F67+ahIIe1yUQVEtma4ro0jgvi
7wsX3BtLjty2dGG1peJAd5vk52WQnBuI4Qx7lshJiBYVqr5KmJSajnZolvHINeUGUotpskWFd8hW
0dJYYWk/K1ZLgtXIrfGzcmSyIyWEJ7+KDYuHMsrvI4j9fLSxa5bJrBreFE7Ld31Wcu1VbjcYkAGA
0MzZPEWHz1qazRvZGw3eZ8ZaFU7hCbTnkTQ76FyyhogQfrKt4e9+bVo3koCtWKzcF9ZeMAduaqCv
9mMfXTYJv7sz/U90HPRfG9+WzEL52sF/vnjxgYQAnR5MdR7ByL/UtqMSBtcLkkLHgEBQBh5WEEx/
pMM+nDF3Y0arcvZzzEgwlHtGQF/A6YYfgM1b8BDZYazv8v0OmveohXXOfqDGtcGdyJ0khey/lLHy
mI1/1ugz0LmXjuGRWVVIU0EBKPQ3Ds+66KwyVOYesKpU8WUsT4v9lon/Y+3/B7hwCLcXryo+jctz
pFoM+Oy4beJMdoeh1R2E0Y4dJzSD6E7EZHiq91kzsqizu6I3iYPLlA+GaPSM1GvldmDK/fOTEKKx
JwXNZ7yAjYaIh0Lec26gh/FpnOgDXrk7p1WrCX2V5cSHHn07AvYP4bJ9oi14XvXxgxdn0NtuWfbz
oZ75jyl48h0g5KEugEcEnE71nNiG23cDvESCIvfi1EjtNYZdkH/89BK76knNd0sM1IaopVyF3A38
W4KcsHaW1+y0SueubVrdBMZq/wzFcofCfn5RfXnmxF6y2auN7uxo4HqjwMqTn1cNSLisC5kcB5Lm
TctgshMOpqFSST9vNd0k8dNF2AMlXuJA4rQlUuwC+QvCQftHjfAuE/EEwIX187HHZPF5r76up1nI
Lqu07Hf4pAhLFVTRc2S3p+CISqlFGglgNxNwZ3DQgYa8d/OWH6C443Bf07CJypkcOuUxEegsM5Cg
I3DYzAwZAq4eA3FOcYcrL6kSLi06d+XJ0jP/mxw4JdgL7+CW0pQhgG3p+tRBitrHBdWIGj5I1N+l
55Yi60bZqJGNWNdXqelWEUW2oGPW7W52gjP/4EtP1hZFT+PkZ0tykJ9ND/GAUwHwnbmvJvD+wIRu
abCgDvdhD5Umgz92u6LykMdbQt4lNBjH/lhrPzLw58863HMO5SwUqJhggZvgCpeN+NiiKMcHFeRO
27wdK4KsU2nHGmoUhExaic3d2uhWr0YTe7WX6B/zn7hLnBlL7m1nqaxbbaWsMX/gwAt86aovlHW7
4gGHJ+YkuTMexdSHwhIVEmFpYWAJNhKSUQ3222+JK2pudMhSrtmWXDuzAcRJu5uHfUDFPJ1bD0ah
i/0zlH1doKBcttcEFi3syW7vRqCWob2jZ6M+ZoWhFd3+cCHAzTlUQGXp/6mZ1Jb60izVQr++wcQ+
sQyUJbik3LeqX4ZoW3Xs7sdR+37FDlaXfWjXpfHxRmTkv36TS/kuv/tpAGBir017SWLWnLaTt6dI
EF0bEQmLFRniWRh+KXZhtWal8mZ3jbM6+ppnRZ3kRxcQL2xgZBd3inPr4ijczSmrzriBl8r1jabV
R41n9UAOYOA7eMAOLRyn6eZwyd4XWMm8Iv0LHiv6EsjlX/uFsn6d1gDK/epmiCpvpf25zlJ1yLXc
2aL60A3lAYImOfGg/8atOXwajUIx3uCso6FaE8FuHK5L52POqAd3TguqhReMoq7ywJ40QowHVxjR
xtwgRcGvQSz5Xkyhc7i1Wq/ZesfFXPTDPscBlJ0MEgDKaAvkRvK5BHfF84J3HFPUZhZTmvmQCAZY
QR6NLIplDI538+l8LtEX0aw3RD+oWUAOWkynPMcbm79NG7q3blxeQsEsG+Z0SbM4jZ5aEN2otTQM
FmwCN4YtcoPXeFYaktezE2uwPY6PtMvVnvtxRM7Qf0cLjkMg/nRl7rMgN3Ez+dDcwbb30Mm3Kvpd
KAuAHBy+37d2XXvPRsmX1zBXgdqL8bMwb6AP6VXIdFixHpZ+2Pjk39CdbxN1y+BOFQHMMovhJKLE
2/CVI5HV1Dg8uy8YoVyLU62VAIS0aS6M2sl3zyVMyxh61su4bzWsVaYi4Z+1FXZduiixGolvpPQ0
8QO13WaXX4fIgt0Xj25+yutKnLTf5Bx7B4SGw/spXPSVROLCG0Cmf6j+KjCQwdAGXP3Sc3CAmGzN
IfJbj1fdRMwvaTNzdvux9kw+guFORlB3oI5yCZPKTLirkWSJhz77L9DsHZfIs36i9M7ZtbA/Ni6V
iOgXGlkf7edD3ErJIXKMeSejfS/N3EUY35L+x82h4/qqTd67u4+Cn2oayy1gcTckup6EPEql8G2y
mDX9jhISnNic5tMeKAfds37i8Lfs4UBau1JJMghEeRZPKnFcbZ5Zg5kN7stV6aa2urQnOge5RPeS
jj+ScI0ewaCNDhJzRCBLtUiSlbjrh/msUgah5ylSH3/HY9B8g6A04PyqXkcYh5QdfI1ffUydF2gj
0F9ES/PKpLWjrVwhWi1KuX3r7O+tj7L3nDxjHq/Oe4plqpJE5vO0Igvz94XwFfuX3M8ItTo4kv6o
RYKWeJKU8Rd0xYia5EUjgQx1wv+hI48JOF57NBEanZRc0Vhu/VxPQ+A3fzZ9rsW2gib0Ox0L1KsI
1BsWE4Bdxcv9zx50NlJ4i6V41anjUZ+m04rY5NEs8E98c0lUZtjr/0+WiDhcfPKDW4dzM115kdeo
FfhM5LHkylyIegmZRymmYNjJ9E7BFnvKkANsS+WNZip7nxLnppn0u2Z6iqIzd3AwdFNSBntwmLWr
QxUaYcA37TwS3brtT4SDInaE0X284VKNjAeBk3/ghm2cS2/J4sac3O6sMaRdVw1RM1DxO0IdZikA
l6IDcsgbq64GwTdrk8f+gZfd0+fGhKk2jcKEPiOdsx3XQbKoXDBH7tz6Zp617tUuCmw+VhPeb2mY
h3Tgtzg5RXyrQMYy3Qalf4DP/aAv/qPyjqdG7K72aB1k53KePBgeHd0cPGXDNZgZbPgCkmUo1Akr
Hy6tIHqoPBpvkXVr0L6KDrlWWsDbuL07i9+NPlNX/MWjO0g34QdAqI6FnXws0I+ARg6e5vXifnwD
okOGZw3ghGDmpZJLVejsuYzyt3Su5LVYka6mMFNkJoCuqOecpB2M6zakIlLEk/aJVFVHeD5J1wRQ
wCb6tsBh2vnSsekBp8895mz/jMM6IP8HbGkWVmTHkiAO8rYptG3UTYYiZts+rg8wM9GjI4dEK5k4
mc2XxLNO9tJUXnOd66V8Lq2AnhXH56IXTlxKNsXRk5kMgtLSxBn2kJOfuvu+jVilsC7YOcxi22Om
dz2M5kARupXiEM98sbwGnPVuvsduGjcYj+9bhWBd/bLnQIcxYM/ppwUYgelwkbQ3Nou4HJORryK8
75FypRYjL6vj59OY/yNm/GPBo3IILm7SADvB/t8TS0XmT+oK5diPaT8nXSCaH+x1rYHGaO3y+o2q
1SnO3B3SKLedABqouNyPEdcEWe+3k448hGk5LswR8dTseSoLexKAy4//A2UL9tadSNTDXF5OQuqr
uC1+wwYURmDV8NIoXYrytaYZ5/M6vLRgAXyEdSbtgHzu/Cz6CUjrICyEiTjt5dGBwNvzW/qOE7Gl
40CVCVvAVKta2Zi0BCQg1jN00C+pXvkDIg6psBDlEYW5aAdNOQQR0bEz1FBA56WY1wa+ywaJG5Qv
nqLtiLVT+9GS8S09fvD2oZvf96W0mFGuSs7I7tNdFZk0T+CvLAJ0nWWZgHF7iVpP20ZbqYAnsi3f
4pux1HDZzJuZfswPs7IgFONexpRKD9ijzFClBFmCyH4SvzP/EQn35khuJGYwUE/3d6MAdqKVtNXp
TSeRyg+9FpVOa6cd5lRGyYpRfy6GVJNCg1qvPikhgp9/xqC23Uq7+QpikOp7TCEVH0ImrCwFQQ4g
JohiKzPOhsKDy1xWRD/MFXpGOQH/RbeYkeuU4NmXtO+/sv3IPgItLiMzzoo7+mA6G30oRuzumdsx
KMgVfxoEzBIydy2DKI21NqoQw1vDEpwI2BEAa6LN/t7dozEZ7OR+9IFQ2HrYMIbjfxgRoPx1t5hQ
wr01TsxX4x1cr5uBXItvp4F9+3rhUx1UWSiOwFTBOnI+HS8nkWxrSi6aoUzpWFP7gfWJXtmiVIBe
wB76llr50KDmNpv6VmuZlIx4hYdcJiHL4c8Z5IdreZitbry1V1a+ObVI7r9SqRrHhhbfHQ5oPstA
3S/BxQblIYzXUM2MTZrxQvGfVzxOdaRJ8tzOLmBEvAeWyLMO+/bsQF8v1GZYixXFb+SO+D3GPN6P
EOSnSf9oicbT/Y2LT12piNN0d9Nou22mnWsWzKxPJNW6yG+1oR91cBvALzv7pDbXOLCA2v0D6mK3
8zyZYJ0CBdgHJHu2/8W5cBPdf/qzWpAqK3fiR8Tj5rqX2uUF+Ze10SJWD+q8gBBHhXawSpmgONtz
Fw0xdRbGVqJhvRQ7rtPr5pLeH/7U6rPRtcQ+JeTEnZTC1cRJJW4GF7waK8O7/AunJiMUTzDZ0VPl
GdsHLEb2ybFuvjT5ZyDZPkY+7yB0pgc/H3il36TDAcnR5m+y1ALNlqjHi8G+X71PrrDtkl6NNX2D
iXnfYMgyEzWp3+tDSx5lYCIV04QUySM49o7genm/bu3tXYag2OrddZOkg7yg6GZ+2GzDvVm/Xurl
oQrTBpNolyRKwAa0YjDqj1FWaI0JA68VBHQMcpt1d38ymG4T7LawMpHCVRMccrjjP3ey64qiQn8n
D2YgCO4ZkcxCEWUzVgugWax+LIpmjOPbuhg5Wl7VToG2XszUEPm9dEcLY5jaYjPlrjqSTYUbNZX3
UDoQhbV6lrEhY3+TE1GDvORYx8VGxTarFBh3w/VyfGLgEPrkh6WMmpkxifTnBWe6Jq6H/frBl+t9
U0+otGZy9Rt6ZI0dWc/4miH5Ivxr0iV8NKOJqTvfkOHbUYcwbMNih5B+gqKsuJzj2NFI8lK85UoW
BgYLh0SaLhqpY7/op0Q0+ToOOe+24dnujaJPriuQ66bOGnJoCHiPD09zw6R8cFJKyL279ZXX2h4E
5Uo/NYmCkiyuJyL0lKL474VgtY4+tri290TH2TRChklp+5CnbVg3c53f7vUqwijcN7EaY0xOZwAb
TVkSNH0CEDXdbzKW1wm0dXrT7DQwBeOQVkMsZy3KjNWhdU1TbvFk4vs9spW01CY5Q52v1Nho564c
YxrFImheXhOKX/PKkW0dMapO+xsTCnAlFbGbtqFnJ6VhMGqYd2GVQ0v4yD99FXp5Ipkd1KieitSw
0gSNa8E0DYFbVNi8R/fTGZjGEKqufEIyABmRe1dQhO73HyXlBVunUSsXMwSAZdPZxiWduzl8Ff++
Qco+3cni7ojGd7rXnjMYxsAtDj/8PEpPN5/Y8lUOUeFnrxDPM5aiNdO/Q1+NVQgxLCo7likz8Hsp
NuidHE+PfrWjd8odlmaEwCmPaImaUaXhmep47vUAfGCAlsi3NYFILB0L8OfanSneHX+YLB0MYivn
Hi7ByT/kyPhypiSop7vb6zBRcEJImEf72Qsp/aSECLmPWVUu52t06k77n/L5CRe/NFts/Ale2kgT
QflOm9UKHMGSkKkEpCrG5YCcyCbOguYmNBWi+ozkAKuL6IwOmNT7OItU5A+3KareHf6GI+wZVc2Q
NT1WA+iuvo2uy9nc/X3+Y2c5BrK90NKpex06aqpS3Mg/QYotEQc1u3nZ1C2h4G4//D0jTT1Mw9O5
kBGXBc60PsQFHeUwNWXMWmGDPxYErrvNOqq3+9YMaxVxpvJ+SLOo6qomzsC+1LsEocXhzlB0MUbp
6ab3vp83iw1ONVgCKqhKqBccN5/uNzIzWNdHufxA4RwZLMHAtkV5QXUuDE5oWPOmPmTC6Y9rEs64
Lg38sEPzMBUmuDsr1ikVk2T5dY5oKaCota0mEECh0dPWWKZtp13GO5vKrUb8VSWzpKBSjOb71Kq9
yyrMOiA+mOgdXF0KYkwjaUe2dDhl4AuMBEA0GM3wT8d9UHwXXVY7HlS+0P6UW5m0LmR+JtxCVoEG
Sxv/aI5ZNsT6gS+9pptcW50XeEPY5vh3Q5I6+EOt2f0k4Kx9hFcugM0ulyzncxb2uXcyJ689PFpi
R6XSKZQ+66hPuDWpQR2w+kgFOZ2iF0rv+YQcjEFPGPyIdi4f5D3BuXMW9eaYLnjWsKW187/v4T+2
DgbgfH/20h7CGae+zsru02Ru+nHv3WnFdlL2x/WQb7tqZEyJrmralavVvYM918Y76gRwupZjFadJ
AKa1yLfR7tsKlEE0PykCmCjzrby7SlAaTzfir6YHTsnEcsvmGL9Oa7TYiDISkdGUqIb5SakvYRNI
BvUdPFNDra/o4rep9IqCiktTZIMZHuPFJzOa+rPRO1Kc8lL4wtCVSSS2pWZ/dR7a9wZuLJOZpzqg
E1M4jWwbkEodjePSDT4w1gEozslWfn3JeoG1gxiJ+P+EmXSvF4bMba/n6NtEi3DWJbc07YPUV2fJ
lQ/lr+u/AcPv/DGRffm+bImjDRFCF0C5acNS8Lbl1huesD1u5uEqUnGfqamyaNB6U68aXz7f/U2v
ZPoFgSoNTSVQZvs+iu3G/iNo2m1kT9qQ2ENQWtf1SfhQ9KRzwRpDUBqzl/tuBA3EfnLBQu0ocBM4
Y7hTmjp/jmPus1ks3D0OI2oTZvKM/Xw8Zw4c8RErJdOwWJbeVsXGwqp0j7hFNsfKZWYwxFtQ1t8H
VbF9d1pfwEpGAqjQbIMr9TNz5/EQwH8wEqEkWcdxWICvuxvrxUyCbbiesogLXdFbCszDo2rfuweW
AcOZrbHWL/nMdK+LgrKj6ML5bs1fI/WfrYm7BJ+7oaeD+CaEHsS93nQNFoarxhlKolvqYhVYUwXO
FLhhF2GZLgvd7IRfXXc6EgVzCIs4AnX+Dab7NlWkmWI0ssrrwOIeRxVdoKsEYJ0wrF4+p2kWdhg5
lfSxaxaTIWmrbcpHOJFsf/tDwcvrGokNNIcVdJvWKckfuWqTzgk991DivLdqaLmwmkEBRbSFMvN8
vu/Jdzq/RAUYF4Z6OSlJxY3yzI5FYL2xU/aM623nU5F4TUBUZ1XlGpjLlW8LCv1YjbEm9lM1t3we
tSEWXhdESgveoSvwgomNRPLwITFHmqIVcBSpRZpR7tULeyvCG8nMsjNDJUpIN9xcxVYR2DjaGISq
+2My3aI4KsciLv6yOCFw6eSxNn9wXpikmWEXaWckqNtEjVlxLju7+yEzdq3WFf3cHkIAkuzMyZxz
El+/luP+ZWoHN5sg5ucOGlY78058hbCFAndUp5dx/GN+KppJHeKlC045TH8T4xQNobp3Qhfdnxl/
XLq46c1POvsLdy6ovdgJ5fU33x0BZ138XT/R3BSHU5kT1Foit2vlwTcqg/iG638osUkjL/TJWtr8
t0KSNnzszeXNtAdqLqxLHTdBhVGWYrxiyypE3AG6anbYOcW2OZRCkFjLos+jqLv53t6rsjPoHiZz
82TFyeOxvm2hjSEHYk8sIs1KbLCjMC8Qs7psgfZqp/b4W2DKxcDDV0sw+qqsZxThwQMQRO/OHgmE
Ry+t9GFMm4mmhbkP4lVVxs9VQpouYRX9wjd4g8vF2KQdgmErGQ/GYaUHUS7GvNlD4t2pn00clKz3
LTIy48Wle+O5o/n4KIG9o+ngAcFs4wtQQUpzUJOP/Uq6zRuD8qW/6e8Gey/nm4qkNv1q7r5NMot4
Xy4FLgCXO2h9OeLj6pzptTAIsapSbGV96Los2jPlDZEr01mt7VTHxhGdFBlAbovlVnXVRAmvt1sJ
hn8FrR33fS7vF1zWQmgr1lERXi7ctoafjFm3tUQKvKt9O1V+G+glg62bFzS7jku8MDN9mnbUU5Dw
fzFT7dNhu4W3oy60vfixoJLcV1m7vvQgbsooO7s0bVUn9TkkxfVyMf2/Ve7pBLWk4nqkGqfqYECp
+TEvZ62TTiCH2q1jRWhEZDTxioJ/oLtV4HhDt0ZcT6fwKDLhHA4NNfA9dXuBI7zB401vh/N53GuA
eAn0fhxgmGNFsF77RvTPRyVODPDM03Xo7AwNjra5VEaApvMQyH7ILrTUgvdiBPcjusCoom0n34z8
YSlPdusNM7UZ/yUPT6XcHjpmZWpMjePEJBbmr4LU03o326V1iScUnWtPJ+J+XIiObGrtP3rTpZ4s
jz9u0pIvQ32iHh6hAiqSXFSnzxV60DOpgmpWa87BcFXJv/oQECYLtY9NHu86yNWnuCKADTrlec4v
J69OK5C7CDY/Nxgo5tIOaMciOsZCmQJ3ctxK8eV11hBus/b/htCKHbIS99aAdo0K1S85NH3XHBkj
8POksMTRV4/sg69/IY4/0Cd3f1/WpBV6BZgtHIAi71rcbXZClmi6QAGGGLfDjMMMpAAXVFeDFnkR
TwBuSB3ES9EvgPp6K5pNMldiL/l4WHtU7+gAgAaZ3xeivG/l3JTXY0Cju3CThllBQGYuFM9kpS2w
fLMiACHGISn8idAoixHXGS/S5GUP9CfP46cdJ9xfg4coq76VYGAZ3hRIXUCiP6dllWBz7MQvlS01
laTZClUdfT40cHcDfEDjsZ9+sUfKq6vzew0eeYijNgEE27jGYcyZr0g7GU9ukFhx0jiwEk0Z1B1Q
msU2lxLpBs8pgbwxEtJF6pG6DL/q8y1tHvc+W0l16whsUev62qDXrBhewH4+H9lYJakqeHk8Gqio
7lbwiwOEl4olgkw9kgKSkQ9DSkfRW2NAqvEAA8W2vFZPp/hY6rrsMyyfwP86z8KWoPbjux+hJXUl
HJB9joMPohC+PgEBDJzxJd2uCycCPFgtcddCYMFipv2nJxeESL7dAeWjW8qELeSMSl6STcdJniTr
W4P2f4w2Ctt4snUnCCyCWhB4IZTIcJ771KivKF3f2MCegAMEBJNfoAXwQba8+SyhlQN2ep23HUA6
8maAIHEz3TVuefqCM9S1g9tO9G0nEOiDcRQ8+R7jZvSMWVTH63MABETgpoRU5pSi5EOCDrhrr0eK
1sBDfjXduWLkR2dRidC4G4udnsjQUtmc1YrdnN0VGOl8aqqDsEEVOCSR0BN3RxrLN25agf3+aIdr
Ti5nKiS4eFT0uM504mGUjwA3Du9TMCtxqd0fMhtm0NaDTIvS5E3nJFMJLXmOe8kcnWOtnfarC174
paiODIdjrZKsl3XeJq+TIPOQ5qpx2aSyE1QSXEZYbBiCsvsWeGW3Rchv7ZE8kKAY1Ayho2jqHpb9
RSN7/4pDB3OQ6Km18i++RvCLfUis0jBmVmiyY4iK5fvzdXmHkyfhKr4oJ4od6x94CiyLZ8KtOLc3
gb/sDhe0OFGIXXtc0FSnqbfb/ccU45eaEhD/XO65/10dmtsyvVkavx/KwvtmSH4CRR0+4zTk6jvi
CSId78hGDFJfEdNY0TDLBB7ozjipgHUvopcrjkwECYR7GUeuicChOBHe8/65vSEQE/DzUlyvYkIk
u/O7yhGZFsfXL0zpTac1YFMWdsVXh36P94FjHEmvwlCYPUb2jd162T5XyqBOKdrsUgQBUMT7NleW
NR+7zH7cQNsdEERBX+y1UbgTrZaZOhJ0QXPnAgXeFhS8wgoEmvVVSc6IbRujD8ABTXPHLn5pmWHy
TGqX+6k6SdBDgYLILcRgH58No9JalMsTltQhX7BxBDLscq4/4hNmBCTKj7uQSQ5em7Y78xiarlJE
byI8hZh9DvCkazgKGaptaCsuwPv4X0lR7fSVRmaeTNrE/ZDIC33q/0P7uK7+IGXz7z3Qf1Eq1CNl
fu9Dau4dk93InROqyLLc3Lxu9WVdbF2eyeGSJfIovu07FZBmYeY/rTBSpfHcH2Vqx3u5nL+41RtX
LoFqzNIGENnqXdYOrydcg7zhtmOWK/iZLC0ilA9WbjafxFU6pHVOyUHNnY66c1/nybr78C0GYw5q
AfmN9fKYypVEpi+1pUiSE3SXZsTWLW9RcQW/wS82IQK5BC0jIHWwUD8f/9GEHI3qBeEIwJ3zPLzq
sDy1uvIT4eZhc1VujYHMzcaoHtxwdkVDYJADnP3HoF2/yrAuA305dO2eU39/Bg/naC4kPZVeHHCg
LmnGuEjte469CKEZL9r4HBP7Fn+TVIn0uktT+CN9HVmWv8OrU72UvJUfzWlzkEjAi4fGZdY+tVyG
ugp1yhH8tHM9cyW3HGPvsIJ3JOw1YRFrkmjJkkNBZ5IgrHI7zQ61ro/Ii6JpdYsbwDCxy28VDltX
XdAeWU0Wvcuanuow35xjTRBVzkx1CM/RxqOk6i1BpGs8LjxooA/BqnaiB/B7gu+xFLh80QPFH/hG
DyR6FA+iwi3xdpug9LbiT6DcqixXavJhNIvWzLgAlTNA+63a9zYYJRdt6aaCBpcggL6fom9ca/C1
KrfJ/SesSvZGNKWXDWe0Cek8rljclt4kxJgU4JoQeMXxmNAfz1FURmCtol5Vp22txgVcvPlQy3zf
WgqmX4QtrjsUc0WHALtYXXDf9KyB9OmOFMrXdqKkUx4f8TF1r2DsRxjTpqbj/JFcp+4wgnGpIMwk
kFArQId/cYkQ7wlbvqKJ3n208YwdY7io44mZihmoycFmLP3j/FNdhqigLSPfKwbo+TdBFhEzR/LR
fk+0jIc/dJLFJHujvS+bTxVXEy7mLNWsWzc6xkWGFowtiM9N1F0qOU6MosAu0hONbT5cboZjWPBX
jSjNU05aPb7D+W7ALgSMngVKbZekR2TZ5NLZaTMzffcXreU36XcT5ZdEBtJMdkXPe7S7ngVhL/Mc
1ZYfS+pKx36GH/Zf2h6fayHSB7xonzbE4q3dzML5fcM14w7T0Mv5QDK4Ik1/e76DC8FA8Rlfl6u7
nGuS6LDIt2I4oOba8VKnINu3XvOEb/XEehnsuqtio1Q7WtdQ3F+lL/yeB4YOzzD3lZP/scCBFsl3
xFl7Ipo89F9r+Ov1USQUX2A4ULxWcWR01+s4/3ivpSAaAicIfCpp+l3o/uVeDoRmtkNAprwPdYgz
8zXPyl5unZM+Z5/A09Rt+v+HGHx0gC33cIv8i2ggke2R/mSvmYFKqAF8EUPtVFEZaY5P7bd4dqSl
FcHN6PNjChXPMjgQrn8s08TtiwEQN4SvTjsrP88u4vNa4sAklgMA+dWERqe3AjMKKHn2OMdSlqC2
5OKLbEdEMtHqk/Gn4lScrfZRMZh7NvFIpdWFFWSjBv8BpqFS0QGQ+hJ597FRm4uctLHXxiuy+FyF
tUcZpy4HSZY9keYqm8wkHDFQ7/qbpEWpnZ7n1n8+RZgA0+4juJJ3abincmxaF1cm60gj+ylnwICW
iA0ZFZ6BfolrCor722lGflsEUOlv0cdrJxpwkgQI8+COw7XMBbkYDCt+qdZQICXzY0bpP5kj+AKj
h7QQhaOjYFE9zRs44ScA1r5dWzyHYVia/za8ykZtK7IUH7LVP0CnoahX7QK6winw0eS4W/DP6u54
HmVlbaZqkLiVBYPzhFNDCvle+z91sYqrrAR9ULJ5mqKijsjKBC1MI4i802haTzWEREaELZ21Vizc
l1DuwiEw819QJUzg8Ucd5ktdfGwGHeEgvd5bV3uHYzKg54V90Culjl4pktMlL+jGm5hvZlJVqK6/
jBQMhP5mE+4MSon2c7Iq5hQUE6z0SH+yvYuTLvkSoo04yo4Q2gD/4uVy0eMnnFZjuz0qqQEv6+Xh
0/bS/P9lGIOsHP5wL/L+96Urn2sSlc0QTGSXHj43q1YeXr0M8jRglLMd0VmY7G3bK7Wx1UsMqhXP
ZuNPP9ZwrYz2JlHYT65URgDC14EqUJltg1PKXf5w9PXwTkoVicNlFWdOZmU5TVLeysr2bAixxK+R
T8wHDD/AT1NYTlxSGpdBJJ5ChiFqalY6jRBHJWCQiQYGLIXgBr+MOD0zw8R25tqbZUEr2vFX9qYm
H1H56nxcOV60QrflaDjSwYVAVfX6eBEvI2FgP4XkJJSSFwkkC8r2KjxPq4zG5IdRrk5HdKtxXFXk
zYp6Pon/uvrLoUWZVqNZ4TDqPF8cvOqeGUyFHf58Tpu+vpm0/PVaTYft/9KxxnkEsOp0I+JB3/xS
Mi1B5d6j3E1eGYVNt/S+vdG0r8ijqBHUWVKsVegJ1lfPe2ZO9kdHJ5I0tI4MlFDIpJ572gHJ0Hrt
st2C2xjkpcWIucDRnZqfDpsQw2cgyIOGej2fHAWt1qhMDB0e9XTZbWLnHbMBwearNKmFThfUrlA8
6ZjeLxoSjaDf7sf7yO9PcvSDEZML4cHcP6uCLFOAo1ALnek2ehK27LRxb7kvQ7ME+te+Qb0oaTdJ
7OmAc2Vs/cEmR/b2/wIWf0XtHyszNVfioV5sGPmM9nOrdm6mjPPnWjx7OiHAGWJ14LPqnxfJTEo7
rSATVpt5ZoJooQpf8HOtLTMfnnkVz9+Mxr5P1YVKO+1X32wfnmx8R9IEGoTlH/rhnnALTIyPjbav
uVAkJIZwGGMsB+9h5jCfWdjuGyhpQPDLLubLTkUn60dnYu68GWAx2K98Sn+wO1Vl0z4GVF705qgH
mK7gW/oIrSfNVSGnAaHZfEtlJnJ8sCIWj5bPuAR3pfuR2WZAtGgPOxMA/KeIwX1mT9C17KTjV0Af
GY9Zu+lRoD8vhH2mGbVaJCm4zFbExtbUcrw7TMIzq0i1Mcw7zfXxgo9u+9nvFgBPxrPYS1VRfWzu
AnHY8HdHqR7gzh91XJvfnyW+2uKQPOTQ7DevfWA4LqfNanK1GtZJnNiildvGEmgmuMQbrfaovHk2
NeTI7KgkP5hukL1Mim2yfs39MzYurzLAoZa5OIMuULvXpDyu2VsP9JaC+2GMImTGAPDlhZ89W9YY
EhMuBxobtoI5uxyrKtDgf32lBRZ9tNqz1qwzYIgKx23gPcBfsAumupDQNwK3ZYZpjvdGi7vTzcxD
c5Mm3y6RFf3C8VIo/ANbwK+HrRbWsoXnfPwypkmfK4KUUN94fq+tc+87PQ6R72rOSedLDNRWn6Dl
obAZKkTK0vuDscxx9NYo3UW9wUubduO8YPjTPbikryfZPChC8dviVlHqrMOk39CMTpHhdKvoXGxM
abYIr6fQez+jkFH/FPnG59mVQdIggGHJVduqPY33PZZJRSLEGBG/so2fvmiEyT/l0IJN/EKMwSxJ
zk6nbk/GNU/NX/uIbCcuBRlQ2wyW3f71hGwnioCcYO0IMnsjpx9CKsS45Z+0LzsAeDVPI+SCrNZr
V+wVgDZCmISIoxZTSqfJMOZ4xoUvl6orOHDUhuNoIvEcnOeaM678e+MfD8uvFUSSAbMgPWH2FYWr
bEufMY2ULDdLdwdYicjMKdfBPqhcpWs+2YZecGLXp3uswsqFH+Dt4EyX8YP7MQfgy5PJFzEkwCZF
GL0iAd5rLuL2x3lpCcq/T+iEZmu7WPHv+r463oQP4ESPeb6xjgof5veGKrbP+/NcT4W9gOsgvcla
iSq1m/H9iceRwjLhUQ4MkwdYx0k9d9a2/YQaOidhD0jWDffZDBbAQ+prg6+4wtZxNROhsmZXikOf
lBfMpSCdBBOW8jtqxd8JxHcMd0FGsGxW+5Hx9+2L6qh0xngMALHNQCCqi33CIcfF4S9oqYvu+tBS
CQRBCqn2dWV1YqxViYAzbTriSQHDgJiv+lDx+79VMo/qkL3z7KfDFV/FL94Am3tX6ca8GfGHEZ0S
XPmX25rpz0XEecRWoNgmZEAvfnz0yvqCpK7xoDAl2U8CLAPtNIhF9Xmfz65EwpK6CceNWXfIv/Tt
NdJb/NbaiDcKELdaUgkSGpFmCG0Dq8YUKQ+xP3rhCOn/5qvX94VSwn6qAryAHQetfRHBNa+ne9dO
fyS674HKRoujL1G61saI2rXZ/P1W8cvCzF/HStOBAy4h3RN/+NgE8VuZn/CJLVGZN9Zs3lbKfWU7
c4SLrJG/8hLvK95payr2p6F6E25ZHjb1l6cIOeXpuInbLdHbWfPZuSEryK7sbhZw7+iWO+aBTUHN
FGPNVN9ZyZuoeoV6YB3n7OovYyoIPNmmMIPiJO2CYcNBz5yfyru0y2eckwfDBt7I85OBp1/z/WJp
cFJT4lh3cx+ldK2ZxpR+DLeEF0fSoSXAHJiVSMbqKQzTf1I+YPRZXUpAl0ikdIY8NDQidTsyw5DA
XSTOGGOogVXoRw6qfeeubaaH/98ue4kIySD/PYxz+hXX9mpEm/J/EXvUJhEhx2bMpc2am5gHTYop
0dj2iWyEGTh15tjhniKob9egCaRltDDZVkMEj41X3P3yrBWcToAWm/S9HAxy6dEumipp8X9zF9F2
VyRv307Ip3pXDKgXi75eCEteQkyIgJeyecIQQdho+HOouReELanUeod93AzxasZmHv0WMbdgaI7i
g26AbEojbdWVf9o6ashX473hiyP00PnI3ypUUxYxu1UMNo6l7KKH2DCmepsXqFw7yzfA9sQEofNL
xAq33JuaXOgCvd7HT99fJFFmJUWxjlUnUOw7HlYFUG/oHOQHwdkXSULhsaoMj6DYP+8JMBY6+XGn
1wJgLjtXYshsBC52n4c8/TKj/mKU6hZwKNcu/8udhcltIhURk7PsEAJbjO6PgEHgTC/qtEZKhBUQ
JG1HP8neqpkX9ucbVci8MciuU9G71K9BN1S363lEWMdvJmJNOo+3jbgCN0GOGM5ZCwndLgNl2FJi
jDW2VTIcInxEyFX4+OaRpz31MmX/JoO0/356it30ZTmAU8bG5PrzqgFjHqE4cBQn2Lryfhx2Tst7
iE/Mz2z0HDUXE8ezjufZbYvga8UVfrmCo4NKQ9MHHE06Meaa3XS08Jp+sPFebxsXybJ9mrT2KBZ6
c8mNW3o9OMX/ivgpEX8Hiba5J5xZJyJ1SFjzNpUByfK19eHzbOVfk/YpvYHopI7hFY6kyYnhk9NT
4XsZMlcw1cW3ZKtL1Z1j3kVjTbe3xX5ngokVyfmSHir1xopp5UWvdTPXA8M63tpSaP6n/MLiNVhs
tpnoGhdw/IJfuqlOEFTEmNG5B/Bv1Jd6wPFft74FBvlBNQIiaxUgbCGqKIAU21/PMvREdNWNJEcV
WYx7CiD5HKd1If/Nq5coIMPbBnGaROBua5+4qRhTGaBVtEic/pGwsBdHcis9xlHQ8089ozlGqyX7
XJ06opVlQsmEnXlEwzpvGsgL9gawQ0/bAKqQiA+v92B/9tJJ0lhbjQN7PlfQaWDiPf2S4v1Eh7SF
Y6GDnvIwR01frbbhicikmFe5IXB6HhmoVIdnpkRL8j0T+c1d9f78wMOXItRb8fFhQuPJ0CHjCLL7
XBeFVHOeBfmt/MZs9V/DMaKtgGveGI1hnxzJE5bc1+jXOuEqhxv/siCMtHvai2ejXb6lx1rFezkl
NTQgJrmXw5snTc9OmGDD+Fd6hCe9L8kfdMPjTZt7jaerGa80gD5BoWy+0SFECk1400N1FT10fMDp
E0xGs1tkDEYxOYEykskGEuvbX78ytUAYpm2Kj13LyaWykPN3xMXKG1lMFLTprSflYJZG6X6M2SZY
GGQk1XJzPgyFReMupI1IWAL32Ski19delF+rBw7txki8BwjlTBpDpAnE6M8EUtJ7Fdloq26h804P
0zzH84sYGamHvm6y5oHeX5puMi33f0y+4I/zAEs/QpOFAU9p5LEj/8Ee244Ed2eD8nxqSFNyC+au
Y06DP7gpC2V+Qe44YN2i3pYvTV11sJKZ+BHKZ4pNMuL1Ru1jpKpSR0TvZAwRid8x5n5ypUSyUSWy
au5HATgjnRpOpoZ/IoiOpCu7Z1TiVltf1K+8iOUsPUIaLvmqnETGYvKCL0a0oXQzbMMYFN5fRaqc
oIipOgjeEoCtlKSaatIUobxBe037OspdwOGRWo7vSAeqGhE0ziAl0bEpnudswkjsPs8JsGPdQuDZ
KFgKeQnAaF+Muz0JdYlNdKkPkn3Jh/vRouarxzONvg+3k/Nz2IeJ9nzXGrOha9E/k3Sd22xeSmUO
d9VU3gXjNhS87y6TwE91rN4qMYAfvO2+3iwewAwGPc4wq1OWYX9vNf43XjOlFt4OtAk5rZDYgl8A
qXT4AIcP8Mteo6AF4WEleOnpWGjj/KigdFiqnSQOHJIIZHg8HBJLy9aMfMFPmAd/q9KZ8K1cHjgD
1ma2PDPE1E9oOxY+Man2KtSSdkG2FsS7ZHTkQ+WUMmDNqHZ6D7OHiQu6z/atHtmHOaeHyWMqcvPF
zP2OUrK5xNhqZnH12PHDGmzFYqvvFyYFWnmmXsB/cAL36h5YtbL9BcGDNDpV8q154vgeOdP2IlEP
D2pFW+Sy5UMaqHGMUMX5n4vNVcwffockEAoAz0egGtkKPafHgeEez8kdAczTtRWm3RdQxaO3ug5G
a1KT+C5EHFWU9dRndlAvUIkiVE3t8OhYj8xd6ZNWHWT7kMQuuoN00XCYp346VPyKo7IUFetstwox
gO9IOfMuOD0Wb1IYyw6hE3vOAnSZR/Gf3qw4m0iTo45mqUBw5VpRhpCx5O/+jCVQD8HiMTFeDEOY
w/C3c4DLoeDQ22piVVMLcrsi07uP0Y8U6jd4CdB6bTfRitMyViIQP1VGqjbhpVC9pB0vctMASA1h
XZMCIXOC6n0MIEL4rYQ5ta8295yJnk6I1Et1aMAs2ZBDjs9hX+jm3Jn9URbr1v+93b6uQaHQDTSr
kUySSY+b7BlQdapPGdPMuZEW3YHaBdltE1D46ILv488PXDXUtmcKcx32NvtDcfVQeIBcvFYDNhHk
dbCYKuXG5NU3JN9QQ1fP4F42Oc91X70mIGk4jpB5b71BHzWVwk59wHKWAwJwLVxCUgxUam63HSxz
OaApU7XWFzscVLx8pjQTHNDsNG50HwfDp8Xjz4EQG8RBHMc7dsJJeFMsjdJ9r6174KCIgJIO0fgs
oxLQH3LlLYAKYlxa2ErKbDHEEwRS8d5Qm95W8vAXkZmg++Nam7c+4G058Snf1Cc0dqe8wMbUJ0t4
WXmecgJoT1grHlrmX1d+R/UoCzvUB7rSXEoH862R10vdT7UQg7ss3ntHpQAuR3DuAfNf2SE9Uvsl
uZ2KLQi+spCM2k7qcOTdqqcbDjQXUKAdNvoruLKePH6OtYljkf98QPEDVleDemavVOLHrVW4Jr80
vdsfzMgvZ2F6vopjnGyHUNWbHsWA+TP5gcaN0kLGTmmfdfPyLtuF/8TdO1JOQpEjP9BqQ9HLucfq
PRsqC+8IRfy4/LodWJxVnAAEa4X2WTJiePHS9ynXetAfhuBHBDKU5GVipfacx+cjUMRcoUYC57xe
FnRWmx1FHm3siA6WsT4MmLoCm3N+K1LPiGAYne5lTyMnH6vsMk16rKRJpENoqFZ+eHnPhDuzlZnT
U7/9fzkdIf9Im5mSuncbxK3UGDtSJDaL7w0IGv0x6JjD3xlYRTJ+EgVn4gV5EQKEYDXlrOZ3Iap7
hntiC31rgudyLQyPRhZ1lhbjrbyMbJXKZKxFjUGpjhpJyl1+LnWzH+67qlZGax2H9+4sdhkKlqR+
c6qX2kJAxiz4ogBpvLOiUISrZ5z4B1UsI/LpU3p8Nc4UUBrHgCBT9gxHr5Re6gaYoU0L090veri7
9KkJbK1p0uP4WrIH3avhbhYE7U11DKFhuO/mq0YCX7YkP0CtJOhN6MzuDzdNNo9mYK6Q6Id8Wyfv
mpZ/1op/Hdx4Wx+RTVbpfnHG3pQtdm1QrjYc2XSOsWj4N/s5sua9g150vJP3S0ySlBsoebbNB1qu
MVoqmpO+vip1xfxD7HM2Z1eSgAsk0pKSI5dCbEm82wcrB+NVI8dTwE1lqgBMdve6E24ohPqrMgsG
jf2BauoTxNbu5b6WraWeyAbF12SocXW0GWcbhNR58swSwwb5Vgkr8Mc/gxAOXRA4+RA8slPATZyd
0KMyEiaFgdbpDDjOxYyYsd0RwFN5Ckugj0lcPYdTr3STJk5SRCieUhjG5OpKWU76p5lrKrKWFQyg
tQmWtWidt5gVSerG9493uveiDupRqMzBz56d1xxVwC7YhpZItco9qi+A3XScO248u8ObxUxggfHj
tMdKXy3zEOJcJQ+C7pf2+/HN3pBYkLQs4Tc/c8R81ujLRGaAG5kZUdO0/O3XlKrBNnVUKQOzGlNN
HzUpuja4EDXMm26ks/XyHJfknQmCnc34hIBBL8hyXZSUK2KbI3Rdc/q/O9MkHOXEwbLZRkon3PiN
LqOoQGlYJO9yR5SrMFG1DuHQzto0YKTeongN4AeO2EqHUL1S67WPAsGXdMe6cuFDjSKYfYDGZbt5
3Fep/nn32C2g+11360WNMMyCimN6K5vJ5hJhbRc5W+D/0H59yqECuTlYag0gbMcnCvpp8JpV8cFI
3BFQUN1l3TED1JcuojnvmYnquoxhfXYPNf/kdNgaBZymWsA/NmHs60tsot8tTef/tZ9BylvYb4Uz
CTbTdijnxxGYih1LtPPDO0yFCYRJN0VoaZj1qY0VNNYVe+oFISOl1+xLPqPeehXLlOW6cjY/6OIc
WJqX8FEnRVozExBZLgGz5qqyJt3R+fUE33oamprefAGp36wlz8qdeZ1wHKb2inU7CP+Kvj8JsF0I
MUIon23hZVSPxVxRFX3SwE7XQ7IhhC1I+u1VO9JtgLCEa8HdenWS+zOoQHMNFXWyK1GozfaIGcek
VUGR4znHC2r/sKzNZuYB2pnMdJktaNor6wh5aP+vQPkmm74Ora0bEqFvaPcnssbKCMMfCV1UfMOI
9M0TfILnsmRseTRMQ0yB3e/DRdDK7lz0eZ4oP7jfkjxnUU6v44HATOzXQoNBdW7NBbzR4fMlq9Tf
OvhGRpsfVyIlA5PWFP9UiKO1rQpYMox7LFexLw+BEA2PndDIdxFPVgHAxu38SMfuTbAjghypL0bL
WY+JmUEi55TP6GzQz/kLkMrrbjUGIdv0SdlrS9pQRO8rkkpG2B+gBK0URL7GOabHX1EQLwAqfh9M
pKrEZc36D+bU/vFwH5hGh9/9rVUBNvnMQTD0184M4gE5RqQZguSGgmJ2x1ToN9uTj41Ro4g8Uzqb
LHu9kKTm9S8duiXHGjsZvCGGi9pw5xB/8VLmYi0h2e3ngTN0CQ85kH3g3pokfpMcqKHg+m+HtWyE
nxHrz6+3UMFpaWuqUwec9XX3I9lOCTbZtW0wAusEBB1xGso+aByiL5+WCFDaOIJvQo7rW4HeT42G
ZfYLlTW1xhwggY9H00dsz2E7b7FVNYT0y3HALv0b5xe/MfiiUBTNn4XgX1EOVt4o/vZN78L/WTGf
c9j4Zlflfd3QeCg7tVxcgcpPRMVBQEcrw4UKZMoEdmuInsCvDfSLAWq7UztjBS6ZM4jrPfsdVX9m
5R0/8v8drCxr2EEyJK3uMLzQnNucrfxPUzNEz8kt9AefyLl8Y4tT0F/15c2CXslsTPF6duaA5kSd
M7z+yg3af++tl5ssl07M9afOjpjEvB6TUgLKGRWNkmTUewXizaZ5fptO2cQDntbbZL9NwMSZBn4W
7PS00g/K8xf6TYtosKJr/ABhdC/CyYcGrflA/tCuZem51rco2YJXmTQj8LF5zvLQBrRcpXkJeznj
ukmfepWa0v+NvIqX+j8r6i2ozTM2EjmFL8KNkKZAW5QuUbgkoCG8mCgR3i3Fv4C7M1mmbmJ6N4L5
u+TWZUaANYO/Cj6Ni7y7xWzjP00JtXEroFAVC3f0sOgF7IsfSsj3jnyq5fWEExXLkSOwP0KzRq5T
HC/nT3noyDbLq1bsifPUHY1O85O1IQ3ZxWKx65tl1x+6fxF/BkV4w+rmDrZCO1Dx882a8RywPKfa
I0ipIYJDBMitgey9PO2nQ3Ma2Hw4kbmRwBy4H8ZqQQ5dO3DoFxDdKNPSyHSk/vzWGUCVD866mPes
M+N/GWRhVRjFFVyg2bnVr1Gev7wtgAZqUUjKnsT1h6I0yuMN8IK1Cl2d+r1n5dO2Unu92DFSUEVA
qGbgqyhJ5tBo/VvuLa4c/p9m60ENTueh8+WEzqoDaxFKQv7jgI7mOkQ8jpfWLtJ/dRvxw9HY330l
0qHFH+kOENmz03o91hSauEWVz0Gr/8XmgBPgB7d5TaNbBL9BtucB6Z8KNmNOiMjAJZkU+88uJDgU
UKu8fOTiovBGUy3q8T+c+RGmCM/2NS+eCJ2TSvxBqd5LVW8yIxs529kaLXYD6TMxQ0rygibtw3c1
Ut5Gi38GazyKMiG3H7ALk52ErWrHZWCQmnIACGOcznqKReyMyHJ2GYHOVP0V2vRQCNJazE6KKs1N
G8GNDD89WGcrDkAfpn5E/KMfhSNcPPMCrqIAymnfzRlqP6PuMhEpx/lAywVSX9nPHWpz3vqlMwvT
PdIUQo+L0GauEHx9qbb/dy4fGYSDCrp1nctWSwugFk2JnSxM20fB+x1oIcriHASZysj0TqKqbSZ9
PNKt5YnP1xet03Ewpm6dlxwHPS9z+CVQ7wJ0y0ebjfjK9pZrFvCOdJ7b6RStWJLNQxRQSP9zZUxJ
S7fujXrEgcOyk579Ke7mcEHRT8xo9vp+8LisehzUd6pg60Q5TMcxbh+oLWztftW30rWBezoqkg7+
eSbmmLrGXeMpYvRMYkWUW+B69dP4fNAsfTYQvVPCGTQDB5JWtAZmwW2tzAaaxLZ2udOCNdvAowSF
HZ4lXqsCV4f9s6bfq3duSqQen3aaSMIUnHfFc56O3m4k6p0zz8ISE4fxoKpcwTgrhIxAVv+3FL8b
sTWmmXAhNg7lG+trypejJmsCJCQos8KzsARdjq2sq+qSD0u3FmPHaVD/l5w9VDHKL+LtvXuCTSHt
ass1/krSG0eETqcwT73EztNad5MnJS+0hX9dAgBGEV/w5Zmicf2RiBVHM+N+uzQ0WyoP8zISr2+V
x1RcFvTJexuaw7qtwNoKP5iFvlTr0cSW9NUydzgZYG7XCT/HBCKvOyU+xChw+To41w9Gt44MSOK2
N5fHhuZ516I1DB+r1VBAA51m0Y7LQP094NxWOPPLmC+Qff/LIaCL3J8sAgxg8SSG9jt1VZY4rwD3
Z6pkUn4aEB4Gu78Z4sNvDbm+BVg2Fw+mp9uyy47M1Onybb/gjS6BZU/6Qp3h5yphuus6/Xv8u4az
SHiEcnlSgw6QJD1PWJGVpewRVWxrcTW6wOTVidAWiPBCiNho1Mz/IhLr7PTrfnfn1sgnhbvM3fNJ
0K0GDtupP6B2sHJMMF5SqTCfmRUKEnmoxH9hdduCWttFWBH0uViucMYjgX1avFt3PnraRNtjCyIH
OglibJdfpRX8Tbr5EeTkoDBVtUJtcFwVgR/Eb6mzvNLRaM/nAixcbFjREBESHQqcL07s6J+H8FKM
oiIb7t3621HVJQK4NEVMczpUq0d74yIaizHSiOkrXXGyYIrR0Ay7ikifIQNDYSlmDp6r0F3dumSg
muU8Mh46xCx5OsPMd639+nKt9jLUSCrB/uMN0Ja4/zdoYmxZYhF6JB0y3/9asSdtcY24AaO66TDW
iA7LGErIOxqvP63P21q4BkyunW1Amw6KE1LNAo4/y8Dr6MA1Haa2OFvYgEVmtP5mZ2P9L9o8h6uM
6lCvzZij7EWW1oBjywdnReLXreQdMBYtzdHiSn73Ce7djb5BrS0Fjh3FTpKBcQH/BlrjtwzpSAoh
zA8fTussIWdP0wFrtrqRsjTE5htV4k1VrR1xY4nwQF1tqfsN1E6iQVyuz53X8kIAGcGMRm5nVsfg
iEYlxlBY46RRVhnrbshmEbxyc0S8pnL3DjAxZSKYuR3+OSCYJ3mE0jGMY+H6MnjopgIhjJEU2SRz
fYdvJhK6yT/u8JNMfr2DSN8Wm1trDO0YCTKp3YFOxexgICfJPrw6BiGN4gqWrDBW9Aga5SA31lXK
rRWWrV+BSA8Q042my0ekeg0xIbe1W2stMruCadWXKht2GgVTxMEtmaMXNUEhRAU+a7w2qJ/b9zSL
LKjZR8PUjcjikPFexB8uqhmByimy3fprFJBzSNixEBH3pb7GVrX79EN0LLDy4ODIcoFCtd5UiJMo
YxZ5ejjbsyKgquSKLrGcMcl1/jnJpG0Bd97uGwvK8FIDmuvrSsCUqRHC/TPlz0e0ZoUTdV2ousFH
tC6NBgXGmkkbaxL8VFaR0wkOhw85wDoAbS/6qYtpDAHxqDw5Uj/pp5DkaMRx5CprhozDolAual3W
iACCle0Xt2R6oNkFz2tuHeSnM11czMpfN1zu9LwTsHXu0+DYgYsMrVK/N0G62iW/0WE/+jcEaG+w
wjaipDZFnOP3NthMquAuFpgqNuuonN+HslEbFeoS5MP9+OPYQ2j4AWP6Kmet/9eVGfvfkcafNrKm
iciAeCeedfJRy8yjT55WdVfruw8ZWkxQHGwvVkoPHzeZZR0TfZpjRNETKJfUXEPT4cPRmxxcHsCG
07St6+sCBVpawYvdQs7ud+Nb5Yj3n2MTtSVhxLuTMiR1FzoCZm+ICOt8+yV6IT+u1fULhB8xHjZN
wXCwuzp6H2bPIGM0LlC8p8hXgAyNMS2mdUGbEML9KjPraMIY26JTQGunJfR600W3m+xrQY3yJyMA
4zmrCCAhyCjAqwnkNiINs6L7ky2dh690iKYQNqWN3pmMM86QkfNj+aNP0visE6TDE/o/USxPOGbY
X+qyyCweCRv/P0+gofSDYQTqfrpM/wudLe7Z/58lqoqxd1FkPgH4O5jfyRgwdqmnKDNO10qLFO2h
8uUzCoBdefX2DwOToYT+RGW4RvCO8ZhpLvUAV31v087kiigRMbuhX7Gj2xQLoAnquUR5aW0VNQ+0
6xj5TZNNSl6yGNKGV8NqHmvXkfzV3WfF0urSXljuwNq2D8Btos77DwzBxoI2nXXYlHdxj3wHvGEF
dhWBzyjVHn+THIyUCsnAsoV/w8AhmioX8S6EicQPi6lJDSC9pnhJYUhjhomX1VDuOR/n7iPsv8hL
v3gaByUAidKijvaky8qg60SfNU9AnYjBHM+zh4+VAv1RWE9KWbalAotW5DtenmYgvkWYCySReYGf
bsajl4vkLtr6ljnh0MSjQcPoAAMP+gBwpywqIPQsbSdBgkV/HhFYikuOsbwmv24EDziGyOi5+iNo
B27us3z7/Yl8ikMwzppu6uTEX8lLdyOWHRJKLP5pRyhNdyUn3kTg/ALR1IVKShdgAwtwUyGh5L8X
AI/bx93w7Fbwsq9XsFkgZj16AubLJzixi0yhCQ7CdJyKieWqzM9Nq3wRzWtsMuPkIYDcGQBxDNPM
t4gk/1/NZ5Sa1s8y0sUZfMwqIEcGXrzoVl4zozMzC/o9ijUZSJxce8aw7sUGz5I2GqwEj73+jT7y
XKtNL/PzkhRBTYl93dNQM4moMuscs1C2GMBifAG45DvWLRLCqmGPzm3BphqkC7aYna1qDAy8cx4g
EahusC/fG74VQKPb9CnHAuox5dcv+RoSEczN9QCm2tpua4CWT49pk2yRc+7Z/3KpHrlai0nA0jcu
bl/f/HYbkqMCvQk1SP+WOJ/hTiDqj5lDR1M5zLxWgLFWp8aHkripGzY9tBGlv3CRsz18Ext0Zoi2
Jl9/JHkjyk1J8OkhhaoaF9kjemPpnWi3l9174EMxR93Vezu8N/pAp+oAk3NN/dIyKLz/kMr1MNsx
buBgnGw+tBh+ce/tUt4SGBQ2/fY89SzmNlnMEUEoHS89f42Ok34rLAeBZqf+ZnxtiRksu92fDs8I
mNjHoc3cfebtIf0suHF6vkRcnpAJaQYPs6y2/t/vEmyYlASo/HHzgAbhnKI4+gQFZfJpwG0ZWnZf
wpJq6ccjln0bVgL3Niuu6i9VckXzL516e0x9eJz9Gzsu4hKTNI/xnZwR6OMMV4OnCtXI7FDRFS4P
3LurTkC7NeglI/m4xKtU0fOk35btN8I52qIaMJELqqiM8SN8TSx8y5s9pLYetjTbKxeUmATzwJ0s
uaf+uzds3QlhQOzwbxdi20SwAVyvNdC+mM36T+5LaaCIwixzA1u4t7G2Enyj1ipBpWRHYTQi2pu7
kmN7iTxtM8guEZrrmO7p6msTl+6VyPPTLyBpaSZWzcePWmRRiS0MjJYFeKmSjKNoKx4AbSBXKerJ
2yEFLUSNJMTgYOpQVpuowBiY94mzhekz7pdxAa7FkIkoBgdUo4T9CmK+7wCoob5NSIyXwM0vrCbp
DmLeEs2YVUBcLalXG/RfvUduWNGmOWKyqMCf9RFK/o4MwwTgtGFXQsnx3yFQxM64ZbKLOpfMtOPo
am5/E6E5GY33Wh1F6DBuiUDPl/JsVCfOVx2Kf+KOiqZunWDLoS6FIJRPJ8nHfCd5UZxDBoC/KOXo
hgk8jqtEFrH61bQDqaA4ujESTLoHM+tEsRmRh+//5GxsSXfsv1N0skeK6t4GN8swiFcKUS8ddtLV
kq3pRUwKK3eMUBqF2stqMbXtk0Gfa1pjAx8UyPwldT9Oj+CHdnT66Pcwv32FCYDE6DgEaeDKWoQn
3nZxXsUSXPWiYn85D2fNN3f7p6syQeunPnFxK/d+b8nQ4Syt5BaUf8sAweAFnuxI36CKUTGTVEpt
QtXvZcsXwG45HaEZKGz8BqX4fhZvkJ2ebpl+dB7jIadyGFm5RBfoYRt1Utgvv+iNnfTpIzBE90tg
cPcX/6oEZt1I43uoksR7GC4EMYxyPusN31DzMMYl7cWP670QcaYqoW9jA70h5qvPcVBisRMo5SCK
CjnALz/QRYhlrc4++48nOPOpYS/lcpAnBMdH+VaDqpwD72a9ScXOx6UiWdkjVYCC13MLEXPfRvQn
LBKOO8fXFFzL9bPd0g2SV86yyAq3MZNSTXBjm93clVHSzo7CXjyHZVMfOLUGzvYBvnXMr/YSIc8w
4nIAl2YVYP91UTioeT+AisKbn3xH0f3ttEFOHmfgXga+mf9jsphltI4A3o+BpSNM9T1p/AVa/gpN
57zgPhvUYA4R0f0TazDIAADjyl4Lq04GjKmR5Hmp1PIhjhtYDwZNEvxyNKtgavn7a6+ElimwVWDM
UDLkYK4ZLpdQ8aRM+KHHr9bplmA/v4TGONOG9KK1cA7EaABJDuOTyAYntFnRHwBGBHmaZghvC436
bnNwWY06Y9kNgbGTzcG4b6NpVYEcg3kPO71JycKALqFONeEiscEdp63SfO5JN3t9hjimNBcFvhEs
bVk4hHSKMfsNcAHajs2lF5cFjAtUPkXRGUY3y0ktK+6i+bDxUve5jvng/Lpn9uT0Wqo9wpYhZ/LN
PYpDdMl1NM+BAavRTv6riK6xUcFJCZXIV7qwkDRBlwbrPPLyXGFKKDRsUzjM36vRkNSXrmXETbv0
q8JFM7h+Zocer0E6rLfRV5D3+kbfucO4j7fO4NTOFKS/mJHooPmaI33s73o0v3qvBj8kOkuD6nAQ
GDLGq3XKg5vbFRG0KWzrqDUpRyJpejYrksYWPYst/HG99ScKO6MAAIx9rOuqLCVU5W6TNr92x02Q
y+hTIqG82jAGvKPqsghmry3Huo/y6rUfa7j3XGXqpJBGM3Zth+mbHCwjth0EyG7w5/Zx0OzWP37s
no2GGcRik5g3/2v7bop4BwIquKpEADzl/9KCOW/kh8DJw04i14fTRG/MZkqbQlHdCvCXY/R3xUPA
UDn8z7YAwBHhjtUeNXGCHiF+uv7FvRqCAPNH4oaTzDTNS1crvJlhM3QnBdepax8p5jDMgCck+L6A
gWJ+rNpz0uUI01wC62aSAb70J5yOJAu+dL3otNRDQMDGeBLSnFDTLbqzUauuICIINrCngXMDN7FX
0E5H/T8wvblxxcarBA1BkMhtd/6LlhBu0Ii7yJDnW8hYTYNhHYTO3VBVmouvghcEzh/yEEbn0g8O
j8l1oJ8+cB+KmkF2S5MV18m6xI0JjzsKngEvI+wILLM4pYWTX4ss5CSThf2j6hfp4IOlO/aJcGiu
oiyxM03RUcEThovesBjWI8nNlnD1yjVbSniAHXM4Y97mEy9bRBo6YpWHwI1VWL9mOtoTgTgqsKt+
pSb869Y5XzS0cj2d4gGhaZHnbuOWylHEI2Hho/HnHEwSeYFFrIogX6zNCtSpQAffD/QAOCgfR+Ny
DaHQZMrHbaovG70k9jtqlF3xc0+EWg/antNpivJd40jpNjUQFbQsJ+EkQEaCMoQDpNrVdpbpIiuh
XPCn3nwErGLSlMfZg6+hNxarB7diEKgxyLcxoE8vIEjAw9ehKHX2Nj9BPxpgrB3vkA6aIVptWh4h
tGV4C+z8ByeJkX1qKRQhvwWL/Eix+KOy7GVt47SE/WSsslanHKhF98soZI5NKPaPBGgv2yPnuFpj
SVmJFhNjoNU9V5B87ydK5H3tsLcuXgjLtXffjexHG3rg/pNm0WrUMLC1664JQ2NJH9rVGo0K9YU7
PlELtuiPyy3ynIAvwANdfKx/XKpVcc2BepJoTtt6WzujY7X8Qf8IJKAKxJXR7j+GYDMt7xl1WsP5
lA27PTq989JPiPgpS1E6rhcNfZKZeXLGFcqW3na0I8wEsT8uqgbPPy1IFxihr9IJsrBlH3Epo1D+
dmQCW9hQ0pqV1Qgu/p9v5fNhgt3B0f7IWybIZy0NxsyOb/H3dAz5myPtFjc3iqw/XzzewMa2KYUZ
mtOLuEJUrh7n3FnTx+Wz+A2U4s8FTWbxqzBzQXDzodNat0qOtfxNctTeVDoQQ83TyY6sfHt7zSsM
dJGmWW6xaio8uFliF/dDWNMCwKWdHiv1DZmDUicRXKicTiQT4yjCeHjrIV1fL1lAurgz/vAaml3e
xdY9BA+l/PkapJK5n8A9uC/zvXhZkdmZ/jTAJzOvSxfvYTOr0MPIPdaUcMhO5ux2cFAt6uVE+rc9
mmEkEbg9ZqV8Ylfd7C9B9QNn3KZvoGaNORyy/Cl4eQxqyTJnyQvo6FTJP5Xj5Ae8n2ZIkFhqYj8G
/00SD365IEi1M8d32ti5oKR4ETvmd6JBTIUAkzNkw1Lqks0iirOX4o8243eGuKn28UzTiHTj3Ax9
FbKIgJe9mGjSF5AT/WtcHV+FTgr3sMolRZGMJ+B+Kvuao4L9AZtFT+cI5K4OiTuOm5IEU2PG8Cod
MlRiLexM210lvRX9urowyClKtdi5x1ZC4f03IDDVNt2dBX+JookK7EUTW0obWS6jkJ77mJDSwMfJ
TJ60G/xaNd6jxmF/RW28G5uB5nAiL+iDyLpYVUcIsT5bIlMCChEKFx6gnQSp8ScCB29ViTyD+yEP
danXNKxgeLAzbfs6O7d+BLX2TKhQH3CDNw9d03LLIY7L11pw3vo0FDzuaEjWDp+LhymmSzEghX8I
960DGpt4VeY5Rqtknuo+svaY4m+Xn3B2KfsOcSk4vlR+D2s3fEr+WGbzHwIOaV4UVV17Uickmz8s
GwGyqd4ETYbZcTVOSs3flH7mNdHKGr3Ueongx27qiEvWQugte8f+2UilU14eeWhXVTWZAEG5wclR
tM8LsyEEncO9yQTcle/puBXleOHwEoYXTJYCwS6/ObfnfJxd9bnnh7omW2mnnIKT52AqWhZF/mdq
5ofvstvG6ud2xX/FradXyuyy+psYgOT5m6D2Gk22E6P2fFGJu6UK/RTNBKx8CUFj8RMuSn6dzaMq
lXrw8VdlGC0JYmh2M4d4jfbY4mPRKOUhx2kQ4QYEBWUxIa96OwPG4dmPik9eiCPs8Bc91Hn5brWY
K7nCOd7lBSOs+T4XUeZKTrTQDEDlrz+cngDp8VzP21JkgYXbc8KCKVDJa17M430HPAfuFJ2trcKt
w1jlp52EIDke2OgxCHa379AYQizdZsfF527zbButN85X3BOKzpqij06Tw1VM2X7jyiPNjv9F86jY
P01l+ZaGeAJiGe+H2edWaIvi9Y2ic/6llPE72b6aWbFqUPYRN4GoNcwlyhcrScx+3V9wzFExocXt
FhyzRLUxaNbFl0NXX43yOGY7TcyeV4LnJuEMNv1Q5QJiqiYUv2MH5pVGa28SaxWusPkYzcv+5Hre
KQc8+hjXKGAog3tOgooVdQAptQ8zPaPhQ+KKclOpiaSf/XahmBcIYSGSJt5beZ1Yhm5PC9JRV5Xh
1uzVemxdyGeVwn2WQcykWT90f1DWHDo2WP1cwO44i970wl9yKUF4LvZti0Dzu5Da8JwdMjnEATYQ
UfnKo9dWYAadNSsXIWl5x/X2Kb5JEXvt3OLq3WuDEGy5EEWo53tDAsLRdRM4F77KP8oKWoKhW8Hl
RWfC0iSgYAYWulHTH0dRmrWMtQZwNLhrhLWhODpJ2wCDwRNlgPidRSJGngW5azkVpJcV9hV5fOUc
2iN+B4Hrgar+F7W8R9QeQOjuQei6VYoga1gkvueyLlHovKtL8abeXUAT6bVo8J2KIgy2XArU1Q5H
AOoo48BXq+QGc76ZkUt0cLtN72Dxb5hIc5tFMVTVw/AQbEkSWDKacfq1kdSOm1Lu4b2uFCo9UKHy
u5Z0ArDoyCeDoFBLx6w1z8WOcPak++Zpt+it6kB/LCSijc42H5A3eh2UFxKGGPOfysiWBfPslzyU
RnrBsVIgdt7iJgJNxguRtDxSZHQOjBv2CGOdRgF31/gt8EJbu8Hz/C4enLz/3M1J32XOn+0fCcFU
ulMlgpkXQpQAlyg2Du3pYG8mIva0rMkBfFZT6G7sz9PfzmqB0q8F0/FSxTsFtIZGNJEb7eSqe2GV
0NJdiJGEjNZ3djzPfwVtG5EbjhZHTKH44Q2TE08ue9W9V5fqw6F2j2IVQPa+u8R/fU/7wqhoIkyf
Ty/3EDrX0vL5i9Cl5qIOed1XCIk5D+hihfHy3Nmpx4xYTsO7sxPf5rmR5tbmzAhz1CMiVRjkK0UL
znlYHEsk3AzcWNkOU/5eNstc7zQv43tTgYtgbCMJpsoay459ZoBeUqjKDsieicwjNX9nx4W2F21A
9/aDw1j11o7tGAEMIpP10vtNuKDgCkyi230YU4Lg8C/tgVo/iI6qD9lKtKFCkE05ypGA+wDRHeGF
CwMp2a5Jh2Srs19qMay5BQ4nGzfTwnhu80SHv5WKypNHDomFEuF55IxlRdLKwHMoX4HSDoqzDLT+
7NAY4aR2Gy86eaV0zHYvuWp/lrG0iT2VZKsNvbMbZABtfmqWaXX1dbUa3mH9jT//FFy18m+ZR1V0
JmqfCjVQwyCOTbeH8KQcx5FLwCqS2WMkDCEo88orM/8eETgde8Mf3vLpCdkF+5XBhNGU7ipOccbM
9X9oadef99J6yZ1HQoAqoKcaCrxFgvmmu+a9EwHe7+WlvriKb3NCJPxUjJ180FuOutRijGs+SaPS
oO1fduseBX2vUTD05QL8skdyxlxFjvrZBkjkrEH52Sg2ItBS6fPNCyFTxi5YySSparMTmjNva6Rk
xcz+GKB4oRlYNPtwJ1P4KflI+v0PWrynUlw8rTcYCItTr5Hcwd/9C1H69KY8GsYAb2DrI93Tk4Q7
VARAzZyZKAVU4+VOKTQNkSgKmln2EpLoUKVWJG/uH+nJsGCZO0rzNwV4ZHY0Vgc2t87/rH+Gfzcx
NG5V3FFV0zqTTWmMFmBV7ssHbm+BcredBUjhPo4pqlP2VEIJsOg6TPnwyvdDc6BTFjwBjhtDCNu7
MnejZPg0kZX56SozzRUTcBQhr6sgz3zs28o8IY6FIjk8KTtJjcroK+qTAUfHOY34oVSU7fbQTPGq
UeybyXoc14VrJapomErQxdYwn+6ALduA/VY+f5dVT+ClemfFxT/175R8CaDsM7IOzUKB18bacE8N
hjFRwK2D/Z9ZWJtgdN6ZeGGnekB/igRoOkaCrh4HovEkBeuB8WNNh0qtMl5v7PHmOqVtHL1fNxON
fjj655umdF0vnga07lhMCmLYkn6tW6icfiRbogZlAg2MLb+I6kli8QTRhhUDPCkF5mYljzgG1kD2
2CseF3dzYEhI238lopBYfjMQI4oosJi3CsF6508PSbRV/Y47W66N95nMEBjKiW6VlvA0gRKKKSmb
vL+s6kK+U2zwP6dte7dqQkokWFA3pKZBPEiJTIN+l7jd1L8xu+BMI4DFLRF7XqvyKbuDQI5soBUk
pkW6Gfo7DS7QViuoFXHQo7F8ez+dcFxdchznvvc/Oybt194DAN1l+by1qIWF0yBuSWpiwEjZlbSn
hKwCTNGsJqh+0nYxeHIPScYhsQgKV8UcMSwTv8iKy54IT8IpcjLLlfudZ4o5bJDZHrQp73Gt8bvU
QRr0TvrEiTmmSlS8/SDzqn4AtW31iut345l2UzLHVTtP9BdhlB6sI/Js0F59Cz85BRgSTQGHmr9v
0qhPHZNdhbIwaefbs9SwFeP5qZtoujloDerMfJC4g6aVf44nZ7I7YJ/nw+q3GQbJ69AcGDvxZNQG
8oYrB39t7QjoUunIxR+cU2irml/ZZphbxW9BlfiwhnmpunyNZ83WfeUNOhZtrBryPhn3o/BWi+R6
BlkPSMFWw6jPoLE49COblRtgPW9FGfdrwJ3UZB+CHq8iZCMjZpiDkHbGJ07mqKh4wqm3/zL0C4qZ
/KtQEP8DhxAtU37Qc/7Ta9kXWgPbwiR1JBD9WVpGTp9mgYqGc7b7AlEjn8tPZRhPr5TuFA+FXaaY
S5xcdsy9hwDHCC+gAu9Nv8eMkdEvi90Sf+4w9RxvOnVNqSeLw4/un8o7NW+ZNAt1mvRv+OP/g3sN
pwaweTqUJgGFvrOjP7tME9/5bQ19Y/9GnBNwX0LFRP0WUkISGxXsjYNyKAHcnL5j0VavOAHEboYK
hi1P62OK3HClf5YgyS4FwIARsheVEL7BycBoEUp7UwTm8rQIqGrn7iiNXF74hTX7NoAF4x+NjPc0
ke6GC3PvO6d7TVBpjQUDCwYs8j5NEG9G4qVSR6L3a2g9fQAphoDA4gaU+PpYq6pfSnFsRQ7e5DUw
rRxpqmPr2yxqshE3jm2aGARlHLFhFCApwjeu/32er9lhlsYyEfTmLU+JLLjNpX5ch1OQUrlhEMc1
mlUjsSeSTRelqXhBTYYszxk88cjMEQFKaUtZsKRBOdJs7PDIXmJ0maooAS0KtXo761GAOYtQTx56
7SWupHlu8BrH7PgDtkDvyBOtnmKmOtcKCf8Ts7LIFt+ju6HzwzssPySJxBidArhsDxWXGVApCEZX
ohcaV2PN7KMF+7tpGVKczNEPEcNTqfbKQPO6hT6WhlfNZSq3cKuJxb9TBU6G/13vAUZdHuGrf04a
ukEaOFXSxbAw8HFd1/uBqxxraVRVl3mcqGH37fVYP1kaa6Z7f1nZVT3/rXzunDO0Mr3Xjabe7WPJ
S1kEugebmXwE26aRTc29z3Yk8XXxPR8J6GvtdOHcK/e0/BNpiFMo9tOIXSBNBjk9DpnDYOK3aG17
kxhwn5imAi3F7YIseMcRRbcvDh+8ReN7egJE+3VFkOimV0gCVJ08y4ghpgFwYAsYvz0wiKv/dJ+Y
/BGbHAP+lC4wFcS3hJFEeK8QSkXOKQYjKzVmvNodwnf6/M6m8oiRm9JpuAFOevMaSJSK+nN/GGhz
z/pBlhsAea4g07JNtt5pNlD0RxvdZlbxONJVZ4Kc/i07Wf1Kdie8hwQ3ZTvokyEW5aM5ZAomSUCw
icnL7eNG7VEX8GZrAV89ZCdSvh5pTXWgNQ75EpFUuGydP/YFpOvgyWq4d1IlC0wRutAagJmWYGGN
7na8YK3mkCy8zfddBpWlqg6v2w7k3DzJmO94Lo20qUIerGP5vofRYw6iyf1ghKCgO7T4VpLhbD/+
NopTEoRd+MoD13gbjL2QbH9Y5cyFvZgBCz8iySDyxtMuf+xDJLsaxQxgrY8C1ZbOahtalAlhHwED
FvNQ8hrATm4eaDNl1/u7mobNOcU4AYD+80la3/1I3YLjnfQ08ezESajSQG1NmbP08k65y3nRaWfX
FlO9FhtC6uC8uDTHYp1KcymWkCB3RGE6OwJZiMfAV7IW2V3wthMEvnBdriKrBUVTew6Djjh7TT3Z
OVwzzevnrHDRGMnTMiXkYuGaKasB78hvxCKiIAmI6c89657tq4wNphYAE7IRGcn8AFR1dVwiaQtt
tQJL7OFad3YZSEvlM9h9ATRey8SwCr6AGLcSpEfIb9uqoRvo6H9j5381p625Iw80+kdswOqC1tYr
EjD8GVVDbY1pBrkAYTI5AhsSZYg+wqcrNXIBkupuYow/Py2Txbhow0hFsc9GMl42chLfOMSCM43d
U0eS+YVwZ77H28ptlFdW/e6euM7cAX36txL8NezvTDT6vitLfgpRk8RJRrECVDLULyAIrmEWwibE
FCg7203ZtWvNfUHTLDxxE9TiEQhyEO4RD+Q16ZDTR7HO0TES3vNPIVcORhwpYG5uyEBFf/GWa6yK
zYFD8bbslhc2QXtoKFdTghqsp6n1lEAaRGG08QoO6E4JQ4IjuP7IyFmKMR4txyuBVG4JHm5QNjn6
1p1RismnunAfNSwKpbtA1uC+H2YmViMEkikawhK/HSevaUpUs0Xp/hvEQGW7mzDZS2Avw6dCQ9Oz
RQ4h9kk8Pgp8DnKHKRWKKrCRhgP1sx0yy3X6LZHDSQYrv9pQ6w/4jowS65uH0aaRklenMbJYo3ww
CKieeY2XzCZHQKe9UnpbO0JuluD4aoFeBwNbrV/FlQHQ+Rk0gatOoTbGBzlQe4Hn7/t/PomLW69D
uN3Rl0tY6uuNZDAUrZx9qKPCurinsfxNYUdnnMHxoQCBlA+f5AQvuEDUd5mBKRz8eE4x3Gkpub84
rS1pNIvmFo+Pl+AGgEMAE5eqifetEoJAulLnEGpeVaupPLsDvDv9WiyJYZoRUJcxHKzGD6r12l4J
YFdYHlQuYOKumGfm4ct6YOfeR5bw3oukfSV1ldg4KFUyN1lcPpirv1maBKyMn4F+1HjI+YhLh0SR
Ktl+sm2GspCFz0IQzBHd3gwOM6OI3D6iAKfV+Eb4ElI4OK2v5D9scdKiWU6cTD1pjZdP3tjnO5Du
qxmRgAzGzv0SDswAe/VXA4lsGBmKZUI4L/Ylh27QAnCQXTBjA2jBRu47rKWwGEgI8jEM5+pwN/KZ
gdIZXxd4/kC9ht3PCBNxPyELpfWS2hy2FjeRTYyEZmWuqBXnGCX3zPv4UtUtbZZes6epmuD49SBk
jgY9dqgNWvgeejJJbdkwq/IKt0WCMC17y9M3vFVu97fOsAnm9XCgS8jjxnax+nBXuOt1aI0vXAmy
z9NAHyPt/5Caplp4VUN5YaIyXiyiLsA0OSWmsFKvVIShRYPNqtlJd+N4VFgTIiA9sD/Wcf4wI3eR
xj3A0ubSn/aapFntTYne794eDbiYk0aOZr8jrqVaksECXO0Ftvpn7WDXVUVfEKrtcesb6StChLmN
jUFg7Y4GajIRPY6cwW2mAWkA6FWnuwUTXYwLyCTA9sU+JBTncsE5DVr9Ewa1120b+MzKMYhBIpxw
HBY8scMUUIv9RNBrCBwUAxzAIli5+NrLGgyn8yfeUxNFdy0TtPmcArtnASr3up8sI+gSLJCDht+O
loUIHw+SLCbSVkmoxYlCunQoHBlyjY64Lknd2mlAyKoiLrEyz1gq9dBug1IfaF7l0Y3SIkCFX2gr
4lO1k2F5GbINE3k6+bUwBiSnaURxWSPdRfTpZ6YToSMd5L2Qa8WJb7PPsl879eK2q5RliBXxGvq7
Se7K3UI1ouHM6KTfJlYyI1XHFJEevV+vEdHoxy3aHwMpGtGyf8o7e0ZDGJEC3Nm683pL8RMrtaIO
ggBahxhKizAe550UyUJO8uTZX9Yg/LAwbjmqHCAMeR1KkkNH+NtG9Yu73eh4eL0X5g3t8+ebpOzt
AgyyQttFf7tFRMVtIHjYon0MxinQHQSjPiBWhg1xuOSjOYmPUgRJI0lF3HegxxdYaC3Zm0ejMhYI
DzSd9yt4kP68O0ZBKeAxBVLLIEL0gPNgDCmcrZFXUGRFmsXGCeDRSoMASiMEWuigByY9Cxy5ld90
tqDIStuqiHp5jncgEzFIsEIFam3DpLU1F8kT1OvP/GUomWHWXOhnHSdSdRfjKVBSYRbC9DdrN1bB
BWsc8K2PV8pYLjjHXzMfO3Lk2xIMxSfMm54RkaZdJI3+dXqQAjxtC9jXxfJTWkKU/xWq+QQkqzmm
Wwi0tutE4RNeJWndp7edEPMOZDCvijv1QiCQrHvGOq12gjYyOa9pYJCYKO9QJZNLSpBYTPA8wIRW
APtAb7rkmo3obfRXXq7ldEE0bhe7SPRJkEni0ilPjv46Y18ZJZWPN//qqg3i0Dc16cHnwFxHU8Wl
CMT728dkX2W7DUet/G0oDbbBIuSK7/WXQhgIxvp+oS25QFkdNOxfqFL/vfhlqOfOs1/ZH0id5bO/
H8FKBJL24NlcERt57b7dKPv7fC/vgTkOTj/D8/KfI7NPwzr9N6QTh1QSPyfjXH4SmR8MshCJsICL
sTALVeKBUGTxwZ4FFiPz6XL2QC4+B0GuaUouPTwwB1iTyXpf+eiB7x365MULRgqg7GmKT8JDQQh1
yn15JWTyGfXJhG5KFkCY4at19nZf471uJgY+cz+g3BXN9N2weJP2q+USq2/SsbTXnycx1OOaS4bV
y2gHQ33T6Ow1teZ57vJEa/ldAc1JG5ugiwURF3KK9RE508pjFszDA2YXouCOLc625l5x8WG/DXNR
kVHPrtUd5SOIj/qpIsUbzrcNFcqw13h+XIq+zQpUf5NjTQboh3mSHbxfKYcxr/apzAEkC0ZxoT5T
/0ma0K0w0ZVZ55dT5xN5HewiWYP7tKiVJTUA/OvT8ZfVAJ9EycFjFDgH8NHE2qALZe48Y3LRDK6S
kH9OzuQpxqOZ3L9cPIfkuScEETqWRtfItsnWdzei971MTyaJrm2E85a+wg0SriT3tXFccc5Qwyfj
07zgAkT40LCfWRbSibfku57+gALgrtb1YYB/tvkvCaQCzTpO2AhLqRhmJnBZCTYLwzOaPdK7LMQ1
DBUKD1Cw2vkYftJhup+MbmOCORqTfDQ+LKe4sxaW7MavPTsPnZvCCncuQGyO9Xa1OyPW38qk2oxD
BbzJldENI++CSw77zNySCMqg74o5JjSqULZ1unte7vQFBUNaNBW2A+doVpx0VCvhb5eBrA5t+R3A
EsBTi/Gk6YUwMCQFrruLGpN4gryfxXTrn9EG7L/lqMdEeAsvcImLpqNA3MqTvmXqWPnYoHfn8Wdr
ltOvVktZ8Iugd9mfd4q/1VXxnd0emxvT48EtQRI+L1rsLCtaz4LOxh3Gxm/QdgRh+ll06kbUJsA2
lo4SsPBozybSRO/ao+R/mbqu5zTh1au6uGtRdIlge21AGaFxw2ogwTVqJzYRaGodMP7Gx2ZIz8QF
K+U4sWu+e1TrmMIKrsKi05lHHcxv5Bp5mdSSzKNXqxlEna9t9sgON+j7Ulr/D0CDUzqIWnRqivxq
3iDDJtpTrjLGgEvWXEOrKzbwRRiLwM9wjlHjA7P27yNPl39drm1/HdIv3PeMG+2e5vFXRrB3DLlW
c6axN+tLZaD7fXi9DQx+n424Wl2K/bIzUC+TWFPZI8HyKsfuZLjBWEgvtL2QAimDI7LXpJZjRXcY
FMcAW4GpJUboTNXaKk3IF8WGnVC/iGK+vVZYtu8L0xPot4gF9c22KRJNU4dWUbBfk+WOwBrsZsLa
p+QoHmwRZy/OPOMps1xCIwgqJQPS/JBA9yoSVWARtn0JKh9fNFS7eheYI6lG1sc35KNcd3tfTRtS
q+2aH6cHkhyA7d0TY1YvtqAyL+sqjIhr+q+Dd2ophCo+ezAJ/VRktgpYjEZ5hbAWhJtcjNPN/Aop
ak5uGHA0hP784iduDojW6Zq+yWR8SMPDHvAB9anbWinn7Aum0Xj/a1B5h1ecUvYsnxZswSGCNgU8
cdMpESyuvecAVp6lcxekzJ+BkAMljjjCd7GX4nVumMuAXKOlx5fv1UQ0l2jGz7M80j3LbWowXzkP
47+Qw/jHpyB3h5q68mXJcQTlxGWllyCY4jncwoYgO/Rjb16q8YZy921e4UzYLGuR5Bdg10g4T73R
p+0unC2RQjHhQIityQFComDeLLC6kpn2fRtpNSQdDnTI84IUkaaDmG+9ix8bMXrNN8E2u1dXuWF2
jaZXi6D0XwohigPNiTGT97lNG4ir1zZ0+SngdAKQHI7Ex4x98/1zw9qCYvrH1HwAcPz9R7wgHPJ7
dlgsjUwKFZSB2n8NTVybP1UUvrbbnx2NlBuH6oyHh2luwjPQo4DWY9tOOSkAcVzo+6LYp6dBnv7g
BZ4sAzUYxKhgW05jNFgYasvQ1HL2Lc+APuEmKRam+ourqOczEvbSfOorVLzuVMREFtwdWk0hSbxr
w6Ae0DFmYIGUZBW/RLwrlfTiF6vs5fIKjYWnJQnjB/4ocEWrqEI2A+wOjUUDcflm8d1zcidX8VCr
wp8fRvdfbaMcMpCwzEOp7VKT0Xz1fvAh+JYKwiiJ+inXGxArDZ5YL7bid25KdkR1LR9RvXmB4U/Y
ZkGmboPG5krkz98rBV/EMAbNQqFg/2kBVdu8nBfFjlVHWxBzwCDjcRciIQLMkzjuwWyMGfkUTcgr
lshngfiS++ZUjqQbwZyIYEfECcdeNibf7o0kGUs40AyizQ8FTWlu0tVBeV2m3zaR3UszRTobD//z
HJgXVFhyuCRMhvDzwsmkqShPdc+m10xqwt+qTgco6UpmYkIp/+QHjeA26vJSgfzViYy7pqlKjWNI
5uEK6G/zDGajyYuT1IF+uH3oJ0+P1IbfkHEdqRRsBOnaF9L1ulEiT/w3XPQNdDbDoLN43msHn5Wa
ZU2LfPNgIjOyxDIt1E71btkGbT/QCDbmzSVcGImLN+T1o8aeR473K4wceregOZmcXb+3auHkpki7
ryKUPx6zvCBOQ03XHM6TOQq+Tzz0jsm19RGvTfM3DUakips17EIVmviuoy0HIDs28Q/binQUkOKR
tMyTUjz6PxD4TFK9GfsLH+TSszb6Ryf1wd5cdenPiiZmDhFXwUsWRcErk698tcj9SaWo/oua8IO1
c7Np87Ufp6n4xxdm1KZtZQ+wqgwXWU9y6say/fehzXKlXx0zv9EiAzo8J2TNK4Z7urHSEuE4Je4S
vIyCOiQOocIQRNjBg1A4BMr+zb0J/oNeWWbbUNmTTQ04tdkEgf4zJ6l/91Hu4zKb8z0v6p25vqZj
zgS4Zz09C247KsZQ4tOSDxUqMAMpdMTjC5XMVE8v/uPU/meqkrAxgdCixt67X23KHRoG7hqBWawu
JlFjmfvLM6213zBcB8XP3ZAA4eFc9KMG0EYGWrL8JRhaFn7yuC+75kwowjcEsCy+CDjrPeGQKIS2
SH6hZQCHQHV8pfyJNe9vL+T8/8D5EzoF+W4gNrkbbTiXWbi8l9QG4RP/LUhzaLY7DYyNA2l3Lpjb
t8Zfr1Pn2/slZq49Ezj0H/wLfcskJ2o17IO+RwmwpU0pYv/iZOCITYDQ8VP5ng+5henfe+oENQub
j9Y9nSZbtrY0zSdgyfK/CJYx9Ubq+X+1sIsv2VR8TiQiPgPm8l0Go3hfMohsL5LDL+w1IvDp8vO0
GZgKu52zN+XlhFtEdhDb+4kPMpn46dIInTVDogAYiGJrQiGgrIFxTPtXmDeIoNMSva/ag+++cYbP
5ldOGSXYLuIxaXlADam7Wj5zVCHd2b0m3Ku4snm8HEb8LLWmF08Ny3nfl5HNsya47pNtLOLEOvYZ
Dx7sVDZ+UdA+aFDnUjKf3rQI2ZNAXkKGbf1Ckr633yWW1ilzhz23l/cThHHJgwgS/+8GEmoZys0o
7TSzC8xxux0bF7KKVMhg48Vys5f4GByplcsIEaNyw9OUbTmMcdeaSHFBban9XJuKLmbmeJlLFlu7
vaM2obbhzmGUU4LdtioR7S6hqcwfehOvVlRnZbaCaawcy401Tk0V2pNYG/kF6h7GIAynlfyWxkOC
4cC5NOO+LodpapqkZRftgFpRPR8FfTSCDXW2laOlimxhM1R9uDRQmJzqmdaNexTBAyH1oVlw1kdG
VtFhhvisLYbaKO4Rfh5wqDUoDjJKFhCRMSTHqb7qN4OtYzpuRKVuz5ibUDVKmVJshhqYEDmcg8/J
d/o2d6kd5WgKbLd6YoQOEeiMfFA9GTXt3mVvxvbFrQB61I2TDffnpu9mmRWUmyznk+QMgkJYotG/
EtvLmg9LgwJ64ABdw5eu0aKMKZz+dL44JC4sLh5bwZNghiIst0b85zcDxim6kai52bCTLqNDKzB7
ohmX+fzHhiO8twyPY61hXnKocho9RkkCay1K7slBfhzxHZpRe2MLGnlI2nNiYj97h14/GKMMq0as
QFhZ1p8qW2CSkYGlFc/olSZqyDqhETh2TdiOPxX5ssng+b2akALM2zNjPA5yvEkrWwBRCkBnNCUz
3saIClC9xvDwIqmbarn4FviRalnKI9IIvfWRajR/t28/0Kbt6QeQ7EO18qerLXgN3Upq00ehysRt
FVhFsgKARphRMeJbePDdWLDm1aBXKVUU/Z/arcxEY5wrIHamJjnUni8pTa8cAJQzPC170Wy8gsD9
Os7cLipAQSv6DoKR0r/+U+aHeH2ym1SrF8ZzFOYUI4vmwSYCiN+dlf5mQcXCdUsAokNSgKi6IlGe
L7yviXtKZqu3RmRCtox48Fg1/kqcZ7I/0CiIHWAptlh6IfgyJehP/d6CmrlMcV6pBtPiO0cw5noE
WuGVP9kMpPozylm16pTUx5MZ5RuYj/NsMEtA4ORx4B7xN4P9SBPDVFOCxoDmehXmiynC8wQul4uD
QVSWPIB3KaRvNKJO+RE7Ep5oSaSJ7/hvXzEaL5IFSagb5NcMzkEdjjKm+NjAG9o8WbgBgAzKmjaf
tae6TSqp1jjiZOY1YRlK6bzX+f5K6v39+O7Twa90r36AjWnQzXRlTsCF8x1wlrxEvF29Sm2l71la
rKr/e15YgRZV+vSW1iR5vEs+GsP0zF5gDCVuCzLfy5bDMBAE0+5N2CYyRe8LJdqTgpvJHTzqDExw
tkM7o/f5nNEGuXt2tQSwolNnyj3ekaENVP03YUYrIcvKrqLCZNUg9U0t3EK+k6h+wo6HXEL3O2Hs
5ZzYF+C1ariRT5THwDOP49aCMry201oqITz4vwjCK3qSbiHP/ZJnH23/vR1zpGryt2TENasajhRp
TsvrwUmj413z4zwa4PcP6BXUNh5jYCyNo7Y0xaxkNzZ8vW0wEzPsX0sF7tYL8yEMtUGhRuOKSjlO
9vy7Z0OZtlp+6qRmSISpIn6tNaFEnMN4p4TWHFS81yiL87UiAOPoJaHEYq5kAK69wKTiyBJbVlu+
BvoWPTX/Pjfxzx8e4vCVyDi5f/3v8DwWAGnghdcEPZknMZuwy2vWniPVoN9wdp2zUHrjaVxf/KGN
Cqt5LyeN5dJbsyXkgJd61XNfUy/yO94ON53eUVd2hmNKWYzuAb3RCVtizHAp/nd1aIuUbn4iHS2J
jYqwEYbOe96gYm4HenGxHBP8kD6lbw0B4Z6EBg9WIiwPobNQ6XylModIV4aTgFaDjXwbGfrGAind
DLk3vCsZ3azsWpGPftgXxXsaov7IahWB9mZy9yOFVwTHDBQu7F0ebkhgYr7qiK16bQO90nvuo6ch
4j8OJM+tXhpDqXXJ/kdXhyUm+Jjx6mqhWhcykvxpo5DoD2Dyfn0FjEuRhpHZ+YEU0WfRemfVwfyX
tXNbxvqcVcNSqHfaJ0V2BJJhHvdsAAW1KT2YdBvT5O0wY1qeaFlQ5jzFG4OnCbb/GnrCvP8GBvz4
51bepxbd9/eTjWe0vLffntHcNoVpEuybOVPzZpSuNRPTjiMNkszarAmtWrz46ZP1WFrCU1wjuwNV
PZhA5+NLJ/yhgIfDYTNZMb0/MKYQR0JXWprAuAO3YO6NKHzMi3SG4Yk3mXDUic1aeSeAl6F+xl+a
FkJoCWlJo8WkxKBjAWhqlKBoLhLLKWvTOrQ4BAJsCnJRgqLlvbCYo+c5swmhVk7VI1mElTmg1Ydr
rmZgsxXgdpXic9pConH12K7BxKpgRZOUu4wEZc4wgxWcwD2DZEeXuuO+fxGFqybCLdjvqPtA1Wk1
YppexO6R7dXYl6F1bqzCZ1rDMgXjrvUxikj9uTuuGuP82bw4Ev10JWvxLR3RZGU6wM3Y6lOtK+85
MtMQkII8WHqDVXVENVTbvZr/p4vYe/z4YufGVDRSuK/LyFn9hPqGGolvJkYY88OLyTxFJDF4orou
aqGmij30iOmbUv7sTZKKus0EmfQD0i0mXjqb1sIFuE3O/icgCDmC5BP1i+2+AOFsJCKD9dIUDdu6
io1ZhBTGDlNnzNn+6IFDE3bZOtiGzCFqmYRiyxbEj5L3KVF2n3M1kun/WYjLoaZmRgAaqAT37n4l
GRo87zHEVXohxm2vWc6TTQV6TD9jgKzxdp4JUpYtmIKiggci5xPEUnwSWpM9KbMau9hy+guYSpRJ
L0BHkrTymvxmb8c/NI3UC5Gdj/KxF2pc/a3BA1AzyavKfQRtXvMO0sXEl1/mCy+kuMx5OIYTC+8f
kb/9xYpQPCXUJyaPxlxDCx0R0tbppUG9vRJm3CgyfUEMxU+tOprQL410anFTg9a6TkchYzZn25gl
pn3pwC5WBPLHt9EuHIiWrH6/Kd270YNEGc9Ye4rwyzL7R/hrZVJBRUfsDkRQ6qGf4NkjZk/EvCww
UcT5KJOuwYmBhkzKxIrCSrC0qqvCMnms/jLtPVJ/D+6acWYZFHi7fAyqD1rUB/AihEhmFDb5Qtvd
5ay7t4aGAPgJ0XDLKN8XopCckbLMQf5dIpUPzmdxOy/iEM1TcSWOUzfdiRFuPuFQZSbm1vBgMbMI
2MzQwrDA4yaJ2rTjpSZoe82YUEPfXIdPSh9ofxY9hGbXLFdUCmiC8pbIsAMtf8WpyyYwyiOhYJW0
vcNkkWQ/O9MmxTM5o77Wu5AfiJom6JgPHPMJKHffs67tadE/L0y3FunDyObY8docsfUH55EuUhWk
GrRUdiW4pyinbJcJ5UzOXJJP/wMFP9l6yKRnQvYwnrZkWHwLrEi+n/qSVOSMYP6y+nkrphO+6cJO
KF8keUIBy6P5uLLh5QXvOAc7xDkAkfJbv5GIceDlf23NlVLe5HZYNRBVi5SSsGW818a4LIyywFOd
6mfZsJ6K+lrN911CocaL5M2CFKN/TBlvuYIvB2kZY69PR/7yHdtA5+Pyia/RCkvXSL9F/ni428Kw
EsDEkF55RSbItgfHE53yM6f8zS6m2TnBdvrQ4Y9+c7CExFLaNmfQgD0LF9sMTgY5gqJtj0n0fYIf
zotXtkmlca6PtHHCZRbbb4jgJd9di7Wixehw500afmfH0YsZwXVONsostOD/umejCOWaz6m9cCqy
gQufTBGWsw9szdKLdai7Fob0tjalkR+A4ntJppaGKMvWLDvJWxuchfi6XrtnLel4hR866P5ihJ+8
5wWDm4+ZKvYhxrZZDa9OUXjUesE33nu3XeULKTVpT3HwAD/RGH6SQUPoX2sWQtROylem8GtlNeCx
Lf5YHH0kAbpbieqx7oOZD1UsNL8Kgz9UuKPFrPujjvcA8b1dXThwFEOO0kfnMqwbeipoyqtYI3Y0
fod5iATAbKQvurGehRbFlxB1iqSTekvgl94eO7iYLZzHuYJvKuw2f8MltdKDW0gnSUTzC4/+2NQl
mvY+4rAcZnXj/AVAVUmsgkYbYwoHOaFw4tNaMfn8Ssgow/pkjWvkmWtQ9mCOz0XgxN/FAu7Sp2W+
nnwajfGMidMMNsHkJESMK48tygiaRYkcahke1MjajS3AncmGzus8x+Q3rJ2DGoob+i2RNcZm0AL/
cUcVJxrNezQRZuYf8PuUORijzI71JRaSsYwhpwelXeFnnIB1CiSKcosHuy/j+EmOEOhoqw2YwrtX
wVdAilbUhwYeVJ3DGJ7Zif+ws6B2xRSGTjU340IrMG5muiH2cLyqn4XZeiW+rttBiLO3d7D2p5Ld
nQRViNGATuby0arDT7zvSkSmYpr0axbHR8gvU7JFIZquWh2WMLkSKRZKm/PEvs+1BwVFTQDQTX0q
1UG3jSvWlyGyA0LYDgYcDAyyOd3Pi3Ac4fCrfR8opuuZQ0qijxqA6NXS2Gnn9erEDVVmq2/rMTPg
MlXKo+Vqi/ji+xRWBpzBpFhdrPKYyS5/52oeafai1apErGozY9LcjmKiq2H8Ffn9vdDWsiOdhC//
OETUUhtIq0tGfGggFP3si+rX03jqVui+oiwW28ofisv2QXlfoGVV5QN/2mueQT+FDAD56p029rgh
AK5NFnhaFmCYOKAVOdLi05ieOPVzQJpJhGAys6Xg3HYFG4g6iKjSv/6SlFgLH5xskjsCa1jPFyY+
IC/1NI6597hGJdKT1fwikwnCjNfe16JIIjRDCMZUgIxFumFcjltIi0pHZhfutpYy+8xoYdRzVQgs
v1tq46UxozNvrHeUxl6GMszCcF+BcvGOMn4dlmY+6bBbyPPa9de1LFdbtVfOCuMJvO87YIvcwneC
FwtoTZoZWTYOAk2gczm+884/Fw7mVi9eFfw/I56eYPgYnb6U7BY3pNcph6s+4ayZGLQX2jB4xKTT
y3+lrwCF+N+UXQLmCUDsEO6K/W6tr91vUdK0GSOUB/nARhqDoNjQDYnmbqZ7Tbh52/TnCYiIhN/J
2KMu8NQqsdc9+wpZvbFxfrgvl+qAIHSiRzeHenVX1DNkbE7r/wWfmkyflW9QwjrDDB64jBgUQyX0
5m4QK47WAy5tqhuaz87Kq827oJdo7hlSSJqF2Mt+lNBmh45fOdQD7jxcMvlzimPgGlikVyGOyMVa
qECya+JsJZC9MYULPIHAndlN2RgvzucJFGwgLYnM3l7ugMcoOrBxFVMI9hhr76+cjgadKifHHsKN
GOXmW32u9xXgoYR7VnmYvg9s4G63DJ/U+QtcNPaUf7/oYiShVSq0asHk6l4T0Sgdga6oypc9Z/8z
FR98sS8SX7dfqrxq6FL5K7mhhNqiyHdkiY51Ms92Mdd4CPBN20KjKRIixhVZQz/9sFU78qwFYHVQ
itoJvAZDK6hnLq1PZE8OqXs9EsDGk4V566eoaoHHJwvRFrlgZnG5dNbEj0N66BlquYBDSQgkBYTW
GY+ktT8hCsGLiG1K/bzAePFCwA3BnfNgloI5mMYERRfF+CSqx4k/F1TqUa+QD4DscKoYs5GDrsiI
dOwlbY7uyskKbDHPle+O4obYmMubD0D9rwSrJkjfFsMRIurumyq0bh8uRidAsHDlMx85dEqUwj+E
o9Qrp1znivbptMyJObk99Z4zQArp9q2khe4Rc+ASwJtmdOgo8v9Pbzz+kMZCAZKRNtVUBkInF0F5
OGv6Q8jqopkixy1zmaFF88gprRrWQIfRMwqi6s4WCiJwBJf1IAp2m9QmGcIh+oYsjXAR8dMZzYM6
CHDeCEor33fzAq/2BWWhu6qduX1DyWjbEBeCQ+WdHU8q76p/xg6965AYYPQmg4wWDetx3lKKO5ZK
8Glyfh8KRYy4ONryR+WG32aIuSBBKHnJJHyZth/yv9dlEEoLA/y+p59MG/ZArgiW3lbvKi/pNR8k
8HTGoZypx0roHvGTbiLj7Z4fxlfF6EBXJT/ZWNtv5r6Kwi8SeUhw2QXd1Fkkky88M0bL3ztvVwIB
jYPQkwJ4zOl0grpN5VyfLgZJ4MueXDHusu72Z1aoP1XeRTOb2T2JcB/doaKzMWEaoL34KjJNtcz1
3eAX80qzjRfhK+R9o9HzwqGLPnesU0W0INwxIEhOwz4qUR7M93s+qMyPVfz8BPEXE6WqVRZoqute
v/jnLXPWhKcedhT/xFj+YjYjOlOGJHRYK/xlwnEljzgIFScB+GDCtKggid73fKbqm5/1m44Q7GXh
5oJzPbKCyfXFEGb/rX4RaUKFEenLwN+zltAaaC/sxBlYYzD6ZCiWfQtQXr9EVr5ku++equMqILy3
e+aXzbtOXgRTKKyjqw8WKgibqB9ZfGRk0QtmIVb1TEGMjND0a5I9alvuDcYmoi3rFFIkGu8cS1MY
KEIIk4DkGmU9EPnh5qJZaTTQWCrhZ7r0p9j/6vWgs1329dO1wsyer1RpxfV/a9Y/FOqkrGeUhIox
3qMWvbygkKDUfsIP4P5ZjpSlTeNQMTY/GEzvlU9AZFdL5bu5R8e1QE7GFOjZDWjfxruFZpqKXLxg
/tCH9nAlAIBgV74s7s51kO2pViTjahYRXuKHDS76/0L9umo/fghCLS9V4+LzKg/eEpcQkuIfd8M5
fJEiJhfOgoi+ucTytDBN1sw9QP6zmVYVBr+7aZDjlPv3GcBH/sAniI2T2sQtcUD6bj0T/to+fH1z
xfSq0BI1RaJpVRbsQs4xMx12C83lM5xF1+B69uM40Go5i/DFGTMH9nt5wlSurycPbpR7vWluUrZq
k+lywYZe3MFZL1LAVJrL5l6nRTQ4sJrfbQk8/yDvfQuWbFcKp9wo/nO/tHNXQwvEiT9kcuUfF6Wy
Vwhfh/oWamMR3YOdD7mtuIL+ZuGOKMo/UzRZqNgz4eqHw5jCTxHj/uGQ1l4EcgDjQauM00d21xny
EofFAN4BTzAoXOJDjLxwb0dfkitpFhopH8Pk02yoloL8klR3RmuUJ3GGsWGRGxvT3yr+wT9nRZck
4fB3usxX6izCc1FLIyspvgH+nTIUDT3xuKa82V5qU3AnciLeo9TdwFi/e7QZFZSjhe/ERtzJMMFI
aPc2P+sJ+v9paz26oahIo1B+fNe2eDRPKXqX9oO9+40UevWtOqSVDms3Y6KjqXECYFVTncMRSmSi
ODSQXftSv7JOaFBMMR9I9pTdhclwuA3rOUT3E5otBZ08C+hGbPe0qctP/f3mAr7XW0bNMKpC2QRI
8xQjq0599fcE3m6mrnFlVhIBRt2WJD2Q5K6qYV0BUvnOyj9zWQ9rceGlts4StQMhWvsGCNe+Z6cY
aGR0KkImq2Jm2RwhX2oP6+YWlLS2fEow50uCzY+WIM1mL5BVpq5ODJfx6W/keC9Ela8W0130VJiQ
87tHOpJB6UdN0rMM5bElIGDNQJ7RNlhpP6P7qyNBOS4DM3IrKzDfpcX5jDWZKJdciltXHJXfox7i
6OgfFP7KTM1f0d6lLKr6+J9+IBAs8+M7Ss9rDKSn/ouxeO3GaM3xDcPR7jCFPVlLTIpuNDjJMEiE
xYFHFubuAi0yktHDHFbRMJvMKAJFn7/z4GwWPipZqYj28deepeJLSuZgXNq2a77/v2z2gAzi1qo4
7kcIaOOTH9I/83k2GJMQzvfOT2juvlZfXAeKfPxbPN1lYclGtQipHxRLrb5e18fJYT7SCx+U4onb
tuRKOPVoL7kWOEyYWIufXf76Dcwm0Q9ZzIxNeoloKa8NTSe/2xfQ1awPLYqC8k6sJGXQ8ArblklN
DZP1VnZAUWPGxVVmhXFh+gze8RorBVXU7k6PtppFPOldXW1oGi7JVRmcBeNflu3ydp+YasVq5gWz
RNUL2cFLD0lMVfDUnv6mZaqReXzGYnrWOmnmtcy3beo2JCkgxd2AeKqBmdUUMuw6Fxo+06vepwvP
/ryAuvr9Mk1cMPsXeoGb+1LbALIa8qioqPBc8HDth5EFGnD11DALblbMIiTYmfVrkfutf4yXuat2
BdZkxKTEtxoZjOlYL0CSXBOGZxx29zP/Nw49k4tBl9u33F9LXPQxQFoR2JlyBTZidjPq3EsV8oSW
y9klO6xjr/OgrKnyFYPAGs4hiTiyQQ3Z8I2xtC5XAPzlEAS/axpbg8dAwoIUdDRjlJf4BfCWFpT8
NQcCEO/rsc1dsP1/RQqZaY+SXoAzoVKFibGdGcXzrarFsTBVMDAkMShOHmKjJCpr08BYrPt8oPd2
fkQrl7BLiImP1axakRvzqcGB0KNLVksS6Jxlxg2pMffXrZacouqrfjG4O+nkUskaLaE65pH+YbRQ
T6UwYdkdSbiTmS8fNWCxcrp43F9KvSNb5rtwNaYX1hXzNvUr1UEsbEmni9g4q1bmnEZ8R4IR9gJJ
ayVM0WZsyBDWUxDtTcCSYdCOV+9CVyRC5drTplw4tQlN0/ak+esRcRYew2ZTtg4qb1N5+St5p3+O
LFvxE+klNAsLRRMPOm27vn6evGKjTFJFq53gvjD9M2bOA/+cMGXdOpxt6wJaBlPxH3ShGhfd3duc
MCIS5PXQfuq9mlkj5xk4fZ6B7r00JJyaDsSy7wzJ93DSWv5NVagRDYVj/igJmoFM+X5Tc3Q/5r/E
OmataMfkc/U2Emqkd9hu37uJJVKU6+mWTmbe1QUVVgwTvXLMxWx3xY0f3MSvw9f7jcmAu2ymMxRW
a+J1SyD1im1Z+/KLZjZTXTVuJrwBsOFXxYU37o+2+N0l6CRgAVdexPbGOPIUcnDztIRuz9va3XRB
Dt54SnThb4e/Hx87kofk5HndD+DuwBuCS3SsOEt0xY/M6htoen0SK+ZKMPYg8FmTdQUn12w1izJu
Lzwn809Ngi7DcGnZheuadwbncPddTu9/270XuQLmyp2hUXuRxg7D+lMh3mkHQEKao0czRKyg6dZH
+kGgmeWMVdRXc3XesE8W5Ivkgx9X8CK8+AraIBN5fnAaAp2r/ltALjC8GRGYkiA9lFpN2PR1/LTh
BClq3jL85GWlD/EhNc59YUD4lEyLEuzOfixjEsJxRpfN8flpFvY4qLXNscU8tnglWSTi9ML6VK23
AMq3h0UiKtQv/8KxpdMXuFZjaRkWd3uKtkWzMdII4Hd1FVypH5Kym0wW3OV8TdUw2nidDFHsxCuA
mVlDwunuJ6B90olEPNxZYMe+LM9U7WJWFYSYt8BiIuQ744BQ8oYFYVHUN8u43vC8FPpBE52ttpne
gydU+dHkg+u9s0pLNIo2q/PZTaniLD9/3pIfP1NupmVIXWUrOyWtJ2Dx7kTzuPiUKYutoUiAwrin
VO/3fTYNHRfU8Y1WhgKz65niOhgarwdEng0JtX+5IMU/o9WTlRlEFCkffAUrJ4dRPd7Zp1VT0XjZ
mbJoqfW3xgBaUYLc1806stFaoaxVULiLGYCQneuONGgCwKJCeWnPiSpK7IX5dzeiUOyG/slJ6mC5
7URIjRZANoJvle/5aGkyTaLKYT+FgnhgzCo0YVzXyisntq1Ynql3NlCSwGK4y/OfPF7vhNTibLSg
xtoJQYqYTgl47tSFdT0PqcF5o44r+5Tlaxy8lm8LtuUWhZ7Ry+2BsDM/99WRXcByf3gqcHZ/m/OI
xQprf6osu/DEFWvnhhFwROnvZqvN/rLzF0omp9GiLo4Z/IhqaulcaXdyqOLIxOVzlZ5WQyWkpEhY
q4T6O/8E7Rk4IXZCNTdHztcUuUK5AK46cPQR+RP6UEht2JsEZ+Th7nnCL9qAPsLVTPr/n9iWCffX
3dKdsw1izHunaj5qRW45UbllnE/07ofaBCKnR5blfxl/hCJP4L+ijCBuv1xX7LoyvbxLult7xhnS
m+/q2r6jDXnyTaFnLmizAaRsX17bKSapBNtmT8qXgAiElsxPevZEzYmvwjDUvGVYngswgl7qTu2+
kToECdCwQj8nFHV4O0tbak6mXJX213RAMJOV+nEj4CesrWu4oojrX/0lchH0JEVX3LwrFaMmgDlM
hnuw3A+8lnCf6TmnxYUp73Dp2W7QzlcXs1P34PnyLjx4y8hY86jMcAYmbgZiM/pCqq+M3Bvgr6rv
P3K65wd7r9I/laCS5YfX0MywdgQpaMB5yciD8nGOO7IeM6C2f9mEc2N8YXBlJiFJoWbbV4N44HIC
dZP1DgLUpbfesH45RdYm8NhtnrUbSirrkleZXnS24P0tjeAYl+jMyNMZRKYCDNZnw1Tu/nl+yR8w
3ALMmDmMakCx0bttK0Tfy4UYqALfjQGUN7LqAubD+grJEMzLnJdqrbVHNnTRrdoFFSG4X+DKA8Vk
N1q8XZCaIexszZAn2R1HUce4CglIjhhFQKdtgD51Dc5Y7kD793CQ8FcC79rWdNBGMutyHYk6QagH
kcSiXMJfyexGHaNrLbM2O1Y07uNyDNNKgZZfIVS7TFYJIrW5mQvRHc7xsD6KGUQBLRHEOqjJBEzu
V2E/nv6bBNMt4M9UcGErsJdrbwSThS8TOIkNTN0AqP53yEzXH5kKR06tSy1yQN3RkyFvINqzwtaW
35t27zIhWfTAldKiXXWevc49SrAm/1NfBdraQ9UAU2SJE2Q7JzOSjL7UdAxJgCKiD+HMYvpWk1VT
N3j/cLxhig/6Q3WVRzYg2TABq4O3msKxAvEao0m5v+Ml3jb/QYo49FUiUCfuzIhLZD8bfSGU8/p5
GlxGqKAbzlV/TAyxZF9vkLk/uyp6KQ2e1kP5yDYCxS47wgD3M2LXuJ889ROLXuWK24lYOji2kTpj
cBBhdQ9gGGqqOFmwy/oV3pmsDnh6/mx6lJHDGomozdVNeUcJ40pCSQWGuHEYo3zZRZdnGdP7z2t1
VpmuPZKe3I7P+jxhYy1kxtnX08Msgvh09z97F8MzavVcLlERKxXKj6HPMQXcLMHe/SngKQDRuBGM
Y6jPAaYBT1SOicaTa2mm2oBmz2nvfktPREfmDTqL9enG/pfrij8AUAAsx+gAmKzfWWVIP/tAKbx0
EoE/cSQ3Z4ee0YfGqqxPhWzguvae8b43sHOBCZT+SerTuWWjL9H6FZIbj/1K0MeEjFXye9kCXlxP
mmowCb/+BjIVLqv6wQwCr4KUmni2dscM2ueua+UzHNLAc/KiedwaLdZecHmrkPqqv7nHwxxTRjl4
+QTt2c3S1eK6jsxuEa8npAwzZILA/Uikbg/42q2uk/OZISQw4r2U+eUYqQHnK1ijheMMEhs39+eP
jqbrIrEEBrjrevONSTv4jgSK8KI9iBLcjeJV/FVstYAn6RbqOjSfBzEZDW0WDUQtwwL6dqtxIwJW
VwRNED1xV+3lchiqKnQZqN7JT/WiEStrw+xMML+Vw5cxB+tV3s2q6MxXNpzM7p50VAD0Wj231xCn
Y2kbXEY7E5LjwyvnRcxzXBEkPPaQPiDq7asMKUzGnn+tEY+NYwfI3dd7DfmuB1IUTwH6IT0+RR0A
n00nqqN2WSPFyNUB/VgW+b3j+e5sDXFWfDEiC5b/HJ4IM5GvpkIDuERswoinEt40Vsw+gwdJXENh
63COMffxTjcuUSuiY7Z3I7+yX4bwAaSEiv3soH12tHqemPk5RLPRHTV1uzQYeloiwoObEjjzRPPs
HoiP1MaQV6CTuVFAcA1UoRedFnwkDJzWQp06uxfjBfgpApcoON8TdP3v4uZBUuJRrp7RqrBUd5ga
7YQFLS9HKPr85II8A3UOzKrJV9d/BbfsK1/pBeHoG/HW+Gca/xt16uug5F8CDKp/Dk8uzevGzpTU
4NXs62KTcwS49P+r4KNbN8Pa19MvxIE9NkJWrcn61rvWK9qlBZXwlP7ukbX9glQ13qlML8GraTkS
SOtbsyCMCmN9wb6yfQ85PR5R5q3x84eRhPCm7uEkSad731q+7qpmVrYE8iPbJ0x+tU8cZE2pLuo0
K3oYg8Eufuj6Q0iupX2ZliAAOLVbhsj4O+JIF6wF6LI9gyTaQExPsTJGACdIkxp2B2J+6+I7lOT5
9L/7jBygm4QzFCgEywx4SAzcnWxgt7oqrRythr1NkzMy/O66qYyRAwDk45zfZDNl7HCVI3Nlkl4Z
pV7OF4qPnF0750qAFteZ/awklahXMtLzifoHz47NFJCZzVKwxG/B0e4JG0d442slpeIGPsALfMJJ
/5Ytunc/Qgsu+GC80UlfJ6NJ5PXKwcqRc+buTZ4AwwmPB6jA5A6XzlBWOTwdBXtwGWWZxY7icgVR
GR3KjUpSC0FHdoyuxp14x8YZG+T2E4XSExESM3cQ5LWRcwdMMFA9OFLkcHonKHAGrLlKd04XF9NA
khE+LdpxZMSLNpyw5Mt672iYFtjFF8xR35hqkPsh92kFn8NkbdDdACEg44UvMq3HmmWdv2szR8Nn
YhBN3SpTaXxFpCRN0GnA8SYCRqJlEaBjKDLgjCNUcy6rCZKYd4J9lx8/odGcmlQDlrm2qPtC6ffO
Pkk1Wa2IDJSJBGdPQvJEiiZPyeG4+yRvXGHPYPsMv4Pnxmn5nuGbYFkk0vPQl+Ep/Gu7z3j7KPgE
x6B4z9MvUCbQ5Rmq6Ue6iQOsdYnGEX1eo1fKrMWU+vRvOzIW0EZLo1v6vIWXfN/pNUxhrjBx59lh
L3byYoCPgCecblIW0aHaUm+uQZOwdUgRQ4CWp22oXARAfYACL6xFl9kVsZX6lwsj+2EgAeaLdLYg
3u5F1H/mlwbXWhH+0PHYS9/O8SumSaEBpyLr0w0Bu6FKDY1hUNe7RbOWuKBO08njWb+XB3KOuGOp
cWaLoLD5q+s4mELSc+8+NY/651pb9irsjyOrLrsBf28csKh5aId1Aqov29mdpOv5teTCf8z70Mpp
LpbNraTijjm5SU0/8HAxF91ZZaCkzIFe+BJ4cY/yJb8zGIfbahqsARXqaGCh+6cIp2us7r1vtumz
ByoOx+m3R8FuYNHH63KwL7QSI8fsGyyX43REN2iDx4IH6qZiqSDC1ouADTx3VczYI6qp7C68nAwP
ELNwxkLbVhVg0u3zrqHGLCT9QeTxVUjz2q3YIr55xdY//aqS3VERlMq/Dr1nOE9i6IPL1W0V7ACA
zaKwq+TpPSbNlWlIvv97u3sT3BJwUtv1CfFYjomnAa4fHNxW1vKSDy6QnwNehg2x9pAFPyan4w9I
V+LC2Q5Xs5n7QHLD2zsh64l83ucVmfthSGNwMUAtYL5e/wttIbNIsXSeHSaFZC4H+odyA24DapFb
Vw9oMCbo7+QCAd3Dg/X4sLLGdWNNzTuBq4/13ebCf5N4rFSvA8ii4KLN+5pOKZpCF+W+zVlI2g9O
V3y1sxpYhFCyQIG76Vr5Cf2BpQteIHgHz9nVJXsh6JGsLYU2YQKk/MWAueeKKl7LdaVuVX2fezOI
+NOqHl1yLI04Cd4DCj6ietKt3Z7qctTWWPB7hz6XAslR6QUDg5Oy+IGKKtb60+/9V0Ufm3cMIzzY
gyRcU7ni6PU18TDT6qOx+yh7sDGoUbEhs3E1QMIpA3jOcIJnFaM5vOS0ew85uDyotH9kLHKirHjy
cbED6aoKoURIWLityb7bfiA/AKrBiKn6TLsn6ZVk41kFcxt/ziO407562dbsdYsrKcv2DSDzrwl2
Qma9ZIkfkhwEvxtTh3qY+hchgUQQnGjRY0Z1ADiiPQpgOZXPHh2SGuXAnesQKE95E0glPXFwKAZJ
VOprv5zpxANJyPzfo04KvlFVcW7KhFWwypEruvlqU1fm8t8pCD+2tG2IXQ1IF4lWUtg2NHlgiYR6
USxy8lC57C7WhIIt5ArKTcF8Q9T/KE+k+6WhB+wveflKGyosPsjnhm8JaqnTUN+k4AmTKtDpuzEU
yKGUw+iuvur8YPiAjwuSKeAKe5qwE2E1OfWAguOYqbyUEjQsUhxdCXCi9tAEIgwmVIsPvtSZtAip
AGRT9/4fVRnA08h2J9ZJwtIrbtKruPc+JrEe8r/+lZ4yMeCAUE/kh1UULsGjPGXCtXfdFGc2MRjI
Zt5jEv+ienKRGTvM1VzIiIB51EBVA08rtitHrFdjA3Ia8s7NRIfj6uKpr/+rz9EhhV9OQkgtWEr9
iYFGvprXW45Pm3tgpcwbKn6CAV8P9Y/HQG5tQ0n5X4d8A6fO0YRB7oiwWVSMkYWfNSQcdH6jykvU
0agUBt3CVczHuHRSKfrbwpQuwlvjiOx6locQXniM77EmrUN2mY95RDWsEG0UX6Y/fSPVIo52bEki
BbZYB4uEu4XDOt3BwNI/glrvtYag+J3L/+HwG3vlVWYYJUNkcliX/PXwxlePpGSCw1uvloq5IqIC
QDKBSntyUpYX7WZE6aP23Q8DFIROYfSAOteyK9S/626NPXxvP3KMRtg5zoImaKxR4qIQt3IfwS4n
cAkvlB9Y2FZ0Zh5ajMffDSLlwy5D3t0fOITOoe6F3lFMZJsG/1AM/H+dh6YnvF/+7pUzgPCj2JxJ
7fe7C6Nao6BdrlLaOc4d4rx1T7y93eltx83+WoqYputaBqzRYNoavlRhixuh43VKeYIZC4PZagie
mJIw/SNzG9tqNAB013QV7alMArc6aib2ZR8C2ZFlm67ZUy/td0FnaOF3osWEWO4d+ZtUohyGDJN7
jjhPbNabNW90orki0ynL7x6GzoS1Qb0ec1upyeCivZnvRma1AwyBVxoGrg8tKiSMT0Dt+nzX6EDe
uHiru04uIXUyhCyFwvTjDi5yvybXx6fB/cQSb/SOw4me9+gn3pS5hN6XS8JlPF2gw35LVsYlj86f
JgP3tPYQfAnQ3rl5J7C69pJSKcufT78A+pP/QWDCtTpsfbDs7/7J2CV5Al/4/l30a9+Sh1DHVVBQ
a27DAbNcPpz1ilEbZ4CngPnKff5vhVZNjtG6v3Mf9CabVweCEaDbml/dT2tpucLqFCJbRP9976VM
71yXrJqliaSfO8ejDLAyghnOlYpg57goZ3fVeZhP0Pv5Xmx0SQdtsa9rjyRgycb5nHtifWy5yuPA
NfCOynYr0OhG2U74EUln1x7AWJvwGoZcgB1Wyw0PnbaXYuiJ72FT8ggkCnCWMMrJZH9xbHxltmvS
Up3xxWtP/2/Z0h9aUXy5S9YDoN1qgQ2SCXBVrbl8lFgsS8kVpGjYW6Ib+nDmlca5g0IZxEIUcVHW
s5lWARt7E5DRJxPA/c8UEf66lNMOT0IyaOFxUB9fztDtIAEaUxBtHrUBZTFAKRHloXHzjdPNmTBU
LSwTF+1RFsVQs5P38y92hcpqq96xmnDttPY7euAlGQX90xviLVT/NysPLWSa1Z6NJigHpkLd4JFZ
1X0AwsiT79D6sZTVF8xs516Ee31U40bhvSYVjSNtNXaBXll5ucprJNo9oUIBh/Z3FO6rWYA5Oj4U
T315QCsU2YSCtYnY6pd+tEe3tZnD00jD51bq6S2AecSmwvi1TxdGR3TIXtlLXuNHnexxCiMwoqkK
1acgSHZUVTwLOzCpsZr1VorCcxcpy4HjHmoHd/w0zCzAFHLu1nUJA6jzcSiJ/qrkHl+/XCD+TEfM
Joluh709OrQRKU4OeJeIZXhIJ3lfqz6Dce6kRnnLwmQPRmZXZ056OOTbXfu1kbRXuWOftXJf32Lo
BmfonEP6CsAV2GwmSbC+PrdqU4IOvebtySgWaGkL39O/sXdWvPFOEs9zA9nOmhYxv+vSOG2Rsz55
DKJyOCxKNU/qTGs7kXTKZcV/Hh0KK/ken7JvmCSopLRS8DZna7hHhBo4jJ9F2UMR1kA/S3UMj2UI
Q6g6H8IR2Vc0rSnDJf3UxNdeExSfPxkTIdgVAv9FaveOczmmilBxTSsft3/tklm+jYXAqNcOb3gO
zSoc/z0eGDJDVFWPF+v3en1UZONyMjNg//V8Kwx7MC9QaFMPgo1Wi1xi/+hwjVdiimPvU7LB/juk
tEWqsJRSkflYhKZfCSPqpRQqAjktBRCXGN6UuVur5VkoC5QzTWWsmPmzeU934sBtU35lRoKgB4AB
l+j30cVAGFCwCpj7eBILUr82SJkA2pai275CI6XZyoXyLDM7eq3UXCuOMIPv1tRGHTFWUZuW6gF3
yopMvXyvRODPqBExV8qX9hSzPisdLy/2XhAGEIU8XCa69A4sTeNFPh0hiINW2ltpye4OFyuy4I+N
2cRn/d+AqASOsAb8TxtWxwLCduDqhcjFKMRDFE+xcqgxO+uJvPUbwQpcZSwexx/ljsKqwx6Jchka
ZBWbdpBhr1M9GNN9f1duCNuXLOiUeFfGvudjEZI0PwWrjIxV0z+SudmsLrFRWi1Jh/3umCo2H8k4
ZFzuceWYbZwsO0cI54HMHAgm+/I4netrFwUH0/Dc3eXRwDmmyipiPvzQKyvMntdqBAcJiKfjA2HR
KQzB5Mlqq8esevTWPIjqwJTCfXz1q76e1v3D0aVg/vYU468ReFwkoTozBA6IqqJ0RM+zNm7p+SEB
W6TF0ErOEkt9HMLjUv+GGkziD5RvO0gmKnUL7IfvV0yuYcw+ZfFW4/rVGXvz0H54oKNegwuV/O+v
AOEMd9JgbSGuusqBhC7ybmkVW+83hhz322LppdPgKQhzOw3jP9sHYrSPCAzKTQP50nb5s+mwD6a7
yXn1cBqr/J8pax5dV0ine95EgwF2UWo1o8t88A83KZSArUG2AAZstyix9DH1NSkogRUv6Qf7pJfS
bUyHIpjnOJN0Bz4reZYBwhDFMv8gFcfj87gD94rGxTuX4SExLDtBvNyIXUhxOpY5ZuSpAH7Nfn8R
Eg84Bv4nxggpFn+jn9ZWZnUETd/5YzdHvQ0+wzzYBRRwMqjtXIVIyhdpMA8aItFPegRbB4BkWM8R
QooehwCAMX8Na7J75DmV/ePWK0W/UEuQ8jS1cxb9hsDjmtgdDU6XmCUD3Ik6ttbtuyL5K3eY5Pe2
zvsUwZqx9QhQvYK/M3sQFB2sezVb5AipqXxadssrZhH9gIAobv1/AxKOUderzaSVq73xwVXdbUE4
Z+0wHGdxnSJV8xwQj2/1+FZFVZL9oe+pDRCck6/dV39Ml/yH/zJNM1yrE+EIlX4vPaib4SXpujCn
2lKZN00CADxBy8s/zTzH51+r6I57HDykDlVo78vH26unFYokg0PLFhTm2YubHhp0auA+iY1Za8Ls
BRTLTvh1xwlSiebRHVHV/Fq1eqRgIV9TsiUaUyB7BRcedTeRgHXPpWf3extX5mzsgFDgutiED2mV
DvaiOZ31vL1AZQzoLLsmDneMhzFRYqvsM0DyiO98NScMOKeuEl9poqVuXak3Zoc99FFuq9cWmeWW
MvcylcQEn7DBYMEcQ8SXcx86Cq4IeNzJ/TyhSySg8mDawhrhMV759hJuM/enxb2HRYdPpERdoZyn
0oyGo+XA2kPzDhB6eQ1dS0J1F42B5d0BUkjBW8E/yaNLf1y26gdSILpQVQfhX3BqykWOJjnC/zfG
OAXSQcrWFrKPglxKeTe+pLRrhf9JvWWF5McxcY1s9kTv3WZzbaq7XfjsL6bX0DfX7GJf1m2qUjqv
0Jge7OraqFd15QanIU4pn8tL+SjMbI5kq2QYyYd0SE9NTDXMa4Xg1ej0nbaJF+NXOJcARnOnzOiO
xvd9CD5g5cPDMbOK0VPVXqGIBgbDCgegNx8+PEk1ped4v+q/xWxo97nLKQo1ndMKq6Wly4dMhUll
GXWbMsgVz7bmEcX2/ikVQwjUdwZO+tBNJkZb/AznJCHIm3XZ/RTQTpuPldpstyqofIBy2YT0c7Tu
AlpeWoM21WWMwQl9DlCSKL+AKot2iqQgWK124TY/l21wZFMe/KT6d0zn3BB7GXMhElGETlUhxATH
T1CE7i803dr+4shmWDV/oi8A1949Axg/abxqjrddoYenofuOVY38Cinf6ytK/ioGWVmdpHJgWT/z
ZYdvRo/tYYRyupXNq+j8841JPmMmBDJLD/RoRK5wzg7FFB0yfI3tU8onIF5pokUB4knJXYUIEJh0
sT2PJtysjJ2LOb1LavlQx1FN+2CybBJgpHEtylw6ZcTmzeVM5uLAQgAUPzdQtOb9j+2Gvl5+e6RD
zzBSpJ66UVLvAqvAIkHtnOLNxKyJv7C5Fk/7fRCGKxL0+ygsMLKgxo//czABBku8vkKyC3f3vZni
5tHIY2S66RRS9xaCX/M7hgS/exJAa7h4Ub+FuMmtrPUEjsuKWYlFQq4f7TaRO9Z8HmzpQM1e28EL
A1qKlWqIxyqsaz1Rvs0LOOWybjpo/zFMPcrc859uQuZRsqQ8uwiTrc+74A68AQPqaXuvuXrKP2XR
+9BtEQT5/uqjCAXhb6euN5o1nG6zr9MmMGvFDkzTTreE8BRFlLWZLXzJYzsg4qFYheWTn9LITdiB
d78uivyG6vXMa5L+M5A8AD2aYxhdr6dDQ6jkKp3fMp6vAUwltFXtvSQJuIjHk0DTVuhTbbvEDV4L
Yshwb3dH/flN210Gg/Jyq+fxhFAXkV6Re2xMbJxclfvtRVVzoB4YcWyjksRKwubBmcca3zOTbkhk
ZZfVjNut67XjeiXDLNJWKVaynIO1dJZlBKo1QW7NNMmPGG9WB67xaaOpGtYDo5a62n6WxBdUoYtz
EY4juZPWCNu8Gm6u520kY9LebSzNf8RimTGnwLikJcCuM+jVy6CtSXz1ZUDZktgI974voM9nv9+J
oAxqhPnh1llwecnmYelkdNz8kw7KVdMGTFTQBt1bKwVmCzut4p9mbugfcrgQW8v3kwnfDhst8TrA
5Va360FCfAc3L1NDD3s38GuLAfzFFCPoHzc3sxAXdA9PKFvbl7GArL7zTTMhdTX6R4Dho7gpVyHI
qdm669RDGAAipiFp7a3/pvHQZj5LuLxPo2Frpjki+s/9AV+m3YGYuNR793tYHeMDnOdzcvo8Eijm
EyJOxvhTL79BLEfcGu+dol1aAONfWnUYcMWBS1dlGIq6CDPXlLMe30Ka9/RbV0R8fVCJ5Vc1l6bN
d5hnbqJzE+J8BlftAtYK2w56A5NNO38vA39CK6QB5Sh3f39z9cv/eS/B/RbsfvCZ6oE3ziEl4B99
cUIc3mD88v+GdGNvYi2jZqhhTDMaoSxZU1N5Pl9QDbje40anjldQJCcAUbGlUQvlW+KgixcBNvD7
RgnG5kiHas4xiTjE7s1QIA1cL8jV152+6lwytI54f2PhqavxO1Cm4HitqBLGXJxIRtR/wj2ysdc7
z5GTx7pxMddf9C/pC666WaxzMlkZ9JuIOrT8qZ4Cy7KdyI8xY8Vsn1JfMX+n8CDn3k3lf2wVjkC1
2tZM3XY1gAjvar5jx+ew8/kuJPU02gikpoH3kDLu2/cAm+v9LzvuhRB9lGc+FTgb4+PZR4yxuylK
CZAfYYbdKRHKBWKry7XD+2rse8DtolMYxtONE6zr5ywk8+WxfjrEhnegPj/SgMK3p5SLUqjsi+5E
AYZdSJCZ4bKDrafplAb+01QiXlMQn6mrdGIM34ha1nNDanMxLeGj+mUon+FbBnUd2kBBtI0Vv5Xg
Cn4wIr0PVYBvrYhIGWopCEge2h24l/JuNDBa431GQz72eXRJQI3u/pZ2SKhwRcq6hDLMox8Oo5Yo
9hIlXWgXD4gk4k61KxSY1o+591qTUFBTvo2KCuXXDBCaRK4oAZzfZoplm7r/OCGiyTWHd9poj7rc
Sxs2/bA1PxQSqEr5nqg9whyLAB61CO5+yyKFjDKRh0agjbl7rL22oSNns5LqSJEzDpENDRYUZ74Y
7Ibu9vSRwaVpfRhFPUc/woKjYEcGy7gv0zhnpNXoBsY/6Hyuu5iBXYE/wht0nYK423ZsZ855smEY
GBtL0vC8mYohebyLKrVbsFl/MFKl9ZjcKQ+XwBFTvyTl3mIdDGn0zZdsCkhy9l/kvRbgyBU2kiOH
2uHLUat469AruUWlFddXi06cW8dL6fFnYGrxTYOLly2uJmhwUrESUFvEuu/OTK2eLoBfGWv+DbJp
01ck0eI9JhP32QKacbFrEfKNJCW6tl7LtkauLdBhkLzhw/UPcDumZUu1xqxzn+NcO6/rq3nBhLtk
eD6sn3m6A3W4RtPkrVU38syrxFHIUpIVzL3MlHNTuPw3iKU9bBkOnPCKHyteyAeN7uCoHU7v8vu1
baKqmRUp+XnTr7z5GFMCsAim/BggMWFe6M7JWQ6CxSeE5VICWJ+zlF4gO/9n3kJB7GjS0/VtdMf+
f3S4djWarD0nUOveDrpXNBUUqm5k8HtFDmOVXJ1vtseNBeLqmctG2le/rzRQbF+Porgb+J9jwcx6
KW1aoJQwGa07w3ZV2HG/MO7INSX5JBHTAK99vm+By/05vn1rJoueW491Y0IC7hqQEoZbc0fgWubw
CK9kKl+nvgUVr3QF/SEQzj9akm+OOEN1tC6i1SZr9fgqulb2j1C72Zyyt4HxM5qgsic1j1opSbI4
Dt9w0E/jgZr5YQkPdItstR2bjBV01Oa6cIQDMoJGpOcBuGTBFW6E+/Eokk6bGAxdA3mTT0oXA7RW
S5bprDZ7QjSSl0jkEyitAYKs00/nDWwIEGMkYqbxW3BjCzUwAsOThzCD+N9LztiXwx63FxqcSWhj
ylQ3k7o9dXPgtGw5m6VVC1GkKIYawaonwpcuVspblgTI4CeC2vSuV9gbFhWZDvyRN82zSI+l7QHD
lky4rx1RhWxQ7sH/XXhibk60JBA+FM+AUOt9ATvr3l9dkIpU7jRjDmbyMe2rlCVJezSUxmkje9Fc
y0NeGww9aBOJfBBKiJWTdVTIthv+hVyZLkdBLEACB/BPxuzB4TKh/Syn1IIgRWMLo9ERnSPExXGR
BEwVoHURUNZobnGkPGvfj55ri5nCpbrwXQxKVudsavBSIRBAY8EuIM6ppWROgsGFIRtObtc7B/LL
4vm4Pa+SVP2AxstJiKPCzjHz/bNDPWCTR6Hauex2TkL77smfSPiyz+/dMEQiPoN5dbdeMxY4pNvs
PnF5oicyPxltdKjsUaQjnOxR1rK3be56QaPonU7S0pfsTCqEnlDxNu+7q2WRy2CmjIMcKC+ZSBKf
fVRUZZACfsdcmOweUgJSAIrOSVHT/mSLihTcpNBPTlvTURhpFqubLBRNCU04EiNVu2RFVHW32Gqi
cZdSLMTQhVt8xy/BddmuwatSttJfGp6bw43zkkYNdBnh/x8fAM++IFwRIqG+yGGt/HqpAOTrs0Pr
mGWJZocY7yWWhGSqUP+/7P9/1XJ0514YZdv/4SCQe9jypaXeFZyQsnH6w/b0iH8Y9G8Cb/Q1JIAF
CjrNsngVH2UeGFSChGSdjS8ySQALmbaOo5Uwb4i7CH0esf6IFuCam59dw6BRy/F76XMJgyMXlqro
zf3ty5nLZpXjpfO4ESH/xH97IwSB4vHDVTeDLlyCh/m+pmP6ZF/2N4ie8mDDX103zc2NoZY5/FsY
3aPxoc9NQHY+KmVo4V2MJL8V0fsYsyVr6lduIsKwXJg9qbB9/7B1cNhhetnkd/rpLXoxC6IYJ8b1
39RjwNTPz4NE12FDSRz0tL2l1Ei215AMjN0rs/NJqweEU6CotuGoqMpkLE1hpGPsLCflvpBlUTxX
ROpATMDx4zaCh8m/HGCTJsP0dAFNFTuFyToTFU5zfiIyJbJjHEB/uvNBMRmof5dJ+KNKwxi7/T3Q
JUrRatficzBDgYq1ut+GDI5hI7YeruScraU6bGV6MM5IeUJGy9rrb6mb1LB4PG6eOLwmbUZHFO4t
4YwmFDIhxqqHMspzCGYC6cKa7zxSNeVcXovTMI0FWNQ+VubiOE0Uq/j2rcIn5QGbzKWtKYc6jCa0
iDVwvvghLtF2A9PSQ45zUFmFUBew+8xhYYNJWX8tvaRx9JZNP1MdXrGKKi5oguZtfhOjdeZehoeQ
T53Ff16lNGNploWRGYsVDU3YVc70MEGdstbaaTiDHbprR4OVNb41aoEH7VPtNbWkL9Hr4eDC6QI+
xY48seolIOa7J8wnTnQ65ypuIH8XHKq5SKRKBsE3dnr5aXGbDW5dEipuGpD01TsPjkZUAyr+NqKk
mbCs+kPMk2I2W3fYvHS2rzfluOeXtJU+7rUbWYbJeoEBXVxeogRiMoPn9h4GqDji2+BsBt2EEdIb
A23JLvJTEQnWC0yEmm21Cd92MTSd3nALXGXxT5mM+egXXPD0LT/E1B1zQVKtnL1DK8FH+7qykcjs
KQ5uxfeVkonzZGvXtcf3tZ20uLoQi3pJ3VuRljjZ7Q43tWYJDQPaPLM94kxqj4oEDYAqHDbxNuR6
Jv5qtWn8OzhZjkcruv+fCDFXTHBcpht7rOglLWGEL5uocvP5ir07fbZ6oK2LMscO0yHj1j+vbDkX
udLr6fbx350mjFrdXd/c1TrJjtM1iAePlAu6+IjHie//DZUuNq4MdOxpoHq3HMpHuuunMKWGhu11
9QuX+eGVKZFI74MM43sNdJR0/weNX9+x0bRQAMyxSWXqcgbj7ngUZu68tQD8zIC3h9G2Ms/s294/
lcrlC7UG1XR66tfi0sCvbBjsJSxNNlolnNx9hy+9Tjw2nTMGDpho4n69INy2j5mn+2phSVpXIpz9
F/lUZy/waQx6SLxNWaPL+C/npXrdUJNJ1bW0IjwE0qJUD9bmYSStCZeEq5jBNfLqnkjyY4zpIxV0
kgxr4f1lndkt9EoRspsKr2j0vWVWg+15XN/gJHVhDUrk0DB3GjQ2yLdpzefKXLvsdWc5rcFe8jmz
cCcG+KPemh5NgvjYaMh/MXRdFURAHi2ZAZcgKyWb3wStA4MmzfZW0hA9HSwQB0M5/UwkBOe4j807
RTFlRKhd13K5o+u6URs2Fu/FAi5a4t/WRGUeQFDWX+Osggk+Gl91zFhDiYSnHtqosh78MS6N8cKq
1DlXXn4W4Y/r6UocMP22xz0lT9pmYG5oPFDrzoim0YdQUaHsvlbT+yPoyMVp/KeACe5XjuyT9miL
gA/J9xNcweyZdzhFc3q4/xuq4JT5BJcSK3QprxXCTakQwpxPp4sAAohVFnjAi6Yg2kMMuE98zUdS
/JhbCPzwT+UbJclH5nVzNH9PvA9pU+2muJao/0JwKu9hhosWtFZuQT6qi93uzd4LYm/PnbpXGdLt
69oZBKx3c3A/cBBoiMGxs8R4SEWFQ7Cqhuh2XiP3Q1OCtfLX3HxmT36qI9mhy4qOc5tdjua1lYc2
Qy0Du6vxi66iviD68zzBuP+jn59hTRHyPn4EOJfSFgUGoH9JW7L5ydvxTAAUY+lrnfT36ES78FbD
84Oh3Pd9+5WDAOF2kXuCTUa6jLVORsu2cCzk92Sa286VOecYe2DpnMfhUPb8BgLkJsBqQXVfp8V1
fGN7vs4bZHgNQG22OdLOE3Zx5fA0CgCdZ60P5pzGSe/AEtxCQUVezsxxeUHaNvaHI0bvgcSU2Sbe
M2sY1cU3OOULUASqxO3gicO+Fdskj14IRaA+WguPWX5PdGN8liuVUOroLjr0DAJ6Ncstuqm+UU6L
5zaQvCOHWp0epWjKJrbvgR7tn93wUzMbHfzmzrc8/ILuOYzW9dGUOEp+vihTV1esVTDFI72+6Rl6
Prf1g/UnqvvbqCCfcYn+LkobIq7nuuC1DUO9IXeczoBdsqd4qFKi5LCIAHdldBsamu9bf5Azvcsz
UqdDFI33Iusg8LIgjCgHJb5L6kPZ5CroXD0S6cOrd9sTcjNkZRJgPRWWMx5CFCYxXM5y0cAPa/c9
mlP0OqO0hDwKvETH64z4jF9N9jrEy9Qqv2jOC/c8fHbHsiR+S7rEMAG8xnEJOeAuOq/GRPXrFx7n
ZkIrtHdTNZsD5ds3W+SeuPc3Z/Y2Ja1p7DDQgN6SR65+CbmFfBlrS55OMNp8y8yp7JKCGdCh739E
HJCaVGPkJAcV2XfMFN8IhEWJPHyS4U827GeZ83tIGSI8sq6K6wlrTlEdSLAPnfPisIADkR7N4RNd
8xOSSXYu/3yHfEzVoWWvjUU45fKHNwTLoIEMkLA9Su8UCoYgjaw+3OnoJTvx/0/g1NlFmWyXQmUz
o0F++mjMZ7KtwvGexl3DCJDOPf/zEfGXiTGkL8MvN61wClc2CfE0i8KNMS4qXt9vocOdAPNnDfS4
vwfTqfnqpZIvD0F3e5Wt+iNSpyWuZyib1x1e9FZlT0OxUqxx4y0GHsA3RL1940Ypex/k6XZOX6Fg
CVQqhCzwYtuPvyukoWJr0Ci9qYNiV1CNorkLfdoTvg/CbEp+x2Il/GY6pUFqT20yh2NxNVHjPYlL
RyKKTJ/nhNPATPhnr1JvrPF56tAWjCru2LMnMB4KF8sx4GcYrmsS4KSE+WlSSecupItk7tNoj/JV
wy3d2N6I8HryLktBlS2hy1Twg6xk74P12kM6FjnJJEA4owem45eSpYoomK69V6/VMZjg5CYirlUT
UG6yG4+UAEoNiOo3+Th4t0KVwE24lxwAljCY4DF3Bf7YXpVdYM/ctMrMzRJbEZL3G329hklcZicy
NFkvgG56BvThVxxsDnEP77IUW0+esHl9EEc3KQUfAprV3nv77OP79KKkSvNYKez6lPZo4iUyJMIj
zq7aX3xajIeaDlqliH7aRDY/Peqx5azcteHfBo5zjUguPnqF1791bRfKyggQs2x/VmWRlpYYWjby
oPWcWDZ4/moEWuouq1IVl+ABbmjPYr80o//hCV9DISuA228431GVByZZtbJcniebxXg252I4o0mx
NG/huPb3CEsui52fDxsUS8sWgHkUvvotFkO8tpohNHH47OkyRy9kcqFoqCHag9a6xcrYXGQVCuuV
iYk0kXzRyLWvzQxo/wsZIuqH3bQX3fqKk/bSZBvXgiEUQ+sXbdNtqa+7EqqwGRDD6eFh4A+Txknp
Zqkymbs5HmBQOG76zD/beRSgRD3k58faHCOQfYZ0u57pd4m0V5k2Yl7BTJLG5dpyNNLVk/voTPZz
yx67Q2Kd8zlt73RyUTMqKHBkxp9Zz6RAuxsNZ+uZiMK1AuzrgtofP/cnBQBm8Q8GhnlnrxjsOIdH
sF5I57OHta+0kOyFFqJFYZFCGGJzvUPzBX3v6eY0W8XLvJgUs+3DjkYXak7YE1dD2WGJIgS92+8t
Ens7c8m+0+yiZRST9AZxZMcDM9B+lVpoEelNG452g0ahDyzUsPb9oJpvy5CAa8Hk281EocjHftpR
wt7+h967ipRK+4YVbjRZkj9ppPGK8i23981aTmZ14FYMliTo5uVubj0w6QG501MT7VTNy6msuEw4
JdHWYZrdhxAVf511sTzsY0YAXTq/NrsHSD8Sb5H544VQlj0SeZ0b0sfFPb5doCbcr8DDEa1qs/nt
Js8Bs1yQypi8sCf1IxTDQeLwMWVObpKtfgVjaXB/qnB6ZoyqhLlwv/beLieTzsRXs0W+vnX23rAs
HkgnonutYW//Fzs7HU78kKy/ZtS6aD7IKzq3IY/rk9HvSQ6AcKRnphFyiuhtOFjIxMVrTZlJMaZU
Dh3l8hOuuISmefD28L4ChlT7mLgTLYptugS672jnbme7ylo4BZmLTsOpKvZC2Wt/ZLPb4HWmsy4x
THdhZ5al6I0qRg3G3Q6z4bR75e6XH/kbVQZDPMWe/QIz/0whpsrA0Z9qOVsTEtjr5Gyi7LjLUgVM
CPWqeorRei3ru6+3MpSQURkATYog87F7XfVnnEOXbeo66LJRK1G54ThXE3/C3ylU9vuscPuE6Gpy
59fXiICv3CxISKRqkoVICkQKB+DGMKKcB1ZXkzVcWchXO6fCSUc8Z9jz335VE8tw4Bxgym2RAS3A
UMUmGDccVQHzt1YlP9tBtLJKcI1Ge0LMPM/9p7Kio8RzJ989OCs9e/OCYyMjbZX/9QV6oVxnUu9w
MBquhNQ4S5Glfgw5L6+UPKc0ISm9BZnDF5wBwkRJRFxYKWO0NB96GB65gyjxAZUPtjZK/IiqtTfy
5iY1v5xeNZ7X4+z/lbOgb1h/Ulg5B0xzr28byYlYdEbP4xBQxx79WdPF3JhdWVANkNgCuWOet6SC
JMZkvDItdF5TyXmsNKFQAMLuBuJMl/FyKkXDlJMSUlOBHl5+RCDWR/hYZrRCdgHozwcVF6nTpp0U
At1tOwMEqpzKw58B4j6sGodTjuOWwfXFZcDWL+ixMRBhCPAL60tAlALoPPHIEjKCMr7ItKezO5n8
Z5HBdsB4QghFLOddjkSmJFbsjW8xPF4nA/F7m+M8UKsgXGQprYAbvn/i4/4PTxNh0JVy6GdrM6N4
MqaDctxbHo8gSl6iBjnezTJ1HVmOD+xG8z0xtPdLpDoePeHUqfvkJx8hQH8Ucc5qMCIJ/NOgFKT9
mdYidbzeiN87WvpFWjKkudDQQD2yX3Fn0km7eDPDitj9whmDNPXOFyZBxkDxPNwxenM4oXX1soui
QNAEgXJofptXMyBS2TxLn5fbpJJT+7QVDh3OO29fj1rmcxpmK2o7rbGI1blkUq5OIC3QGIft/Ne4
gIVIby1IrM1lFc/xHj7BWHAlHHu5a5zTM1yxHoHlCrLaBhIXJ/BtuE6OheZsaoXG0c+tqYOlZ+Q3
yfNFCqiTkG4hnIj/5M9Qg4oRLQ50tjDOUOp4CXcEpQlX6pyTu6sZtT0eb1dDVyyaLJfr3tlYX4ml
XMgbSGu6ojBMJgdKzMCPpZx0qJDnDAhfORYIfOHKbEYSp/YpoMaD0zuHjKbrs7nYJQsaSXcPqwJc
m0dn/E4crXPHMOxRtoYeB3NbVtP1peYHeVY5wNQz0aYG6zQl6oYSfhs6YgUIcGEHgE8qBGZX15a4
+3oPl5wVht9TRnsGtbkFSUaOZrKNBcs20uFUIvB8SSqDnopvvLGyfFWKNK5sOfuWgBkIef//GPRQ
r0nQNe59oTjo2hnAMHWjAM9NmiYilKxkDbLKsWd+dXpt6Jbv5tTgIKmQbh0MJrBp9WO8fKYxyAGM
Bh17aHUI6nXYT/oIzkrA6s9RZl5MJKEYsUWa3RxCR1MGmLIBWy57KdBmWYv6oGJZaGl2edudbodH
eXbra8GAGneoF46dFW2VQfNM7bn7oSDdAzjsfLMcXjuEt8KzfAcL3fOkgkiFKpdyUqdMYlYAVEDo
3JYJ68l65Mw9qh3DOK8rbxrKZpjPnDIq6HcK71yEsYtXp6N7u1omtWtHFEJKfNRWYqS5V32LxBul
MR04btWwdsELiCJLenXE3ZSBN1PKsoLSV5C57z+EU3flf2w1TdTkUUjnyxQmoIYLMAy20H5SosmN
ombwFOURVmr92iEX/eETu4Hy8qSSOdNsJBSz4kFT2sQnxQ5i/ozOyfgQFzai9GxWdA8nl2CfAQ9S
Yy0psDeA5u1Bkc+fzOg4AuL89/LTjVS/m+RJDUs3LAOubaxXpzRiljuzOokEpHJtiQ9XY7/DrEGj
gqSgQrPwjnhoWH6HByDrrd2O7W0NyPowdyPS4X5bdG/KLI0Be8KJPG7Vhz/ltNFStGyOi3uHIvrl
KBBmMJsdi5eBFwtiopDrluTTQSGifUgRHQJXyEa4eeszdsIkfRg+Ms0eECqsTgbk+nXGHYo6zy8r
NlP9zt7qF4TU7OXAMUgb63qo3u8JZY+aZ4j83F51IYxgn/nU+ONzIN0QxrE8/Ud4JEJIASVdbmWH
NK3MwOswS+L0p+IVnRugwPfAgiSqru7qcopdI+9I0CDZ7iKu7teZS7KfKTxQMkQj1lvyABYyCa6j
nnbtnEEKUJsnkYGNNk3WuI+yMKNTNQGNK4uwUDsf6EHKuH8xkQ88Y8R5ZSGN8qH/FzVNl7M49nhY
KHhwgOty9JNd2SyIREI6YZ7hlTOW8EX/xpPKJQyRHMjqPkbpWYTX+/xq3/qmtFh/dbdBGKyGwH//
UW7p8fSNpTwwvJEsc8d8D71eAM4n76eq/vNZ0w6K6Xqe2mt74hotvonbBcTqHTt4Jlv+P/dnLZ7n
EK4dkHv0z7Gq0qPca2VqwOSkM2NzAH/svZ+9BNIMf1MSOYPYzf8wfRL+H+RInViRPRhpgcZ8HeFY
209vae34XZ1EB93miAKk6gFwkh91YJ7Hy9g/A36KTkDUkyxo8/hJxauBOndizqbrStJHSvzSrtUo
VpeUBqudZOWVtQ1EBZC+xiWOoJou/zgmd1f3Gmt3LXQ5NiAdw3keYxAwfa140J/jnvJQ2L8+S0/o
0nNJpthf1AXZACxn7Dej/oJmpAGsJlyDPXUrRs11O3Ao3qPJyHjUQJNGsYqiAG95pZRExl1XmCI7
UYt8XicwaL5cZ4YWbg7LxwJ7hoHxG8dvtkTE2T2jUOrtWaOVVt5ztLyiWHEi1kwejs2+U+GG1vzj
bAngbz661fq43zYvuOEM7z1Ds3Zh8s1cehVtKFOSkk4KOgitKJeYrHsYtOYgMfNy9LPh1frdtheh
GNQY6VMtse0xvHqbyHMeEg9jeNIXdmttKxeSwIJceyW8vmRCyILq3WfTKJcLy7xk3ES3j2RY/C9j
nRHUO1YOBTTIAmZf/G98shbz8kDLIijSD7w0vvotnh+8wLIHs2oS9PMV14KzEjpjqPmlhBcDBSPq
qvcwWWicxoyI3qq4I+j+imTn1OSNzgpbGfPQmYbCu0AhNgu18m9eIWgqqs7circW39tl3NEcpTTv
dp8MAX+zla/Rx0qTr6F6hPpmCbyBBEPAKfKZvjVNW9YS2ymNLaks+KA91QaqZaS9pQXCKtVtXjSC
OU1vR0c0sOSoW7BGIiBYROV0yloujF10ODkKHS9jMCldaUfqGxEhHCxK7WHbXY7hvoaSQWXGLMi3
oDdMDKrd5W9Ef38BhfHh8t7WUkaXztr2qWt4DTtcSEs0IByxDiN50wXgLUn3UHBCHJk3x8EPqFrl
v2whUbuh9iOth3/GnkJL8tVNfTy1rAWkAAPhWLlifue+0N82g6ZokYMmBEHkw9uWTHEVWEEJ+jpW
aaGfGIx99QCsp86lFC7Q2IQUc/nbJF/OyOFql0C/AWmgcZAYZBtwlrZpDULP0GPC+BeM739IwGqr
bNZHSyBD2gQBmc3Sopuoq1BqaIFToG66J9NRFkVWamSpMZlRPvXtYA8ejJG8+IzGPxE504J45k3s
VJkbTfoDrkfKngpOvejdaJYe6lnCdUX8Nopln4EASPRCyg33eEiZ+G+ybimFGVvskUy4jLy+zeCW
Gkn1ruKOW8o1vqC/q+I4/KCDbPet1Y+eZRqn1iSgysRZMh2XAM68cTNSZwu17IrsZSquiqXEEIsR
UfOHl+MY/IwHnG/sVPn3kda5b6yMV1Jg6zu+tzHe+fNikuBbRrulfXgck5rNDp18NK8vxoGkcNKv
Hyyqmp4n/lFLlPo1B8ynf3a60ryPABHNGOWXg55KFJSRkaRrY2lNA6q3typ1fGH3GHGqz9+JN5G5
69TfQcea2uD34p/CSN2fJ7nO6U07ezYX89ygvIe3P1PGD5om2TsFe6ZTd2iUea/to21GPFJ56O69
B27qO4wi4I7sjSzIQR7mpCIRguh28PML97eOT4a+SVb06mU+4uTu8rQqGZb2q1BQclTZmWQU+vyL
JHGm6+i3qJwW2HC/Pjx0gO38N7IIsEkpC36O6TsKJRF9HvyLkDCoErQTB5G1e2vYlf8NmHeF/8iq
CmYEJMoErx9isnATLUHEwV3B1/xpxTEz9ewv2nTjesSJg95pdzstU8DoaJM3FeT8lmONbqYnz3E5
mxWLFatf0YMefciapALLaM2P5h/v77Fn4PpxO5mkVfw1Zej8leVuNXjLYDN+MOsUYAidQ4zYCgJu
qE7edavWa2s3Z7b275kr8OQEAGNJe08YNcbKs19XIoNIisx3Tb215H2rVT5HvuQj6sxouN3UzGZd
6BfojCdyCAKj+2TS9NCp1ajUpyWFmdRsAPVMKWvvcW6fGE+/i9Em0/VOowmWI5B/5cnhg0eHlPaA
0SLIMjLSY25UEZPvr8+y79nZ7pIEfym2EYIZUuG5YEhdU+r+cvjNNckZ6SH7W3pgA32z2OYyR5dc
d21jpK6u2hiku9Ws5GdLJwFgMCF6ec/tJjhDriORKhPN/NZ53VumvKhVz1rci5VlU5WqKU8PbU52
PBXWQvY9MKbjpbhyubo4m9o63gMt9OvuCPSmW/Ux6JXZfo3b9OOlaxZU7wUHvXyS9T9lYL+BXAEE
pX7P9rPkYHx+osf3S222T00Z7ICHkAycAmK52rgt5PJ6r7kKLSrD4/Y2zS/pv5XmRVkR4Eg1JdlF
UdGpO7hHv8QahOIBSirH04DiOR6kGKLgoVIOrZJU8xZZiNglwoWcqzHC2WV3fpovnmDPUBK4gbZ9
Logx5xIByD3jm4UJClSc1es1OC35ojztUII2pF4+ZZpLSaqkvuaPDdNjpIwl1BstMfXg66ZEudnV
CBh/Gi0oR+dBXGCSKFWS4yQLaD2EMsKalhnmYBNFVydJVLXQz//rMGkEeqOrdjRggOquSZtlTaE4
KT8cWxzFg8CXOw4kL9V+wpjK6DE+56ztUOkDThRykM3wcuMNj5dYNCk5UQdQ6/RDZoXnZ0QGMlEU
+2RS/Y5U1GhaxqjZHSpoRu7hEdRzr+7asmjRvRovwdNzPLNb0QaJxJHHteOUAIPjMw2elBWCoHRr
XATQs64vosCM4RBRg4BvjP3fIUHZErTuVST6qVz689oynI43LwGLCMX1DpLLszl575sRrRy2VEbc
ft/hpbzNofyV1iQjCBp030fRuPpaPF0XBaL6lMeWg1KYv/50eV1ibCJW+uBsYPJq0xPNzALOv4SI
jsG8HpZ+65WkrYZhwJ28NVPtQoDO27VpMvVOVps6sr1uT+mMMOXyKKzyvwaGhFScKcdDqxjMRXhG
XTWDnA9lWIV5Nwa/8n78lXecuD5kOJADtb7gBPXEBRYKw+YJqD7PdiolcQIBNVuwF6wbOanR1Xif
RAv/2X/nbYKCJ0Ig9i8TEgBBCh95R61uSN6VSPYmmXiCbL+5X4xNCsonkQXN34v7JBx8nO3V2/It
fr5hKt20L88hu4FcyMtW39IsGfNKYXPoEwya/8GB0av8hWmYmCl0fl2y5TTQQVhK3NKI2lEuyg7Y
SfjVS4mvqgd1NMlxxg1M4IyeqA+7CK46+wYhfFM9FqO3s7sh5feH3wDaA8DHDkipVRK7kl/5Stum
7CGe20Z5pxyfyioyXyKDMIZm6VBisX5O9wgJsoYhNZKioESyXA5NMa4Wv8zwI3Tj5LNcpPCm4M7P
NT1CoUj96sjOYguKMmpEe5V0bAYmGNUWqF/KQABnYHDHS8V+FMv/mLjuTtoNH1vDt07tVT6OD75c
OjEYATxZ08IevOd2wCd0Jv9JJ+IRS0PMklWQcttwDAVxg5TRRiLROiriXhuSrGKl0yIJoiY7gmAv
f/H7RTXetFG94qb0iGVEqwZcSu+1PsehHgnXT6J+VvlOTh+sr+Vm+249t3FXXtMfh51nhphyPf8e
8DI55kHbtMOwIlJUkHyf3CvpoN6GUavVb0EOwHJrn6ISpl7IP8bDF1RtkPbiaKgGo8awzHo0Xgxf
2NndYX9RBBGd1vYWb9TwTpluKVlCmXPUDLaVgTY8N5+mIblWiqWh+TNHh76Y10+sOkCAHCJKUxau
7UMjLgspVcu8s7tos2n9GlHYxoTnKOT+arLBatok4SPJ53nKw5ilYVuXZw5EQ3/KyyVXTlO8l5GE
0XyzSoSyrRmtaWqnLPR/5O0ijcIp4grYDmGcPnwfB6kQsvwv5djhv6H0ohCbsdB6a1aN7YkIqSB2
136ZJT/DTtL1q/HG1129SrTIYNQaOiC5lSiFgTbahLB+k1Oksczh5Y1DVGIRyyQn4u9Ag6Z2PQCv
n9drXFepcjqRzlBW6kT98MoRzLveeLX9XgOTXS+xMax2yr1fuSXlbxzqXd18ZeVR9Ur2anfkm5Qa
xImSzxFOfVrSXkIlz4D7K0K1+m0Gr3eUZwapkGgFfDBB4Ke+OZukgWJc+qRtyn+0YCCZwfXRlkrZ
PdxGZGQIpsUtiNI0BK4qg4MztaciTFnAV7JgL3do1zDweTqVM5JV9GzMjDMmap/wejY12teTGFFY
1fP0zfN1Pywux4DCVaqN1gxNOBChAMBEJ5Kous8isjrWrqL9xnb8oN5ZtY3mYUYlsPCgVpaET31A
njab7RP958QAnIVrreUmaPaVm6Q82K4KegQ7jte3c0CmoLnWSvwt/CGWXfUwy4ENqGd6gDrlTkzy
yYWDuxhjiwIH4jpKGB1x8InzBKvqt7w2PWXMYF+/r89zD1dffTXs8walfljbb3D1cITDgnZ7OSrB
2nKD/qejjttZK9rWgAKWuc1Sh/x//5O70uVo4/6QQKA0nRwpmEODCrdpMjN4VkzPSbi//QrwUYZk
Wr1JSVc55um+ZkOQONrjzpfz3jXE/IotEtnqhwFWL7yTuehPGwBLfsAzlvpP6b3VqKVcnGOGJ1e9
DG/AGETkUbzim8zacINB6UHSVxh2wSrZZE4Cb5amCd6rtZFi7Tf51QSs0bvwbSuqfuCvnswG9tOl
BMQAAW/w45w964evuzMu0Zo4BIHAc6wX5RTjfvx6Yr5XOI0a2bgTUR2gOhBL7apOjUSSy9I5XCwD
v20ZJ5MZbyfUyAabsVlLGYaZjzX3JXkx1H9otuI/wavsCb74+jHUNsT2RiDIWWOlLYjQky6LUIVp
UvBAW85AQ/eqmKfp4COYPoR+yVI51F0u5jyz4Yvh44O6ObeNRkh0DHev0AYzl8vtnHaClvB4hHVl
uTtuXqOKUn3v243X81zZtKEo1UjRXlJS7m0OHaflYrf0g+ooYK4EJw1TxlKXdI6+YgdSePhtVIQj
/jgRopo9aTy0q34i7Y8PWg7/cZm0LbEVgGroj9Jqke8nf4qAdPU3hu0v/pWBHIQsAcXAN5/YSRId
w/8iJFdsuAQmcaM8jq+ZOGksbrBHP7+O94wt9elmqPfuv2b/aWaztR+4uYoabR/GM2nuVnNKD02w
BBjPRvPNqyQzvCrPnGbXUferoBObPo36OhapnbferDqbJvM5VkOZy6CXlz8BSD83KVzCRxvE5ZCe
giGBBRpNv5CaBR+cJ8bg7SHORFbdLev8rsBarOURi9Q7d2DrquKdm5D/iWdMZCDTOeBO6M5x78Fi
4iabhmb31Ur3BDD/hYIdgwbDLSaBEQxoORTP0S6BABHVfRk2WK6icTfzcVefAYkPN5JkXvD16o+9
nkeAgjBqtnwqZ5cDSXKFTgnGYtFyrxdicQ8Ueut4OojyYJBdO7m7xtY0wMmpyZ+HFyjCo+d7HcFg
fzrJhQDQ9c9WogmPO7I6sRIxQ/8dwrVAy/d0GLULfvrtVGxEzv/S+d/5SsBtjteeKBIBwLSG/3zE
OJFmLbzSqdaYpLihCsnYvSjRwmPLXOI6RBbCM6Y+WcuEHNT48VQO3qWV+gkapHb+XyP99znAY2wk
R/fsrsW2OtUusl9b2Y5TAw262mHmtKg/F3hRAI5fqM4mS7T88JNFqnrz7vNjuKJgV08GcVIF0eBq
Rw06Q1Ka1YOSEKogvAKFoeNjrdjANvOLFWtBKlxmercajgZCAJt/zll+bSfNpveExWiLCKa5k7Ny
wiqcQoh+OoSrNzI+X5ZJrYWWi44vYpB0O67YHOQB1OCVJNrfuA2xne0DhpO0FpW6pVAxLIZpCvx3
bkwr70BFY/HXQqphw2VNBJF4TGtW6GKn3AvGKr+0NEysQZnSvI1ta4doEQ1eyhWxieZObEeUu6Nf
0CtOmKPNrZ2JfI/iTIlNmKPzEsstIERHyS31/G31PA8h6fdcNqRS/yVhCvHTdSExbwE8sUoRixRz
C9MDK0WWOHW/Xk9Yh/b5Bjadfb/5npnivbQilhDy0P3z7zrJz8L4sLpaTszWazQWQ9CGxlnq6ZKB
H7awfXt53IMistqHxgX2VFj9x+lQZTSS5KtDSDuXTbPjPyUiYwOOoxEMltviqCtbHio8r5S+fbLP
rmKnFsfMCNnV86nfC//BdsguU32ZEIyOWXiXJJZDPDOQvMM444IlkqGHXEqhsTp5XbtoX3mpyatu
AABSbTQTw/0Fwp+8Td23poef+//XYpZZ8UpyMgSmRLEMz9zM7/K9x7Sp7Q/Hcw3214iTQH1aGKlv
ByXwVZp2yJWo/1X6GhKw0SZoRsM7m7RNhZ+109Nt56uW3Xf0wtNpz2cVo9gYapvfis/giaXazxdR
pUkK0b4X77gVjDcoXsyWM0AoaMglxZGDWyKX5ZgxTN9YK4URELiDcc/8jWnD6A9vlO2H3KmTuNSD
jF495/ljl4VQW1v1kuapF0URhkLxvLm9Bi4iYO1TZn081MlfltRlTZFf/r0L2AA1x0BNfWyFlx10
N5nnEb9UfJ22sPwez5Ba6aLL1RNhevKtjzxeTGBEAFV8uhiclBnKExruTfV5d+03+gkhtbfWjUp4
W8cstS51CO80gRwWZF1/uWa1CNTPwQRns+xr6CLMzz2gQXqLQtDC+MjNpSmdn73pGL46gTJz7UBp
npnYhaM8MXrgaOCqPfp4Aa53PjII5gTRVVQakaFy/0FbEzEE2rlS3oozyrwG93B0oPkYGhKHhvPO
RthwQEzslJwcubNiOPA5oAxclCdKziGAPOBONqhjnyfR73ujggjm0184XcNZz3ctxl/TslLabC7V
YZYUpJbHIjL/J/8mn0Eyqv+HnDJbfgSi1WHLrzUZoMb91ECYtFupVDi5t8ScARSTDwKv22BgwGXK
XS/+vkxoDMegER9hKJXemUNazl7gEA+dvo9wAUCZ8y/OOgv0pBC4YPDI3uSw5BRkSsW9NXYgpg6L
X3zdSuocnyF891pBlBsQxvBQEmuCIXF80o9lq734kdQ+Z18A1sycoRf0jRODKzWNn4g7YKv8dRUO
To6Yk0sY0XmLiOxLc0/N04iwbFttxLlomPCgaEP/8OYZ1wRW+XNGUoT0uB4gcbpiElmXH+4TXVCC
Mi0kExoavLCj9uIagY8rjiq/zUdD5gpmE833PK/yOm7eTkr2okBUbAw/RAEFY91oBZo1zosEFWA+
+lw8PfHyZfMSifZl7RTYuRJWCCE94Bfs8CgDgzJUXhMHY3U4dVPfGp2yPXNyzyATmIDIM134QxTX
lBEfHn3ZjZDKzveLBlIBsjoAtSekLu5qHrUGgTnNpqfiMoQ77cHZ0wkkuTYrWUscm28y+K2Ej23t
lW+rxUlQ6fmJOLE6AbpUxgwXYtorBxsdfaDAGoSqjVdY9A0vZtOVuiHznXvQdjSQQ+5lIuXQe2Ad
HSehNwT0TssKynTSyfVVQO5ORDEA1pUqSwj6JrpqzLhpL1L7d1YI5syN7OrE0jvyLDRQ7hRX+GaS
UA/Zxuf6ps2wTz4HwhoxfUoQuMamfkTWf9tIgtmCztRrl7OgVeSz+FWS9s6y34D9a7epzGHSEXbe
bV9yKbsk9bH7Y+vckcrPSCrYVL79HVegmS1RIn/b34+lKhQTYk9H8/IkhNNV9cvI3Vf1GDO1TuW8
/NJjm6dlTkEyL4Ad35IiZeyk93Ug5SazH+ScXyyPRsP4itqllw1MxkhLzKYkTb0mbV4NUYn2AzAn
LbSRMVx7FXD2bFNMfd940304A5sx+RNrTQS0+xdRoCxcJ+0ewJSD2f/n9lWd8WK0eYT99xt9QY65
ehUP/ylOsI8ibbJ+wbTuf6krAxvrgn19MZfq9Wfc8HGMJ7gIz66DBdICNEnYvg4v3VSzq3HX7LY2
y6TsxCFuNLOWIglG5C99qpdyuA9RKs1kLAj5DSfikO6YYNa7kkJfnhzR6wj0uqgvYRdAX38F+6De
lzFSAhD9rW2JuKCUtr2P6MHhO1ym9EYzc491uYF+OGpjwwEXbu9GW42kOZFwsFblNnx8jC1sArO7
BxLlnqeJtRdLEnFiMrcdfMJHzQH+IR2FiYYuvG1o3LnVI+Is3PORYLqbisjpYW/YIZ3E3o86N9I6
yzijsb4aziqIDc9VK7ISvRgMDZRwLvlkS7Wme6kXGTvqRPoR3MS+vqVByNfvId27S378OyWff9vr
bDETnOTdC/64dawcI2KEluiMCHpMOizPruoikFRPQ2K8Qhz/RO4ZFUyY7I6c4klD3unx2apfsLrs
Z20bW5mYemNiGjinTyrnI528eiKDBS6BhjUyAFsj2lAD93dty696wjDZkE2s7ZI7vh6wRw6m2lt+
MIUvjGGVRT3nxx73WKTW7DDrJ1QWquQyDz1/5UbA1eW57eNUMNswrq1BAwB8NQtQQ8l2ADIvcS6z
j8ITTZICVhGcPa7OA5eu5nq4xp71Zg8wVlx4lS0lhXQvR5eQrPYh7ZmhmiPBZEk6KfnGUN+4qaaD
HVB37tZeb0nS9EncTgoPV5ViC5QdYZ0KL44BudRkVI4s1vZL6xGU1Pds8SrF6NjK/ULgi6QPwNJJ
XGCY1xqx4LQwG4eEp5IF5A2GhzyG+axIvDjXC+/iGI+7W4blIxQN0Mw2/U4Bi0NOLGlHCl5VTtuS
77AFJ8MbwOxbJ9zTXSpbj/v7Zy8WQEOGf+pB9Gn4AVuDJkSMiZil6btf9Xmy/Omh3ZC6+n36qm2x
v3kQNYHWLUxHHFpu1GPUSKFsvVgrJh3tNTwCp+QVp8CA2f8ZldpQpvlYl7jOBebWKTN9eyI5hX9f
GDL90mJW6Po2nHpuH0NoyD4b3ja4lnJVdzZOHZff54vPK7HpSUVaJBozRO2f7ibLeMoJeuMLj2EY
FmpXirzZ3w4u0V2bXsdSfk5eQ0Ih15c+Roc0QtsxCIm9geNMUoMKq6RVp5eoOB8QlPAhHNlgSP7I
zdNhEj3mT4SPAq4SaAlvXfVoAfar1arP15tCY9IZF6P52YOORkNkaLm0fcdAbVzKWkN3PYJ4e8I5
2dXy6/TvRgebgSasRTRzSij9HRJNfXP4mWsW3ABKEJPsTS0mCJ6QKJU4tydlPAzjAdrSvIb2csf/
t/6M1lKcKXQ2+2N0mYK4VU1e9PhwUz5CdmRmwgAGsNED/lMFld8tlXSg5wCbZx3SsuzLqV/tfyUi
E1ZUHTMxJJPltDlVB63xl17pSflvWC2jsp3k/ix2vg2aWPoALLBHwoyri3MhDB3TR6CuuwHyYsHu
7qdGLbh1i16fXTxQtTXgK9uOwwhVrBf84sPD90b5YBslm8pY1WHIgmntm+eaP4G/RQmQS/NaIIwi
/kCt+udvpzP4IhUtwve/8VhFFRNN7NRj7HpSVVnV+mdjAWruAsq7KOfX3R228lwnD+ZSPtalOAqf
BWxgGVV12cPAI93C79Muw2DIsqYzhVkQTaz55TIpnZ/+8iXuxCKIpAJz3sgC1jWpjZbC5b6LNVk+
zKir2Rkhpl1yIsdTtIGv91VWUl7/pcLM/pzoJfoEJwfyPW86wjU7QlJDGXzIOeHijRcccarnaMAF
6QhxWFtkKs/khy4Py33/yPKv7bAyjKAcDdkrziDPEhL8RvcGBXV5loolBjbVwKQn/LgL+GGIamGQ
XnvVuM7HEwZWc+oh91DRA/jwCORV5LOA5Ce3NktSyQyWWPmLm+j0f70YAYGPU/IM2F+q55iD099f
LNRqhCLfDcfV+U4ap2cV8+nflT21TB6g5h2xQPqbQTRYyS9t1+qq0aP5FTHRAc7lTrFKEPcGS/rH
Bx9txsz5z1akr8GGfINJYYdGzv5cKzDOamXX/7NHDPA+AaeULjIYkU8hMeUhXw/UdUOdEwToVwNs
3abDNJmHk/euUz7sfUG7kd+v2l3uZQnSUQpvcfuEN/XWkd96znM0HwfHylpxhdq/v04rml5u+6NK
jybNMEIJwh/lJcXbqn186tPbFw/YRPHyf/PJtfnGQjkPtlBOAwkztR9axSTXMtQR8xwrZcfNv3d2
+5kr5WKmcbheIlpsoGeBDvPSupxbwGIeJNEuMvX/3UC7UmrKNgbgQNzXSfJIGf9p9k0SDXzfAgAS
DdB/Bojs4RHwBntsrh3PTcp5viW8J3+FIkXzX/ZvKI9GyUhJB5MPkbHLb8IjemXE8Cmn1M3/JHXK
+T7KPWrkJ8o1hlB6gakqPJLWeMjKyOgmStOQHsre2QCu9pRz4KMj5BgjtDopSCE/xGn0l4fpABDz
fgJ+n8SpbPYrm4cMu4FZzl4CB3Z6UUm9p/gNOGOS/+asdS5VtCdk95C/2hVfPr4TlDcA23ue6Tn0
0F8yX50zVGjZHrtHMs5OY2cfbjQIyu+TcaUzVZF/sl7bkwa0uHj7NOB7hr6vDKfSTWP5wswQekBm
Gjw2bqnc7YHzWMoeLc3AWM1fLDcbnsmHl+YpJb4RzZpnwswcFA+tnqUjKZIso5yttJPETVfKzqDa
KGLqenrKJVXgyBepNByjIv8jP4j8G7yXjrn/hXvQLtVqcBQ054mAf5GlnrHLKUnqUjJKG42hAqqO
jGGCQ530nnk+cZjZSqG7IIAg3/+xu9KyIFwsqNyqD3JrS1DPI9AczkRVrdhKujwSrkIpSOAFwhhk
jybC5b/M3nIFgmmZWk35REpNjCLuDDqbTIOn6fIOEEnghu7sC0RvaQ8F2i0giYC+9TXhU2ENzJ2R
KqOxus1arWVhsUO/hlrOlp0SUkpBvK+TNpceoZ2NlKojBvO48enisejAuervgb4aASZDM5dkF74q
Bi8rUE3dW77fRNbT9Sggz2vHA/QfaveFtH0LakHovI7n5GYulCSiET+wwwMMCB3LtcUuuraBYUsz
xT2q0c1ACMYOM0n6Kc8A/3bRi4GbtKPLTOIqT3QpThZdubMs3QCMU2JcSpju1xnfJZK2A8UuzUM8
S2xqUFCF02R9pFqPoDsvS7EvLqzTF09wA688Ibw/QXtjWaKf/eXeEZcGKm112DWAxGyWoBb0Acwb
LCcST7DYkoQpyNNTkYzC84AcyX9/m+DOspxd8vXmgayZacmfV4EZLc2b7cV7G7y9bpspuL1IfxbZ
aCYRhdz8QGnUc46g+npad8i8sbJjcNZWtQoFltrYLweH00n7y5wvXplMvVRV6DJv4EcJtnx2GxiW
52xb1XOG82cyktvnJ/KHazqine17U7aPIa+ja6kQJFqs4FCxrmS1mapR5/lNkG3U5eS8PM8zgkwu
w6Ub9U6zsAdc2Z8G7Ptz8fVfHLMH48vkKRVFBFNgk4vy3h9PynSPb57T+74MbELNyYv843cy5lph
SYbaID+OYqQ/TCokZ+xcBwNkJ6y5bFJGX7dmzFx1AEG96ffhJsSjip7maiO6Pc8mO/Kxu11uaF0d
EebXKzyY9A+DeDlFgcOZNE0k2Xk/eV8F3xjaZWJDSVLL5VHYHNNincgOYd2JiYDhupaOgy4fIp6j
sH5WzXO/MCtAusyEMAfgiMGmFiXluUOZAsrTi/248RWr2lENfR/3k2ZugSq2mMeqO9IMMIjx99j6
5HY7DBowTQa7tsGFhYCqexEy+320lhBQNvCel7OkNtj3fyZzCLUUCTG6ZiJEoDBPcUnOPapTfLTe
ivW2rCRyXrdNR/nVCfCMnQIgKdjqBr+6O4IPngTyLZYH+d3mx3nJYW/jlYdAQ3mluzkU+3ND6ewQ
7fhi6QLyF8uNPevghxIpdtYGPBoWSka2Ddf+a8e1JVzxYJnqdRKVPthTyalDHFP1+HawQ5SUNn60
oLOzVCmBsrrajWeE7C6zJG9Fd0pAtVGQbMgS8bTw8gXAPjUGnHrL8qqPSUaLrYZinQZ5lx9Zd759
jHVvCZMKMzBXCSqEGIj0i4Cw0vS4GVTp+LHNV9BgKtFRH+zCgaKvupm72upOtmGmM4ZuXAB4P987
3NETSZhYr/umNg+6fY+MBcFGwBJm3K3drqNGX3OQzvgicp5Vkljmha+F9gk7X8cBdcUfChDnJ/vQ
O3VNQaaXw4igT5ip3NoY7jj2bOkk8fPXLVCNGzl4D8rRNmZ1M7FXCI44LOMzxAVMW0hfV7IHhIi7
z3lUQFw5OrtYSr0xtY+AUmD2/QNADyqEJ1A2ZJfTxMZOaj9GvNGF15vNFntXuDCWsIfxUPgaRA0V
rYVqduvwDkdPAOcPkYsr9rfMC3BXU+YdAWZOk2nsO6mTahgA7eY/gtEvhyHFRcg8mdpciYcsQxQF
BeDLmBdyabZ6k1S0JoT+GcI6C59xHZprdeAxWbh7DfuTLRMmVpKxXNTZgxiM7lF633WZA7XopLR/
0itykLXLrcWQd5L1fdJI3Gcq++vuvOw7oHvOYlGQNdh6reqAKdni+6HRoMDxPzH49WlSh1NvXCae
vxrgTLSG8neaXJMHSKYqxnmDimO/E+ekJy+uHvsRe5GbTym5RhlRckzydgyquXmGK1NVx77acqGt
bV/3ho7HwyMt3jh+6Szbndf4wx7ymAcHYO7vQmzfYae4VaFSwecxuQ+zfodU2DQ+jyPzDqgnbMTP
89I3QdT6kDYVz3RNyxSF9L3hfDcFLm6m/LOpuGTwlyI9aj5ME/NFwFbpLnjFHQIBZflYc78SVRGe
1f2aoPtoeXqeFyDt0wP49WImBEauaw8vA93xnIqS6vtLwzez+6PO0NlE7gMLGdHgoRa5EyevmfK1
pDac6NxSbQyvNguLu2Usnno1ubP6WEXX21f5Q3maV00n7ogDtwUAoKWXC/F0rUNqK9NaFydye9Jn
fdrT+3nTF2kOrQsd8pa9MGxzySTCdXTJZQz2IXwNhmLNslgtA3FmveE4/pSgFCsEePFRYpIad+BX
Hm3V8APLGTHCVr0zdVXrPsa7M+6vfsn0sykMKVqlCxwSMSX3bMvnNiGTysmANs48TW0Gm+ft4EUm
V0Dn7pAVejX1/8sSSLTkrmJ4N+jIl6YTNb+9WtOFszjdTOZpm5+EfFq5CQGdGwkMRqOKt7gu1LTn
f+grIyxHGsOqNaqcVROW2S19o6LAi/pOUAD02LO0VX4h7qTAV351SyY7TQWj7ZvhfkibHJ8ZGdWV
1XhrsNnynWIp2cHMjofcEwDepC8gy/Z5Z4Zj7iLAImqGCfpgHPItIKsa+KhWrX1yx8XrR2TEXZVz
E/PrnwleF8c6YptGYALpwXsQg3UaHHvUYg8ZXjrh0JDSsa0mREEHedZdTdPaUkeukHP1ToFKzhp2
pJZJrEb360NEPCOWbL5I1AFEaGoOZtiOSXHiUNnRndbK6RYKzTRzs4r5YW88s+DSrOALwQ9jcjqo
ptuC4211X9DZs8NlkfckqwM3rdnvEfOWucs3/GnfeDF7iTiNA/UjUiQe4PxCEVHAiuwwBph9Zx2k
+beE1wJ8DFuKmF1AOCckqQhJFvhkll3Aj1mMOLxy/fduKQrPF7+jWhgg73+A8KtoDe5rSaVU+KZ3
4HnPwOYkD5TZo1jAZFttOxFjZPdfMpYuXHGDX4Zl4KNxVGRldAVZdodmSCyNYgmM+6TkJnxKg4O1
aEFLdKue7syI2DLHTxhIlJxutOqEmmYOc9i4xRdm9yENf+eIX8TvhGTqHyWybx3mPvzf4djSgst+
kQWXBpr1wjJnXrMmYhyG9r9MogICojWomYotzHH1eITIkKAgvByWM9y+EbfBpwf2HlGNR8yzpGN8
7r92BTyZoYucRphRfxkc+rPFIu9FmWMHZ1QL7m7JnsMbhU9gOvKrLa9tGnO3XmfcMzxN2VgiC3V1
izMTc+OSq9lBnWKj0AKjpX9C5HBXa/W+RO/h6M3ByYUNhLAR2/J8KKRLT/5s1XsDXDBHWGJHIcEn
8fStMg4Jnosx2aCc+D2sQts+gV/x1cbafz4c/NLqABuvi7Wt7A2VT/qdfzuN2MVr9pZzy3kLiZju
cCsSCsj3jHcJSe4i6HSZPqXQb+hfiubJM7UYK5PZL/kyXFZDX+oCL4ttMSj7KR8hO9NQNOp8t4Xy
PJ9HeLDpBsOFR+qKy3TEb7B6BBXQ+6c1eAPx2JHymM2QSGT6AowtaJWD/kZL6Jns8z+7kwExNRZF
7rEd42IyKcZCwM/NCRshheWrV5JUaBs5GNqikA+Y5QWxHmDO0lpv2I9YrxQEM5x/grh9c76nnUxL
gLZph6HC2tzEKVQu6mqOs8/q/QyvI1+xD+V3XCjnHXzY6nCBBvnYDRk3i73DSECxLni0SldA/Hpo
Gzkkm3HhUdFuzeI48lyK8q1a6p9fcry2YlR1wcqIAP67J2rVX710mR5CtZy8UA8oX8iRCBUcCwJV
dqBER8m1XVMUAkRWZrIaRBTc0nKKUCgzLJIDybPe37uD0ZZz02iZg5hgDPxdHZ7a/GoNXNmhib3+
H3tgIkfhrx/rjND923eexb/X/d39vnhFN+tRKaieQNbplfCFzZXnD/5LRMJh6pUqmdnaQflfPunA
mCU0bLD1ZVywUFjv6O8wQJwqXUvDhtfgLHfrWHUN/Pje/9rN8FagIZsBzGCL5HR5Kbzhhspo/nga
Sy+D0+kHng1bX/UYNYrwkWSBuz1srTA8RQmU/KDw6M6E/L7Ox35jN7sL5qaCL5fB2QTyj70HcDP7
7JGlT6teaJ+qGit9OC5eE5xE20mGKkhaS54ZrZ41RglKHl67lmCO+UjPxvJFwc+tnx+l2Wl3WXQQ
AxPEZPNu1WIOf+FddSXgdbLNZ7AblKCzZ3pkD7GRgeqmvI2pk0PLKOmN3pnvcG3DWPj/nJhWlhzE
HGyAIYkQRJZ4Jqf7g+VMALyiYP0jCFAw3seh+q+6auUE2QDvzhWVgvZrey43QbAz9cH/YGg3pjmT
03izhrs0w1oUNXuOiGjqW+OHsCGT82y+PscqfPw4sfuv8rb01CpeUYu8f80yvMW0f3oWMTN9AJVh
ZTJLNg73+RYvSoRuWLxdWHpekF9Jr/6TPIyp3WA6KNTzNUx6ie2fRiOjYMbyevPbrRzqz+iWsCyq
Z4/sZuAxT+LbQCikrnxDSVyfT2+cBA+yYf9WO/BX1ks/DaILJBrMUfe0REcg5SgiE4+GB54cslNg
Qvov/vnGiObbyyh54p2MGieYa8sytJWxovAu5Ii3WwppextNARZZEWutp2IWgfdFDZibAf8QaPUV
JHMpTbAwg0dJfAmyNyp/zu2/tKBZXQqqSA8JLlNWM/BHpTce480y5cES1VVkWYluRGYCJxpG8/tY
BblmMMPPUIqSe4TuozTZxgtROZY4GB50Pyj65JMR01mZCDyffb1iU/MClA26N4ryDiUWB/qQ41Xy
vujMeHpesXPnh/actg6Il8UuE93nE27edmc/GnSdJfkMIWK5caUE7/lJzrqv16qOJwYK66J4d/zK
2i9S0vTP0yh3bIXKFJnmt7QuasP8/1HJ5O2QUVr5RhL/qXAl9rbXHl9Lcg6DLYX5lyAs7FCNkXLO
vd6C56JSEu3R22Wv3211kSqC8Fuk8gj20kJcLeTySGYx2CqeIREuDnkRL/pjy9o9kfx51YN7F1bM
eW/E89l/08QNmXzhqD4jhwnsKlNe+I4smrpH/Xjr9mhLasGnu1Y2q6n+u76urV6FXXt1eb3V8/tX
6ZYve9XOf7CPn8puNkiooDbldgpmHSF9rFn6W96ONI4My4Tf2D72P/q0lVv3qWa8rzpnW+La5nJs
F9/w8NiUyTQXZX47BIugikx9UGgm7plMaHzT+uP4kll7TOQgWlNbuPXeAJIaj8byRBMeEY8qVX4X
1AmeS8YKypAWETv7uXpqkzO9H1/y6TkXz66ZSSxQ/wPDZIHvGo29c4xJOqRE/6V0eVVC5Ke8R2Js
ZCyggfGnq6+28T4wuWnE5d8vtFDvCn7AHiTVaZ23cV+pBOfucPtXbpsA4PryeOAITZHSEcensBZp
rBR62yVj55dSJvU60Pn+09v+LcikbVdL0wb7owkEWk4bQR+GCWWqyEcascgEA6UzOv/UjMXce26L
F7Rs3r7z0CndnCiSYCJgS39ynUF0Rd0UpSBxFbVkhL7Irnrq1KfrNywS9C//cfK1wOhwA4gvoneT
3dAIOooOVWGaQOpNc3ZPW4eS54SNpN37YeoGO/6zprvRSvcrm4oyDX6cn0VswFbSHSJdCesLAKnL
zbgTOg4rqS2FjBuVtSGsSALgjvd4L/WJzFGY1/VzLNtoSricVGsRWXHcYBo35YC++ZUWgILBFMTz
e7y09yDprUXVLD203+w/VQ1cjcNhneh0t/Z9QwNMn28DZM+59Y3h0902PpFhsB4YyiME324CwyEO
b96n4rx8Z96zs3FQARcZ9L4MLFOrkKWqZX8LiIlsVVzNx8cOspF7SEZ7tqxggNRu/OtIxdecBfWm
jWoqvmrFsqRjc6w0AD2OKth977Lr1vkMymdxxUayRnSimLYppO8Wp5Uy444K9HiLOKJKwA/hmfab
QVtlwzEaOc7psIy9/kuX3NL4nHV65e0FMY2DIyo+EP8yhgFmGOGOeC3Fer2oHSjDhuC+Bl7cESUu
p+uz5wkWBAH5soBUfvaGXi0GCDvH0Y1iSD7gszBVSCkSrMSAfBcjar4ydyEn21ra+DHerg/zNqOC
SBkWPL8q5zBEDvdKWH8SxBJJ90gprNx0sMJjL4PH0+HdjZkGY2vkh6Yr/xUu/vNsz+RdCw7U2wGl
DLJNeoKVXK5oH2vq4+2pWVbqhXSaDc0qo87WC31d+j4Ymip0L9MrFK1bl8TEhlaO60GS2f5zHK6S
oCXWjR5VfWXxDxkojmz7PN//eKxfqdJ4T1fDNItLBs9/6VdrMALp+uQc5/wCWxZ3XSa0Vb0ODj8U
zd+/yIu8m//PfIiA61aCL42rH5JWbI7WBSK77fKVcXslWluSJ3WXroekHnyj7LH3kenaD2aSBMvO
Y2zfv3CmzXmyERLvrfyrLWk4xkScUEjsCgXy+a0Bp8loL98ObxzjZZFFW676NsI5VsmB2B4R8IEa
SKYGh7miMKbbANh4uhv2TY7icQyc9V6DGx8B91Tpz8Puw1vkrmE+KZlVdzrV03fteZAFdpIbAYTR
heH4K9hy3yjt9ac8OfJPYbU6qh5cyoY8Z53BYOEa6ZcgpCpb001aw2LGCXLA5rFfxcmZ1E8xp2rY
131zFk+Uv18HAYkrBMNjA6v6s+n3NIQX7l8QcVh9YN8M1pL4HRIicM+3QwH4b9sTqs8KN7msdvvK
4HR4NQvAshWOF8erQFWQ47YoIc0T32BJ2JSpMFJjyM8qtc7VF1Ycz2M0bAib4NnQ1M6tIu8g34e+
R+snFSaVRvhrlHedCB4pmb88S4t+GZuG8MdO+lVwaQIyNoZMbdQPi+gyBmAweNLojbT8MA+9S8b/
QHLpd9+ITzQFG+/cBZxPyJvxKN1mZ9210VkdmvwlP6KbCN8nNCi3rkxwUCwxqNxbE/T3H0NjeFnF
wEAeKGOpHrE3091mc/BT6zIr/vra7lMxWFWwPUcx+Juxg2DN02pArgYV/iw66kON107elLbsLmaa
W1q8tNl81D/Un4/lTi+1oLIiC/yZFyjcpHZT8V4tORyEmDU4ubI0Y0w1E3vdKH8U7E4VSMWYXzqP
4k8NuoQIGOjFepB0VxEGMhLQdahOU2TxGo6Z9/6EMm6C8uklLPDa18jVf1eceODhNb161Mcpyplp
7fGq4e7KH0Hy5ateg5D+6Kt1ZMGz61IQSBa/RBzC+pySPhKQG8Pl1gtbK3oZN2EhmUNTDK9QXa+r
HUF3Pqhefq7R+4eBA0LHVU3JqQUOxsK2mPhH2haDwiJlX0nrXQS1B7kIrAFPT6H/VonEF6LdwVje
FNBNbXgZU+r/4mDm2vHETdlBNvq9LtdC4pwiVJK7A9wB8BlP8AWkmnwpKs9yddmJtm0Q4Nq9Fm/f
TwsI/n/t9hJP6DP4mjdx/XWAibzU3nyd2YTcS0ZRMADpSx6S462d1AMaldB2CM0SxqYrFYdXYyVb
JzTfrx+By19WNOAl4KAP9XhIG8kYJo04qh3bwsHK1f7L/EzpJjoG4vJVuoa01WaoLbclxXj8ITE9
iH05owguGOd39TJlmthxtiROh+/WJCDtYgkP3ulUrgUHlxC+2onn2IaNJfmIg2iHrJH3LF+mJfPf
OQAX3eCElINrNQNvphb65TmUPmdhfVD4UKZXL18wgNxFt/EUbpPhT2mYw13OORZm3nivSDuZGX+N
HPGSv2fkCC78nY4+ZdV3N3BpohY2UhnlKEq3CQGji/DfmqbM9w3chM6W+KQahZSN7aS9HmgyH8aK
jVhB3eiWhAmKzyqObQtFzbvPgOFiuylVIWtuAqqcptjCXbo4YxJzbnvYtnbahDcRqMbXxRLqsKfK
qKWhAkRbMoWGmTAiu5u2N+Fi0Ui7hKXqPbJAedRrSs9RHMn4m8kv1Qrun403Yq6n905PoCY9obGW
cRuIG/uNMMIGcreZ3BzK3//tApGAu+RtKQoPR4HtazGbbTRZ7DmrumgA6ErAGUKnIJGv7wUzbIB6
lSbQ+VornIfRwvui52G+zNqyscRtD50zg4+rp/w+8sU51H0XtXly665LuyYHnK8OI7HSxuj2Hitz
Z4ffo/Nh7oVKVVKTnzzxUact3Ve5GHZ0fxchX6Ark/c0s1a7gID1Wiw3RckBroU/ULA2F/4xBPN0
TM5g446HOILqVGCm8rp8rhk2WTC/LtTGQw3Ihkag/uW6zCrMEL5/Q7AQaCM9qyiWuacLFTK5MN7I
Be0nYndyEmVYB4t2DWimjWPCSdHFlC89Vy9C8uwrGVngFuCxjBp1b027n0st2F2W+A1DyJVMYM6t
EnQ5/VskLnG2hwUOB0oMGDgjYLOqBegGAGXSry2ZYm90mDKIeAZT3x8n0PhCdN2o2KORbh1E5dxn
5N/rjVfAlFSYuO0dBuKlWLRf6a6oYA0IqWc5LmnyMH+j4PBhf7ZLoUQXB32JtodTWAKoHk8YCoyo
EiX9TR44u7cA/vKsXSNFUqhLtIW4WTisA3N06UrPa4sRueZbgzGhYTAmwTGgHgL2VQfVjME1Cjy8
CntqIllU2Pi26sMArn5txtP6QOsExSUmRiaGPMcUDnfBfK/eEK0hTFS14Gv2STk61puy/Q85EFSo
RCxwERSP4DC55tWo+u/+q9g1apZ/KG+rtCEfy6urr8ga6neh3aZNxl90Tm0qaIyjPThmlxZK0XE9
2rVq7FfsPyAd9yj3u4AQ94IJOJE3uzlxzTEuob94eUwzIvjrF/+qPYPNaJQx63nKmRAzyamXAbSG
xXqOyPOoFksU3B4sDBSWz2754KnfbSAZpSZzgHwGt88nsIe2T5O1O6zbB6HFSnIbytOmNDvH9vkW
s7Ga3Ql3hqCnMiZyKGpgZRe4L4UGKLlzbmysJFpdLESOSveAXWYjAmdwZ3UW15V11Ujr+W3EOzu7
jpk7CT9y05r039x5dDOJ3IuNal944PnbnR3DPk5RfoKnVTEhPeawUi23Wj1FlNMV23ciyuWH5hrH
d8CHGX6EPwtGEcMjKknLqvovt3T85OpBtcGycCcnVHhlHi/GsODXcSOQj7WjgLPzykDCDHBnwNHS
W2p65IzYQAPlb6fbYLepJw3A1hg1f6chwXHSbxLEzkbPdpTPTiT9ut86QY6c9+5T2dhj7Ujvh12U
flYvBWDjm74R7aEWEchYtWYoZOqysmlJpbjzS6xwDxrciVKlRQ578pDVsVpAmTPDzpRQidoqbX/C
aLiKd++aysh6gs9ShJMoyuFBPBmi1pZXzzUupBqXX1Nt7MY4Cn6xatj0asGci4+NJJvwxHLhuGnS
LJtczprmX2z+MkpIW3RxfxCxnPIDyIWwaZ+LYy6dO29NkVUDrrgGK/JtC2DdZ6Hqv6RmEtMVi/V1
ht+GMgUD+241R6FaEoOZJuOEoQuvCvVxtK2TGV5LgSuJus9jz3v+88kJBAoh9Wt/DGY2XuUxKF6h
303sq6wtaI/9UwZAUwP58LQtXzTrFpvfZwLC95FVxVnZSqmstNqOEtCJBgyT+fdUjPdsnmMXXrhS
vZNruMrbRQaJjqu9gq1f2IQOG5e7yTKrAsLEQafFGOjohsd6treogshS0QH43DF18yb78UBewk+/
3FDYI3O3Rk+DgK/YZl4cXkhnpw13wmQxlf9PDz4WNGz0EVYmJz8pGUdN77xZN3OKYR/eQBMjPA0t
Vt6bMjIq1ZmAiirU5FoAirygtRVNMPSXg6aoja3q6pDNnKq2BLYkZ4ZDSo9N4KXYVsPqNISxrYRW
G1TzBRi0+0heY+fBA+n9qFpz7OppgllLuKImiNJnYKJPZPBqjesHZtpGDfVQXrBmuPFdkxaYb6oK
1v2UEaP3JUFWch/pO5yttroaZlQL2yVID27gDJ0gcUQxmv4rg8p4SSvC++COm98KL0GDvcGNLgwN
rCwj6B62V/iaqlBPWMY732YIfC7elvN310BB6A5ivRM1xH8pkALehh92koHbv+9gwlGmRYqqSrws
x0KBxwTFg1LFsK5RlmaceXwWSG2AICabX+N0gsT5huEqrRYgFCu17jCT8oQCay/RN4p2Qe6uGI4/
1OHNPC9YpQ7mjeVaW9dHs4pVfLL3SofqalCSbbBYPLU6DuqOBzyNKPp/C5I/VpeRXqqJqU6DkmRo
BNz4TrOiRYT2BNsPFbzi2MAGQvZzzs+CSVmlSGzcsC6nfs1614R91rQW+xuUKhOtJkBZIx0fCgqG
rhG5klBTMgWRdhwj2SWt3pACeKAsMD0y/UEclVNQaSBUga+VH2Lp51bkdjx0/vvOyQItXjQjZuky
cii6WW6SGD5aKfiPSX0JgMEKjYi8dQgYJu3WVf7APBimhy3RWQtsA5UjbDZBlyiCbFZSsTrGzSa0
NCWXS03hxfXwZy+4L8NENSYKv+5yExUVatSytG0HT8/81UnL1oSq4KskgG05PZ2FKYz0di8ZsAw0
Pn9mbUzJ1njdQL7wsYuwJo+aI9f7lgX4cyfstXs6WegEGP6dAb58+jv0smqsfTZ5OyXeJN59Dyfu
2LiWGnI4Q2w5wfZMNi8hRYpPPNLc4UMt4ZkJ4HfKLa1VfBSl/fmNrRtlwykWrg1+hWL0g1TDyO+A
Bo2UsvL4pZHY5Ji9hoRRnZiGGnn+fE1iiQcilIwptkuXsbTzGlvk4+vpx9jGoKGxCMqJhRriba3M
2ER/rMqGFT+YhAuHhJae6XqvB3A/4YyHRRARBfcUlew/M7KAcRJqUK2hkCyIUTComkUSiV5/M3ht
zefO0MB3zgAuU2V891VC1P8mP6du0+MKMg/Gl6gp2hpsNJCJa9UOYgPAqxyeFn3tVtuli5XqOPRm
Ir28FSb62bBhBAkrWZYzumok9o3WZ2WWFx9xA3BjJHxl+XC3aOr9rqIFxMXf1k4nEfXn4H7cps3O
cMmUYbWDvcIL6YfznEywzCYUj6FSsVKKg923ll6LXN4iM/Dz6Dfv9WuYW9Xph7wyQYYdFUvJXae4
ynEPMBNlQpFV/3ADoRfpPLsTwSOmowDkyGUw02yT0zA5o2YzVa8qoZoHdyhY9NeWzkJf91xQajFj
64oWcIlCwX2ppqWYVLPLF9PC3PEeNgPcR1asEu4zU7x2UFgYeIR5BDAfXNFDFkLkbQ56Ra/53tua
4v0UgAUqEhGRB8uQqLMPmiN1AkgsSVvQDzU0wJPyk8lZO3eZEKvt5OmYoSZDJdd8G67pzgfWLbDR
JGLnw3aiZUtMwWtmsh4Sp2QzO7Ilm/kz2qj9OW9aLFXrImZi6brWkwcRbOUEL22myJBcGgJX0DYR
tc/tvTltcfu+FA03qSqvN0Uxp1R6VvywCLe6IiPxTE9gWs12qkoGYHvCKSq7AlbbmlIRFbTqRxxF
dd4fj2mf8vDNGmQzvpcrkIE8BvB7vbwWQtRmAVg1oNU6DGqI3I8LAlGKJLTpbh3yaHYSkUiThJXV
qd/NcCxcBQK+lC487cHi2JL8hcEoSiJyX6XzoogH+SiUbFF/lbPYvywzctDxmo7VR0oo+Ht1FzwD
WZkolkemkjA0kmcqi4dwJmrWVK/rFSY2XhV5q6uE5BO9Fgaw09/O8D5RrUvZTqJEVCEB+cDI5mOs
RXg8RnhIqGF+pQo1z31H3onH6k9hq9EWehEREQx1CR/4+4FTQq2UW86dosh7P6F3SIaZfn5q2e7I
Iu0CLLpTOlIJUBV5fTwtq/wDu74YThv64Wh92tYY3ZM3m0d80xRiWqjrFLs+RJ+OCLT1UgT/CkoH
fv9JwZzraMb8YYeYbefC60wKKdKtMAXlULCr7zx9Wiv0y2zGo7HEuZ0ER3Cy75juqOF12JTJYry3
MFkp9OrFfss6WprrvssnziGnPDIHSKESEAwvgiVM9ncr74YxRdy7PZDY6Z5XyEU3K3OR66kAM8/B
56jdBf17RmqUfnrmaK33CLfNrrIv8huMb1CsHZe9AOoD2EL3Dq/NQO2Hlq2NntjwAoslZW1oS6CH
MBCB2FzfIfxp4cYcbPntmsSUe9VsN3SJgVLcMIycbuVkFoX7vYvHLeLgek+Za68xyr/F3MNdxcfD
hKk+UAAg1+m4i+R+KSJ/1kct7AWOTS1K48/Zdq765vLwloc+oGBI6DWXS7hfKvA+L4X8zALv+gGh
hn0E7uXndMzSpTsdB2k29cc/k3OpykqsY8jPI3VUypEAOPm//VP7daakCb5o1uI3cwafj6LydSiU
5cIDTEDTNRPvFVnoQ2kDSFpd/uu6MYfBYTJSF0/E5atFw5u7fneJnBCcKF44msqAJQmZeZqh/RnH
Z8sP99NtgFNC3glp7+tdTE11j7BcVh/tVQrw1CXTFBB6JNCYXCIOAVxCJL3Jjus7lDbt/zo9/f3o
SjvI+rHSCdHWDYX2Q9CvPndSECmdKNneJ2FC8TM2JsTiNHc9enW4Yiz4FR45zeyToo6IQdFKtgjL
GkSRKrRQsmI+w2cuk+LafwQuTaGbSet3wvUCzsLQ7DzCCcXgkvumZtde0YfoczIJ8vRdcDV4OyuJ
h9iKTu5NkbMEQhefteDtKNt7u4+56yXJcS+cfHy2qUQQ30Bz8MNhfoSSaw8t8LkB54XHDBVKLKDI
kLu2ZTL+6vJ+X2e2Qq2UOnzPgZQu9FXL8MCm+23sNvIeupMpGka49nKcE56E/df+hN1tasfpAYBL
sUJcEld/jUdlNx7btM5b1fTY02vG2vbfKoUXC9oONQ9gsJZOvpP9aED5j4E7JdjrMP69pbAYvc6J
BOcU2xByHPD/8RfDXNf7QcfWwAOGXDinmgwE2uX0/CqDwuq6X4Q8GhLqIL7hLkvHeNj80HoxE8A4
xrL6k7Z1+1hF1zO65Npq1UN22Ab+kLv23GR6wulwBI2hER2OawzOgOrpHwzI6fGAyHH45SLA+NgJ
7PzIUYhnV/3/2Gl0awifw/l1R2oAI7IWUMK++bjoekMGJG8J1iXP5in3RqwVXyrRtwZTx7zDA+YM
t8xK4BXs64TWQ0JA7fMuwZ7egqUUrC4mG6CwZ2GhuRdGj1vRwnKQv5hHNZI5Qv30qN18ic0UaD0T
40TNXu9TQiymHlPJlYgj47aw5PVzIWNL+o58AFEtrt942ZNhP8Q2U3Fh0S/UmFY9zAtMxf3WQl0N
ctx3E6S6nSAzfnXv3C55lhjvNkLGZjfwqTcG3y3DCCP3xuEmgCXGTuS9aEiHUyx0D/hp5cfidW8D
1lai3XOx43mGjezvVDzpHm19hBZ0MtgyZ34DcEd3/YKzIegWQSTkkA9FBzR/cQPWQjYcUlaAOaFM
mFmH2d2Dfqje14wYP1ALePlwYb1BkecKsNH7WsKMEZJPALdbrqJjcijBzIiJK3OUwgXimODRRTOc
JUw17yy1VqZ42o7WG8VeqvElBrOPe6PAFSwBJ18SHqW4ENWN3yD2ms66FdCSFYqZeUc9YEBy5x2E
4+idkJihTAzpW/JhQrHd3g3O5NTps7yS1m8hYDsG6sGBfwGLE/UhRECsUSGbmy1/ulQ6RQC8B+cs
l/325Bp0icTLSym56LPBRU0sStqH6hq48OxErALT2C8ECPTOAOTsyT3OZ+cg1TPA3nH81BpaoUdM
lMuXAK4eSu4yb/6GrBlpTzAAlZe6R1uMKMWntduXXWeOmnPfa8k0ZIaYW4eWWNdqnihd625GShE5
zlsGqwUCKa41QUK4GfULggipx49WOu0d/dZwvNXsvnqHeRGfglFo1tyaW/MYFfQKjdDu/8bpSJ/C
Sb9hwFmyHqJIQJET9IGHOnxfsjyRB6DVO2yaitmEA/g4+Tfs9ycC/eH1+S3H5UAs5lpKcm26Hxcu
76INiZx0dRX0aNft2pXy120iUjyjZffdHooQ9OfZlZmwXigMc/BqkzvH4hquKEVv8A85dzrmYb3Y
A62qN/rJ9RMSbz52vo8W80i8i/foU15x6JIxR3hHXaIgsDTG2D/8OSYGK/Y6BhWg0qP2gjD17+iV
ER2p9kpmaeKLvyQRNRuQfgB2+kuOKh56A20q0RN8EKz6+nxXEPqYSXJZnzQuNzeK6l1ZraWCvHZ9
Rw6N9w1WVf+ktiewDkB4qX4KKHjk32kNbce+9GS5VpgFpkB+ulDg8+SEbWGA740vOOj+Mt7VOdeK
DrR75eHrcoCt4e0eeVaR/SIKsJP7xs3Ayx63hr51qcwbvqAAKgUWUqiI3dMHHeyo1a/y0kGLjcC4
x2XrBw1gSKqhDMiGG7NFcsmj129Z88Y87Ueonc4GoufKn+BVdLdg+yvMLA9BCjHRPk1D3b7N3tv0
rgFyCnBbkf8NTI2mLi+LeDrIosa57Rj4qfw3BTZ9ih7VwPssrkY70cH5asDrC1gDy+qPQGiRIWc9
y9VJ6z1IYWCUSHQIJWS2Zdc55YHT2V5UWnNoDVPC1j1yVhIXKQ37WPcZldoTC0HBNUX4YYMWhkEU
54PucQ35ESy2mfVeWknmGmdImTKclqmpKuzJC4IryGDQEDz4YrEuz4QH02RNDl4GpqQFteGiifmp
e8kX3Z5j2MhdRYwnqoisimfa8HDtPFue4uSzKSHlJXjYH4F2Yf/Ur7n9xT7fPu4nhSsToHo2KjkL
0iMhRY5uZDZ935evbTQEIbyl7IEMHgZQlgofW8nAKaANcnb02uSHv6JiL29E9VahMlDSurrtm3zy
NmdhhF5fiZ67jNc1gfASg+jVWBA86YZRhZo++uke6XzL7vpdpTd1GScJ8mVT0BdxSTPjCTeEnVIM
mf9O5Ces7jvA4tsVAs3SptAhDjLjVw+oNMvaHtHBjvSE6ROFy/g2K7oXlSfEM8lwaZnmshqzOQjT
wReo5hxdVt7neiD8dSXSf3BzBedCcY376dlGHEroP/mQ2tHstKahfYeCZqVjrHvSh4cID0puL12U
tQdA9PzPVE2vYZj/sGlvaSfSZGAjLhYf+Vw0YaTbtKx9AjDrPNnAdAXZH0ER4nS9omKSLc+ixg+l
9ddjff1PRj68Zti82EZAlGbNIAN69VGZR10wcmB/I1Phu4OZxlTHgm5PudtcQWHr5MZhOQrWtfCx
Xn6j0dVsqgPtrZnqpy3PR6VcHh8Ne7kBsoo9ERrFInhMQj8nCjezI0QHka94o7xTPwVm2ph0OAQT
/qQzwv0a/AzQ+m9DvKigk+YNKSCAbZK9BNLbW1NRnq8056QvsU3Lyp54WZ+s2snMvHw8Dx4o4A0o
Da9Bowchf6+U7UdLJeewgeSdUyrvCDfUM9spjfPt/ooaMu79/nfwPjltICB+rTeG9GeNU6uJ4eZv
dlWUta119En/25SPIatNgbcAcJVzm8bDvh4meFm9h+8WRzPU+KyZkpBSccu5hzbvM5U6h30IE4r5
CWnbjrdLAZ2KH/NPRS6hK+GwyjvKJ95qudfymazKUw7/ewObe7d0HS6RWsgvvxnGB8tp+gCTb7wC
wrgRyZvmdc6dc7Ap6DvorEPq88MG8N9WYO8uMdNAjvC3GriOc4vvMPtbeKotfY01CXXBMVBOOOSn
zo7GsSzqMD5wmML3WN9RJDkT+pqKGKYIcW+JiSUC4phORqaeCPLLB/CpXaPEPPGg6mu7Mp1608Uq
GS806E0Q5YevWBMEqbK+aMW6gbtV2QGOv/uSneBrLOgxaSZOosMpmneDH36M7fS6ZRkg0nnqDdfS
m5RbRZVvrcNO+WjY6UG5rXbzJjv+c623X7Sq0sb9nur7KhG5VWundIyN7eNB2Q1J2V0V5LhHb8J2
o5CUcMimbq90Ddfp6eVurSEqZm6PZhda2D9Lcq5P2BO6ZRZtKmWovYGEa7uOIJYfu3+1niiTrb0k
3AArmqKUH1TYmORkPGuQlHVrMUVCot9OhcFSNowISl9XuKUVsz/cucwudu3YcMT5HmzX5LyJsbPA
X/QZazH77mC5tsHl3pwks/0gf0tYWG9cwcAsvhaBJ5J59kuA5xmKCeiEKv0hMrSdm4kAFP1XmzTQ
nrtEgSKMqgG6Np1mszhtfwV4bJjzdxXbH0vFExQiahktxCZYR1fzZ5Ap38EoIIzrG2+D3rF8f2yG
fCdSM8uRhwNekVEIxx5gfjJzL7khnDf3loeHNm4sqytlHqu433/uOPIXosetGjn/smPuYsHCYCPI
9R5Rb5S7GI7ArOrgJuBgNhQNuljxQH3QMettnC3EavNY6MtsvhgnxKBkIvI0+f17+MeHAFPN0rGn
ucMoZdlQEhAY/Yf8ThWRAtpj02yfwirBpiUsWN3yqBWBsbGqokeDTR437F18YWBbPcHTYGL8L4CM
s06zcPGQyYgSk5zT0/TSWGjoN9Ll0ur6sWjG89Ot76o7oCf/6kYIw2xMwKUhoZeybKyttuIRez7u
ULZSjWOskbp5Z179368NZ9Tcmi6k81mcP1T4ESz2ppjAE5QsN2uoTNyzmTSicSnOtwSe+acL37dv
KEQ6KvNW1EUrC68FpfddSMc98PJUV8etKPQLDw7jXF+ziQCe5An7tbtQhWcugIruxnx5zCc/8juo
wEYmh3HDf8zYV/JS8L4OOSH7XEFMonqqylLvIRfH9BpcR877DgeIHGb/ebVmPkmBiPDRCXwy0bcx
ogTu3YFH3O6CZbQBoqnX/8ctNFSTbwk7N7iVdl8hCAPnFOrOnV69TYq37oG+OktVhHCX/gsdoU2q
8lkdVbG3xSkkrmGKDyjofWe7+kVXZPydeojL65x8iZ1+TEFoN3GQUeTI/XHToRqa2es/4EBvRSXa
suAswbTy0wts3B+1wR9nCq/KUrX7t6pBOA8hfWiFdzKS6ER6peNRFEhqB+KJfA6IY8Ks4giYa3GI
c7lZB1gwGaTy5wAp6XEwVqAs5epkfW4fjy++ASsnC1dgAPjgKBibb/3N7F3miQ+E+opHiqGfmurS
Npj+1fhXwGDcw3LMoGcSCsQC9vK4ANVq/I+ZovCWTzNf7/BgPscxGS6/mVMGFF6QO+bxe29oITHk
oNbPyJd7BRfUhSbGOgIVVix6fRRZBChPyjczyIAy80577fzmwv2CrMUSlfx3e98JVTP9C1epTOKt
JSKpY+M2fe8tZlHPyMTrvpc6KuRrAf12unmkJcgz+rHo91o7tW4gWBym4UqvjhYdKuCnJhNe/fzg
iWno+hZCY/+wz9PRebrDRJUt7bf0ULt+RDCgLkM5XUWC0CE/G1P9i7Hn6GWwT/alfQm0mD3c+yaP
VAIDeWKa61abAwIwticpgu/zol3WSNub5v4yzcyEH33YH49Jylb1wNqP7A5uxREpBCen/4n8EJ1x
wgRJDfSZHq2U+6DsRQVJMLcMiJkzqWlvCxI4EtmRsTYDCDBOeOT3HS+s+opsJBZzltjlKO2tRJh+
z4bHpS4p8y5RodCBi4raovN/kVPEjzvqdG6PeSZiJJJEGNkiq4nTW4bqWXyF2YFOhYne1U+xXQwJ
kOCX0iDiLjLxSt4Auo91tjFOZ0n5lwFlFWSd2vSf4xY06urUqzy1qg0bs6VJN2MNxARR4P8V+nLD
2nwRDs/VlZfjmoykSvr16C07K/dqDPKYE2HFl+gpLau89NM7KYQ+5SkpLB7PAmVYCRKWn3U6RVM5
P18Pg3kXaZOewE6YSXq1MjtKyg/bCmfxBZVEZdJoizypmHP2RUkxWtIuZhksuv0fYpbY/b+wc1nL
F7145BO3tdN5VZZOvxwL2D5wx+bj/IQ+GwQ4ul+nPWykBg4G/tckZLBAXkVXZvLw90QQwYej3yaG
02Dx2go0OWyQouuMTswmfDFmlVKim8CIy7iU6JFhNq9a2UaEqLu80OIJGfDT7PbnprWHOSOpe3Yn
VjGPZ7sQIfsdTat+ZJ34Xr2mDOBn5xHqbeMxV19bCs4zaRE/BZmkAXeUXwhn5bsW4TLGiHI4Fa0L
kO52z9x66DmdLIsmV1kPl97FQV7U0yasiM3XKigxs3E8o4dwpf0leUKtl4jURvnZgrL19NpXW/5r
i+Z+15bX6JxlhyfUvhYIb+ZnT0B2T5oY7bzyD/BUuByPoG5W13WYn5oMoIIcrbCY5PB/26L5Wuta
joRU4cgJcaxErsA9KmX9T3B9RAzAzSoXGJPbquHB+gPhrzZJugsqXoX4yA5xwdXygnbcnATd5+J9
KKdXnMajQRr9LDtgmoKuGCiJkmTB8t92VEh0KUjgZwm3O2ylISo9LzW5svKvs0q/18ETVTaWUhBS
9RWnn+66xLmBrhCANOm6UVp+8jDZXC6fhZ26e2tOMDDtiNrs507lcNxxhwrffSM+Wo05k36ZPDBD
6lFS7s3TS3PdL4oA2fDJefoek6cqsWF+TNTRL3080905E7lozLFrmoYAzGGKyrhP6OmHRWqX8hZo
jhNBtuJdTcUEK+FRCcHV2z09zmaQEjxDnH9WHxvHMIaC7ZsfzkgLG9SkMmeXFqV+c2pwRJjJhC4B
cw1BbHwCvbX49LnrsQWJSDJ9u1iEdtBGwIuIAJXx3dIhV9j27CU9lIEZY+kYEgZpVAG3trL6cKv9
8nq5kyQlblEbkOj+Q4B2pn2GOvY3e2GrrJmn3H3opfoCMXqD/Y+1hg/ktO6LP/D4uCQSwvaGOiWh
AtDsVVZqTz01eayrAtOqehAEnp4iejGpEwUL9vXiOS9KnXMbcxlvW+/P2yKF7QMm1hwir+5iaKuR
DqDYR+TT99tg2WGSVnY6EdWcxJEVY/GpuSM9uLuPuZmoRIJwsoULpieBg/J4Rr/HkWrzYDrFL/W+
IqDeTbf6u6GI1rnvyhUTqHJzvHSIYSoZBNQhRylXhI6Afy0SJDdCfUvx24pYVfFzfF0qjebNUgi8
ZlASc8Nm2Ucj71zJLu7RQr2mi4wzKuQsMfXNvBaaVY7dt8JlkfLLy278Nh1yv2scMmYAlIshEwee
LpGYYL9q+OS9IBpOicueo1/W6tbWMIrSC48QiiUBovCKDafW8nP0p+0e/zSClVYbt70uw3WdLP+U
TphLNhowBD+MYB4D1xib3QzUDH0xIH04n7bMCYxAq8HG/KPQT0eFz6PbtM7xQwDypiFH7cCXVbzg
f7rW4ZfElEa8vPi+Hv16kzuk5tiBnjnWwkWKNti7Y32IZRMV32wueidx6qke6UOoO2qKWkL2fykS
vR5mel4kXvo0gp/xPl1DzlNF3G+joGPjiENzs0OL2YlGXcBULJjbkRO30Jn4a8K8ACuvPAHkrJWT
Bz+xqWcygT0z7cSSWAPbOEtsjKQb320HHUngKs29rthtrVhLt0hA+UVUD7lcIccEtJ6YJ6dqM4wU
SJuODU2hdFL1YYwXE/4p3b2V2ixAUKOA3orLBWEnQ5SQD0Q6PVQKzUcWn7oc3h67VXlO4M9gqPsF
T1RTkmlIsGCLVllyLZ1NZ8bDM0T4kY5H3yDIc8+sEWVhMdhFNEVvlIAK+/yx2Xa+YvE2zyfj8DW2
t7PIcmGg40u8gw20nmExPyF7P0Fy72sAKtWujTULn/bhAXH3OLXdNg1KePhbs4d+szLL6ROTyWAD
1dn/JKayRO4eZTK7V6ReLJCw0gcSbxI4AUvnEWAs+HbtBHJDTxPwq6NSqcT+OFYFDFyO2n/3oUFL
6ntd5aQyq/92iDfDve4u3y7hxpOTGohbLnZR9ZbCUZpQh0b6Ug309OBWYsQ8oOw9sA+368Dezwbc
Ka6HPm9oSz98uPg9vJ0KBV90JdmY5UAXYV48ezWG6zcOxv4sleOWgJx8bOjsetXvi1DaFy+VXSTo
MG2/m4FpIRek3D6hTnJNqYVUcrcwvkMIHbrQr0HOIryKyZWNOgDr/kPFxMylRrLDlTC3fWJHgp0G
d3Cnp5GtzG8snd964iB2/ZoJ1FH3BqfNnPaVddEmVwK2iwKPtXuzp03f4qTIEf+gRM6gu0XOYj/y
nkp67eUIZTKDXd6LCk7DmPkt/QRSIGhRznRSFKzj3Yn5aIDx/T0KPeNz29enk+vNZHzUyz3jpef1
GGmJJBOeiVPAd9u1fs6/pVsaW6BMS1VFTQj56Ix+Xa1iF5ZELBRCVeWWgQm1wqTO36vyDaoxfuzv
3BDANYPap2q62BqRSiCZ6oXwRJ6Fl6j38xJ0zk9XMsCQvG0CZ3+NK7EnYU2PETF4k9E7hM09PQ8U
HYzew6S+Sk/sp8a3fPx/1L27SxL9/IgbrJRaG9eNGy1GLxVQQIqLzRy5ZFf1KwRT9Zr3TzDJtURW
LnqP4X3k8aNF55zYGYKt2f2QNyjok/lUUunrzGRFN5+MjA0qvJCCdZ3Tzshh9rckfZHiWEdQ8G/u
edyiI8t4hoRjBx2WCUv8BplQXCAd7/M99K3l0qcQKpa6CNtu/7jEByyFwu3AoLbcJD8Q5AKR10YD
9sUwqf2+8M9xrt+uCdT0VjkM8VwJ/l9I69EcrWQtINcaFrqJIVdDpeLQNEuBAVqL9cw5TnMN0PdZ
4S2oegBbiq2/K1zLw2FOg1bgmvF3xBFcs1s2/bQG3Z8BHor1QuL3lajgqR5Y1zZ4t3pSubeO8xQZ
YWtONOBaT8bvvT43ljschqxVJWHoVXtRD8Hv0xL4qxOz969Cry69tJtYWQddkQtSmAEwjETthgx0
jGXB7OVdEd5nvw9wNnngAG84DmZ1LPYxNgbtWjch4dGn0rMS3FP7FXBVW7s4YgGcho7QK76TYYr1
n1jGb7xNLzC1SUVGmPOiAujD4JAQEXkMxX4Py3pI5TM4TxBcVhfsbopZCvtrtpltburGg7ekOwsU
Ecwvt2Duxcf9n3vCA8a/e8iekcfz1R+Ka3ovkHNn9qf8aj6mkdJzZb2MT5hjGXsMV//0HYgFz3Ol
mysvG0elJ1YobwBJUjULItLUODiOBFJ/jGBZgi5wSo3wmokLZwj1g1TTdta8iGFQ8omnDm9Bfn90
UnWx6lqtvjK6orgh5Kb1FSY70NlGXLVVXqLb9YlhxX4pnnAcH50Pg5QBV9bBOhKueMtUA9ejoBv0
tQ2S5knxrq/UtOvgjFOhnL3k3SU+MYsPSj9u49rmGySyU3q+jaVwm329IEC8vqtfEJAeG5Rmx7VE
fMm40TwF/5BOIO/tIywTgcVQJnwIM1kUq0TborCn6eD+Ebvdtr7cKSnJKDpGbwe4dw5zJgH3Grp5
bDXVFwcfxpM6NKaGDugzJ1O5Ijr9TrsvkDdCmi0nGfX0bSKtfrhni+a3Lj3eV3Cseh330TfNx50y
fQKmBP8ZirDmVIl3qbOmKSvFg+goGxWmCejG+8n8VbPpCk1FjcpaN2iuhcmULycTd56eMavEzcGF
pDa4PoZ0EZ9rKIp683ig9rCFw1HhMVLA6EtXhHIZM1yhqxO8QIGZrdzVeZtyrQRDHNq8boGCDAD6
qiQb34OYuIrNQcZT4alABpMxL91Eqe18n6CMyfdkX4r8MYEiT7qC2B0uAGBFzMvneLuvisG0eH2W
rS3CH4qMu9vPigfHuIp+fPtH9wl4ToAZ+AIgDjGT8dRzk8S95KrU7RAq+omapgd5RKqRdTZ2YPVR
+qFRVtAaQ8VT9LC8zfWFRhS50dCDc0Sq+zkcE0wbZdoVIe4FDn847HZYg15g+PUoyAUaq7TomZfl
2L8t3GUa2gktwxI3QEY6Fd3UviYKf6V8bbEg4JcZfaarF0b6zu0I8u8stgxUO0FpR3gCN/7WbibJ
rGRZAlli5xfGykcg/0zWdwhAeDZpHD4ebCbuXdEkXsHSZZDfSZIkhdroTs2XtFIXGl9v1VNCMZtm
LQBm4d3742RVOfgGzrotIqU7pbi0M4SQmU/GPKx6vrysrYHxdopVyE6HdnsXfe/OMWfyrGIt/YVC
wLr4rqFr/gko0UkrXtk6C6TmGR2CsNM+19EvCk/4EkeJklAAAKsTq4JA3SGqAu9g+l8Gc74BdDhG
60WEDmpfuAGxLF3fHo74rgrFK7TrHB8IOE3AGV5CMwcI1b0HXCGzpuwAtUs+MGEp7qZA1nA5akE2
zOsXTnPOH7IATPl/l/YM1uRqzROUDGwN2CsTk9uzdyjnTGdStJmhlj822gujXdVh965K5zsIKfIw
3eoXn5XmEwgYWVcdMh0Bvjs5dIEpnEtXKTrUHSHrtj0/39Uwa6xYoyKNYQs13ICzOQF9Pdgkr5ih
/roMQv2ZGlQf2j/fd/09zxt/EbA1CSn+4myQcB1i5wfV/e4xKQxSjpSJ/3WDrQjeEk6qGYY5DtpF
m+FO44WVCeNTIjl8xKcQn8+hD89WT6jXdJYDaENpbxoKBH9MCStoQpzjrji4YMVqizMKVhQVN+G/
I90y3hDQ6eL4wT3CugcxA62f6JxFVB2AvMDmA/SCW/k26Gdpo8yHbVVenupJvGr/9WnewINECkTq
9P0JOIQzWK6yJoV2S/7MB80MT+8l2hxC4nNrFGbblDVyuBphQrTQY+On8G06IDmIaNX46ioJDt06
xaQ7eI+ohG5kizLYrHxynFnzpQgy5DSgyoXWWSf0rGAgIhJLhQqwaNozbUBRdM6/gQ83IX0/KeO0
SxY62l68v7k5PPjdW5a09tJPUYLM9zJB8zYEUnQqZzS7KjF8AeSBFwG32jWsFQ339NQ9rFfXimid
Oa9AMPPAd2kejd/aWzflnxoHGB0ROypzo1FRD/ZYd6T0pFwgjaIU2H04s8i2jZK8HDIRxu15xQE8
DPqgxXwnYD4sz42btQWE3WsMXzLy1qCKUYmZ5l2B0L26hDlg0UlOk9uly2P8QpMCVzQ4gS8YRwvd
NBlrTT5LAijEHI2NhMgkdvD1XYDHmaTD5hy2wnk2YI/hh4THI+AxymJdKwpBOcf7EQpAY9ag9NRG
AEZz2A1xWmmPI3FDZBMu26P8YlIU6tE3bSwevKo1lBJH2DWH+ueGQc1ustZGqVpbdMC3C0IpEe64
waVlFoPzgId92XMrr/Kyu3wf1Y/TLrZMRyrRViXteTxw1Y+DstVw9HNpFv03SDZkHKEr/Im2Q14n
sZQBmrNBZHJdy4S7f1PTopkwBikvg01SY2bfGYjfGsW/4ft7bT3H5hwZrNQwEclzeqdn+e0Y0mar
TkBRVJ2NSC9NCXeJBoxBNc32mA9fUM4GM69qT/Jm4ymIODbhTjHwdMQ1tYKGq6oD2p4vphj6s50x
BhLFEXCI+JOeopmPbionPQHYTQLP93I9Z3f2itXcZqrOHO38MamF0UDtjs9ZsBcHM9n8XO9IAydK
+VV/TgkVqVASH5fmXKKXHE3A1i7iW5HM1aLD+lyESt2x0a7tNOQOoZCfJBfGZ9iPl7TDruOgC6tp
HojxbxpSCN7F33Sud5I3z0rfKsAmBCza/WW1SWSSPn/FBrt+VplCq/qhC8exB+u1H8pqvsa8Y4R/
W0d26RxbnX/BC91PHWX8vTcCW1EQZTQdDBlGex/hg+EUOjwdL1ql02VQENfk0wfBFsqU3J1/l/FW
qDUEpJgQA3Qh3QXYuFblJ1pDN8DZPjIiEVrEQ4+NS2hpx5yW9GIcqlT5uSbc/yO2B154X6b3AoiV
ttXVw1zfLMtWl8qXN90BSmVs8qeE8bu4RfxTKUEbYlAianuCoI/VrzF/6r+Lz0BUVjx7I7uPOW+1
GO84Jvyh7jbk5C1uLoFveuoGU7OssuB6uWAdkl+jaFpsgq09RurkRldvtnb9hrDd4vpVg+w+1+10
KYc660HduxPhM+uykkYrbpRx4aJ4jtdbR4CZsw4AJud+DtJNrsi+xV8nu7IbkrELYr5bUF4dKYVT
dNCQDeiMTl0VQ5avqZaZbdSuGkdeDjbi/GYXXS54JxrGZVgxuVt6dU/bpdOZxHvvag4iaoj2L2RM
Yy8+V6cODz3z71QdVVNDJp3Mf9hB5Pu8OeoZne5xrifuGGUgxAgdHxrtAlBif1neIpmSqydU8CFH
jwTU+Wyr237RqeanPbrlu1jxsfMXoad6knW1FtwKm0Lb5OWFcvNH2uz8/3vHxmvNg6t8wjWtMDMM
BtXYq9j/ZFO5wpitlGAo02sCVAKk/aTnxc1rm6sQu4nP4vYLLCprSyIYaaZjrcDwL9wDQBOEAbS0
KiPl69BySty3ijf2D093iB0DxeDLO91SH/2dvWsh5W7iElYIERI6IH49xJaFlQt43n2adxK/sJO5
DzZiAB5wprWT1jeAtf/Qd+FinHe8tGF/09VWuCPfotjjgmpH86Hye6pFOPRiZurPTfIdotJG0Iqk
150zQdXV6mIJwykjNSrNuWMPs0Eh2KHtt0/JNEgWV0refV08UCRvgZArMvQ+u7gMSw/Zy7AKBPgN
006rCuIAhgktDCmBXUm61MWam/5TMY7L+cGHDlvjTIkf4siSmWcxb7fOpzhhS/nWA8V37uJhJonU
YB6KYywniPaN8vBkBJkLPbteXcRbcHNYd2ZYlmsMH9kl4FLGLGDbEDzbz8uF56kHo8woaC+CHV/Z
38Sh7K9tZZ5yENi3Cn0AU+7rPQkxT49as9sPNNPvg6upCA29X+hk1gphOFx/7AiSk0/qidZM/yjY
2o/y/Dg1mNaoaTEkY2DWXmmQU0EqgQNbVvpE3bV5H6DKJA/C58wfcBQCHx8ugLiMkaKr+lOtP0Pu
f+0p+HHBO6nmW+Gj9Yh8jZkyeZgvgtKioUW5JYVsiCzoBBF0nwUN3f5u9lMXmt1LuAMLFKAYe+kk
jAulXIOA6mSZYEtfG6lSfrkB3MNJxqKZ9pgBAIPnGZL+eWNypMtJB6CtajlC9Lm3NXdyZ4FZZCXF
2kCGK0Xbk5n9pMA+P+vJKMjp77/nYKArPj2lJ7e6NYvPXWJo9tZvntWzTZqCUh7ubCf/J2PYxERP
/nsY/9SWOeIgRYNosE1VUI9Y9OnyDdIB41zHQflPsE+uziKEc5+w3MsNCM2tA6Ojb4iIi9Y3tVus
PARIo3Fpqi0kvIhZUwP4IlouON76582P6MPY3S75HZf5wr55IRLz7/YyE1rylDLh+4f2KDt94dIg
gpjSlqTaHXDCq19DYuLmMuwoaQkJfDfJW+3KB2OZKVbNZ9D931GUQYsc7wJu1Kke0JBBlyhMJGI/
bT47aH5hNjPUrL3DaK/KlFbEpPR/ZThPXsqPt5hmlqFCCe0ZFtIeIsZ9We2S4V3XgIDmPVlVahA+
7kaSErgCsoWQHcOmmkFfQyifD/yEvdZ2NKuQBF3em3rftEjj7/Bhh0E4y5+rQlgkfEpK79xNxBpg
fb9m1lh/mVImfZKo8ANziTBi5c45L9KdKNWhGyDo9o/Ds1RYqie+ZcPDjVSF7I19swZPeLxFXBaj
f8wEKLCxnWzys2b0cLqECx440VHJEdwjPuTuzs4GUGg4CDdgxx7tMi0Pgdk3aDTz0bd6Fwg5aaLq
8LvA4rmyLJtlyYHSIRSKEiz1Tmr7Wxs8FKKqAxGGsub5Fl4GYYVTfO8UkIfWVruM8PJaQBSEB6y/
E2jkXcCMXPvcG/bhFo7JfHGoq6ag1BvKnA6cius+vcin2bixlXXCGHXeUNIdAjVTp6uuDdtmtxFc
sa7P1q/nNCNjunAJmEWYWMqNEm8LucEuACJxfAXCSMCfj/uF2G/FxMjYg+aSv+QcQs5d/04Cl1o2
A/gWP/PdNQBdqXTdIcl+lBR5oy/QZy5pIdbtGvw0g/YreX9zW/cBcP9P2hyvsd5ZutCMFuUDku+2
NUlhv7rgvMqMgWnmlG4lrq5d4htXGqTcBS8YgSTXOCabsad9KbKUbWskjWQhfH2WlAB3sNQ6TQ6g
dXv5J6nJbxTlpif2vjjeaycp1iemuy/FO/EV/DP/XU2ZOgEitU/gFj7O6/lrClmIOxNE33IA9PTx
OZDvaRtNwPEtbxybRPluQfYLbboq8JOs8s0SJ21nM+i1pv0r5g9gSBH/CSbwMsTxnsOajlgXvJ6Q
9f2ljLljC4GYn4BO9KTLQD9Ok/t/QSCpd561OWHpvxRmFWlJoMOejUjB8RJ/gT6wZDcemGOXgC/0
xdRhgJ9X5j+yVW2L4NS3Th47BFeI3MINgdMDj3c5HQHXaaAXbFUrYDemQGKYQfs/sNZqiA4pbjUA
+6P+aj47jkbwJgblsQ/Na9UHJGl3Z0/obzefblmqYxhRgnjVElzREM6Rel2Cs0QT1cr1RlCT2MGM
8l6M4LhYYEjs63PiqtexMcUiRRDAAiD1r6wxmsfp+nbDna8HL9ReLoQx9S930HPZXd/82eeP4iXp
sSCyI1eCJdrZQqQfvgvqI2pV/TBmMUEbMS4rMym7wQw5Fk6nEJynHQg8bi9BKRORxVArjUKr1AyL
jh8vShxQjWV02oMXt4mrT2qQfkQTzuEYr7POyYfjaYn8Utng3o7sLkK/K8J8kg9igTibO+iGizmc
IiMzxyn2QCrsjQ4Wv3XWp+eLW5u4k1JGzL0hXTihMthDeAWJMUk0fR3ie8vN06uHjzDEsBeJqb4M
ThGuhs+5GdkSuH4VZmO2495ZqqMi6mXKoo5MBjkiP7BJhtH0/GMYJxry7Fu3fxINqm0Ano+VbLtS
/pjOKx3OruRLbVtUkUYnjrVzUo5eClxzAPhcrJhnO8COpk2d/hHOKdJMBvLVby94///DC5DwGFDb
SgxhugJTtR3FG0cUBU+bxmn/KSqRYJMml7SA35Ebco10McRRQQ+C5R9eMcW9khaQNzKAodmpf/gu
4zUHteyPvr5p5HOjYobD46EdtG6UfhfQww8sRcWHG1m2Rt68agNwZc5dgwAHGr77v1MTLGmJrIGr
leIcwntn0sNcAlMV6tumteeVUfEbKuGh56pOamLn0RUSMAjEgeUn5BQzDe2WGK2pMGOuc7cUiwHp
5eZdv/h5GoIGLGgmUK4ABFjsZ3vOoleK8Kg/rOHV5JJQ60P8TJMoSP0esQMz8O1OSSlLmDgQGyW/
F4WGcIqYEPssGwxLjPYaS6Ssh4cXPjqO1VBoRYkx4V/j2KbXTW4qk/BH0EMw53kTQAHl63MmogiQ
Ce7DYdXRRHVLqjlr+8Jls5jzeYnrmseQYP68vG6on4UjojAhlf2eOhJQRuH7P9muwOUWmBMyImKs
bl1HDPoJ5Yk8+WTt9p/P0w3+7CHxG9Lh6Hr4caA7mcWGsD1Fxuc4oS4IYwpvhBsCVkDtotiyJIq1
tDICzn/gdu1FVJwHNBTD9DZ2P0Xem7/yjBJhgknXha6F0nuYvo8wmNPHsDnEx30PZQtPi4y+2F8F
p2pmJVVhofUiBlVadu03Gjffv4UKz8zzXJKhc/relpy7ygiMhXxioSlFyxrVwWBMU4b1TA6xGaTB
2uoOifMcdiFOePPokTSD/80UX6kZvjMGBFe87z4GY8EjYvB/daB1xk8BCtpGE7LIYKp4b6oO9OxT
mzB4Gk6DYGi98UafBptkFSvXLL7bZt7qOczMtjUt3evWiOGhTODVLG41VDMCqJPADDTBDAAx+IQv
B44r4cz8H+nidEyJKtNUkASkpPp/lDU/Ryi2JLtFawgPlNLe6KYuWtq9p9S06a1cY6ZjGdjf516w
vLzK2zF19OuRhjSLtFC1Pr4ghsSVxWeXgtgVnipHM4taS7c+auf+SoamnUlDMQnByl/49pFAe/yX
krLDspuOw35eqW40ZPCnbGNcDX0OSclO9PkKvaph4vk31t+iRpYju4o86q8zC07OK7wAYbiexGtP
uT9z1iitDzn8hYxGD1VDNxus35aGUlomiZmBEj7G3FgvyRi7uNOfYHBEhRjQ4tkNlHtziZpVeO7R
+hoR0/YjbF4+SSX7jOxp6CDlDzwGOH+l4QERiGrtsTIpk82+yjC2CGDCcsxIhCYw7FXFy4cI2L1x
iYZagrhvqP9TnZw4bazd62zNFQDbx8a54pPEDGlyp5Sn3WO36zJrya53w0rx7Y2KorCZmtCDZLhM
toq//dRL1VQkchW7eKKfKNeYQSVomibRKGB6roXc3k/+VYMkzygYH8qtWyh0NbC1FSHECs8Mdcs7
+nhX4n0WAD96nopBRoajbymQKrDp03IFutkZpVCKcc5Ax+LYx4xVt4Njs9QitGgfThgSmPTg8nYz
08u00fcngqVF92z9NqOWh2OkfuilIjfh8QlaplAqNPyYw58URGwaGGp+SPhz9wGym4JG74BUjKI0
uEze52CpLAHYrgb5udUZRCvU4Kil/PPajhpAohotg8uPg1/i1zmRsBWeGLcDCNAt8n59CSiWjlWo
oJBtwh6Qix44noduN8/MUFOmdOL5qgSPIOqx4BS+LDj45qEgExrDnPCixhQ8HIzPhvOAZepB0rS9
zrh+6kOERVzIs7joJAaTpTFd2VpWx3eWX4vveadK/PWT1pTRey782/c9dXfqKdvvcJKJNmE+YSk+
ij4NMcmGk2SGyyfyBktY1ClyQ1IRXooBzUd6D768j935XXvuNhaWVenmRFDOnzTHweiH6qzkCaaH
6FZ6LfYiaoXSew42Zj/Iqy3RcLLinftNIwlhlpyO121TxcmQadp4LiDt6R/BQXt8FGdeqj8sM7n+
80AyQc+3fcV1W0HD0xRjZXpP5fTF/dbI8HA5eAHizUrfTd7PBu0XNmXp8+4+B8CUprrPgwXYMYYy
6e0lm3+nts9dCHdZTIh8v/mVKrz4Qh/HdgxpmYuC4lHK73xNNPyFn9ugJqx+bqhPO0riFyW/62Tf
qy/7O4K9c7OJOf2mxE/eCcp2lcBKgDf02LF5JnCknAKRpwQUQETZ2hiQG4dKvpeALBrK4W10DIOG
PMk6XyYM52cN3im+uTtlHsfVA0Glmg4P0uv7QH5wOX2juidkGe1ZM2X2F1VyTx9dvLrT64PMycfw
seLF2UWu9aYQP0BTEw1j6JXU7feylQRuAHDIWfJgtvjWdcTFTuHwPYXPHyP9Ja9EwN9k9pQNMXVv
3D/KmRBci3AmMwtJHOuNV7++vaMsAo5UzWS5r0twLoi/MXJrHRFf3WOHjEt3ECmriIkj/0qlshVe
MWQw5026WP4AcDSln78CxXEXVMTETCMrHn+WiP91DJy9vMKyNnWhyG89F3d9GsGF/gWXJ72fdmBd
EZlRTs227N9yRFW6psLJrBycL8lFXksfk3NfJJ3aJqcYBb6kGsrKBPtOpNMvnG13vJE9KQWSQ63S
MF1JX41Wp/z6og6BWOXz0Jrsp6F8lftuFvxQtEGMDXJMf3xr1nAZnv989APuh67U57DlVz5KXC3Q
oJuGwBKELmHMUn/3pjlZfHfE5rU1d3FzwTaGWPpZZHy5iTiq5AipJuQxfV58dEh+MhZ5gpVnzY3w
CquNDRUzE9eskFwjGzu1xSRYw53kfwtEfiP6r+Rbl7b3DdAxm0fYdaTKadS0O/DlFlK2+V3J8yHW
Gftwj5odDKt38MvS+wktxAJDmQuvhe3HuMzzLQ9Qo1e1981h8wh8nBvy89QGCG2JGNJHf3V42FZY
/HhC8quso+sJlawkUqZJdKGyzkV3ubknB7JUVej2ai/q37fZN7STSd0gGhqWoyzkQdpqExvRnONZ
Kt3+c4vF55y0WilxY5gje1dLjVEFI9vc2OFFjeYOOCSOCsklXHwUDn9DM5pmypmTEirhp8M/6Zx6
3SdEmGNt4V/4qyjDe6PmrGIcz4yFpPZvUJqwOppnfTudrCVIN5BSPkwghrQpw1LgTkB1JDD6x2ou
i/894ms0pet2nTDB/F6J/xKE4QnUZ67Dc9VH5czl73ZbyPq/AGpQKi/8NSNJ4lFF5Drmp4LkwAE1
XaiFEGxWVIYesOWrKqc671z7fXPVlANyLNmuKuQytE++o7dHLBYbIL5qU6WWJ0G24dEiiMdFrlou
rB9Rl28j7nS1mQl5qZeSNeBodlD8UqSSq06lRwFGTNDqlIZ+IlSwyvrUO0zn7cB8RdkCI7nsedHa
/ZnPdGpE1s+Hepd38vJBezwMajL1NCvMWiifruCDwsbfVOm8dzmb+JfeuwObmLBOtXiver8/CVzq
tdS4JPPZIk6aTiV5eJIyaW4AMj12yCO1ULhXtKrdvUSG3SZzUGFmNzUPGwP3j90zFMV5UZdqAVi6
W+ZrxJRgSHin1FaMguYJsW+cg0T0N1KUZC8I0M5NLzey6RjMqY3kJjtKNpk5frB27SX6UiIBLZIN
F5hrRfwG/BOKeHMeO1lbv5y6f9GqkWWnoiLwCgYH4/ewI99sYX5/LJV71Zc/MT34TVP5qH6yPWOt
iw8cht+JIrcsoj02MobBgCrgxsnrWpE6/+TLap0Ppp/5GlF9Q9mkDQQ2v9P/5TZLjZJzFgGvuMro
Oq4/V2LGF1kuS+qU+T+XlqxiVZpfHL6j10hBNjGFekn5HXZ0EQgrKymvvnxllkid6ItQFxWsGwhp
txDFchtB9DCclMaZG2saz8q2pMZncjxZxEYRhq/EfdLl2dgfviT6vszEfYUuxDBBnNL3Cyfv/I7H
JGERVosXVo/TWVL/iSEBXSnxVzUPiSJHmIEhNhH800rp+SD7/ZARnrbTmKKNm8oQJygIsF83AL2h
YsRyF1ZiVcPXyof7EwnMuHljXIvu3zbZpkoIdSufVo3Jw2obZH8sMp9TYR3H5XGuErwVhqmPy9Ni
vlC90LXHCJpFIJjrirrV6hyXe004ue0DLpHvHZ6PGkXL70YdUqt7SYtWDeLLU8PSafeJu5FI+Bg3
nITv5YPEiVpuRm/eGtBBajt7OPp0mmpjwCCEWL3oVnYBThnisFF/oLxF1/qEiRuGST1fsv0CwfwS
ax/7g2Ee0+ttfkM7bMovxOXox0H9gXX3f00l3GXsfu62C/KvA9Q/BUS0BH9KjytvdyQzidEZ+2in
WCo4SwBDFUOy9xmgh2xIFVE7qKoDm/Xw2YvRN41Gs+1+BzenXhNcIUUwfIzf7R1qkaAQLaHqrcjm
7MmVtnggkLmMWH4kuo1F5/FEdYkwVeXPG+WHFQfA1Nt9Xg/0PgkVEwId5IB7zs6sf3sLt6w8ZMis
Ac9gyIYDGzZcBmn9t+7OeLSmCXO8cysP+zXvvtPJAjqAo/SnA0AOK7Bz0dkDroHOfep1oKLaaafk
cq+8gBrDFFRXiWAp1OdhntVPkqXs8wMZN9lSguH/ykfrmdEdH2oQo9k/qYilk/WumU7XjW+Yvyto
/BPKgRV4UqS4qiyM8lLDYnYanVmaTzaKtmUkE9yHonHrlz+77f8FPXAaYz2NBHdLpIhbQ1dmsGnM
CPbQ30EUbkktvBmtxwcWYL0DrpQ8K0+FBmsEvzkWVziZSgNiQJtv7Q7n8l9ohAoJSG+ZCzUEInjn
0BpdIfR/0hgFgixqLTqMGU0MZbZ93PNhyZZpzNh7MJC1oDE41ojp1up6ybLvZtXWNt1MOnGkPcFk
DMbygJTzcFkZKILLHy9XwN0Gr04Wv+YUVP+D2J/G31FtOTEJBRlCUDgPwosAbTyMHa1KqqFDV/ma
QNu/njy/ExA1zFeb1DbEtL4qSPDKfZ/ehLCO7KqeHq0kaAL+ubw88qQlLfovUpUIsc4fHI7Wvc3g
eWfKD8obs6EpkehzlXKbcMwcGeZ2e3/v5edk5/bgU9NJvNaaD5yyD8Q1ubWrFaoK6HvhH2uvEoRI
zfXd2K1wVJVRM34l7Br3tgpgeFkw48rEFq76S9Z6vzRPZ7isa37u4gvp5PEkf2mS1hepgY1s1wIL
pGZ+GfV86GzGKOWG+Tb6zGAjTsJqqaKpwgwWs/oMXJg/AhbCVdH6CSWpLcHY0KnDeSyKZiJDTK7P
7DObK2sDlTjJLUAi+1F6IQglXJLKhDiodT/iVbGlBLDdj7ZHFi4bpXAolL09DzqGIoyF4p8MLCxZ
TPyvAmWh+/8uAmaQolUq9EtrwFRQtzI0EAv5Om/uFSKWLMpL8Q9430Yy0EK/mfEzBZ+YjWwwWx/n
hYK3yClNUm2NtEi9+C7MfbDb9XRxYef3IHN78Vlmm0b/o2eTuvGGcshAg3xkgTML8XHJl2jUJqGT
eiVkwxUGnCkLEYodmG7UiKTPO8Vp5062FbGhTXBn/RbMQHnYwUlNzFZYHaKbpOmXg+tFf3i2JtLM
Rn0d75/BrR59vU8xsT3e20JpxS9tC3BZKwL2+ywCzn40Ao6N1kG4piMVGjZZjkpxUj4X46NHSRNY
KPCt1P5OcE+bt4Ub7OS/D/YB43e/aDoDtUgFw8CL4pGPCZobfQvsvFp3Hd+YosFeVaM3mk9XdGvY
vQM6IVepggmcR3Ltdc2ratDvjcfWbTnB/QJyoxh3nD1nHAwk5ZVgPGY++ges+bRiBez80RcfI+1r
YarAxRrOAQjPAsWYETQgPfcKJTFxSqBmi9vYDZYTArO6uOJQ7vdpftOTeWoM2K4CNqSOp6uvFl3u
P22/ar/FEHkRCmB5iITwaJ85cylkNTaMmJyCYEU6hU5CWO6GSrC/7TJrzmEdGDLB6/x6Hnw2r56o
EsVuQTv9E8I4P1+Rs23x+BAKi1egE6iMoerXGSFPBxp74ExelwWsQMlHt+192NSqpvGgeP5sN1BR
ovJzzfk1cbgGp9XzkLKeQD9dJq6BeXO7wYpzHA7TTSWBpzeJ4jUDZKG2qCyNskuWNcO+C5U4UwUR
c+5ILmbWD+1OLqbnNNhrTy47dyqxp3SUsOnwVoNFwQp8E35QBac47LAzd7evSU3AKg4kbsU9/fuH
B98SqWwWXo7C+BzWK74dm3VGWfObVDPFhZkmpJWkBaOrJVhRVBYEMHB6LaccKJm/2JNT4LtOPpQZ
RSl1kMD1Y0pvB9rqeVOU/lOvorh+4BGRf5SWhUZ1hA/7EqwTqeYhho30bOoCQkj87fuMyzXMuu3q
KTi5/nKTT3tRkgxENYR6oLv2t/2KSFomW4gzOHraf4/I0q2XJIZ8DcNEgYI90qOlwEy1XeAsFXba
U+76oQ0MIK9EVRNdAKaZIFRxM6/dd5oEG8N3mChkuPFgnxlUlVgoP2jIMrZq/ERkclWqq/yOknSL
Jw1BRtkUZEtVcQpt6jTPGgDrVvpRvg20LZiQnjcB60IzeHGFXehwxBuE2vt2B4dCuKimfGpUI99R
YW2924HdWbu177RAym3kgXrZNaev5Ett0jSHA5aLZvAx5al88ho8NrAp8LTUCb6EQ0+ARfDg57l+
+MacNcMWLLpK0CYovU+aPmhaZWNXERlOgVVCx4jrSMemUYpz9DcGMpcyV4GoNe+38ImCSbKarYS1
AJ/Xrb4aYf4c8DFszSBwRN68+PAu/y4oeq8dzOmqsC2O5IeA9YkxxxzGWhELBDH4SFpbeQw7oUWa
0OGQ7t7sG3lnbAn1ovkjnqwQWs8V0ZpV5m2Z4UQYBlmZ4/oNrNmlMwwSdpSjMtxAiLkxa42fJDHN
2bZdldkwI32p1R4uNoUpQvh11eEAF/BU5LvoOFBtPN+2oIYD+Ak+FKuuPA05DeEabChO7UVC6C5x
nwrUOtBN/c+kiYN1yfQMJUW98IlWhfyJZipxewBrToTdt7uoZ/KAG8GYHDSn6saFmfZh3yObyHjJ
n/PJvK0POodN3IbzUbdDpOh1RMKtRGwrnIeEv63XQMtQhGPLtdk0jrowPxPW0hvAFp80nRdlCkjI
+D62iHwu45/gCmwsyAV0StSn/39DyIaaQbetSjIn6VVjmMd3QI/JLouSpzvMJv8Q/6AJ8YNSsyhZ
vIFUJc1wNVB4xGqPUI8gZjdbOXDggqbQLsPKiwnrZl680rxfIGGsspCUvfESNpxaqFxFeVzHsdAT
PeOi15fARDEca6uCEmJHwT2z1e3PA8pVMxrWzWDwv2xp6WdzYZ0ih9piM9l//wYM0H4uT/jM6Lmc
812lNvhe8HI+GkOvM9NLxjITNuHUBc1wxaLBixwnL8vl+JclLQ5HfEnobZgyVjrD1Dfa5ZTTCRiI
9lNwNrKCvwsMWzah6Jstah+q3sY6hStL9nG5V74CdYnxqAyWe6LURxLo03FYoQEN+4Smyhb3OcS7
FBmpg229iHGF7c+RxRZxuDtBZCHSlFO7xbCv4knZYo9gZ/Vi6xHayYvCnUtwHmDtlNQgfUEfGw+P
pmgR0RrYvaFgrpmWaqDkLNG+LL5neYSeImn9ThIZZFBziYccqn51jxlXmOINeU7MI4DsiIzVEeT4
uzEqxXQW/VsIiFmzXp7DanhUaAqJL/NEhnestOVvsMlUCol/NQwzRqvoferIcP/VqMwINx8hdMiG
aXLVJO8wzJdLN0gSeboyWrFBno2JhKAMNdj/wViR9nwdVclM07O2AIxNCPn3DapimYPFs7L2o4s+
O7/IBvl+6BJCbCJyj+lhWV3Iu+0HMTDd/g5ghUZORJrrHgdjsw/zt5aD4OUWDKy4BLv0zDIg3oDm
rSb119SwDsxVmHH11v9ZLFk/wRBMVxbQurYhUQKK7lKxlKqs20jBLrduReWCiF+EqfuHnWEIXa6p
v03dU5pIB6CD1YEpoyU8nsSlbiDbiv9gRzIc0jt0/xl+6+r9FeMwSh641hoB4pYHybuYfy1UG7rj
aFG+rQDpecPSc7kFI0Lk66fC/M3cDU+ugPat9Ud9PhA3xrcMDcY4s8JoBA3Q4oWixTL2mkUioCm7
XCd2Z/0wDDQc/lDMsEq1q8z3v593AU+uJGcOQRkBFE+3NpWojvHjyjkk0Vs9RdnFiyaCAoFl6V9E
2gv5tUwT+qUCwnAteXWvUE0dNNm7HOxf3GXdbwMsanG4c0xctgcksi3fSlDxUSVQaAGOGF3LWDNM
ig6wS0HMdP5phIQHqYPlQlUaakvBmAS+xcvFOQyJ5Zjp+QuQNji6eFlL9OddMvY/vuIoizhDXBin
7vzfUvRVxaXUqCnoA4GN/RB2XMyx5cFspIqnCXuxFXtdwUDZQuUnlt+GW3xj6m2XtHJESDtPI/VF
GI1bUGaODX5iNsQIQBL5jdmWAVY74yx0uX3mL7xvfxqnjIEN/8DZP2iq3YqkvGVlLqGtZ9F4sHV7
sVJ1gDGBvp3YTdJq4cMqKmebYqzYy47Xif146fC2nCEqzO6TIpaynm94Qf2xNgNAcp62cEmdedzd
wLGogHAQiz8wGr398YVFy3pGaGDl5ClPWblKnbVRXEWNxNtCnLomANfn1ir4+dm5A55HWBqleRtM
R+UxKcS8qQv5Ewv9ESWKBiIGCoTudFdpjgdX2hPo7dNad2SpLC5Hvj+gMDc9I9bLK+xY7GM8k1VV
WbsAHHZMwt24dmSRd6+I93nnJ2VPa71T2XaSRX1+BOYPoH80EeXc7HNUvcmT3eq6xNrBRXpsyWT4
lPaekpmE2Yx6ZPi0CES2WC+XmuzrsssQwVm5RkYO7g5M74q9Hvw/m17XIWFrCETmuxTFiSqLo+57
Kf2PcPlhyU51j9gzAtsT3U3PIcvFExvdo9suv1bvx6i7vu6SmET+9uUKxcT0w1kKOJxzlmYmmFwr
bQT0xgUfE3Y/aIG+m0UhD9INNEfHjz7FI1blpkNdexYXLLT6YEqwdBlFJWd97uVrbpmyEhCErtVZ
XubTyRvDectsjFW02IkCs9NavLQcyjTrAh98fa91F5VMfEoR58ijBOWnz+fOqZs5C/OPp9E/wUIl
fDGAVNuwM0Yh/HZOybEhgAQvwV32IBTRNc9AiNwR6BK9JYreqiB9sHaiF5PS8ia0Rz+cq2To/y4M
L8WuhnItzo6RkCvyjyyDHlaWMDWRtiXlMbn6Vlp7yS1kbQHX9eN5b5+ApTJ9vuSLhLw56q5TOtVa
xIMu/fEq2fQKUpVxLzOfyXtXfbrBjrNvCdUrcvxioXu/CU80lh4rGU7Cyr6YQS8tQA+00dqwJfIz
HMiKHWo6O+MIP9DejvXQUkL22B3hBJ3Jrc0bzqNppEYwB/pLV/poZ1VMrl9lVOuEfPRwzQfgzgBB
QEm9u+xJ0rVZ+EHMk5lATgfbsruYGPqjzQe2k7QEyW3rB93UHWXkkb5VwcO593ILkWcbMzK8gEGz
2JgVgmgG/T96+20V8px4ld5FRn49Z/2e8zh5Zbj4w1QIW0Xq7PxsTVtl6Bz5O4fZqIc7gV188RBq
DCFKKRuolTLa4yAKJnsG8ozoUQCgLCu0XlnkRt/WNp+s70mDLq1M6umMHhtGapMwkcEwKRUQwPi3
TwS6BpB4FenfpHG6KwQJrJgeXnWPa9RhWGQb/QcWkCLzpJGww+4XYcakuAc2vjKVeVd1Vv59nDey
kgeKMhQpH/Qh7vfzzwL0eDy6UsOQTExvhTJ5Q2yrOfmlvbiRJn+YGohheliliMpM9FqGDpbipWze
Y3cUZYSW8sUKphiZa5YIhbX9Efh92IdZ1ERx6h9hEw/njZvqFZbBWcV6FucQmrdvAHmJko2BGxsq
ER1LC8dBM+ezzpECPPr0wWYaqGR4T9/8N4fXc09jrEDwjcPQy5fpStZbstWGbJl5nxpDwjkS4Usy
kwvbQA3PRWamtbCvwT8BnjKZeJCBVYiAfnJ8x8Q10JvGsIptL8MFMEiynjysC30LeTR0Jqho1ZMO
CX9PoxibYZ7ih9W+BeSvsxXPKKJLwiM/THa7aNzuFjYNG3L6xx56eRzizeMjPVx00i1sydQFrb+b
57qj9R2XKl8TGaDWpPHlLSlxZK15JVmMbrHuLa0VqyNJxKcCe/NcM4EyZJsrUAyJC40IyRF7CQpI
zGLHtcNFa37B37Unbwv/ukRM+qhwzLF3i/XF7yaDunWK1qMs1JVZD8IwghJ4Jy9TDlH7ACLvYNy3
PAR0avkKT5S54WIVjGbe+OTWGJr0Zw9mBNFR4Xy1aSTRIC3tguqLW49pzx0HSzGnDJ14ryudZtYF
GcC+jJwAc3pyKNBqQ+21Gn+3hW+F4dfN/Kme4u//dQ4XbHleWdTNwBo93M1CaCj6UQOXtyarzV0H
0yVh0yeQbnOFaQfTOQ2deYYHrYpY4HV2HSwB1CLKZ8ytT9NA/Wqdi+zORSzH87Sn14bfwU1abFtW
WFyxWKSEUoVhYziVS2dqcmc9bCKwjBlh4sh7M1wxTZzSesXkhA+1ysEJ8+cUWXI8PFqDsCsCsmSh
FNeCCGoLSkuYEz29dBMdEeWhyg//PUPnTQztwosabBAaLDbieZC3Vq3riBTVgsAxrZEnvruIkqxV
63U3QKQp4u3BFoPRxnpe1Vk+j8/mMxXzlRRpoQOBDHdVCdQ2/zTzNYYIXJESZsyJF3DH3nWNevge
Y14e3ScI25hHvU57JquUAbuk8hz4eBTMSyJLUHMFqe6WgAmygd1D6ywuo4A6UlatXOnkFNUm8M33
6ndUTWcFnc5jIiVyoZ9FiYO9mA3MR2nOGz2U1+JA6mmUNk3yHt0OaluIOunSFxY634xlVpQYS+BG
Q+06+M6sCBmZoNY9rIgtxOLzwUca0ckQoHlrwYP+vrqU58x0X6CphQJ8oUmBjX4YfdZ6ix7xpGbZ
DNT4j3Il16hERY63Ihp1XjlpEeYSYeN1PRC/RkFUmC4clbHFcTQr2NRjWmOF4j+5Hr/iEEfpZcuQ
BAxW0lez/3uvnn8JqTrkdsorgsBgqyZcrpBaGTQjRHtmhWh47UeFC+9azQlmbq44uZ+kfj1Dlmy9
4A6yBGJgubsPfzyhsgD3FRY1q55/FQ5am954k/CVojm+L10f71BATXvHS6dVJtVpW6QzzlgAEYHZ
APtrd3AkK/ZW2rZTf5FSiJDfFoAgw+V3/qvTTw6TVV6dgjeUuQMC5fYrm6galc0dk+xGCp88767Z
WZXN63gauxnCZMfDyro0MmV5WERzNpvbCiz2tYMy20JiXnM5OFajHe7AzLyx5DgajvnibmSe8HQz
+UIR4TdFijIScVbBZ9rILRSdWgsk4w52QWEXSX358H6yVDAj3RLPJ1D01BoQvRDy/uCvkDuAUcQp
3Dric02kAGOXa1E4HBrd1423M+FM2FeyvQd5TPpc/JVmTjt71et/fqT3pk3vs2k/FkX/JL6sBbmQ
EoqA8U2N42G4yP00EXImIp83st5TWy5wg8fP/LpsW5i1faCT4bf9hz+XwJuMNORcLFdiwcddoG7L
NUIuiFBymXDd+uAGvAtvOT6vNixSaizafLazGAbcAkzKji+Sj0vq0ed/hD3FAMjWrnu+elqIm9DW
gjBrHdjSle3pQbIVgSIwwM9a811b3YpvAu12TBjbI8oST1O8PK4Q6z/eLJRNvTBpxglbrsY26/X4
aLDEiRHYBi9pOOuKcC39cESCjphJasLz4/uwowZSAM4vLz4X6IEcJGjm5uQfaST9w095nB/Csj8N
xUsxLv8xq92yI41NEQpbKADYwaCoZh4p0aG77xY7mH8eJZEsV9N0npNRQBw9j4JIEwjwl9hBcKEW
MFBej7LdFOKZkIHWslxPpIaamBqsgu3kmyaUlAmHQ1IuBvkJqgOn1v3+OpozVfw0D5u21dyv4U3D
Bj58K65VoksOu3imuDMokD9hAVi6vYKn9vO7K2Kxcs0Ils6UrvuA26sD5wS4dBSL0htKJRf9YYA/
goOa6huNbBSgBYuStb2MIyykBf6nRz9pAg1WbqcgUZ7YoiFwb19PZ1zcKYQMyUWeySm33wjuZ9KX
9FwWiBufhjEVZKh2SqZVuiRnfZlZfJhvoEthVGvdKousSMa5Qlz2oyi2I1Z5M+g1TpkZp8qvVqKo
+oQ7cHq7z/ogyW42nm/pvlloWHCD5XqyOO3zkE2WqX/xy7sncnnC3QUU90UFIgKSgNPY1TcKY+8k
6iUHu7eidFSz4YeuMbwiyh4aNdCrfgj++JEEqts9zPLUGKbKS2oN01YAMtE6RSYpk1v3yxCjMfBq
elKfOhgL3/Bv6bgPKhz8Tz07dUtUR76tXEkJyhR/ifmYlZDXYs43zMVEfR0Eb49wySYdPoPqyR42
mpGtkmA++hcSMwfGmvdFAIG8uDOenkAW792DN3NU7IUXipOHID6nYfQqaqOhRzmCyTntXo+C4vMh
FyC1ag8nxJnYaDCmQbMiA9V5n80W7JLcQGUMzNNwSWRXLiMHJFtyKO4mJtO6OhUhukSSut1BYAkL
urxTrb+p1bCtp3F3EG0iYoiYgmxGOC5dU4rifaK2v5qpPKfy0dkFq/VEqdVNkO7bZJSxQFPp8HeP
QeUHn9iPMWLAbgTtQpUMz6YXXqnkxgJicHkr97yK0DsiCt4x+XEuMDXalarX8EdZpi6vCYHeJlND
meolTu+4hjk/69LWG4MXZ+rw52tKkJZ9l7gabZcj2UL4C9TAkuZd4bMZfbnco2lH6BrDx6PY+e/l
PwritFRfwT5abUr/WkaIU1lL8QRb4XTEnlVhe5G6M9ERRNXvfX/9drtHwd2VDqUlAZKzpQ2PkS1P
gu0KtLNMvD1JEZmxrogsBUMhHg2QstQccURxsT5Kg2t/Y6WE0NK9QSrq/DimPfvmDu+Rh4BW8zzf
WlcdhEyFBr31iBtiLeSJEclCPqD7H2I97a8qqqu6QQFMong2/MuDwqNqF3+vgdg2cISSDQix6Pog
eDPwN6oudEI5Uu4JYNOYERsN59ie7oMJolaPIGVtzTipFu4+1bz/Y3eC9Vk/zEz/DdrTlnfDWxHo
OUIHGJ7hVZ874gB1PjW7uBetqhGDheuUpyp+ViHmY6T5606f2T4qBntFNIZBwiJMQgtj0NZFvW1j
PGI6S/j1cPUkcmPuPj88GpX4BKQsjJyhDDRacqjh7qrpt2JjVx6ar5N8fixBcMAPHEBV9QMrhHgB
WBqSXSY0/RfBbFDzn9dzKNvcq2XwGHP52txORXRd1ZEewhvTl6rvaiquoYFTub6WIMBj7C8dAYH0
ZEZATRjArt6eZJe/xpVxqqnrVtQ0SgOxNXhxHUtyd3onM3bLarz1O0UvUj0YgBMoPQelOcrtAmvt
EdobIN587SqK10djTT9d6lcXrv2XAIx+fB4yAnS+odw/vXySSG6LSrn68gBnddiYWPKIZsi0A2hQ
mlDGj0AHo/fIgGE4uagQE1KTLvfsUD0jwyU0jII6C07S9a9IEHzOAH4sJpTjPD+x8PCQ/122rWsc
R8WsxAahzSBK8TcE3yKiSpyicpNccwxLwLmQHQuLpszeJQvIc/u2ZsNUrCYfKGzF8K9eZ+av6+++
TdP6NV4ImBBzX31Rej3fxvqIap4getaCU1WPbYFjMaZD7lD9UZsVeCgtxfNqCg4z9L2tyInC2lPt
QbW6S9Pz0Btz9fGwrVV3xXDNnRf8yWvvSZMn8xRJbxFEqFZpv6zNn1lXmkPpTcQDBhbqQeqMf9DR
7YAEifkiKC8o1jhDXSuP6rNApaWESjDCY3gxMFUZuw2+azb0Z9uxCFWl7jkEZ+1qkfVhgJc0Vq3F
Q02gH5j6YXH2pYr4RIGDF5uXqa/kdFBNyQmzPvoHw+EQaevc54iQUN65qLh+/4Rub6D/+PlaAf9e
jw0IDPCREDtDBCTnBEfhUmEWFTNN3GuJ13mUWUVlBmEr/YiQIFilr+3y8A9IqF2eQJOO2Ot57KpL
iHZwiAXINEnTlxIwl4Nj15uT4lhfrR7HjmWumqrRyQedWM0mlW32/lXT2/5inaX/OZQjO7p3iq33
0RFh5U4LGTV4t3eI3GMSVd+ugiMOFMMepy8CwokjkVhZwQ50pFWUWO2SNyaD/giiZrP7iUKlJzSu
oCHEfE5zlIKwor1JXB5GRliue5sAs4tsyV+yGPBTZnDJKJN4OmEAyoUiQpY/n9pweJDpIPlu2XPW
6V3Ney4etzOCQYUYb7e2sRXCSAFYZhy+GtSB2oz0YVf075WMNhxiBKE3aA8+04z/jYJRkeuVfj52
ThDD7hsWT0zAqV9QeHzZqIRiPASnhg+VkBIzAx2OvPDrdZ9ZRdwt3tJjrNfEY85axvOY2lR/WWVT
vz3PD53VFHJdhBAMYWLoDLelB9i2j55HDhz4+trd7ewku4czVgSk0PeFkn9ISUrMv/X2TfxH38Qv
pTkymJLoeL/zd3RWBn/2sg9U3F/J6M3U93OwBsVG6CyFWbMQWrvPLxNKaRx3Biq0QBChQpyT4f5L
iVSG8i9hVs9Rz5/CtT8OqFgpNj0aZWx3xbiU+lHUFWQVD7crgCdFXB9BIrHdoWIEQ1xtLrLBwUYu
h1VkV9XqpqyEAkjVuKoCtIv8TJXECXfGfVEHiX0gc9IEfwbWQfN+/v+Rd5mGenh2Rnf7iRvSUQmh
Xv8lPw6vwODQ15KB1Ax47oOg1BWCQgXrH962qwVbUYA/BdpaqSHhP6oN3y4VeFKX9JA1IpmJpP/T
LleAUKGWapOCg+mx0k9AzNeuzDyk9l4W1Bz+9tZojjHs73tJN2XY3pFVOALKHaA6I/MH6NjSV4b5
moGuR+U0k/f4P+v07OsD7F0XEfYUEIi8I8tSEPPO5KTB1vckRRfJerSeLgP0uqA8JxPpw/aUd8T6
/Y6WkC3cqqgcbsevHn3p9JnWgJz0v8sNXVjXhmGdh3Dp6hbOxv6uBHKkQZeBDnPdxHCnCzxbIwAo
+hf9pn49kqHtD6x98Lc6nIqYdwASP44FaWUq2gnbNMcXyu5FHrPjCtufkw24HHJjycCYHUilyCMc
ZYH43zKlCjUZNhFoc72RvRVmoiQdNzoptB3U0nTdxQ+6+xmztf4d+G0CmFCceuxU75BxCuEbuNbS
kah6FRNFQ0Kjy3j3iXWAZVs1GDXmL2wM21WbkaOuZDFIy0cWPml5fjCPsQet2DY81mDcY+RCYrWG
evBr+nYiaMKTh3fjrwO7+4zILagGITQIU9YOhR0jaJfSfUPj1r5sK5nhW/ty+RUFzzeCzFj34Y4I
fxV5rqWTh70iKkekD0Zy+7QhSbNt7GtFW8uG9i4Ng+QIIK6pBad/fQoLwK7L5Gu/iiVnMnn5HLup
89NZ1kW+iHZ4NO+tWr1O90U2RCdwxT8TThYexBUMjbOnnNRF0SKaTwTBT0nJaq5xuRZEZVbjyH5X
E00DFkjMjXYMDLTFxhDJpI5wOM8epmXlIE9eDAsw5AqTw0u2d90yaXD1S26LDDCE8vCILiISfUHQ
5im8q5BHeSQ4B3k0V6fe3gDZRJFyhhitVz75GktPnT5NzB+MbisNIkXD1vNzjr4lM+n22wAIJQ/B
rpyBGgqC5l3Cp04DNInRAj3fGsGP9zreNFSGHg5+fJ75bdaAzrSclGBlJB3JN3ktCq91rC+cSBp3
vs6PBXt5PK30adwQ8GHjIOqyucFHMuayUgAqOofUeZCwVxKv5wOVLWDg+lwgMjKTLag/nb5N0Ewx
mBUUhdlxwKa36tEPBrPVRaQ9ciBOweRzzbNtkzhEeAjmJ5WuCLlQ59nCjhYruy++UdyT2d7YLW36
R9gdMMJEYQRLPWv5RGrFfZdQ72KKaVZ1Y9Q7leSdiaFoU2/KPVNuIIYugTtXQ5zB+JwBZs90b+tn
+RJARIl29A06sL2rL/MQ5VG1A0uPBGIenKmGfRmbVoQPj9KphLb5D8/LRKEae8JcmcQyitQ8B0mW
LmBx4D30Az5E5EqFfd0DUeoNR/1BM/yq+6mKMfuoomxwpKsOKDH6f5gY1YwfrbqOcp8NRl2tHrwZ
RI/pxoGpxbWS/r5Cqk2A6JP0ALJfB5vqju3I9iZ1fsVXXd1SGIbc3DeSrX57frLIJSw5FYU1zjwJ
J32pes2rdbyksfwCzqJGfx9huOQQu2nSmxmc1TsNo/w6/lLdDEf+EtkK3eOW8BZntD9QIgxohfO3
3lyp6Q0QsUS89bAgUxwPeb99ikWJkPDjwmEjC+2tdoJBvJqdJBQtvuydRaBL/a03QY5+DLOdhmno
z1Oeynlxaet6PdQMTqcPjIbUk8mSjw5MTalksZGxE9KUNbGuxsyYnmiOCnpcr9D0f5/cqQlw6jCq
vamd5vNC0GiGwY5LZa1+uET45vatzuSjF8CTSjQluBaaFhB8OhsgPIEwlEDtGGeyqH0tVYxxwgam
+K7VqN8XeM8kHqWDTCUUPT/n0Yo3PqYGQ2sQZKtRRbtObsUpn0UBXmuOWjghXdGQqo7RMN1TZvqo
HObEdhqcfmQf70HbJ71dxxYA4NXLSbnTMvAqQSpTE4DROrVdHZziPKVOOAWR2agoL2h4zAb442MB
tkW+OlyXRG27p0qSA9MpPJwlKYbz0COOvYeY5sG1vRJTg3s+cfkkxynK3D5tVp58dk19DGdYTf0C
76yub8MHu9ATDyAEBkSen+yOYpwJU7PZUB0d0uvVNs0RbeGs7nGI50N0z6/GWS9U4lK0U6WvGL1N
6p7W55VVDMq/B9GRuvF1+XDxRUbzSAFKK1cVh2QhqMYsQyQi7BF+D4W//eSQKWpVCSsfqQODg5PM
NVjZOdydv6lDLhm75qwOygn79zB/4wnJwWF1eDFHdpgkQKB+Ymrwjskv0d+ltFLrqwEKF2sI8tCt
L53EmUUQyp4qjNDZtW523Vj38KTqskaOVnMKaH8Pte3tUPrjUZOrqOXcKs153+d27rID+BmG0qxj
XVambwQdSuJD6jNd7+yQPLv6Eh9GANKnuHn++vjH3GuEJLjF2pp0+e16EXXFTtp/Kmhv2IArqSGL
EP+TdICSgoqkU7PPnc2Xw8Ts/0r9KvKSZf6gekSKLy1/LAktxGVQcWq7L5Opl5Arja6uaIpEQAQ0
lBIWzYK1vnuknZ6ntIYyJOy2TvqjiGkevtrDh3DIJA21RTO9gEzKIPqUjG+7K0vb4ksDskKUMWi5
zsPiGcqhiSGubuxhzcJ8Ll2FUC5DcX04W/bMns2Ctr26WC8mT7sC+p7Of9Tut9zTiURkp7L8zU9E
PKAL1yYaLymh5riDMq8WIgTRlvAt/+YlMPgi94D/XrZwbdBosB6V48wGPM/s1Ba8eXGCb+59ri1c
ELzWEWuAMWc4JFETBl/HRfLVDznRnUJttF3z6cwgFiS0sifyTGPwATdkXKZujZ0RIGbXU36BWb2n
q8nj56SOazWvH1CVEio7/vyOosPUU2Du+FEa6CYoHLVckGTGY8dYflUAnfMq10YgDsohusjSKBBb
FLnxnF4k4Y5N+CDPW6QtMJAhFZHlOwJsxAIozlylAfqdTCEEYVvLaktXFTIML9bbQUWAnhS9dVnn
R+0j/WMW9aOTWS0tdCt17oTj78mFqJEzKxdafFG2YvqA8QGAIlI+Zbn6Elq7s/Jk8ZiGhCw3Khze
3z7ZCyVlsHZ7HZp/RayeqWlwis7m7JnBgwzU3pvG+OB7M/qpMvkeqL6aWal+LJj0E68RgMcelfs+
JI/f4Z5dHFINL5A1mA71WInhjimesLJ3QzbVKzEsw8qbInBe3UZivV62MKLXkSg53qw/P6mr/aKs
AWPoLASwhBI2uIEncSOlAPjst1pCvdkZj+ZQKMHtnOC9ao3VdDlsccLZK4acgy8GnDKPGaDycRLh
dMSUorCd1L45GhB7dCU06ijKcgxnKprLIUH1NLDeA6WgVkCAN2HcxwQf+CTpm6h3Ih/vJ6EBuABj
ULk8/SHyU33suCZbdJrxWkiwAjEX6bn/M5rRZxUsqGgdnmdfk1XOYuhSc1Za4Z9/VxhO9rSanTm2
OwT4BxSgdFrbyg9lYCMXSb3eVMO2OarfcoQ+5zrTksdzOoJEqNs0FtfreGSf+hRdgHyWb7osjJgy
A/h7Gifi4k6XqQINNVYjxRIzHXmk0tUO9BmoCWwpPXkf4iKQ/vHGpZZXNe5MN3XTRpLE+1wF7qXS
CnzPciIajX+oCZx59CcIDkW1HQL5IlLN+adpr9YiJU1iksBWO9JQs7lhpRAcEzRnpeMD00QcY6lZ
HZQfyDy26SyYQKl9pcFtHEFEmX3jE8jfpdhr1rs7JDI67QKqv8x20YLq7aoRoD2YGNVFlJ/4XB5B
rHh5eceQa4STqY/4YmRgK1tDUDE9nj2D5G6yhYWUA0n4c5meEIk/u3IRBn1Lj+CsA4OIDOJVZIaD
YlO5W8/3HtZDKaUXkp5tuiKRPgDhlGXQIUUxLHCiqPZRUimvwQKKFJS0rLkgXGlXdsc46Ru52e6Y
GKY+Jl1pZ1mHsFppwIDN7JHo0ZloLzDMwml2kTCpKBBZTjj7IfPAfPSp2RZ4raKXmv/oQSrtmYCR
XiO/Yjzi3rQ5xe4jO2hTw5Ggwh8xCzr5bj62L4psBCQo+TWhxkS5jwRSz6Tr61zIKFBjaZmTpgc+
iXpsGS9gUAzIpMk90o9hhnskM63u9jEiJw153YT99bBRrNrTF2Ge4kBYKzV/ZYiFBT3vjZS/Ypv+
iIoKbzCh+9k6sgRm65pzm0qC2iZ4s3o/COlhUAva/QofSMdVJId7g5oCbUX2mYeUbwU/YIbRWicx
TDkhRFnxA3Spxc6bvh1rKRPXSBaeHY8pmHEPa7FmUWs+4Jix3C+vpN9vvJubU0Lb7I9coKHhW2lZ
W2WRcPamTOQsYB1b1IHrphUYpHTbZOA/Mi8kWcT6ncnPUrlF0RqictyrGZpVETXyL6eYwwOS2htd
nINo22U/CfV/6wZbPiToG4tr6aVQ1ARaxqxFYxlJdWqbnRPwsl43Oxsg7p1NXWKgRCeVP/60YfDZ
IhsWhHf/SSXDhKMtoel/6itxYLGo6lvyqKM+FD3yD5NpxNol4sDwO03GfoGamNmdjotMjA/04vVD
iM8YzZSTId4qGq4FesZukOMQmg/tJtngA4/TPIJzpt96g+qxAb4TfLWuozOOU9VHwfFqgHWflm0G
bSAHIgZrkH+IL60fq+KeHWOviwLfw9W0inD1/r2IfbXQqy69ySJKPtNuczRAhm4EXIyddAX9n7Uq
V9PfUNxwSK5Ire1k94PFqlc+VjwG3xZa/LlEp337Q/rDgNTK2eWaBtUGY3KajphFqexiY6ikgL++
/uRkEx0qj1HsTVG3ebcHTS7xLcTEjZ+70Bl12o5YPZ2joTtT9KVXMPxK2aay59ijEo41FmmsOFUF
TPti1OzpLn8sJ+oEurQozpONafV/bzB2RwMdSojHqmnpCWeEF7DNiwVLghOQOl8afXy1UofffhaH
s1JsWBgajEwZ/doPU09pm9Ha+Jx8pUC3csuZzjkCPNb/LY+FJlLPGK5/7tkJmSobpYd3KONG462a
1tSiVQdVh2A6FRU0F74WBOuRYKuzdinxNa785FbKr2oNc5YAhspNsFoSl1fCREIxUbe1igszIIJQ
YB7VvjORxFAVg7C71hKANcTb51rJf24dFpCRkQdeiwgRtOc3NYNOvmvIPfOBoa1Za2YljBawNNun
JLFgVQqGA3NdB3jFfejXa3y/SWlsmj1YowvAwIB+m5vZI8CVs7RPeti+lxONFbCITNxczi7g7utR
WNuJSk2Um9w5v96ni8cdmbvQ7ctQRsESxQ7j1mq9sGy4StyhlRNKKDawhvB1usAd/sHP2Gr0UG24
IDHKwelZI4/PD6Z77K1OG5fOx68kK1TH0uOIritliLOr0G0leCsQz8WP+PakkGGY6xngwqe7SXu0
OZd6Bime+qDOkNM/EeCnIWJnRmMY2y4OZc4phkXQ1iP2j7R77GHjPk8PtNkLdJAUZWytasv4Hyhx
KZh4CACDObflSPg72/XKEVbv8WbGdEEz6FwI6Os0zBuQuZ8gjhFuDyjs8WBHwTFS/NujGgU3sxTK
jCv9oOfhNFOa+6bmpn3giolRWyGOZQNV9298b1VnVDUVlRcv0QpkQjmrbf6cby9EP7NK76zmia/J
czOAra7x9bI+qtFwi7sIYWqMtU6NE+WbnuWRzEr9A5v/g+nJqinOh7SDTHKjiyw9gk0htjbqtlkG
iTGQ+LrjaqzssBMFwP5bx2nR4Kja9SbuoaNhENAKnkkDNjXUmWxAdo4VSGT0Ki4S3zgxDp7jnp5X
eOZ2KWfKteMhGIcfazD4TM/eQbSZX1Lcn6pdcPb8I40p+3ZsJiCsRBxsXyFdRc+rRUrPxCwAMxy+
BS+Ze71nZz9Vj0omcKG0nNLRR/iaBHe30Mxra4Mwv1GvK6QbNFHu+0gtLdM+IEGF7g7hBGunYYDZ
a1QhMfuZU2b0ajaQkfJkWitaZBbzbXTD3A+MVxx0Y6RELoiJ/fAtkGusZaUHGS2pgdvadV5pmfiu
5Xk7xtbb2khmfX5GCCgGNB86TF6wjGp9hJpTW7TZkk//OwxykErCJ1zlZJP6fPkVMeEIVQOaQRgt
S0xf7/T/QeZVmepvnt/GUp8nh7UCnm9Wo1fROQslM4hy596VKInzwdgbe8FmuSfzqnDK0b1DF91E
lakZupjC/YDkqSr2fdUhpP/S7kvUFsgQFETWXKLYPrIANqr1JqJx5RSyaq5je2eJ1O1wVogaqd32
u267xEGGBrOQPtFDQLW7IMXuIb/PEa95zP+aJ3sYGdptrzmiSgmdC95+M2OWtFrhRFWe7+m71OnV
4IhhRb4TOh7EZIsVLDQcb+f9szeJJPJOy1SEz4RtcfehA4mesoVp7/55xF+SRvDDaUqHpJ9KwvNE
fnmI4aOiVsxf+qTrhdhitvorV83DuzKL6AiMG1yTHLljC0ERIDWIGh8MbD8P42dfSdiF98YKZrIS
/RDv/GMc4439UDjAENy07IY1yFU3emLh811Ef7J2cSkYyn2lApgzQhzOYu3SuWRmlEJUDQ0AxRZL
BFeLPbQBNE2dtCKBt44vPEcRAlKCSuVJPKyz/luMWY7Dg154DULwh6By08VAOxLXUAjh6q9mZmxg
udgsapqncRkSKMUqkWDUeid1FtsbE088RCFUZR5C5Ao7a3d/J5h6Ssz6SIWgDIAAJi2HOFkl6OsO
+EU8kIKvNwJdTiu3CLNfFh7B52uCPsv0s4Qbgj6uBhNbtczFVNrfqbWIZWFovTxz7ucqS0NiP/od
pAq1G6tOn4Xi8AMotS0CEISTfzlNruKE8zeOyCVO+++4SkM0tVcwCNOURo20OiEixxlN1rVVLpV8
VYGej7QWzkbzrquaap21GnyNefQcjnIcV4QLbQYwUoK/KZOSxIglKpKMX2GL/RSllDE10eZkQn9K
eVXzyVbocZFx2lSYJBhoDRVvW/PYcaygqvlGu2OmE2lyh7hlGd1QvxSXlY55A70AuBXQXgZTkNZk
q3mJQA9LNg35cIc7yAFza9yVRUA3UCvIwphIB2BA1WyxqGIwu0RgJMiiW4PlG6ZRzXO2y6FHYLUW
shco/gXdOfedhqQpKkNTfoapzHY0V81LdBcsMShdhuROjckVX8rVzMkrlo2DoMKg5IWDyzRP3Dfb
rXLzAqMex/TxA/21u2D5G2KxMwQ541o4Wyb0LNNccliU3+D6jQmdFgz3aeuJ1xZBfLR5JrxA+6BV
67P9btVUQ8Qh5Wql4x1wE43Hg81RoNDttd82mga4BREMCQCmDnrcS1/qkaltjrRdsAvwSa/US+1c
BMxbxey9UNSCoQV70dOCTXuz3sS1WPBFejhjs3VR8e/NPq2tLWF77vI4dx6OVRGe2clQzgHi/nSn
cHTIre+TR9Or/G0NmAmq6mOusYkZEwK3kYdzc8p3J8l0sqneHDptO7bjDquKF7Jub1RjDaRNk8Cg
iHhmJkD7O6p8XjCnIou0BYVs8+KbvhoqPn0L5PMpSoixnxoSNpjQfiaz0WVfcUQHeO+0D2AGwRB7
xHab0ejUcmSgROdzcrz1AqtpOFHoZKTxhpvOOH3Vhz6LFW6D33LSJA9vRviYyBjZ6eD0sWrqe4bu
EM8Ge5GghBsTGof1qkJ4FAN9qVWinWAQllH3pzT8MxfJk7QBwv1WuXNZhHWmEm4UyF0rk81Tt4ni
ojE7xBjIoge/2sukpb/Ww/aoHlQ0yYhRDCKBxU7QQA9AmBiGbsGh26nMmv3IANqd6H97PotZSweL
yPcbxIMailKPQ8BQ8d4Mf64wjEQIIv17sTqOYUn7v8hkBcoLDIaoszT00+Vy2npIaVlO3ZXlRzbY
cOsarGYkN31ZOuOLbV39a9MCiHmuHox2V/zquyIaZakQgmiMe9bXvWye834OaDY7vKfkZE8HXhOb
cKMHonz6pfhzNi3VZGkD01S/l7XJnssggXB1NM626mdtm8B2sVkoVaVbcleJanwW0t3Fw7Jjgai/
FIaaRlJvb+gS9VTj//MSHMhx5hPh+PXPcBJjA6IO5XG3p8l90rRttyVSxRAQVOtWhphlCBlzS/pW
5dsEUWri7YO/ZCEZmiQlOZQyfPWdbdEY3n9GUol4VG36yudtD2/hf1xiI8NhfLFPKoerFfsAuaJa
MhCovE9hh2SoxyDOsJPnz9BFzwOgpUEfDJktDoyxqacibwOVQJbgxjxLTRzHR87b5AZL9B9M9M7v
Sfzf2HDpGomg8a4To1v/YykstoUBnWzmQGFjmLUPc2nJD9AfEAxdG6QpsTK8O/8vJ1pEDLEE4cnb
i0h9Evmf4696FItFAAPflcu/8dumaSBLilcf2aOo9PCRCRvXyV8WLY5E7+NhpCYj4tvt0E1WwhMc
IiHvRGPUoE4+g6TxInPnOp/sv5b2N11NDKOsKOQFQUXXPZDVWVKLXTyW7YH1Qf2l0HmoQOg0Yzff
BTr3h8gJAlqukwxSoXR6rZn0ZkXrUVqVFr1eAIC3g+dY3iUf13z/dp/o+iorEYHlg+uH8ibsP5h9
qofRwxgsXS9JOBb0gwmOFe12RPReizgRcqMD0Q2rvMaCWKp/a4oTTGag1EMtvjLyONCNCU66cqbf
0xl/Nmr0y4oJ8dmvjIzAtttzD0Akle5XMTrD9fZQx8o+btArjvZHeLBAPifoyxl3VHJI2K5AfuNY
AKYE2ZejeZuzuVCpNbR64J5HI1UFqrzKmImOkNtTIL+q0NSgYPQBT6YyLQtLFqfHJgEdTUKRfWIq
/ottRomj9SSViaOfEspbtHALO0Mxor0IO7TlnaijdZ0M5oUlV+wMjf23mCeU3HgWgBwOusrVOz0f
xjao+s0qkirX1tqrLF5NDMbrXRmmRRB+8TyAnn8smNH5L2p2HagfKPxW/ghcEElkhDs/vOQ+D7pk
bR+gq9tz4iS6LYKS2t72Kt9A+hDu9+R2HuSC3JMuUmiG4mf6OnHpXkwcOa554iC/VHM4gpTQv5t3
FewZ0DbE8lPysa+6Uj/eDpP5Efz3uRkaGI2RrEWMAp0YEmAbPR2Hb4R4WpVd07EsA7j37S5qIMaP
YCSEHvooehSgDTMScVP18+BpsgHZcZhyBenfni261vpf1MGlfy8Y/h4lEJyBfyTSHJ4Q95XL3Jfe
U/yGhwzJxcKf5IMmkw2rau8035dFM6ovzgBEoL2hMcsZNl515kfcfg0FH6sWjOhTOG4uuqxx2te/
x6jyyJpSPYbQLtyLMkfVEAhIIdklP+3kmPFi2m4l+8+lpIvrpXGluuxV8zhqIn+1tfPbpTLzgq+x
DKEprh+Se8nurf9ZJH5Gvj+nbg31y+z21RS4DRsrBpJQAKGQsr6K+FMdtoSmhVYeqZOqJARdijcM
yj1JaYGVJpBMgfopBNBY39LyR3nbImBndDmGPEE7nEmP1mixE4T1qGx+3ve03cw1fnR3XtwzRluY
XBAsiwOZRfIbg4aKaSJWix4UgE795GKfCsfxE6V+BvlMorLSWGkP8mZviCTye8Ldd83aO4stYY2O
YEBcGTtLDmN1bJrJr1wReJB00tSChZGPhyZbfaajz8yLVfX/xNfMW5wzbcdRTaP9Jn4LULXiljLs
s5HNOHdVXyBmls/vc3pvX4a+rOCoevhTshXknEK/NYBIawiSeA/LJdtiWO/qIo/ihjjq95MGKk4X
T2Mgnx/ga4VmPsUJ5ZmK33z3V6gInPPPszt1JfBH6bMSZeccExmxLWoGg4LW6Aiv2NIL+LI1j4oY
BYYOmaxnYYW+RhVeoJoxCT+6PUS2a0UGPUm24MRwmSpzvJLK+S5NhzgQ+ur3j67BiG4bCCZaYsnY
txkXIXj7Re0k/t4u1CSxsYmPighzNsXTiurNhc440GXCB1r0KUWsBjlG6bE+qYBzRWYB74vPIXLY
88XUOzNDR+pz2eQEzlEAXVoxCr4hKLxTbsrDOGPmuytt+vte6xFJ+ubml3YbkBr+wFfYXkLdHnOV
8h1vtUVxdg3m16rYG6u6M6rTC5o5T32l2sZokMhfOF05pUve55huPfUg8q+oi25l3BFYCneZ8D8/
VjJNOZkYhOTKilb5suWq7rqFr2kWvUoxee9NDIL/C+AoeRtGl/EDzeWbzS3UuUly5QezBzL6Uxrw
ZxT4g3YloTv1K5yYyffRJLKyzQ7qZp4jFPD1h9FizrvfUwmsOu2AMmxqO322zWaxbTMqovM7gR/+
B1jrcUYa0vB1xzEbQTC1YDQoaQXh/1WYifeQe2XJBqLHtUy8M0VkFnpf/HOkUtrDDAy8C+hngXhx
BFH9M+STv+LZrbkAXwbNXAER3EIRZZPZw2iPM5Loswx6FahgwLsG5k6h6HxgCKjcXNW/zCc1B45D
/3M1BXopjkaEub2b6z9EXmsRC/YYdgJXC99S/8keSuzwdFtlaLn20jb4trIqsNiekMyBJ/722mnB
7i1TOTRv251Aiu3LZPwzOmn2uPbei7KjotKx0LV5CXm2wtUZnqwM+FzTVmjDGXodh739RshRB5qo
Dbc8EmWuErR+jnD3nU9ltRhtHhH4o0r12Q8nLWZ1zvmXKvvJ4gmX9PZIITelcPTSzyghQJ55eV2N
JWETxh+WXA+gHeNtOzKpHq6rj246wI3Kan4doJRqPtuILqrhDv/fx68auYabS19JtcoEipCQTBgW
whtia9br7rvdLkgFDBRE+38LXp0IYEJGxB8rrgpJJ+q7ZXcl+EjFnxHtYGE7MUtkUfkS+/ezSeXc
ZIhOy/6uyThftEjtKkEktRhrqOEMz68a8/1eVAUp1DtOQjwDA40rYqhtPGxXxKdOajq6DJRspqHm
VWpENXjqifqpunVUFaHhwTYT58SetgmunfuAICiyyqpcByXtySBbqR35e9+4qnsXeWa2v+2KHaK+
6AjdbUXAGeQKa02+hNP56C1tEQEWNQ92Gp0pYv552whfGYi3IFxcU2aeF19Ykx7tiKUkzX3234Y5
yoZanWjw6wEmDrsdUZJXlcl5UmNh1RUMPdw3xVWyidPjrFCQfUSAwc11NQYvs/KmxhUXty6sZxW2
MlMpmx5FLwrMR9Z7I3H93LctxvhjW8vjCeDX7CCarjPcRpRCoKExP5cxtbxo95QQUnBLlR+ftfbO
dlAJ8LH5zvXSExFDmfn6WnTXb8H0EPAA4ez4V4+YAXBj0FxwmpCkaXmR3UcE6a8h0pXRT5UMndjy
FktpTUxHhoavJAbW6I6DmO6w17jKgBUkRk4XlAkw7jHkLDJSLe10TYtdOJBZCd0CEXu8r3pbS/3c
Uvk6eDpJaAcIOYLdyZoBW+EeJlPOYSDH/TPOW4cR4cl2cMcJIObUJXraeTYqeRHwepValKPKQ7FW
LBYypS9lsIDJ/oi54MXKo4Q6celYvoaLOErSy9rGay3pJQkKyTrZDTYt/ec3byD72cKrmu8b6wdH
aY+G0Tiuko6yCXIytdJDDAtTZij9lbggsksQvAhx/A9MD42bfSlR+66cHZBwpWHrHyUAuPf6+lAM
N0aKzu0UsKxcf4MH6H1w7iUf9XrDlIawXM5uo+iiGQ6r/JkC7Qcninf/fsxt86AgLo8KnDw1sTOB
CyjCwh/4ND43z5NbK0nLlslcf87TnQ1oMXdsWgFFzAYS5LvFjJxdT+15GUSGS3zA712JvufHfqyH
S+aZUIeJkBtNFVLOuKaCWUhpsTY7ikPIKPViCrcTa8ralEHZvCo7tfKepba8qAQOZzaVOohcugZ7
fUA+CNl4/4Czq8hE5/H19xjkVRQ44IBGoSnS/vBP5awDJsn4T9htpHLV3JnfBGUyfKV5pF02TdH1
IT9IAzwWRCglwaFdIu/iDRmmb92Xg5HiA88hUbwvR6+o4TQbuTRTUMqPGr3KoTnIesfCQ+es52xz
go6WwFpwMnH6pSecYGKnNWq324JJ87Xm9J3DCGseMMCrdbr0w193LxVPy6KzdJv7G3qKN2Rg0cBr
iR3Ts9hlg85YnkGypjn//KN64srFaEKfOICqViwSc4FDcqXm+skwe1pY2ak5+nNBSZvAmXiODB4z
2/je0COT+/abqwvTgSQ54KW8q9t2XIizqzYucwjE4MS1yxZGwMc5bkdqBpXx/zwUnyKg0TWpxLSa
h/DMrrpSQX3qttPDxjvhlaCfcXJfRthttwUhAC+dQuqJnRDXfZZS2EquAQ7gGn7RD0rcBwWKwlBV
FmxvJXkft3Rgh7xc7k3dxdjT7aK9jz199gpg6c0KGdnShWSwI63W7NnQXSqIOLGmfVic5mwrAulz
HMmSSe4oIvmMboRhqaigEPMLfh+HDXDwSsYmYA3YMdLoHxdMtMtAydWgLcxd3p8JrrOEzIz9Oeeb
Of71Hb3/keyLn/0XddURHlhnMNkIh0diaD8pUygpHW1lwtrHkI7RYYg9nihjapCWQaAdGjt0POkI
zuIUAesQDe97uzUhJQkR+fADgVwSn+Bi8c5oBXu7KGeLQywgI+zzY8CCXINCNppQtlC/WD5sfmax
J54ukHHHvzDmUI3CtP8PUKTwYUJHE3HMRAcqfGfXgLZh9Ew+clhqRDtfMIcXcHjFlBdh5Pvhl6Fx
iKfjLUFXYn2xHjd/JA/m5l0j5V/3OCYNNL3Lh6kAeqr9YwYkguVTiwm8kD0bbkTzGe3pxwDKn53l
a3EQGH+H8Pba19m7YAdz8KkQoDqGsKkEFiqiQSso2eqoWWivgL0YWq+5NOXWOeOrRvSq8eyiSamf
quYopewgH69glll7FIF+9NhQlEtQOpdlqedJhPpb4JExXfzLTA6yhtJjMlXunHK6WkUH5njvuEp8
2SXG0E91TBfIFbgcgD7SAr0G3u4epmFUBrrGpftleH2hZF+xhj02rtXHVNFzbqgBncEKmRaw31Av
3YD1zcT0dEcZe0pHrqo4E2dOx7+A/qy9hz9o9y+nytxzOseomxUSncfG56zwMWbiX21ViIVlXvRY
05Ywueb/YfZjLk4kW/AWEIOrVKFvrYDDI2diGw/ZS3bkBO7Kd0i1vH5T2okzaVEa1dm+6Gk1guEf
2CO7HZJs8I21PhwUDJG9uPPb9AHFeRa5ixGDvrmzMfjfW2LvgUl6jtssbpbPV6KKWcdrbZ6v4F2Z
0yfWtTy9zX3EnCvQ2pMtqCbyB1ghEBazXNzski939u1SKoPKxQvJO5xSQq5f6Vjfa3NSU6sVUeEE
kq/zir0vNg78nX8/4ZeTCGTYWcPY4QKkUow4Za+T8Ai+EdCB9XB/L/unAKCEr2M8PO0M2re5pra2
Bsc1KpR/yOGn1x7UJ8GRVjx8F3VvM8plCBUSZiXP2GRWPVU5IwVEjZ3dvDK+Cyzf/1TH3/FSJ2ov
V4TR4ZeAAFohkNrZVrAB5Ip7m9g1jMYeZtqrCe5SIu3orG/m+I3luro3GDGErHbS9mwGbltCWl9Q
nT//cLX8e1bcmHiGzR8WEEQ89Da9W8lkxOGnTnE9u3FNaU9/qTregAlnO4yrDA3h9OMUtPQ2Y9sb
y/w+nBHjy1R5rDwn4m4N1BL4qBCR6Th33hlAwOpHZNoJXq3SoRXJ6BcbUXLkHPGGBzY9ITAWxG1H
XI3+Dzg+e+/6GiK1Dkrv12tft/iAKgS/AwIXuNQ60gVgcC23HW7Ql/xkGePmRhRkKZAW7zMnon0t
16wokzaA2JkJRNKEdptNMGiPkJ7PiKCsw00Lgf9f6oNEkdgMOaHNSPSQbnaR/DMCtKJN4yyyaFfa
GDbFgRrTuPQZS/GBPPh3K5Tl+bTYaC8cns1+yW07NNUWChBz9MgUHs6VcDA9NFQGX+RuR9B99qRV
YaSgYoRiAcy77lXPYaoSNQmjF5eqTmQ8vqksEI7q8S6BOuTMpkIkNeEMZko/An9qs/v1pt8V5QEX
V9KlMcC51+6WE1yGhX5xJvGQQbew5BA2FJpVO8AysG0Upg/1TEvIV82OTZQZ7miqUlqoWkXYZVLu
I65CTld/4puKkiMPpYYf8x15+PIrCkT9vWHFBmu1jOnlG6FYDo5XTE8wXAu6A1Gy+f/Fogo8ojYC
b8CFkIGh/e1sd2QDRLqDOf075CGTTtjjfOx9zs0kZ3vBj0OPSh5VZ+LzRPqcHWOhhRwQ3tXVn5wb
KnQzSvakp2dMifPl/6b3pcEviRhK+Biu2oJix/YHYdhscSHoeHdxzhBpqgAzzPeFI48UUVJ3v1lY
OgLDowWwV2qKK44xBcBO3JL+6yzQJY252T4XySF50AwWPz6Ui1sxxnaeViukZovqSG4z0faUGP6S
vLsHueoEk3VJLS+thmyQW/V7vMWsOgEazTgwJrFcQ+RLy5iqkAnKCoqJ5Ljot95jqMLsbW6XKknA
QKZjyvZX8ijY6giIP8AZX8JdNgK+myGNcNFFg0WiE+ZHWSzVvsci5xTRgvLCF8EVjgZWgsG+15J3
/rrp6jBnZJwYbcmlffhpHjcLkcKGljAuPqpfCTvqe4Jr/9A6QnQQdNWavFu7vpMHvP2BUI7VnQcw
EIgUBtcJ8tKq9A8ia5cV5+RjMaYg/RQ57KuQqygWt0TjtVSknIFjJUFGhefrUw4ZOO81YqSIw4a+
0p9kFH0eS61n1ZLzxBP7fXIBEMSR4f4sfFfFuLa/MnmpWWTAG1OdEK6j8muY1Qv8dtuupcK52jWi
GGDat1G20NwYx7kKl26ccR7AGA5T89ZXvsUWHnu0Sy/NpsDXWDYoNKgFS/nZxeNWIZKRlxM/rBr1
jauCMgvfKoMXLNlusJ+TbGsyzRg8OU4RV3evyeIctrkJS9F+4fpPTaRtglq4jznnuPe2janXWANA
95CJ3dpyLN6Sv4IK2bjN5yJ5+LsAivgv3z/4yRe8O+vlzyjFCS2Bf44HzeknYH9BUkKYp1yf5Zfu
iRyQv81JD5OgT6tBviWoJLmc9hH7p2OgBLJbiID5r9E1wgpiOOl2GemGRnfIiI4PhBXYBEwtbAC5
paYEtaLFKO0L1yRvDzFXJxSPD8b6dvSISX4xwdH0AWrp9BrOU0DinO2Bz0HIaL3rpZwjBY2UFHn3
iZupcvUw+kHajQDuHNeHB1OIiPtosiR39CS8EBdfakdsDaQsxikTw9nJRvD5M7L57lyFK0m1nQqa
P9kSdf6DGcXW4eTF2v0Iqtc9mfgos+xK+8ACqwDx6/JEZHJMtQ4uHSH9aVER0Qy0YIQQj7ZgzHzm
91ffS7wbpts5vfTgM5PPxjp2kFeqsI2oY3WzcYWoIrbjh+JWWnCOAF88FR9wj5Tt0CsrDQ83Gzg3
avge4XGF8U12CuW+QCeEcRuw4wd5GG7CuBNJjNSpBwDiatbNtJEa3266K4BQanCkr1GNN3zh8oDc
UsMTZHm+2LuhY5hwXaTVbhxaJ3BisstH6S8218vUjuSfyn1++sm1TfCOVBHX5ScN8GdrPqLFrw+J
aBLPo09JJV2PpynvL0JafTrz9jLyt2ifB1xaWv2EGJwLSZEB+2rDVSjKpKESFDzk90UcBLq07vyT
w34ExDX5Pi7ziIXdfwWLxSaNEvpoy6VLuxIpS66pGNNqHTddzrytfLStRR7nX+ZT0QREzdzSDtnF
wNuhBHv0ZR73s9UuLlS6hPSgyveja8wEpn2MW1Cb9sNnx5yfJ0a9Ot9zQCvbx/Fdo7Q0fCY566iS
DlazaHmtyg1Ks4evuhHK9dzg3ed+30tnAvNhEhAyPIeVI2/qefVfYK8XvcXrNWFyZjNtcQ9MUg9t
UATtH0IrIHLY6wVXjrlgXQ89jF/SojS49pQ5RzCZgkCTpJU2N2KApCUSYwViOcZfhihxVEpU4FL2
QzsbkP/4YzkWFRNlbuiVOTgFLzFKY36G90W17BOsDr0xrN7FwzzdO0pM6z2QVL10N2K99rq6CdPf
0XihkCg6Lb7q+2bKtitCrGZDXecU5T2YIjn7UHij/LV/gKe6eOfehdwC7QoYuv0PeUriPx/g9MzX
sapsPKEn90qgbj6OFm86vpiJXAz6hSlWZuR/4ppyFHfJybQVrcX2ez6u3/R9QIApNA+sfC4+gs59
il93xvkTaYAI7cNFUsADwR/b1+2O55or019tKRi7YwGwQniBOrZwpc01EPHPWrg2kUDwzAsDPJB6
8DPbg3MT6AQyAvJI5nKQV0apeEvZODEO5nW2E4iU2valAFUtkDKA+bOAu47uCgrXPMZuSemU5+R/
WtaiWOUV/0AcTgb5sw19ZRwxEIc/aYvKpdHO8qTwG5c2U60UZ/Kc+Kp6uYfYD2fLvSTVkCLgyBXh
p/i9KsEiUyc3GNen9SmJJhPo+uxMfrYJMDaG9QtbNUVnAW3sRMH4UX7kDxQZBVbcVdKfBVlYfzi2
aFK5VUsJNQO8dh/FKnDf5xSQvdHPsyh0F6X9Wq1iWm8Fo3xJPlORWi0SRrHVWCbaXfYkcXenfHgC
hB/3/vY5oGuIcWDp5SmeDI8w7FZwY/S+aX55CIU+IX73NdfPvWa+EN6JsXwtB6NNDtYCKrSeMVlh
4E4zniJJZ4xlEchVnlMP7nZRMCu+pw7nwDnGg4LqCIGIeEF73xFCifCpcBqzcYgMAfacpwLm+HuG
rsIGEwcdvzEG+ZR+6aB0sbb/he1E1Smojpd/26Dnbn0ZRqRN5FFaQStAu0OqvxmDNnkhYPi8YL/F
1Np2ATBqhtxDfi64OzJ21+k3NqAVZhtuTE3F68/ox6H0Bi5UscMvO0nHRn1cWmK75bCkjC/pMRHI
p5qOb9xZG2vZWUHxgV7bKk3xJWRPNWVIqeG4egzaMUOnmHzBiljnH9MpnKnWHV+bjpmCi15/IlZ7
FXf81MaVOQvGmUTAU/YwtcibEAn/H415La6NHI3N+ziWHf/2UBtlTARfVyrBKT/nZF/Zohn2X9Mp
OTvbTbVTbn4ipKcQr95Iy/DXxnhpQS+3H8UpUYI6YAN1f0xVnY9uODPInHDlerex4VuKZcTFfN5q
nzfU3T3ZPoZui6yFnc5JgP2Ok0JtKWVPchFv4GMHHE5MQQ8TfJvAVqlm1Obbb1KE29KYIbj00G3P
xr6Q6CkVR0E5lJTdE1lsI0FhrfWguwkTbupbA6aSGB4yeO/2QsdzVIvfL69IuFd4nl/jJC5qLrN3
XXEbzTJrOAQKohQR10GEyieo0UEX35/WWjL8zzyFeaj+Fc+//XsBI4Sdx+GCcrUOsDQMf/QJkHzA
IXCPUSQCLIBqx7b5LsvxI2WTiclGQQGAnX3WXgjjnMS6op2va2fmd05vz2j2P4miWzyleBkww/HO
HsdrK78azz9B0Umxs9oF89t3ysuXcafgD1aVjg6xBVyYMib0L6zlzJFP/M2iuwlN3/7N6tdlU5in
F0HgHaWRvMZJfEopf1KeNmxzpjEERnvFrHbC/MUTDmVnlQ2sJWBMj3szC1ezDsN1MlIYbdgaQmHe
bo3VvXZTcQnlZhpEMHPJpR/m/PQHCcuBshbwFJPrrOSvzJFWESSB7qcAxUMUbqg/eXTKZ2kBk87e
mhkoCcV0/dQ61B6R3ZPHqPii77eNL7saKVlLXscbxzoPlm9oOV3TgqyDZOztRMm9yw3jLxF6dQfP
U3mnQkHdkGJ0NewIloS6eD5OdDWk5vcH7Tw7ZG6MQHXN5SaUsXSMLKL2Q+PQFLLAcFzoTKmq+iIX
WgPvsdwcwLC8+GGTFEx3xW0UPTJKf9eBTBw+8YG4yN8Cs/vl9pNrudzSQsUtTh7V0yz76MBwK685
8TEmqBRSNnuj5LLldIRLMR1bpYriESD4mLz+rXkvvio/lJB6H8pP0kVu1dHqPJx+ojPfUlQjJbJh
4DQSvCKvq0o4YCQh2O8rZxV4B64H0lSEZCvKUPc/YyaoClXHHO9PCvaaUNhvDLgftzYFtaxEBYdx
oKFNiGVvWxIoynLkIRgKLedVewQrm/BclB8EoJnUWVM2MGDF0H94OzNEsCPXoea1OOYBSdbg9Pbm
3miCFsoAt3y9dLmlgzrRG1RSlIr6a9fz2lhutHHago/exjur4AEqkFvtv1UsFBjAfYGWzS339rmy
hiH0l/Kkak82bTvFH/XFLKR0MIZgxha13FXdB2V6XVa8kmH5XG8AmyhDTznzQ2fi/t+JEEZjag17
ucacRM3W2l/4PBHuP0+YFjzja+Nn4kwSFJ76WZg1e6Dj79g5Hn4338BbPf7yssL70GxfrGR19P8/
GtlTFQ6xu2EEHvv07bNHdGNlEupMTjvC3CSwhKjH18ToS7EyNrZheMxk5i/90VyIg+tXFB/6s4z3
RzWx2Xg7uUnZIIVhsoyasbnL0JjPhnxP6P7plg6H5BskkknCtlI4PgutJY9l5H8t/fxknlz1IVyb
07d+kT28KehYd7CS1952+Dsl2lkbhGrAw5L7pa4J7/MhFoIlQA5slEPun8juAMRIwzKYt32ZV0wp
7/gBeaqxpycvLrZNItFqdBRN1Q/MvYWfiE9o6NOxEBI9XQnJ1pXLHRSOJt4W8fGZ5xJBDryE/rA1
Ld5enj8pJhF6VHfWox5tkPdRkqoqefPygriL6AMpcB89j+SnxK7fDqBXU2tM1KVyjpBq/LL/ilAi
iuVgO/nkC+wawSnbSqD7e+jQ/M2FNyzWE5pby24FIk5kzmMsi7bqCcqb7sE0w6//8NVjIkCMG/eZ
vPJm9Wf+mvpuSjKNTgyRCzfsBYOCLExoac4SzDDtVCURaMfKJjlAldW6YE2k6Fk47w/0JpmwJdSh
YxbHs37NNfUsxG+RUp8UtdRfxmNhJ1el/5pbhANLq9R3bpc3nj2hqTJiFS2BpoQc7V+8iBXfdAgN
+tNRvArfwSEnOfYVzYLwkVFHvicTm1BURERe7BycVX/QhMf9dbTGgeUBfm7IuvIuajtirSJqfB60
wuoSjGdKQQKpeQbRs5yH2ZOmLUv7igsc++wDVJfNBUwzo+zd8IzkA2tG/JNLrkFlk6K8qmXMzFHm
5r44KmWfAa/G4yMI41MTcOHm9TkXDw/JPR4RtYOQ8ofE/2PUFYOOE+Kf7kMuvlHfCUcytEaBlBd/
5M3vJ7qNd319fL25ubFQy4OFORJlsArgW3Jr45sbc0KfGxUowEZguOVwFpz5Hg8mqqhopXFCAxIi
D/wrPWoCJfocTLfsNxDQIt2XSfvJB72WO2cuzM1sEa/qPwEqt+k+H4F6IPAHb4NjxD9zZHZo/xlh
IK0WJsxTwyfZUz/6P7OcYn2qBHPMzJllC0KA2VcUDACu4qvIohVLw3D7UgGWrHcVG2n+w4z1uME1
W32342BGgmMn/ju603da5DNbbUQyTx4+C3h2nIm3ft1d4uZaxVTGGr/c/GY73EMo9fYl4X8of2YQ
v7ZyAYNGrY+PccZzDYdXuCgprrls1e8HLgA3eXnY6Q/oa2uF0JhOl3SnoinkRtr8tyhldlW3vcNM
Urf6jkixrChXEn3jEAbIhwIgaJvM5VO30MPiU1CB8mrqBIfBFzDB/6qwM8APLkX7RUFYQ7fDenbg
X/8O/MchAIBUQQWmxzQMf3G/T0NsQO5++r/YWUIyFFrmOV38iPXuBoH4YpbakVa4j950t5ZVmbBW
6IafC6xW98ro0zjFIZdKK4MOaa9WBIqxQIRR3HJnLHdBUA7qfxMAdQPWOFozXK7kfjDvHipVQa5+
Vdfo+qVH1JL2TWVP1RsdLivYPohv5KrnJ/JBqD429TveG0M7PeOJAvip84mDwabjy2/ypdUALgQ6
tBxyo3HirRLfHgzXuq+OjSh4k7Gir51CRhb8GbO1NHZzGULDV7WXKNpHtesZAFis/y52xGI6u+Oc
WFXxAOTgSHMmuhDup9rrt3TgQ5jUWYd3TO0LUqlks86JLaLxinoL5GxMEJb9CudFwDi/Hi1HNbwV
Vc6/XZWg2+rj0r7N+u7arj3YvxQuBYR5nIvUiAYSCxk8qYjqVEnBLgwmHZlUK3VZOQZahi0SYYs9
Ycsi6z0GpVLEbYRL7MCWOOQvkD1woxmM2Bjx/4cGO7yaV4bGTbO3FeOgLiPor1+FAp/cr3a8TznD
C3gN2S3gqEKFYEyO1ueqK5hjDUE467UAGTDyASjetVPFVjNBtEyNqXKiz8EbPyujxjg0E045H3Hx
qpFbghZxg/lC5FPK/eTNK/1QeRSALegn29ukAHv/Aomw9UR91vXBEdAo90YA/UE+fkDmif7Fyo6z
+CN4YomvRlaeZFGkjfgdJ88lRwlIvPZVQEcEHgiwBp6DMjsxWY1RCqrWd6SV5Itri7kuHUXhMUGA
0XRP9JCWFYX29smDDNGx1gK6Dga08g+3L/xNJgoRqkz89VfERxiCaJXOL/ycywUC5qaw5DUlQZZu
u9DkpruN4ImLKAmx3O1j5JGtY5HtbIkjWZZhNGqzeuyjET4w6WasIwlNqCTrz3NwAXYGvZK0q7oM
o7mfIGCmA+cGOrJfBS7CmoMqVzKDlrt+JxYdTmoZEWUm0Bq49qPtvQ1X8mgOtV/2ejDOlh7Te266
j+wB1OukowEaezcv9vpUdaD31vNzzAhtVcXxzHRwcQSx0oSigAnFX2zXlMdadIK/7J1MVFD2P/7M
oDuMCVRrK2XMArUmayLPRUFLwQ0DlNZqJ94xFemf7KnZsZvgZr+bxjRdDYWP88TExdmRiVYfSTXO
EqCR+lGJKy99dJy7Ort+ai9IRWz79yrYmpD6fIAxGIDx8IT58DXfhHj5bSFRJqco+ATWihKP17KI
IyWFoOZdLL7c+q2Xyu9K3CdEDn/9txuhFZ7KLDRbh3LFUQB+Qm1u1u/Xc4bYj8mIMKtEPZNQBfzA
WYNy4RQS5JIsknEe1mHh0yNBW8csKhXxlVaZBC4jaLVo8LDTDMudceoHD3MMDYh06UGG90uwJRh3
Wx469JPPjmkh445gR79tOVWuINUhbrX08H/mcYY5b95wOa4IZ/JSatH2CEYi0QxjLv3yuUV0y1X/
jJ9kiKhaVntQ1WWIX6k2SthkX6n6vBwBpFP+n/cdABT9JfSefQqGQ0rcaaE8QKtSwHHg+Lr3Tcys
WeXV5MCYM7t2urTPYmP0Bmybv977Kc1wiomlrmuCyKsaoth8mCsfCMz9wq6HQUfIHHp5ngeZed3O
KyQErEIU0IC2JqhERdDiZ12jJmGlyX2cfW9cEJU7Kp/a6BfTmuDHnJs1iGGv9FVKDQHx0BwgWzT/
Tke1Ki3sjaH1XnDejljDfW/V1Us6q8G0zkBGaxNKNhJSY0ex8itkOQ+tFU7t2ymJhQciYhCPhxhn
xvgJxcHRWVF2Dr5dwAt/1543gIT9luGCcQSinCjXf5uCQQ6WR1LUrEIZgYdHXI0yeSXdQqJm5W41
bF7a1G4ehesuSOrVvyQW6yrbqqMHAPIsXQqg3RaTrrcwCqHgRLdPdkrdNobq1LbH0sgDcWM6bzRW
Xz2KfYutIs+PMvTlZdsnveo6k9++uCG+Rv2Q3M3mjas867H4dsubYE75GaFeYeTS44Wy95b4OA4t
TdVa0nexONiXYoZVnyXel+qkqD7LgtlaHAPJXQ9sDqb/UMLOhlfhGayJ69+ufbr2la4akQNNG+LN
o7Hyj0rpZW0QLIz6NhBuhzTWYhXEkjLcxr0QYUNBnohygN1CIrLGDXTS9kQJSjI5bZc16iBqo1WT
4LpD8zi6wjBYxrGTThfEYfdtAsIrcbbjWETe/u/e1y/lx0CajPsIvcTAzwh4SHmyF9JHbJHI6jXv
lG6RrmcSmsMn1zxcvaKrl+osFdo9sT3S9tHkRwaoptpOWRO+yMBVKAhdIkhuDxSPF+vquIx2zDPp
3Ae0hAqccNAMKWB1LO//6V/kZxtQYJOaCAuAu27liw1+FfLAmySmF5CD+wx02yVKhxQpqtKOZMpl
dRXhypl+AHvpAid4KWo3qNuue9P36Ug4hxoxp//c++lvhQy4FLsT9mJaVa7ea+T+6S4RP0s14jnc
4/yEIQlHSDE2xcQZXlzC4YyUO5icMz5l5X4+j4BCBt7ucWhLYklrSiisOIurEyBR8Fvif8aBwDUn
B1c6T/AhJmppBBvSEIEuJXowj3flGv0nULCFzWYnfjBVdEOPKmFTZh4N+yzi8RhwPr52SoQikSBT
+0s8PpZMc30Beh4flJ6tbj/+P1eR2bx0dgSzXfL8JqAp4bQuqGjKa1JIJyegZ+EbPATVjio36nWj
t+We5eSXcidM+6CibPXnvK5UU6OuQCf7Qui/O8E9/WpL6FT3E/CBTkQxS00xeU/1aTyXUcbLyqF5
Nhe2qsiD2j9LNXv805rIyiBGtDIIMOXUC4zrdDQZ2iJil5Uz63ojug/4OxFnNZS22gposUe39vGH
w/yqMQCx5278Jv+EftSFwDQoyDJjgyu3yMMBwjbuoeeBMTSMWBQ0F/LC+6M6pGN6Q27gEtZK/5BQ
Zc59QB32ThkmibRuhjtTNjT5LRsQ5dtGGnLPNmhcIPFz0Mp+Uw0/yqeZRyyD1BFtPSxTkjyfSpes
+JJX0l6KcpemF2nnaHil+8lVhELPZG2TtokRnJH91nsFyAT9vLvJPy/WmSuro+Hcb9yvCpdfWs9z
cR7SRS6yfO5k0PJtqlbPq/olRpw5/d3fB5Bx12xRM+cMKIyUtrFNyZhSzNyWfjji5PSw11/ApdIF
wkN7b4W1z1Ryle1yksaJfrLJ8RKpp6qzwhNmqTuEJudtBa1KoarznDVniXsXcMm3tAnCSkDoD9jB
dFxz2otX5LjS2WjZS/grHCBWpwFIfwakfMixIi5o9sIihZo8zLATttZAiST5rK+yme4R/cLzCfRJ
cm7huXYjaoDzwxWirv5QxfA8gHe0/FvsNZf+IArgoo/wgMO4EoJi+fXaxn9pI/L/3Cjnv+tA0wvm
O66l3WS31iLpOvN4K23rIZZ7hGbNs591kSsWEj/Y/CqewoCHE4am7ue6Hy8pq4s4LAzhSJOWDC6P
13tTxQJ+wFzQu4kHV6D8iy56HhDDA2jChpu9iy9mVE0aVojL0NRMdyYQLVMGEEvoDf/SwxFjUrHu
jlh9pEg5vxA6JBGvDShgyNJxjYyaAFaZakSUWgOf06nOikdbapcZrHmG+GGdBM93SxDHaum+iYyB
lYopgBz/HqQczcHFqL9cXWHITAfk4OhrLjAyTfEO97EWI2z70xc2UwP6lkL//3QSfWDHn/omFNad
OI96CzqB3hG4DSHEfb5pvVHHyVygzGM1kgwPMNE0J44p+zYmjHJoj3a0RfkgeFRUHq1nkgQNa9DL
GIn2sKb4UmBbc/s46rMmnJiHkdGPeageUfS5CIBpnIX+vKbTldzCMv/G9qIlV9vuGTd8Q5SJRyKQ
PLlIvK3GAq01yypHGIIC+UUoEIzg2+C18po6ycuMbLW20y9soHyPcmkvsDuLNTCdu745LQUV/y91
DVklaWfLo+0nsoKUzkXIpFrL5hHx7+GpBm9tJBW6qAyZD75W+HZ0fpLKuG76QwjqcYOEj3UJPW+8
oms7eeU/lPuQTiwhppo2R7tNf66ySgc1xSP0AIdLhEoAX7UTdq+2376y1jy25gMY0p9AIJaVV34T
tHZWdBMnYOaf6rZQcO5GhLod76gtbLE/vVwRNDdTqXWZJDuthOjisgvCBYbUiMEtCHG4Iqf+rKXA
HnnvKCEOi20pT8pF/b1Q6qVvmVd3mX/F39MQJ5dmyHcOr0Beiu1VS1oerq2SHL6X3qR8C6TlkIRw
d7J4OxNwYzgt0isfW/LRRjfWIU8DkdTKdA3SR5iMmhLRND4BiLCtLgzCNiLt+PP9bODPcN4/Ylyp
dAKQ00lRsW58EbxiflDLWn11SP5N1BT5Nt7kqdGNXihTFTwOuGz8lMId0fwtEsTdh16PivuGgk2N
ic2RYvoIq4gnEaPfx29jjgNY+b70XxEFUQ2YHmP0clHpLf8PoFu7B0Q0q5aPp6PgKBWK2pvUMtyg
EcxOF7cQszmZwwh3XiBOFNU7DVCu+Ho08ai4/Mk+2xN++TvGKiVPkqOdIJzjGRAYDVwVA8V59dNq
xVI5wGA7aRlVLaeOxKrj4RXrdKNrEPg35/tLMtrTh5v9CUI4hTPi6OuhcJ2FT1NgydoPKv8aqYq5
RLv5CCBTn6TKnhDXB8MYJ61z41D75Xoadq0FEjiT71SbikEoVsVEksxeXlA3DoqiAylgEdGpya9F
T4EnW0+eKnayFak6xw1TuCuR1JjPIJZIuZZcF9lbNmk4TVz2cCqG9gD0RTLOYBXla1dNbGxXhvc7
camhpRlLp/uqkyKCx1XDhnHKeax5kpNo7xaGUJMoc6iGd1tl+V8wImdrrZQMlf9K9h8UUfUwd1FY
WHAgP0Ja33FvRuhwZkklHmExppHSj+Njlcw1QUAU2nzpf3Bp8C9bPIc6TdOpW5EoAKY6pWpo7ExA
ON2rd7wxIU7tmOeTFTj/nSGe25YJD7XahbmvqrB5g0KsR4iZn/xeJ1mYIJo+37FgNg4x5WQYl2NZ
R4GBB8kl7GVShd0TKVAKPz2J+FfhhNUIRKCMeB0qOirHxCJS7RekVthGcPF7yr7xjbk9FXaZpRaQ
T+GSR8fpVSinnDE/EDyBSP2+Z57A0dMs7c2YlTwZHSMAaEjKOIlamftD6HraEtr/YHPfmJBIzrNE
gnUo/SHu9geEm/Sr+9/yx+cCxLlluHbtnRe8NLz2EV1WfkbwGwBkIpzXMaIcHVyIlBTBYGCCeRAl
SNOXsS9mylIL12cyQZ0RbTtvsxJhRbfZ1XueQRE9ZlqPvwZ7LzlxAo6uXaNXkqSraEMLwpmGPhXU
9HOHGQjkl4f+MYIDJtEXW3U8wa0oIF4FQoBGi8IADXi9ZrfToWUnz1vvFZ0HtopFHjq3E50RP0fo
lxQ7b7rkn3Thfg8s9A47wsvb5Za4xCXUKeHybOywmNTLAvS5Dbs2aDaepeIb7o1EcSfMtLxD3kTJ
2etpUnJX8IbDheIhl2TmbzhJ0TA/Gl/obKfeIH6NZ2Dp3R+8xOBvYHh0AD4YmFihCP3CLC3bdu6W
qqKTYCYDPimozdPBVntNb8H56fKC0neZDSRb7CDgT+i9S2PWXKJxgF3r9ZLNOfa6KAusUz5fUiK3
nucON9vkpXt3MxtCV0JA0mhU59PWK6kshgif1Q8Srz18OfvkOPJ3BDovPIrbCS3GZVzqKAfBEu9m
+z+CoZ2xSXLY1BIm7Mfpn9xcFRPE4SYsdSrXLRuBWtDf5LQYoTWlPIFavbdhdVrtdZFHAxvOz6Rt
ue11e5re0xZQVngONu6TKdBefqWKYl1kzStYyzjDza+kfahHFzRB98SGwQfqFJhU17Oufk5MyEu4
DqyIS+WrKGjASE40EAY9XOyuykFvD1BGdSpfOsl+2uA1ATIru+VpS2YjK3hWVbNunekVJ8gqLELV
Kk38cB2WMLHYH2dn8+TdPE0I1iJFvaS64hWqBwMdejipiuDzqIrwo748BClPmNSmmIC7pn70r7Fy
byffg3qdyNQ5eil4BjrvbPxYDrqXYkN32loY9mDPazcybd0Is7SyGOOydAHNA8zk4UORwJ0v+veu
0xAGJOdpX9ooBAyHe8tpxr/7fH6OzoAGULg4afAaU74gXCuGarRH5+J4YNJzNgKkAfDWc489BWkW
tytJ/+W110zv9dmXS5ukk8VQD5NwdZ5Vm2sdFbpb0Jww+5yktrknHbJps/Ji3pC7dcxBTfszzPVk
4mQl/HWRjrCaIv2JlTIemHU898atA4JnGpFZmiwUAaBXZ6T07P8DOTqQZ0c6WIEr50BXtHIVD7zW
E+jRIBRsEPceFPVdF3521JnmAw/WRgmoHIWjijOpJbouzKGfEAL25XhNauBe7iMkiqA17BTRcc88
7VdXlN0Fyme5RgNo2JISpKQioE+9IutzSFFTRGv46Q/Pu0G7r/RybQMD6Fq00aT9Oq7lAosWARQG
Y9AuUQW6ZbeB/FfWJahb+WIQBCNP1524pfGI3pCf7N7HYeuGuaWJ3wGXJtXhhdl8RkUaK+ois9ZW
HPsfWLqejsyb53fwzNmXhJxmZGrigrY/ph1qDi8EvQc4+o/aEKeqCrMjrOMGORfLWZlsvUvQQLVg
YL+x4yIndftLkiFQ0DJWWcJ3qaNSb7+0UQ9vUbQAhab0I+YIg/+oOYcyPE6a/OZW3S7zL0SV4EIi
iDxPdEgiBIAzXRPfqqBSW/Rz1kMiM8YWdmsjlSXI21SyXkMgKBXdSGB/RPdSIkbnd2aBQt9F8eXY
4Ei7SejgA1h0hWC9h1BqaoV7OlcjYKk099qfYonboD+unUDaFUbKG35qaCxKMA1p1iX98xoKLPRt
Z/Ijbsp803M2nRd7GYIozRscdXcltarT0qN80/E1hgiVAorKld2uOUAle62g0EpElA+w+ZwQGP1F
P03BIJIssttjN11XVq/hewZVIkz/LtRObEraeDB5H1ClSVMdUBDFI4ppGPo55YmLKx/CBRMaP+zD
w0qWJ3I90aaIUPvvaIrru+arOtW+DxC5+OcXAEekasxASc4BiGgeWFGIcLMwqoawvB2JsaJQeswf
dXEZJXjemgLOBNxV44HrX2G3jmBtQCSZwD1AFsKKjf90/Gy4E1yBGZ9MRpnSb3oR6SsSiaOmgMqW
I3yAs3Q431RFPwPZamAllI1j1rJswz7IPvg1m1u/pqD3fzx3ImgwSTceSTaDXo8xEl415PcDs4J4
F7L1iXRyAFwynlxmDTE9ZmnXhbWhA0pLK+kWoiql+Uh5rfWs3tlhfaCv/4unky9Ce14Gl0wpURcV
rtIFPpHA2xe8+3UdYcudeqLHZBhoJaaB5fxniPRil0o1HCDYRKUFRUYGUHb62GQYPTbEsdoBvcYS
RwlxT7IKuuFIgygVC5Hmqwz5bZen/t0M4Trkfc06UhWimycskHqC1SVk5RfYrIduWUKNW/rb8Z/j
C08k8nWSK6IT8u3on3nZxg9Rn7Hj9aYK6j72gE/5zRjw9J9fIFOYAJylj4x8o/B4f5pvbR36OL3X
RBUkWuNqnPQs2jY1uPHdjsVTscBRfIzQ2uN+TQes8znx942BLAkHxA9NgJoVjbF5B6u7djeXXxRX
GEpXHXpGk9Gy74rkgifznz4AHDMf7RQR7LthO1mRbf4+g4ujfe+vG7XpbrBoUQ5JWxXFJGCNVA/H
/Rd2zrIuk9xz98bwOQ58WfHkKNMbRWi3cvPm0jdcl2Z2t4NPOOIZLUbVfLW1RelabGX/XDDMFvKy
ZVzDtpIk9k314fr4/wmHxJAI8/oax3ZPdYhYQYvmkOHj7LSBgnHxvvEIhfmR/1N7PxfmNX6xzfRH
KCm9pHmqdqxrMHTeSbDAk5BOa9cDoV9c216fOGQYGPikxywPLlg+WW0Q2/8qtu3r5Dv7kzEDU2Jc
shNi93f/Gia7TrdDUuLSPFHaCz2CD4dKzvIHKB/kuX7PZ0v5VfvOno3dMHHrRRb4O4D50Zr4W/ks
wfwrcxt7naERyz+WXBTB6nPOvuqDYyeRUwYAR2O6dCvna+GKy75+NXDItYZJBXm8inBLb2B3XlNo
ZYNmPcMNiE31rtaZWBiA1d3O3QemYFCdvhTy1S3ucC3g422iM3K1HQ8A/0tvKnBjkxQAQaA/pEC+
foHpA88IC/o6ssn0igm8syMEznVWgcKcJruNI0XlaWwOhnxIk0+fbqCXT37ECzS1K+yAKgLtG3Jm
rmbBlUXz8Jl9d+Btg7pjUhFvIOCgSJDqiOufCFj6FsyJsYIlUPRPhmRMMmkaUXRZ6C4vQYcKko9y
enOEEDGdAc66eI2jrFGsjoXTvDdEELTuyzXSPDly7Kn1P7edoWq2WOcC8p0RIROD/UKxmsKPP3ZC
BoW9wcSXkilpyQuOpNtLqiyIRyCztSSnWXuvky0IdYwnS5NQ/R4Ykgf8XDQ2exsuvKW/fwAKm/TR
W93w37jdf2Mi6PqMKFZTvqdV1GyxKYaItKRAgKTvY5+KVHIPoSSYq7XWfvBZat+emQlsiNBPGxhQ
gWCEpeZSOGaOMdWw4gbBfePMx6clpi+g3mj50Svrp0StP9T7/av0eYel8L5frJGqMemR2hjkiC9X
kUZQz2duxRIdyUVhaNae/qoR8oVRo1v6aIMd/KbXLpimoNtj6m6SrBJ2xWnKIU5xV4SbhR8Z3kOz
mVpQlSuCEVPAxx281l+xRSbSgSjjzpS0T0ZMu/dV98hP9bkXjm4AyMnwdlsjF0WvvZrUTLfGaiaM
7NiDE7caVhx4nVBixxKjvJU1GVY3gen/K/ZVdPiKJ46jGHrePlsdR3r1h/k5RIxMUSgx5HCD2MHy
xMQ6mZNNQ1rZVnHCVYqHD57yMPaoKS7beoYZQbveCseTmab6F09uXJnSZW1pLjIKu2bDmYgPZotM
tk8gZiDOBD+BUV6s++osBuoScy2BsTQ/4GIhuzLQT0iSZ19nqUZYLi7bCq+lLu3W7fu33Ulz+nsQ
hKMnN0hjXTITt4oZwk02YlUN5DIBA5r5qRgvQIxKz9i8czIDx6Q6w5H95fEjkdI0F8hKVVvZA+nR
DWM6Fv35omhSuX4Tts0/veyt5dkWVh8TwxyIANcwAkcgd/w0mAss+tRrKsQGLN2leZANCv5oC8X9
nY6DvkYx/HxyuyMz9rJIWOTdjIrennLoTJl2cw+n0RNVeOE0rqrEYABpy1looGAj8Y2MNevSe5uT
JkD4i0Ct/iJgc7fNHBeV7rSj51UWrGiAAE7inYAMhFCqRcnVsUrU7Mn13SzY3hEo63NCAsiVUqvw
UZwue5wdsaZMuu1IRkgfKX14Ko98rKk3UxlzxDrs9eeFmrZhO22ZLiOgzSqhXkzSqSgnRPv0yvPF
GNOXAgtt22jXVBWW3d17zpOQ9ifAsf3XMchodtFnDgcLTDUqDE1Agdxq7jTfeNggqFE/eSDOQeQz
IwnTLnrIQpIprEfEqEYK4IcT0HLdJy0ueAZ+zYHrdusAVFmQtRmuc2xXFAIX1QPXcwkLPc1w+KUv
+4hdVl0YcGHjFXdm6zd03Pfb8PGEe9KWg2y+4h82wIcimtwD0RPiKKwSzYDkF2Bhb1CrZfR4KxGY
2j+UJPYGO6Avii43GZxhSfezshUsqNFOjoY2qVMf5GU7JRb28YDWTODXYgr2M/ZuYkEIrtlcotRd
1dHzZSKK9rFvW1YtL05DxIq1cWPtvxXlGyuAwDu6y3ngSUXZPBqdWBnZwHaZSIlmHwWwoueL3RDR
MLClMwId97Ocsxrr1NSrDeiALqxUSIeNV1ONWijNYWAhaFSgVslfuhmUmXrUgYyUd2lndhpYkeBz
lamEF9fACf0PD/XdTBWFzSgV8eB9VK+erg9Jd80QgyhI+/3viw8yQqZn4V8uc5UNz175bTmWJUTN
2W+Ne/i1HD1BlKRUJOFkZAtPU6Q9/QeNoxtbFIWwl5uyLcH4ysuOlZi1meylzjVGybKj6PymAG1C
Gh4pZy9sgseQJ6D6Da+kgRfPkT1fvOVzxcodpC9LOW2Ugc2+waHa91aB5g4WOPTkRpGdrPUJeCqu
oFs1BVPaJHrGjActfQonnMIan0hZ7/uSs69gFnctzKlxkvBT7mmosU32GodthMTnIjimaXxsHi3v
UHKnVHgpPx0pnE5UTdiaLXq8wkHApwFIueZxWK4Bdus8oiIbCWSHkhtJfBG4HuElzzev/r5f1W+Y
a4Lu6ZjBqofw+ntSn/RpJly2HThaD8ma8lvuQnMPorXa15Ja5813LTXykAkvX2vabc5NNlKkWr97
QubM2QMWzpnvbysOOo7nyAq2R9U84UE5MRv1oYAlPAPcIydu3pxHZ2mG9IhlKlaynQYmbmFL8DT3
w97JzAmn+ryBjtRS8iOBrFV6qh9l/ZlwW2dSKHr2IV3gZ1FMJRDf9fKQ56PZkLyaAplcYMszZisK
oIF4X0akSBY2nIKZSEYjN1B82lzhZ07OromY3jbOsXHdIrASHhq3KtXbqF3wFEIStLjhwqJv9dIK
2zOUiFwVvwsqf/hJ5qxJqLITOFi6Mypi1agdxTeL32pTiDMDkSMNQQ9eEw7vLf3Pg+nrMd0GMsKR
9CF3XGpZD2oXXGQd+NAOJBw8U636SUbhMn+uSJANvaZ17GUCExJt2ykk5Ht/snfOts6suZzQV8Yt
X6FQFCumjuCW2Qzp0lkQvg7XWFFjRbAGbgSz+0cQ/wizBecNnDfjKSlpuW/cMj9v7sW6jMRWf+ak
9dFKphyAgLk+yAu4cIJTn7aKx30gLsQ8RaCd6YWn8x6eeN7URX07TmX2GJKpjxGCKLyuIfXHogRF
xuygb3s/uE7vO6oGyw400+cDB1Kd1qaDVlHz+wdvmNsvm2D12iQEKdw43WZiZXM5Yn1VpRZEIAIE
QZVj3JQNYVYeFIW+vpa+oUdSSXWxaBZiUOOO+S9aAJASWPlcsuyZuJylJFFh8IhjKAy+b+FO9Jtk
KQFgNvY5CPyiu87UxSLmqhye0+RSjUO7vb8sVcsfVPC0bKDNbXdeSpZJZix3VYW3IeT+jyEGCFPr
CimPrFDAvTwx82VRWr9Xi2OIoJtwf65yXBPL+0SmgU9RE1rKTJkzpBYQb5IHuCUnyh77wpVGxKEo
E9aNZisdjZQpAxyOl6amd0y0CTqZUPSTQMZexIpmCE6/i5TRl7tVs5IGpIsJGW1OOdYz6irXAs33
0Il7op9RxAjiA/hVhGshuyRC5wXehDBaSxnHmQGRs8pyCpDm+DQ9QTOL0PZazJdfP7//gh51Jtbh
zYT+h8V8h0gDUZVbbpILSa6nCPR8IQidin1mI1huaA3GKwbO5ZqBcwdapYvOrVUl0r1UVocLU/Wn
A2S6jGGzUdXkzzy80lkeojDHtnhvM3GDKLrqgjmtL1RMbQ/KH6QwofTykacIorlnKlayNuluNV8O
RucY/GX+9W4FiZMlMsWKkqksrPt/ifuO/XOyOjL/86OlYw1RnjVw14UMz3yBSGaARcY7blTFS88a
8DUnDaRk6bAAjnMU/ZFwuYhltMDHJrZhpYutUqf2z6A65Cilb6QGU9s/Osk/+LrgBneNHNlJ78pa
+Ky8cL+o7YmoyIfD826RGbkz4Irjf9XCUJ5OFy+Qb6mJeAdvIbtqYUmUYEFEIbLKVG13RA14bVly
bRpBSF/kwNfwrJVNJv1E9FOTOTWgKm/FMG9AKisk3PpAezWI5ZRN5NvxzKEQf/fvjCZQPO95uNjs
pMm/musHcAIQkz4pEudckvfJuu6G9fWYgDCQTwrpy5c16Jh/2r7E7K0GU8KU7t8Tet1THcvgHfDi
Rb9zijNk3wnqYqZfmjgMFh/P03kUnyDiTSv40JPIpvb2lKdu7DqeG3MQ3j8NF0vIJBWmb9WIeTy7
K9t3VFYc0+mSYjlD28CZdFpixg0JD22XOT5doYVbGzBo3x+KLRBj1jiKlRWNbBz2fVP/MGtZr9/r
ZkUmPYIlAoi5thAGeNE2Ufu4taDk0lcaBJDqB/nQytjnVWxtmx8K//7tvQDbpyfoa6X+emlpa3BI
4R3hRBGuR4noL8PejqxbJV8zZBOnBPcGd7nbxe9i2YfCbgIDVTq+clLciTXbzodyTWKE3zYNXJOD
oxXUWF7gp7rC3hLxKKn/mDwpS0nzgRkzKE4dK+PGjgByYP9TjyxZOl6vq0hrw679JJ1JmFWcdLp2
Hykh8WWdKaAdLjV3WdM1WwSTNmmNJknPMMyPsxlPvNRKK0Prd/x9zQkXFj6UJxMgCTDYWUxkSZbz
yUFOLoGI9gk7VH4oWFc2w/F513bifx4ZSkvjQ3W7ikOQPhMQjUuHB1qZyBM1EWNH3zWkBabkkhaI
RYU4EJR7rzdsOdpZ9W6few5mSKcA4Q2S9tmz//mfqZ4NUk/jkCAwzFd0RaK/CT0vcSahyGCl4360
alfeKhUi7yLs6fg5WzOaz/p0Gw1T6aIujweTLuL58ISkZXgz+ffTClvrj7p4bYPz3HiCeRZv44M2
P77nozMEAKLiM9QjkPa4uSqL4VQ57g2eEkQD8oJVcZQufQ9h8oMpv1Td7s0Tffg3FIawRo86DIA4
A9rENpuVkJKouRgA2/oq7OAjLXXFGSyEIkVWKPY0KvcbFh25+STpF3SxmwTi8tin1I7ZYFkvage0
ADNAjYCr7UUqbxenYZ5HsF/1LZjf6fZ4IjMgfzzVyanzmOTvTCkNrA9i1+W3ox/rdk9C2shAJJzp
SUA0t7T6UhXAsyFQOMYx+FAXMXKE5iEdHc6tY4JoVWG5h/9tmrrT8HqMqbfD49oJ0pJgOUmd6t8G
djfpVzU4FX/2lNcIp0El+d8RmE9oCKYemHcQ6lWOVp1YtOR/fj3i078FisICRsS5Qd/nS/QpkKFw
1XDsvFKucf3tm6Lvmy5beOA8MRCnnKJYb5WKupkAVtZDcpeWgbCyOxZF7z8xv2NuZIJmshevr9A8
zZnPWZueJM7Nlc4DQ1UhYqHGiXJ/U2Peo/HADuMEAqOFwA9bMTjIsKoFgjD76RYTvQKGzaAfQ6PZ
nqwHm2gaGTL63R4NdWv74xbHewSoWu8sk+ccwjk88oVOZajUPvGwI30uSG1WHYmhWMpQu3Gi+7XM
6MY/h+VLd6r+N9KnZ4fX3nAkOabe7fCZridy5VpOMw0vebF1gjc9oGMXtuA3EffeIqrvMZtsxKy9
VKrk15KoiqHSimbMdO2K3xMXNMAh8T82Ay+ALi3gyFMyezvhBv256/yklLPq950DONfle3QGLhN3
zrwQnVvIQ4WwPJv8a6CCtHWtzSasW6dobWnrEMmIzd7l/sl90M9LZqrTJPPEnC3IdSNX0ZWJ1LoJ
JqUP9L4u2mrMN8N5FQgcy0pePF8yxnQx1VBLAVGst9rPWsUEoN2TGzBzUG5hbvT4Ht7JQKU4WCHI
/m7QIxpAzfScHEvm1QlexL2pGEFRUQiergx5PvfAK2XaCwyojlU8M+kTT55SoPlIyic3UWsL+Tw/
+ZtWBBoNSR+kk+p0kDWqFkrIBvZG2qvJTF+phUrkBgoqmImLV7sioa3NrGwQ81YixsGfZdUGBCw2
9Ib/N4Y16uHqqYxKyLmGSWTI5KbUNUa9uOWLwI1Jn9f7QJCslDblDp2WvxLsKCSM0WlAYTyYD/fK
r9rw/8O9Mb1DPS209af9vprV6mG9um9auLrg8E5Cw7z+SUtEOxh1DBGEO3asC8Kogo55+qLabP4q
fgE5L3m5h9EYkcws17FZqyOYbcPhL1YUGyj9wQG+S9cFOq3nyhs+j9gD+tusOeuji6b1w+t3/F+r
zVVmKBMH9byxwW/7eF1S7STHlkE/QaMjPzWi5IMKbuOMmdXYxYij4Pt08mItUVPADJG6PY0c1lNy
Awo/qLXCroNzEUbBydwikwLlEjSPl/FwBT+aaiFtwSpYAXsogCLRwizpHgaT+mcK6yCc98CA8sMD
ItwUtUz/6EncIbQA1sPrENeysWgxM+x/19sSrq8JkTRQKZ6V63GQt/8Rb/QLm4GVL1X6npwMRdYP
WJK2xlv3iNt+q2b5yHlNVdlWLLUY2lnUdLnJlfIetwRCvwxsE4rSOeP8apSkvfT79TFQJs1ixmHD
x0WZ18exCv4a6fl1K5xqiUtvCHxG4T7+OjUBX/V6ZUzZ4iWihF1cRCAkUbjA3bf5Rdhtw9e4WwxA
Un/4Rctbcg3LPeqc4hgSRm+4y05xSLrvvHLZwNfYEDnFcLbqO1niMy12Sv3clTCdbXc0YZIegi5m
E5CHiXg14MkCiIltUXOLrOntSg4z2GGOxfSwJeLbindJmbSwCjYZFMvSZhd0cTP+F9QHpfzzdLIQ
/Gch3GviCgWqu/07yQgejtzU80nY44orfAU0/e62Ue3OGgsEDrEF8MtclKsLOyfP1/JDa8GGQBRa
qRu6K3aiZ4sSnuSHtVPEuDSigbo6/x5KDS1v6Sd1I3HoHLMUYUDzVP60zuvZ/CONT1VdbPFdkgq8
5ZvOaW27qXiB8sHmi+e71rpVdGOM9BzuJgxmnH51X9v73aqCsJL0db69AL2taRPuBY8BXVvevSxh
14N7ngKeJoHEGrzNpa2Uk46bgb5bJGEnUpVEDz97V2oqcbRiE3qdGEuvI5fS9rDLWrqsbN/M1DOY
Cp6vkREKyiImxTmGzt+doi3AVvdJZiKkAD8sIr3LpfHU9S4rkdpuwSZfUzPA391oFvDJ81bSbOVE
PbZYZEvJo1HVBvRsonYSkeGLZBE4/rXM3luwuSxji3pOVR8FRPLi0m9htZd22WXQi5H5xYvab7tQ
5DPlAlrHbvysOkH2Fx5U8GEtXoenWWxKgCVV7/b5vVRTTEiqoaPNJNh3R6/YbpJ1yxio3aBQ57io
qktYMbJTs8xyLeGS1bGUg0kMZhcWLIyv4xTpIVwNeLyuz+3Eisoi4Nh3+ogqdtDGB20n/gMriJeF
g+1sSzX+mUoX0vvoEipRHAZ30Xt6MTej45u9yQNozAmPqrPOo7Qsy5C1SSblP3lwGN3EZl7ojGC7
ZNGVBmGlLfO6MiqoYmsz3KSqXFp9CMZVUQQskydESlA7H1i01KZ8UYYlK8HGVqBYMNPcfUmnGMUV
bQgmebBQ0ZIqEGaZQMm6ZCN2NxDman/GssLyacpLPXdQyedpztScnXrpMkrxYymdwBa92j6nQyQa
XFvFqk2his4GuNDQmPkw2CMMQu1ixLiosmg0ZheyxIKKNlsDTI9m9J10I5dd6LLBbI+6rkvTF/Qo
zsmKF4UXajLEHfNM7m/B6GChnx2Na+AsHYNWd0HTzpP0f7D57ShqiCOtUwSutQajJXW0wRxSD0+B
gQw7ANWJKF0SBbY9fc8SH4QagxVihJYnS7Z79r1MszATfAyeDrQY4Z8FlxZwuc70G/o01SE3c7LE
hilu5ZFbSmmMNKCJITvwVinr6GZlDRPNVSEDRQIm2CInkep9878fZzt2vJGA91Dz0NHwiQHSyBaY
pXrHgnH9k655wiBT/GOblEOMjjZCgLz6PlPl8bTdkVVu2lywtQW2cKurWrypXqOFvcj1R0cVKal0
IIMfBYSVR5x2R6wJNS/ixRlX8Bo8iipfjHVNuTpXScAL+p//IQY1WhIzgif+X8ZH7lJQMNaClMu5
BSt9uOrM+IwNa0qVcnIG9T3MGWCGTPb44Owzo5BgCyZrugdULixMy5wUdowCFgC8pZ74nM0mjAD8
8E/c/h0SgjFJESXBGCx5oTV+VrH7wiMKT6H4FK7/wj8VAwcsEFlwe4sB/4qp8Mbqr9jExoOMvPWP
rXTFcxTrKBWi5zLNjb3TXVdzisUw1mF4q4EUfqGDSlEOf5Vbb9f6K3q4rpRsREnFGD8uaFiNrNx4
95UWnfCW+4bAaeXt6yg2nCEpSt225/UKkOVApu+RnBRKVcZJ2JOkhdbNKRLjA10qZIP/kwTzoXjZ
mnjGSyTXr+9EOy8I/Gu7P8XBniChKG1tPj/C7p/l9alF1bfjyJulVPSfbmZZIjnltuiPCJxn8Dzp
fs2HtuCOQ533Yh7XW9s3Ee6PKuK4tD2V6SLJ4K/jXtO5YdUMuyyNe65WHNKKw8BwEYBm2iKfuHhc
fvtvLBLmz2xJop1gVy85MF/1GL7FA3s0FSSTb3eq6oOScru8XamZ63nkOOtcjoN3TfCv4KTZcpHu
iG565lCx0BV/pO1yezCiJqAU/nNumDreU7YpZfywtV0rMP9uwr4/pyb+lvOc79/4zsb0hxRT1ugt
y7CevQ2xH6mtSC5tYrKTN3ox/KP+Tc8pBig+7JcACiKiOb4TQd/QwonS+E2x9pPv3sThGjC+SN8P
az6qoM1kBsC6r7n76KFEoNGOk6MU9qtUvENhjPhVyp/kPsMUaY4/imoNd8rV05nXluy/IuEs4qB2
xzK0wUWaAZRLCgogMqoIsBj42J8zC9fSxKOQJyAaNhtZyKl7s7R7ggrfPwO5C3u4QLurMhUg0EnN
DJt84dhbPVGRjvQomuT28Ei1jI0Cq5lajpe3SnHF9ZvForxUYy7e97FDUJAwpC6LRG5EwmQTBmrB
v1wSEoSCH79oyi4Z14sGaoOiBqAa7Ar4WLm1sX4noCYYlZ1/aOojyiCw7zVoduEQ5aN2Cg2NZa7z
3LY8Ag22n06wbmFKW9/K+jpD847a2yjTItrTIe6ROkHvHMigKuwehUYzbePGgHHbhr79inW3ytg6
80Uq9Z1TF5At95BlXbFNDCf4qgemiOubZSvIzWb5Wrj2euTr8Z2ndnOIBRNRBJKQCywnEju3Wnh3
R4b8Iu2ipbrj23DcJO4cyIHD40jygexTAQNX0ax2HSMeFBDF3pCrMdqHk/hPDaop8lCoSrt5zoCA
0KZaF1MfFFJslPJljzbV5prW3EReIQo27d1k7SATS0tZjHEVwr69mv7ZOuHKrbxV4BVyjcC8vdVc
m7Kh1XnyO4KRI9JALU+GXxRR+SWHENDPGpHS2tF9bAUUXxFXLSXiNpdjRgfH6I+hiyzYvDaFFOE6
qrZFmIUp86Sv8e4iQPcywQP80K8KkjmZCoABUlDzh7F38EHu+DJqsEMnfgoaoV7kMf2No0ty7BMe
wj3imbQOPtHkqeW/SlvIil3qEu2fu/XLshrVEUk2899iLrmkR2tf7/zprkaItzWNlML8SJ4W8xey
EgXvwIGA7F3Sz53xaVtWI2YXDi+JYT91YCUEOkOZB0QGYMw+390lwkZPOwGbWkA3CALzE8X+IHOj
ANm6KOUtUppUZ0is7q2sSHLZ0MLoFwvTvV6c8IXZHYSxmAO6TI7pKxLcrcnFQoqEwVOS/y0UiiuG
biWJwLzViozdpKWyfrqbusCO2JjVhQPCQqvEAwLKt6AMh93byO8itSqr3yit3xcnx/zNJ9yI6djD
ZRv9KoCvijqaBHSAX9lnJJAFzJ8UYF7DGtiy7EGKwTAOEpQUOtrIDKsIcDHpgiJGJtueo+rD3LDY
jMV0A73kd3Da+oRtLzj/eSm2Vbzv/xwtriB8bJwU2sMO6Z8vTnJr3H6yBmo2NuzO+fAbplH7Vejm
U2PW6pttLsj9g7YVezHCVBTNH+bBMB0qa1H3RufQ0XNpLGO9OCXSmCgtvqJzwd7yCmT3ENN+p70z
3ctOhfhBSndPChRVbsEr2Ax3JJbyKcT0R0oSKVGkmkXhQgOXrim033e8+FiTOgW+W5WYZIAHOxEa
sgxmABuVcNJ285jllI8jkntkAK6GMIDLNpXMl6WiU2WolKkksAB4CV5mfC0c6ttMI0nx4ub5/TEd
mbToolxS9iIqTvSJQAmv2fq3D2C4e+EOpm9XbHvnCmBQNoo0j7tZGYLzdSY3rcE3Fu+lg/psa2hZ
Z9uXpQcXKNexPsv3hVjlbH7US0dbnLWbQiKm3+pXTcUDbB7bdQyBK00gPpFpsxJt/3rZVYDEirsg
6sqvYoAnCqOXiblukoKVH3QUMXIIKquGksYMdanfibPU2MM3LLQ/Y042assQ+XSe+r+DOHUgEE9l
usFmTMlMSRK1UudCblrkVKgP92O/R5NlFkjqt+kGq+QvLIpJrv5Z5RZ1p9muLhgOrtpRMwfZJ7KL
nQjHnT4bBg1bX3eR5GV1NELYxAUE9tqcF0USM2EHPJJa0kxjLVk2vQXLtrAeSlHO+FJTcFJnI6Vl
ZQT1qbsLFlIekZeZaw2h2cDYszaJDXeWaqTeaLiW1l2/RG9qSuOjXWKmyM6gU6eE4Q8Ha7OOZaCT
VLBd7FOAH7wBfpxqxRKmaCgQfV8HvSRjbEm88CSywfrfemwSUruc/a/7ieWgUp6Ae9Fgzlhu4Y9d
+OJchUIZt/Ni6u6DUHVi7VTQTM2iAZzW1VDKWW5iNe+7TnClxe1myMoze3srEw1B3rcuzvfsE/c/
HyduDcerC5eWRpwuqGW4YM3RRKrIRyOxonx+ZCYTMW8LNJ7ORO2UddZ8dGbHuESf6CE9DXKDMlqc
i23GWaCvCbtmW4nspBOHB2k2xoLTI0Y85qTCPQ0+b8hSukGNFgONYP2l1iX6hTG+fFuR5+wv/EVJ
6YiS1QDHmu5PbmOpuWGu4EsmxsvDncWKck8QOxbqp56LMhyLTU6pf2I+m+iC5S1Njn/blSS5IWfp
FVHtxRxCgIGO64EmxWSbW8MJlqDJLRTa7EW12HjJXvstYaPqcP25ygMWXdFeWagBhs2+wEaNBGwM
ObRkS/wr2hq8MRFcfLhtABvIDH7BEBgi8IZjnLvaTsYpNR1T83M/RTvhXhwkle1RvInJ84XBFCw8
EOJuCCCf7PHGC2SfgonwlzDh2yijq84m2FtCqdgb7M7j5A7Xvm92ZjxQArR3wss5RPoqDOGDadTW
CMZMge1SpIg1O312u6eco7/MVt9krrtqGAk9/GARexPXMQF1Wu657G4x7x/FcDiQlLA2+1RPLIAz
O2TGuNTCK1xQ6tSNqtf5sKcPoK352icxgBwmzxBG63l7xaObNpAMbDlSx1mtH/h8xIoCuCxlWAZL
S5CAGmTPQ3B7sUMIld6Jv+6+3nsy7a4mlQIw8Ox4OCwMyitrizeQzwlqpzVN34Nvm3VHPHAj+byO
iyjyiTOYrt6zUskYVoR8zD6xyALn2XCWozN7lmJNzWbnmVHjNFLDlhdI0j80bl5zGRNq9Z8JEptc
K7qBJoUDlAJy0ZcgopVM0a6vIAmZNjaq9pXkeApFRGWYTQntqQ8/bo4DI/FMqne0jAQb1pg3MuAO
oGtui8ivSbpBeJ8Avy9kq94VECRkXg3JO2ClizDP2ulRTmpYKRYj16bggmz68DyfFVz+K6Zm9nkb
EE8nhpmgg4sE9nIeRMUz+Ih4ePyjY6Bihze4tnZ5r9we1+z7MJhgdljzPafAyT00SmbqN7yKMXNR
0GUGSe2ZOBylQI/+c8BjNB8K2I6Xr3IRmOxrSFjPGamBUHoMtYjO9y1liDi7kXI6J7QNoSeJ81i/
yk6Cla98WJuWH5yai5sjJ12JCseH1JcyFGsodzAaGe380oGa7juEE0zQvugISXVb74Kuq8oUOKAd
wDFRWjbz1hp3Rbdzfx2D1MeLftf7zqnvcE938QNFSzh80H8Q4QJIjDvE4rG8yOeirL4rtNwupdJk
hMkI4pUEqkWIgQbFvbtyL3DjmZJIrcLlZ5mkPN9AXXEH7K0RKLXEm8jwWXF5orHgFy6tK640LfwI
UHVqRydLnw+agh4Dqemxl1kbPZCCSrGKCGdvpQ/imBf2+RGLMIEs1m0ZoNY1gbG2wZQatxBwan/q
9WawZmydBFSLBeF1bNLFbw4VgBZhf4tBKqSH4ZD6yI973/PT81qhGFocfrlboek4a/km/H1I0hvX
+H4UfAhooLWPJTTP2freM6LoKr6M8GZqTRRyQb1AALl5egope7MQwCM1NMJQLYop66jHGH3MUxZP
V/iGqcGLIuYyayVSXJZNMNf1UrTGXvRr+rqphhiy7g6lmsR1GxJjTjvz6+8GUqmdXCSbkVv3qbBm
Lt46t1/2RG5IK3BDK8VIe4meqrSDbg2NYuidp/XZgzfdQoM80isGOTpCmCYPKgNycNIX8iLxxKq+
6770ro+VqWTksBlDMsFq6MbRIyDOX4JuitFgsJHa5c9HHuJCmezmbQnseZOPJIsxDRJUHKrU/o10
pX5VjztJxAqCXUopV4nAD3IRrhvO7rMpWkFJwIOT+g0Oi2+EN9Ai+Z5kkLYZ3PcO97M0ljAnBu+5
fQDX0Ukk2SK3GvSMUK/G+DD9W/wblZ97AIjmBrlrFWUx6CZSL6MHrtMaDXmUjFRM1oRIULMMspMq
vOpuL2ayFiHfmEZpeX9xqleeBmsCy511ynBSuLchqUx0WvU5wtHIHduPPkgpZwJ5bALu45FOuz04
EPcvhvE/lpIJ/9GpBpNrdsLkvGLNextqs7ZU2ASAJYNVrJwy57Tw2zkqVLPScg1IyNa+nS+bH8Nk
lSvlWX5Y0W5Fgfmq8BlFFs/sp/vjvP/vNsbctkmUPYpdj1Iyab3oTaq6O+P15exXcMP5noKV/ilQ
ORfr4yqFrqYoVSRRrjQP1UxHDryn6cEHdC1CstgkCXn275sr4fmkmL0lfy6z88vpTpSZIhBAYyg6
/6MlTkuOTe2pUgPmj0Jk4NrXD6g3vBryk9Hqc3bBdHcAZmz0ISURACoPfLPfgd7HDhcspQGP9L5a
cwL0nA8Ydh81KfNSdoPBydImOlh/Epo27AbmiVhNE2NVqaO1tkXkO4EUHW4UmRbaImAkE1wqRAAz
xVQkROBHhVbZnUchTbViGHATVEDFRw/Suqr6HLbP/Pln/xtRCQ6zp9kGe0ngtpQ1Zths4Pwv57ef
MC/ZphrdxhH3CbfIR3E9AXjfSPubYyWxWFlEIMxB8+qJFLNZDzHyWdAn7wY+hixQWG0ZqTwLZDBA
G74shSXMR3ptZ5Qrelru2nFRk6LNdQHc3DY2DSzhFEOAl+2NfiDhIh56Y5i8x+GTMCX4SqSdrGO3
XY4G8n5nRqX+eJRCt6twBrAhhCUa3ornyITEKjzHHjFIK4N66fFJmg9Oa/fg5aWwoxrLVEzyHlBP
Z0/PtFdr9DPDCAqt7jYGiht0YDwHqiFFe5UstWULQJ0CRnOhPes+J1w65rh+fRSdkMkQG+MNKT0v
XGNwB9dwS1k8RVwlF34gFg1lmDo5v9/VLVfcYRx2EYnxKR0OHAHcY45dmzq6zILUSQ4DMfW62y8f
1oiSg9UJsyNzWCTc/1c+r/ZYa1+FdMg98wSFu0AcWs98inInr8rgkmFlB0mZzfVS+0O8afJ04k8V
tjhLCisEdXISlSo9zJ6ZgUHo1dgKZ/raNlBlZoFyDOPb1redMZU2hwWE6Nyxpgr9w8NoJq9URFai
ZIPJB62ZrnpFIxH8ByqYSMpAWhO7v+OwEQdqeF5OHPNbiLNuR0bj7aoUE3ynasdvRQSkFgX2XY8W
DJIlHo1endh4JJtdX9KblJbjzN3UFIcA4LhFgMNIeh+hQ8BMf1LOMje7FFIkL1cz8tbz0Sp08ybR
ML7H8X2gYdwYQtW/2XmnD6RMI3PcFptI7xVNs61FpTshTkoBUo1Mg5ee74r9SUtgdrDOsYug/K/b
2emE2vk5hEV4czGkaoh6zSqKg3AgXj+aCzrOVOm3MzHU0jgJGT/42jxEhp1+EU1axnaReauTpxP+
74XgoNZJ3qWAXduACb16Qd9aAwSTzSTA8szCf8kdcAUulRSaSKkkANsM+X0IO0eL6hhoNiHo24bd
twmiw6v/iRd31NJ8qEAryTKediHlBk42KE27yob+gwf/ptb+JqD0XGp33GKjP30oxRdlZjP/7Pze
aNraZzc0Q9h/PoVmUSdZovAExVTNool2acryREUW04A+swR/d+ndcrBaWrdbI2HhaMxwb77zklz2
lgs9899xt73Uezy0FVE/N6dFPgk/GXBoGUPqETQZwYPHKUNgZh0/NPPLDMWQUATDx2tDJsdes61Q
diG8yOzDI3pAM8dI8YIIVQkyI8W+flYNYozTTmAA21Fb+/zsR4OGiTjevo6gQL6BJK/I3J8QfkZR
h1axCCrWPYlFfVKVFG4gIpM5WVjaYDSBgh6T44OV2y7FQtDb5Jr3qbu9eBvk2/Gu8ByP5rdlzllG
lBA66NGYJ+v1fNaYIyqMnucLPJV6FYnxXn6jumNqrShtcnit8SzSvHzU4X9WO2MQqwaGeX08wG/E
82D/rNDHzA0cNv5aHLiPIcPt4dOfDWx1rFTBxSLulGvuPT/d8G/Khd3BoFvNOPVhv+y2UkRoFlvx
1+yu98mU+EDDopQ71gKYWh3EYqCTFRwdHnyYKeW0lJQUiSUm+sGxMjHh0a1zeIvI6UPlQkoAawJT
e9XwPndFsP1bZ9eA3BsP8Yg7aGpNz8DJJOdUGVzzEs/eF8Wqnk9lPPehgl9/67j3++axrSoTi4+a
OTOqOPCEoMcsUafuMcZNAW9Y1/iPNcdB1pIeDWPw6f/HE5hRamfwYFAwHenn/RoQmDc8LurlNR6v
oMgnVaxXP/9hRsni8nzEQxd++ROQVpCqhH++gs59S0zWzqP/h50WzBh2rR7ehww1XSNQAQ0TGxFP
SNuLfolAzqTdII6Jd9V9OZfdLcIH6xWimCkQfhWxBBAb/QiuoUNE7ntRpLxi/dnySMF2+GiIAjJm
ccNAtK0HZ8GZgfnXfD5WRS/wh3CAvH2mLzqQDVviPFrVwiCYrkjDq4FsCN06h5rqD1XUzFyOdKs/
JQbNrVwESXinneaoUp/TzfaxEMVWcYcG2uNh9bwsKAiFW5edQrwIHTl7tliMuIAcFfNSw82xRWUR
0J0XGGhrtqQwXbfKC7pCNpOXy6BwZb56G2wgoeKd5HBti5egNeJ/y8F+EZwF8yrQhg3GGi57HZZ1
QL1J5w10UY349iXsafORO5+US1lonqD1Z26ckp2ounRRzq+D1alXbi+DFiTsZIU/8fMSBARNsbRW
i8X9immqqo6zyx+6BzMHW6EQOoZP+IlpVJo8185EugnmKPZuuGd+WneIqBdehUnSXsZBqZ/IDwqN
O1ycyjOonEhhOTX5ep06Sr7NRFJLf2NtLV/CyZDCYsbXJXD78d5dvcgas43FzPraNqfyMHUjKOyV
/2JbXswmcvGLESPPXdhFKQPRQ6o1VbuZvXM9HUoD0jnS+Lopnr27nVNp2OSyfM/LtOJP+4UFge0z
qGbxXwu4oN/JPJhYtuTrLCobcICpAQU6e7+4n9Tae+lzhiz5D++d6SoWLsLRKX0Fhv4awLSshyvB
UEGLYak/e6HcXKAbVNONyLEiKfM8HJNAHgbyYLhhlsWAuXVJadBeZF8gtT6ywsswktgbLwk7h0V+
pa+CYxljZUIYYCDQSo+3bsDTcl3Ybtyva1knrpYckMg07L4vrmzVGoF160wm6xBg3MCqFPkQ5wKd
qCs5mgCtyQqhlWl7z3OaXZ4sq7d7pDMMt93y1k/m/G8qdpQKVWpg0wcfrEpEcag8G+wJYDi1nQFy
cMErIk7W3R+DyQHvy9kzpDCm9g6i36kbxjSdGHoV4JYyL3Q75dHhtUte0mCTIA+5Vu61JDNTi7Ui
f3qxe35JV1rRml9tCYkF5O6jchDaGHqK2aez3fPO78oQPqIpRCmE1UIxjGVUxZaAjjDZaOfiF2di
cOXWpIsXdDnJmFg7l57+7Bf8NaI5iWbLriEWfecWeDdt73Uq9NpiuoG2NNDhaxmoNqlcBPF2j2O2
TC3D2Gk2fjclZltJceqMLhmco/rmQu86uEcBHeUUR1bu/NMWV+JZ4wvCd4iF2se7KqQZuOLZ2x/E
+WX6nid4PJGCuWLUTe5f8ePOhK7tvrYZCPoqtZRNDTItk1zOcASK+qa59PBKmVfOKU4cZh8QvGFi
Xdai9yfwNYYLaMrfPoFXg+Wdis1PpJnT1mhl6ksdPFU1vy+z3OKSVX/eTNazcJu2wJfyPY8svc9Y
b94jdLizBomYYcLiCHy3vkROw4cv50e9oov9qjayX6K6ImNOx9RLaPcz1xWU8WEvANxoTHPJW5sf
uj7gPJk05rpNa6GZ5/qmPCyKPye3kj1KZsT1uQPnEIlVYvDbqGSlkH2BxO/5PZPOy8N/5eO/A7RY
ZcQnthElJx0UK9srV1txXSPrZ+rxxZU1sMjJVHjrQ/z0kfQVJQzNGE4sgWx+AflLQkgjV5sTXbSt
HFYmp4GyjYU+VKWxv3eezuTa+olLDGb9gl++W1y0GOdy8o/TwcYFnDdk2SFnew7tYYr+CBIPZz+t
3qbGHF3OjsB3zvQ4DfhlUqgSV/FrnMWLUCM+TMdDNJHUNJIKvscZaoRd4avVMeLrwD+UAnemQey0
oMyjOxDJYv5v18ZxrcUNgg7RAkXd5aBHRy/311n31rgCotyljOazpckMYUMoIjXtjr2KNq3OnkLU
g6Cv/JeitnQblkTEkWmbTSgFa4XlWoFky52FPIK/GNl5g0Qzckdh7JwDApZ5nsaEaaSzsu/ICPaz
8ms/M7WftCayqXb1h02I40voNu9JFRWC9AXOHQe0yT17KzA3Zms/s4cF42gi8B8qkG+cHHz0A1V2
ha6BoX7qevhkKYuZuyzf1HQ/YvU9QqA2gAfMd0qd7RciWtUKU9eJwSOqcosDcbEVZTxGx8MvxgZA
UFk9eOE4YSoQ40/FKOaEiIimfgb5b5+zMMnjZV6qTvxGwF0a3diKMcdJ2zEzQM92U0XdwVbQrVki
BULaNAZfFRRoIT9/WlOUjIr8wsSgdaavk8JkOyO4EQHdlWJp2axc4dILeZ5G0oXGuj+D1moxrzNh
MOQ1bGvSrwiJl4C7xE4u6hMBpbHCHDYftlWlsGxPP1S0Z8YgOc+Wy3CJS3WKLy3hUHLSD3PDLZTE
qKMLuBPboxypWQi0DTWem0hZGiaSCXZVpu6Gbnpqnk8VF4DhT6AjkDKdNodSYmsX9MDhTvlqMw5b
coqT/5CpzPHdhzbtz9BpQkNx6WMFEEejUwI39jmG0gRuOnXDkn9WArCwwMJg6R1p3r13Rg4o8MJl
CAdM0edkt+mYWfrPQNNDhByAN3qc5UlvbP5frnQtAlUMrCKlN0LH/zqvw85ZvjLzcHchfYXoZW5k
j9QiMxP/NqWKspji+NsqP/datqMgxq471ttZxmSgW1ZCNcukO6JpVbhC/gn2PckRBpYg+3PFdF9R
kEqAY6OPowIERnZ4x95vsvdg+l8nLI59gS09ZVxSUhIObypRmgivON4I/4DhrwtdzR+ONcBRKVbc
GTq8ZZiXV1hgeQ6v1uL1Mo2n7kH5XeNSU2Aa/4HaNIRReMspJH55KFLka0ZXZqgvYRxyvUx9VxAr
P8Datr8Ujw1TSWV6ud4xfkONliRpw3pPGgiF8cL/GX4tO3XKBVeePI0JcncFxpQngz40tLrrRZmZ
ea26daRvd/JcR+kTihT9in9Ab+G8wmRr4s5bDBVNuDX9D7h+h5oQv3pzLO9Qu2zr3Aewm6v3nMqA
7Xm14mzckJhUGOl4xPRL8zKuQoxNUEifbck6h3MfxAwm7xtnHd/dwILMTPPWcyK1rSR9BGznuPh4
3Zjt7FF6Sm0+KW6dleEPOba/kRa2ltKd8kADez2Evrh08QSdbymLEzTvr+DXi30P+F836fBuw5Zd
iVLbIP3kb3se/thOzan0JQ5ASmPjzBf4/3CZNdfeh+VMQEBHuYDo6o30XKeHcuIdgzDah2DRF4JD
izGfnFDmm/qi7pHf1VM7Fu5elj/XUtqwlPELnBgnEOQeAV2hGhzYurOQmAek/3WfOsTNcDUZwuWm
jL5c/EOCqCRLv95pH3y4QeItgPAReo6LiDveY1Sadss9TcJGw7NHBSJScAZn6ZcoFhs4yGDJcxxD
P2Vh9jgL0DYdKML0FU1+rOm6hjxv+bKcvrMgo95m2RpJgVIWBZckVRsVbYTx3W/6R1cyMIyj6W9x
koxGNNIorsKXAPygCLeErV1wuRNyAxGG3ZEVu8LO7v0ul4y5A31bBz9cu27vtwLkhq5FtivdUufC
6UQtjiF/wIKqgmVVnUyWCqTLiIZc65f3yadoQwhazi0CIQYNmoi4XAyZqRllKZRdOSn2xoC3MZx5
RpoykQDHqMRX1KqGsht9hNRPW0KFRLWkYZBEewA8Qsm0yJKp+wK+Tb+grOBICD16ZCxI9rqFr1YB
hrlBCEZQixgaIK11gh/Fzrnccg6CYhoRawpbshk7jCIJ0w+tM1hcF9KDEkfuaRFQX12PdHPi7Qlg
iWX9hBr2tXjmY/9n1nKnBVAF8D/YueKuY1wwWjBgwlTW/9bTwLMc8MmOZJeM6TstPTOMDyixVbE3
Wl+X6OB1kjy89OrsJ5od11AGif72lwYeUy4CJB+JF4NOYZr3eIKOU+hNX8a/E+BZ0/1lJMMTvFBf
gnEKiXklkzxQ33rm3bXg7M2/ClYCjAIl/EPUjthgZjMOs1cgZ24wLHYRrZylzlRASGi5KrpR2CNU
gLxyeA+6vh065xdhYyFFkDjKVT/rOsPVmlK1G/hrEgwAH1nm+623LgKoNn1v9Dm/BgJMoQ6mQ6BD
ygHbvFmt1ZHUmwhDr7ZoxLhP896RqIeSJQdyR7DD0RYreHH+LVeBPLp5Rvfs13J0jsof2dsTszYu
/jfXKhrO9Rs7RFbpxOvX0l9YQ2weB39u3hK6N++twQkC5Ig2MTT/4iC9PBkSagW0JZWjSd5tKmu+
ocJm5PUdrTPB0a7HXtxUATRAUiofF1dtDKvz4ge3jPm6tZC/atVS/VPUBCGILT5O20EzXAnicjuw
jStK6nfJgMM+pISGObTanUyWQZhNMoRJLfomRkK/6m6EcobyVF8CVAR8XS6NAtj/ioxuT9duMxOp
le4QQuPoITVXGJjWkkIASTrUpzDV7GwIKkag/paEWVZjUprvMkI4Vy3xpM16X3hEwmFbp4bAjQgE
eaHtJDAxp0mpHv5QDD/CL5Kh0/Z8iNB1m5KWKqDOdeX8izDopxjN0auJhqXXj0THjwEJuS1gbBBn
9uj/pZlb1MJw53gQMGIpqmfvExLQEZvZ4bgLMBbc2jTAIIkGNoYZqngljKtxAted3GhuPY+Qoake
r2ViIsHaK4bkv1STAsq7f9cEtXjQUeN5xSfWBfdJ74MVcnXX0VaAPvzhrBIGSS2RvwuC2uJxlL5z
Ay66oJO6c9oYeUnOxA3xT1eG/NLnLMJzU729dV80q1XYfGiIsPVFvCtPjGae1WCENbBnGYNFBk2K
iDOc9zYAQkY9M16sJJduFnm0tOe4v0AulxG19iU8hHnVSCPn8/TBnlftuH534JbDO/jc9fwqV5A7
YSm8cGHLO9gMiIHFt3CNCT/EH6RP2urTqmPAe5bPAukbC8/xifoppcrjORt2lOuIgL+Rh010mS2a
JPxt4eF5USvknKoARLl5GupIxAuVHIuBzuTRSk0f1prcupx4i09W4nxY+cHbU8DO1ec5GywdxPQK
3+SPuxt7CPMai4olyXmriqlpN9UKe45eG1QwBacERW+b/AbF96i35OQoGw4URBRmhJKMo8lvj6TZ
q6/NsC+l/G7+i5t9OSKKVZmhz9lcD464MepJ/cYLZLb1tlTD/CFMGu0tssxhNeinVItRJHpzIDop
uJ11Qi3xtJMQF95eoEXk/RnutzgKDTXMLD6t4J0qr6dpME3wNyfwjIkaUrQtDoMNocX1KjJAW9BT
cUuTQKItaS3fnbXtk3Wxn+x5ppFAMUWY9K1bzl0Kgsv8p7SzzHAH7rho5Mg2PhCBP9qUMeqnpVRu
tgCf8AXrvSkub/l+fc8Js9L93JUJQnRbDeQCBUDG53flp+AaVbyazgY5u9x+53a0Q23JPss/0ssP
XNgvK7m5hYvvTNN2l4VQN4tZCqJiWfuSIcw8f8CNH494gz1Pwi1o6TmgeOlSh7tWRUAIirzc2wUy
CQ9wE2bySL5VM9R1hXBrWdWdvrOch/0NorhD+HP22wzeuozaVhUVycudpP0lf+7NkWj8tYKUoMpe
1ZpJ1VvqDZEYtHaRPF9s0sGjzf5lRjtAROFm8vYeK4KX4sRAobP7Q9yaazPRxdWfCXQQ3V25vAY+
lWCyROXFBFd5fSuoP+wyfc8pujDXq7+QUR00n7u+uSYPMtWmSeUSFOfnUbhNYnj60EGcGqQ303UP
iIjvJphpR/7MJlYQhBrZrvVCDrbdQ5nOgu/2qj5R8AF+8PElunm0tnwrUa2wwQTa997n9mKBtUYz
r7WxdQmuLfIcDUG7LcRgCzr/IXQxIiSDpki/OTcY8e/Zn9W1nWxQcROl0qn3Cer9I/0oruXkNYPw
swBSNhL+M5nrFCYupXGLNYTKF0LY7+6dPHiNrJ9OkFN0su393glZP1sq67RUtzYgTcDja7FlTtWp
7DOgA9+9LVQ37zqfbvmPKg6hBGje3wDNxuZnJqRicn0Kovcc/+Oyoj/tzdcYAcugJiYu4NYtTcIs
+BdEG/u9iDd9pvkFsIejXIwM00naX1YnvUKcy6gIPcUECf/g2Xa3aOEwcIFaMe20ymJdPVFeLr1m
3+0dWW6WXih8PaawVN/MvDFmaMbBQe2Rt4JPz3XkkgzRwkFwD1kkOrgvCLfCLzZRgmPmTAGBqHR7
/AFT0kH0rY8JF3K805CrQR9Pp893y9osM7nE3EikdeF/RxKXIbmN5bNfmLao5SMLFWYWgwpfkKqV
s2NxIcP9D2zLs76X6AqXd8hd728H3rXxJvD9QTVx5ZFdzgJre5fchAzeoy6kkTmxAkk0BegNwmqD
zDO56a46Kx20y9IqWCqZUExPpIL8HMj7+l6TeEYFGtb54IIFqXTKbsAXBgGF7CtcL+eudUOXnnl1
JiSGG4Iswl03Afygc4lYE3jziD4YzGqNnm7GdwcFxMyog+H/GK66T/6OT+E9+EllBnJCWfMHwcFD
b01C3jDIhicag48KPM7okaZHBSuyJxxh5zn/vgn0kGFxUVJY+7y0DNwAYWIVbnQIEiDldhCzk5/R
v63fNliJShL4gSUyBM7zPWpdQ1ORoF3fGqJ2YzgafVXU0RARYj3PvoRrkJ6l5ubSorsWdrXg9U2j
ZMgkQF7NnAipV4gGhrGIVvACZFx/7RJiTZsLqYDt56DwDfvrSzNDW+uruQu7qi3RWTHL01N4bG05
E1COq0Gp1nO5X9xSKxiDx0jS/zq55UHXi28bZtuv5JnlpFuH8rK9XL2i3/ZiTAJ7lfDxyaHInAZI
bkBiOU3HwDp5rvxe36VHc1YKsA4ZbPPUMzmqsvDFt4zS0wKNB2aBPrDbicwfwKog0ytc07P+WHcg
jFSbMNVciwDNMJZci6QLNQOZiGVNmmo5uywhayTdw2ere/LJPgY6mkKB9zG2vrgrJGCp2xts8qG/
7D+LSEz64HXY9eGl1PBSsp2/E37HgPM8ETeH3afKMWYsEmK9y8aIo0GwVWkDmdaiH9DcdlrAL2uF
vlcZDvMZ6d0rN4N2OpRUSb0DTKvY0slEQwsq1xYRvKa07tLYMoVWfczDnAP6d6x8P3irR22A6sLY
4reiS7WHoIHsrTj3F/KV2Y8ozex7uoQ5HQHtJ6vvR+rV8TJokPk3RGP4nVDTQq839cRncZYRtNeG
zQCuMf8Eb7kqTmBhdA9DLN/wmXhl7gT+CeEd9ZD5Gfn7l7iaZ/fyTRJK7LS72wc05RurzZIeMmwG
Mp3trq5s0cotosVEbJ2nGIiA+8QocrKM6ri7CBCJuObX0ohGp8ENTdUut02n2FDTQ0EQkinOci3Z
L/l1WOmUkbsPghtWlJO9Nd8TGv2n8ieD8eFZeWjSmdCQJ5lEFAdNEPpT8W7aO490kjgEOhaLKK1d
us/AhHenfTxul1sh5AH3os7WYJ3+DtZ01Q3PsR2f+S1FT7zEKv15AYc5jyyhRMtpo+8aXJNI1LS6
agDlUFovRoFxTFfTWNlGBlgmBa324utq7/nKInp9nnAvU7KXLd/H1EMa5WRhDnjPBkN+8MkGp+xH
OTCBndHc88WaWWX5jCiQnXgNe1acNZykz1m6MHBiaqbJeef5qAdfEcXwOHhIBmklDkcEZkv8x4/0
HszzNwDM6jCW4+VJ6uu0w1/MEvb04d5gvfyeNAaiGnFKACgW2waUNb1QZqQVXRLCIeaGDC6Npabb
ex2pt5O7njXRkoNzCVH1EUmgo4bI1+WQ716F2nRDc1EKNOkHqT76twcR4MWbxmxUBPQM7b4kyHNQ
rsA52mKgmXzjYj1Yico4nveVxp5igDtgIMOtU/Ey7LCEpOcgV2x1llmixg7jkxaIuNv3gIc+QZR2
/YSUUbqhzW5qbPL6jHdPeESRzDL+SPL+8CDVFxg++CObrGR3vS88T4IwD+lgXbjxwxGJ7o+3xKDN
AFlo1oPK23UqOr9Ok5yWDy5112SnS2/BDmLsMt9dehim+2hd3rmWzbWC/YTun4d9qDl+RNwIfuEi
TmLo21VwYPnqHqmJCRiuOp11CB2falVFwky13GK0QzlirEsy9dgzKb9IF9mr6oJi1Qavf4dMA1R7
xpCpcDUCjetb7JekjANvnFdYF3RIdEjUq/A6++Dq87Ck1iZOsjz3/x+cFiGNxZeB+jvIpUsvkzi+
KAqX+1oLCgfiwjoRhPJJBItIelo6Pr9/RdcXTbdJcOwu5lqJ5ZzIOLsd8E6A31puMsYlFc2zznPB
Wh63GADQZ3FyBI6ByvmpVYFWsEeKPB8YTemBd1VPfjy1dI/dJ+fLiF1OkwSdouYF1GoEjsvGdjPa
eljwv+Y8ka+xnR4tkggjmEwAboaUUKHqN+HATVDYOhf8y5IYY2eJzZVgsD1qQy7U2LfolXzaDT5x
AKEuzRXXQ11q1fSykePfrN9PJt9oYH8lZUwAn03IYHLHZSQgBl2Y7PwNY/p5bBXAuneBQwrWd7fZ
UgyHzWBresoKLQATI9z4tA2CIG7BSc8bwYAOqW+0bIY4eO9eJpn6zbE8QJ/RQllgieLlTdOlAjJ0
fCxFlBUwgHdbQywCg0q4vEZ1hx/jcbBayvvBAN0xWqD+qrLkHO4Z0a5gAlxqZDZNdV+8oir7US3H
t09GwOJgdDg1dKwrqaIpw/NndAhSLn3r8bhL8l5CjOk5LcXbsXiwfww5UxPI/mzzVQEc2AoKq8Lf
0OF5MMugC+0UbstXyIMWOHZh+u4LDYfoVn1r97W5JApNBs01ojizniy5iPe84V6DE91mmZNoQ5/R
FHxANLdVxeuQS2Dc0r3cFZV/4QbgtmFF7m4Rqjfyx3W6upHYebDQRadp1EIcM1jsvr/8Uo8+M9ie
kpVdBhwCPo7r6y9tNSjZpJ2nJBgT+T27IZP/VYGUkZ4eq0zRdiq65dFgcWxFJzuA2CePFH3eoqj5
0JumKVkfOEZRxeYpoatUrxEiyR8qYdxFMCqjZKnB5ieLxt9DqUyYEFZ5frs77uAmKmmK19k6SvsI
aPFAilTrYxX02si1gJctpKVzPmUoHjs5p6Bt33CBMUdQr8oQhbIHi+Fe4R/wH3+ULJX5OX8DJx+3
KUwnFYQVSfyysrRWzpvV2E7Zpv2lpW8kLmr+Lh99slmkjNqgN2h+QFyHNFa60Epa4a+QO4NhySZm
84HF3KDvZ0FJ2fHR8rASYlLdbGeukRXPxhY0NlzuIUTVCzobu2QnqgT94wGkuMdUY/snKgyzQ1dh
jGt1DHBoXRlmJ0GF8pCmdDUJNPGei+3Xpv64Wj187k6eS4WjByiAZ6jcThzW0B3EvVmjz0Yd6Wbc
lzQ2ji5tOz1VaD6y1jcv2rM+f4zMnT3iODL0znogtFdcTe3V5sqw6dzAMlVbQgs8FbAfB26OGV5f
Xm2q9EKL6t/05pFKGUq2evteBVCadb+wFDwUzZpsrQi5Xx7JEb7M/R7ygpc7WIt4NmICCkXoSbj4
nenYhE5OKd/cjoU7Hr339txGRzP1zOqQ1lQT1E/xu/Dk6LVhNRSn97YFJfvCC9bRKGUfxxyQ5FXg
Axfq9H4d99ImxHKb4UlJ6bbqutyrsIudOP4NJwGNAXWpxCvPrKhbJoJsDW8uLGrnn6DtB9fMhF5m
6Bg1agKf+RkMG6BrqZeXk88CKilk3rg4E7bh7roZIynzk+mN0Iqd8qKebeIHRAknBX4zzIFkKJC5
o0fQv/URqAhmBzEzjrlv41YMXolvfaxBYDPa7IlrqOKypOkbM9oAa1Xw7A3ztgEfOmAm7rXtbI70
6VuzyDSYNKNPGtopivjhZ8++4pgp1OjkN2JKP7D5tgHOcsMEgyivsIq/LSve2eioGPgVNkhgT9D4
vnUsqxN8idsXIjKgdaoir20dbyJtriX5oLywFAdD7HwiYe6DwRuc18WIWXTkQk3kdn3XAQViG0oi
+hMAS6UQnHv/EkBtGBCoHLAvnYiU1AEyz0fKFqI4BQ83jARqN9N718rmZ+7kojmU6AGM02ppNiaB
C0XLwtkLhapX/lowmY+wvK1S2dWv/5GeskoPebSRIt3tclcwPWqrtLJbWKP893dA9WSdKaHUSrlx
x33vDWl3fFWcEc8PXx1c3O3gpR9fYc/7jvmTwPhqeRhnZq2Useqmvpew8+q2zwf6ZWavKWUW7DVA
ShmGYpB0rx8ctJm9aAPY2pBLg28ivZy/hEZjj8AiVEGQQfheEt2V1cz/hxEwkA4PwbzWifpkZyEz
p4h2EM5Z87j8VWfzjFtpubUrKPZbEHVCqshDcEWz6jyGHciQdNkdqTxse5Q4eEDNEcCUhOhE3SPf
C9GhUcfO4bX6F1iNpBlJqouuV0O8mbpFDb/3mr9yxcqswaT6T/UiVyVpkghiEFJD6nHi4fTxszmJ
IDlhR4adWWdStI6nqdQI0mVIS/2k6WSSvg0roNIHcQ+ZPnrLo+H5lA3tU/iKsYG6zo36WJYoMJYU
nyqenJTqxX0QPedK8QOuMcuMHCB53Yku08DmY2AnYMgmYwUuOyyFxDwQTPzv0Aowrh+A4j7rwI15
R9wV8T+/+vYArVLEDsCedJ8qOx95eP3rKoU+kmYEyAAz3boWlGkyBA7PF3tQzhC+Rtf1dz0+p8Us
e0H/CypNvQOMH1ZdJbCYAxkYgINjkgiBaVRn/a/TuBzvMxKXiNXWxMAQ7ILHm+yufIlCGZCoBThZ
4DdTKsMA/o0HoBC8pQFzHszQs0awqulK9m9L8TR+zARRwiwZhXjs+EcwdJwg0Jy2miM4lNWUhHE9
bdrb93soK/kMBM63UCCsP6eMM91VkVscbp2IjL87xH8kkhIEj+rktMV7BmjrcLm4I3eaj+Fkb0XO
rQbx/KdJvJ1S1JNj7Lf0cHddawO3ZOD9plSeXoI4eu6UWSy1gui2kWF0ceqKeN+daqkRkl6dPkSs
NIJ/DIkuEmDhTgIIHBdqi/JFx9cGoS+ut7ozoe8jgKHJIboK6WZptx29HKhL+JQXECSbYuzwchvK
O4lfBQsmCbNppV4dLK5UyCAGG8FSl1Bn1HZAvKUb3sTQ37Ez9gWzAXnYiHDePBBkdks/ls8HoTBZ
N3ZIQRKK1DWMPWfYtNRsYv2RCOJTIcfd2Uv3sm8U2gnCh/wp5fkEGu/bGrmFFq+GCDfHQ11ltfQu
ZZy3bCF6nIgdwiYqTboMlS8npVZmow4L9c8//fkxbXu0zLaQHwadCvJzDogYbFxsvDyq+4KIfNgA
Xrl57Sjpkv7e33Ya0hfbbbBgD9ICNE4Fs4stvuGUMaXZvegBV8dGobjpJkoFZFZIw4p83ZQ9o5/x
6sPxFeztuo/PGGOPYJm0zX5w/aUh4GqUY9JcS/Hbp/c6S24+118Ep2WweWY8uYLdHiTEg4xfhMSR
EprB9IkI5nCs+oSJXplCuyZh6KsXIgPEd63KiB9BFy5AxoL6HD+N4x57O1UqS8ADQWMEl9Q6UnxF
z5kUHLB8n5A3AQNuqtePrf2T9wA7924w9/iaaPns1b0cYtgHdF1RZ7RZ91hlCnwhp+rxMtHz+lrk
EEjC3JBIFPgdNbLhZ6Ne9FzeOTjAsRVbUsrt7LGeP/j52gsqZlT7Ra6CIQQ1/ulOwBOXq36HsI2p
UpTEQ1PGI5ayKq/nmh3VYLmU+7RgVhccA41NKM95RV9971/a0cvoMxeIo/gfWk5QVPavEGOU/H3V
X/WoivS/DQUClbSfo1a28zO16jEYX41JlCBu4AiYxNG8dQqK267PGaqW7I6NI0ptSMi4SGjdzi08
95WHesadOdRGK1himZ6OYIyLtpUsYsOVa0bnRMVIZxWbP+QcB/spsowLPQ8tLP6VP5Y+NwLhk+4Y
T+t9lpJQ2cPSR25kD/zb+KQXlO8cVL2CYu1VIHd7yd74bGrBFUljrV0dSpJ8Gjct33Gn+sSgnLfC
c3Y4PT3xra2LJvewJ/Sv+gu+uVdBkaFLUJqm+a/chWQhirx6Yezj4EYWWnmlNtHQmGLfI2nUW3A9
N/4zC4Zhn3x28q9aeXyUHklSoibP//ZW23jIJcUIYPsgJV8VW7s5hu5v2J4mTjtZhweqI0Negm2/
uURsmPBv3mg3swoTDF/ehAzd+uMvQz2YsP2jfjctSfH3oXRC20Ypk2Ku+niZ0pMsgq4r2/LxN3a2
MNwvso1SOs969XSxUfn22tLNpobgvxDtwiY0PFwjXzbF93gzQesSzS5CQTEghL4lI5m83nKelvbz
FGe1mTmLIpMQkb/TmnzcbVA1X32C+MGKvYXmmohl8R6NZa0Ikr5TUYhIwX6odfi+4v/fz0PGvqmW
X3Epwj+iNclBhR4sFCwZZi3blIpT2r3rnzGpLMF8XbzShg6ZEWz67A2jH3whYD+1QjRATSZa7Y/B
7QEbETh115GzcTSJrwrbfloziJ+S7hfMeaNnCwnr7F/tgp9Zu3bGgKhkBYvU0RLIHwUxnzgFn7XJ
9uWQ4F9DV8Dn1SovVfyRpBmnVmrum26qNpijpGYtReaVw3Q5ykrTTGdkwcPUsI5HX+BVll+Eb1gI
s/Q3o2CQ96805scburbPtV/Va7qyKH6jh/9oF5blGEousYMba6+hoMXmcSdf3IwA4l0SQU3wteB8
MWMnLmgpcHKtms1U+Q/NoOc5ZZ2604S36T2GVaOfPGVKj4dWuIXvnu3rXeaVymcoQ0RV9qbbBMje
1kLb1I4zOKmqu7AOLMQf9RTdBzxKDX2L/g4iKrW8c9hqLO1DnWKpbEj+CSLouRmc72Fan4P0OQaS
kcMT3LILxJy3sfaMzQWwAihqVEnFcYKk7vb04UdHKmk5wxdHM1hc2fjPOGSwSn6Z+Vo7gZyAciK6
fRSuMWnztQB9KUARM/LR/ekmPn/S0cK+qj4swBcNp8Ly5SlpRoB4iz3iol4fQIKDESEPY0w4ThTh
3aY/FeRiGsMQrgdgqkMQ6WC+vFeERvz8tKltk+Q9OhuKxr0v7rzNGdf3VYsrsR9uVetYkAy4zrRD
+y1mNsi9oUPmsiO+GmmY8erkiH47sfQw9SFMMAmvIg+GSIaw6ExaC4kL/XMMiZcwze36Liq+hY9k
ARfeQYAakp29+T/1jUIMTlbYhUhNrWj+YpENSXebJqzsFseykBSRAb1Zy9tBeNc1+5R9MLlVdSNB
TaRtiu3Egwkg+Y4zgGCDGHib096WmxrnZAdU8wMBtCtSG+FRDriJkSRiMjMu2IqprnzqDJimRdai
DimJrDdNF92/28p7SvsIRlPDc/rXw1mXexBhLDaJPHRoM5WkyuFSu+hVgJMAxnSr6R7J+dWBfoUK
f8UjkjeXd6IMymzk0BjHkQjOux9K5LbYwo+Wrbb9ybvpDhtrwzrXtC0RJOQZ2kR6GFHjbTg2WGId
dW5JE0C/K6CDEA4VboJ7m6x0uOWRDh3JPRp8A+7GFtcx49WffStxHX/ECFbSx6qZ3GTh1dG4ylKS
4bb8DMkaO8IbMpzR39ky/l1Iv19d6lRc9j3XwelfyA9cMnq84Z5HW2EmkBwbNCMBoUTPWXkJPWNb
UyPcLmrqsjzfhgITzFC6KIfQ7dOU2YWUWSm+h02ViNEzxgggiR1YSXgJKLaAaJHyxFfRO6wuxn3q
HXTHg3KyzCQFgF//vJoRq4zsZ+w4Lmo+BkqUau6RrMH62k5j0t9+PG2CIBuQXel2CB9p1YxYaAS8
3EIJZYpzNtZhGYrrxoQVOc93Xke+qWOYH4fA/FPjoD4feOyX0zU5gfY114hamx99hT7cSskbKMXw
tGzMLIPsTdxy3dCIJ+835yutkuzN7Eeb1oe1PTT4dzIi3b5n7D194I1sA+Ymw+X3c3GzWk0NcD6s
6zkIPCxTpyo8STlfaj50uUfIxbrs9C+6RyhVm/2A9cilJtCwVjQndPImEKnzS1b4hLh2+HH+vvgM
DDVcLUJ7NLC6r2azjHv/zO/eLgMKf387YTDpvBHWhZltEOXlfCZprW9J3mHr6UgGNel+3TIIwb58
RW7qcyvulXwMPeDD4AiHLZ8qCLhKCG/tJYTJbHVca+Vw7XOPcx5Mhv3ZrNasFhLLqiEPs0oO/ST9
iU3lDDbZ/z3iQknoy19Qsq+baMVfXPbXLhusIl5GLyQYkqPvjtkaMxf5xocvJVSj4Np5Jj9FSWO+
6xqHzsgVgvGzOoiyogUfaYvZsP0uxFPIizGrAAllDd8uQocGkd5q7PsSFm+5Q72gE8c391JcirkT
QoVE/eNpNh2S5oCycmwMppVx08WpEVmO0Zzy2hS98D9EqzWyGkZASqEu4iFttztysmKYTihdNNAT
rAotYpRnKlIFmpsa38k+TPxfl2FzCoB/x79X7ddyW1C5bLkxvHlo4+IEhZ37KrivXIGBl8K6Xdp7
I1KMD3IWVMSdbiFglowOzGzJB2kxnGrAmAr8tCujplQrATe9ASOvH9FeqbRt8CSE3Y/yEYC+JDYp
J1k8PGk4uWC2Eac0nLd3yVXDdGSXawD5dVapbaupqUUJn9OkwAn9lEZpe1VsAzJPe4Uo3KrSnRYB
EnNkVTXHB1DCnsgUuSJOdrSi/vxCP5RAaJjOTR/J7Bqb25TKqF9/0zy3lasiecVIUAvwdgmvEtB1
/mugmqnyCCKKLChL23FEXQqIn4o/rZ0IKXav63EN4sBEBKGcO1oC1Y+jHCenVicG1ZzGzzzHwjX6
ZyOsNp7KxarN2W9l+Tl+ZSDFwOUXWLofyTlTHxR+m83xlGB8n7ER8M6olPUevXGs3E5zL2Rwwi0o
ecXdcz4chonuXVyzFGnt1GK5GMFIY0QD3eg3VvlaCAhbv3agsf46aaO7BCeP6XeHNpOEzmjToCi4
V4G94ii+h6OS3anmp5XgPd3QafR1aXY04CNoSigWk9UbAEegeCk2wUa3oZi+w/rTvFJnJ+I42UBe
7Robd5DIPcvzvd7kfiRdm4ywULP2mTicx0YmVGF1ml8hvN4NV/jc321t1fPEd8hD0ZM1LiO3b4N/
ov0ZH0M47WHRI9RWJI6dHtz7ebZu1KSidFfvbjZoucTWjfQXZmLoZH+b0xe9hj997g08zUld2l1/
SD5jvzBxfDWfpfnSfNQ1w22sxi0eCTJAbZ+sgZl1fVhsLsKei5utVYakuXtl02nn3uuvZn6JHMa2
3D8tPlTJ5SmqWgPXQ1ga2gIPN+KzYHUf5XMbyL4/0ymfjsZ4p1a1rKaRch8kfC+TaWqC+/NOCYIg
nFfZCyQPp1cLiJQX5UiNsjKu0BaOkckVajjXdUqtaJlKXu5HJSWAWiL7u0P74Hq5NPyKIqhiohPL
mci7zbNn7RuMSBv6W3fOcLImYKZNvZaWol4gpeY57te2TUwyO22dvmG75QOjE5H+Dn0ZxReM1EjI
DrD26SHr47oWwA1VSC+zr799jEc5vd3lGnJFO3eRwXvqxtsLe0s3bTbZKI5QkoNvLIVd/hKetzZC
m2cqFWoHRYCUA75unYp+/bky2HRtKVAqUOqd1sxr95zNw1eTcMkWTwRTHwGCT/kXK0hKalleC8HZ
/bhwQF4SZC6SCMWmtkcEGhjoWCbS1sHlM9AQO7/bU2iYB6pzVZ2N+jj+B/mZsdPUSOMRT0Yvtvtz
EtRVtAkSdN4tOXWIhRQCUreRlbtJ2aX3BNKJDyESd6lgh8HPJf/KeSegOJW4HV+KEIx3qsYNC8Wi
LBaraoXeoONb3Id8FXBG+fcLq0TcMAViMKvWwfgH1vsZK9siwhVggWqdYRHWlFSgG83D8mLrFugz
LG1+55+a8/+DZ58QMK3WHRl77mW54PuitF59eV1Jlh/0XuP9ngJwyXtMSjR9rPDfdB8pi97ItvVY
tt3FvCkYPS3e4wNZwy9zxtg3Tb5QKcW2PW+T1o85X8tJ2OnpaKdCCJ93m63vVW7OorGZ2wLZlNjz
1hy2d+o1K7tHzmuijlqaYscCvlj9Zb/xYpYeMrEpWnqueUMV0wY4+lJjawaFptDFPuCRuKiI6H9z
5UiNrIyjZ+oq9TSBP5hgT/hk6NRlOCeHed4cWqCC6vc5DGclmHB4fcZKZXnfhAAzZQEwy15khm3p
7R2crU6kqeXxYu6lW83RcRccoR8QWDqAlEaXIEblbizaQ1pw/YqLZW7y0G5CwqfViGk6Au2a9n2K
GPjrd40Q3Vzy2EhCZbUHdOPCPMXgPBvqVEGV1E/Y7oyXfued69eva2ciBT7+mX1gDzVYS5y1VOOh
hrvRHlQVQNFXNOXma2BXeWxVhf86l7rUhl1yGIkpmHNYUZIYWiH5/KO/Ezd8sQIxoLaF6WPw87VF
+c+zaLmgANywuZp8vclaY7UFe8KIFJLBHHJLIj2lZTQNa3B7qW4PM8ucPpWKxkKliZzZfSyjOtuB
JwP2tLqt9pQ0VYtHzhCtPRYXeDUXtoFxQlKawqGeQxdiTSacZDa+8pdiHg27thCWrYwuSacrcuqk
K5VKC0TesNachwEL5yPVsbItdSrwp338ftejhPNMJ6wOfNmFZCzKFQCe6EgFcfl4f71BgZhnWmTG
PO9hC9UGweWuuN8pT2unoGAF5pM3fiaQRumwzTZmA4xGI7jIrZMZesJZwsVgoTlpw9kI4cAH8eoS
snFcO8bRq442kf8QbM74k83CHiNKCdMogAowqbqZ+8G5xjj+ZWMX5xeWaRBfBCs+reY6Twb5xPcQ
sZ1nHg6VPH7VV/l70MvOMYlfWa3VyQD1ws5ZzVhIA6RRjw2Xvk/lociAkkJN0sRueJfqjfE2laWL
A0cYQFonZFSQ1O+YSEXSYQcQ1Loj3DeUlPR5friSyfok9TRLrWAZvCKH7NOgGM2hZ9/FfYQWnKhV
eQHSkqVcPN7jXMbbUS4yMX1gVOrUuRvraKATMR7AnCoCxtH8LjJZBaF+IB7FCCQX9kMYD0yBHCUW
7cNsiQn8gtaNmogQzEOYoESvUGGZL3onNNsEekwlc+6FbxUK64VxpvlARTyPeJMFtXk0Gh3gdRHO
S2Yxa2s1sRBiNHLqYas3A7HZOXCrkNC+aBnVdmVZQqx4ShPt+gkta61TZiKUai9v1xe6Ox+/cKJS
gipXxi0c612IwW4m5gyyWzejxOWCv0mmeI67cCK635xHraxbJvJ2uANJT/4+zPhzNRch21CmpMY9
rmqnUJHwk0NQKqPA8fWPaYVEds9iYMFi617fM0SgjAJNSHI/5kI7VIDZg2cPaOtP2O9n2YIsbv6l
UuOC2W8fCu61u+dhr27C8Fa3Z/wlWcATp04vnBC5J3BI6gDKnbwFsnTIYwAcOT4s0K93ClOcDyW+
oBNrYQRDKT3sCTCcO5kWyL+4j2kgqJ2puTxLvRZaUXYJPVenGk9m6HtluJo4BXXPfWzIQ3HHkRMo
u9v2CkDcU0kOG2pmGWXP1Vfl8sGyL+n5bcylRjEsN1gnLzlGJR9TrHYigeedUROPvEDcIsNzIm8h
Y6DWgs4g/VBODqQf64QRfAahmgIWHyboa1X+xvciKj9+tQIb1jOCZuPNZ4zH/PEBQ8nwlAe54iNg
6ANIhCFBEhAceyS00cJih5Uijh/14b17rv4mkdc4YnH+GqHNGh09fRnGUxEFivlI8acH36rgrzAq
I/aNXB0fxqCIdyh00ajwc9hWEJOjvzJ7RNQdSQvbN7U98mqZPmCk052/m10Q6sHlrV4oDDGKSDDl
dQMNPo2KMgGB8PeGxyx+myjb6IRwrKdUq4vcEpakfuo53Br27yp72YUKSkWzU/lQFKKeiY+3WPCl
M+BCaS3C6Lp+0A3FGykgsrKXQ4W60nwU1b9VnBwxb5PLuZuvFjT1raYcPU1ZShXBpvzGr1+fFVC5
ECU9omBTonZQT5gPz4LS3Ds6PFxZVSCWyPbSpx4GCcVM42As2jPd0a6309oltQy4JYdxKVOfMx0s
WphMVT70ubYZv1wz1+5giKyzVI38HZyZovEJXKc0pQjc3p9YI4gHWPcVVegq3ApqqRbeAg0UbqnZ
oG4ASSPfsrnZWBvVksnbMdeeOqBoirHOxl+LwmcgqGUW8YfgCpgL7TXQ7jARWX2V9JN2MslIBUd9
rYgy52otuhzPd7pYLMp0A80ujSJJ0fd7fMjSYiSWtaX6tPHvI5bSNOP2PiTWRvH+ZkSPOgAJGRf6
jJB5n/+wuE4+TWjf03i68PAtYolFoLS4Tr5/EXMd94gsXAPDq2KHSZ6HXtSSJ8noh/41OPlD2VDU
COSiUcn49Ogy8sEmY3jo3EkSDfF9MOtioBPI3T8h3zT61h7sFCn+vvUV6q6PO5tv1diXR0leEL9h
SwP28f6WlNWSynJBFjy9oXywqKu88gPKlf74r0kJs3ZQA/49g4MCCQtvUYA9Vnla/lC2dYuZDSIV
6iCsN3sf0M+0tDOCSOOckb2USO7fIsG1tyP7onJ5V+aet2QujLDNxHgAyhGinHjbGUyMdRMFwMwO
LPwwBf+sPwGgs45Cju/Fic2bgc+F/sDpvl0WR8TkNEkfy+Foco38JH2WVsV5fdhEC6DWi03UlHh2
QzE0o/8tvbV7WuUrFYNqgDSfp+IyoV96YDoUOZdysp+Kw3AqEAVly1HCK+zCXDH/jC+brCTDaORr
NBwIHXbsup455x1FSrQ2qRrJEyYfV1+Fpjo7P6cXbWFkswakJuQu0keaOnU45VZRe5OZwL6EN3ox
CjuYJYYG5bO+QJcB2YwBM8Ouo4SwmgXqJz24Gc2hKM208N8U15/ZdcZ9B+WJZioT96/LrAIPJQqG
bBmTbLx43NkpM2/qKTa5BeeInL33R52qHmVUXvLd84bwHKYQs9hkny0cVWVngeEg1rnU/ria+ZaL
9u1BcnJ1AEq+EcJVvAzsnfrbVLI7q/M6wWgXDme8WTGvkng0IPCi89DKYmYcN6Bo5phdLdhXGmqx
Wm8ysEk+fxO2uEsrfewendaqsM4WIuukTiX0lvss9pWyiwAJI1L3/FVG8QsDQss5eSj3nvMMKTIF
3Pxq7cWtWh8n3zLgPgtG/QsAE4uWMKxz/oT/5gycbUtfxoX4qxxcJPwwuakOHi9jbBTC4k+oUvjH
JHADVjPc4Dz8E56xBAoKikbvg3aeayYQNMBpbtwLyJyArJeK7+Fog3vppTuB6MlgtZ1+8raj1z/G
B641aQSNVMWNj6AW9rcy4Qhg3x01oAUuRrN592IkSGye3sELqS/DQKnW/48enRnqs8K4NrWsJY5m
xh9/HIo8z0l7iKQYIRmtF+BUpFxR9Ec3wpx4jNqu+VqJ0bN2Rqw3eWK3JO3ld3m2QYFZwsau5494
PgbUgI12MgWlqb76sCBhvs61uYoQP4gyHPYiZjw3oxmWFHWH0DA6ZeydFNxN/+do5sP6GfIcQQp3
Djptzy+SJ9s5tO0teQWRa1rd9NchE5nxL84U0OzkUG0LZSJ4CZeRxSRvnY18zPADLfzqMHOBoRRr
h4G7cdFFPWDA7pjQSG+/zkilzM0uijnDZNv3NtWpmE3LLWSNMXOmihuwQLyKXio9LeGF5602KCHB
1YsP30Y3Cf8fT0IMlMeUyPUZlhrEOqN2FiWiPG7R5KCTMGbvWqmdNEXBK8yJO3YYA1l9Kl8C0z/H
wT3n7FCHK3EN9ErIbjsB7YfuOXrNk6XwsAiEc3hXXiptWHyfMzufeXBks5+NI/OPyLsJhcHOiNy4
TvQvrT/bM0lrk1n/95F0uSLGGoE8v0d9W8EgcDvAQXGrherME4uSFsUGp9EOxhi7IZILTpgNXke0
1b3fi8zenEOSZeR2qdH7Gy/xIgfwemEhzENBxgLiLh/2yJOCkqOZQtyz6+RAJcz73XqXW+zReKra
NX5GE9bvQK28SC7R7Y3R7Kmq+e232lHXUraMGWo2CecMSiruPUYicODIJSkYBVZvhOxABbBvUImF
p+NkJBIWgoE1KYTIfn5tImHqvcxIY22tSlcchS3M/rEncBc+IYVD5JWDu2J/vDz2AinyrlxuZojy
fF7JkSnrKRTQxUu0iFXwR0p5WVOfQD0aBVrzYG/4St0BLqVnnL52hfUJG+aQrVTX0A8xXMFHsxPb
KhkJt5c6Yd9czUpGegDQrGYI+S1qm1xpPFR7E3ySqDmFsjf/BuCmroKkm1yj7U+bzDTT2KS5BDFL
BF7RPbg9y6jDjXWyli0iqnNLh/ambuYll8y8E7fKZEaPOphZoF+c24FuLDaSw5H+qo2H3SXj0NQe
QHJZX/n3wa7DZsWYFwwpTzXP9vd1MqhvzLlM4dL/r9ZjKf8wVpD8AngIenVl6YFsgdflPoSxU4Fm
CJrW5gFX5aQTEfskr8QACu+gxKNHsTZAMfS4VzqPgEs9gK1x25KSkS2YqUbSxeV9Dsc7cne+tERg
WMwEp+sRHZfM6uiSia3kzAiSmVFCbqjSVBF0eVeV5IpFuM60t5dRHGor8xti4ObW+3769XmQrjfz
sP7eP0M5MLnUQbk/WuxeN6FnVduNm7rbTHEfRd/ljaZ3Kq1fGkrT9D2WShTY6+e3A4OAcOvQEI/t
lAxekq7TAjY5G9KuPrhcu5s4Xvk+u6WbO6C1aYll7e1vQajtNZkZAMbXvfg/Db9gmgJHqAaxaSM2
9erUG++n1JV+edRba7/FymFFTUQNFmE7wiUY3mHGQQ/Xg/1fDtGaeU3HRNEPHS08k48ylfhXZ+Uv
XKQDbrY0SclwC+XloC0hlAFWm8sxJmq3fpVTQTmuQoFXsdV0kxkAoHfpkxAVDhHivV2kRct6uwkq
HfP2C7s26W/uBFeUzqhaWTQyZ9Bou7yuuN4moD9mI00yi7B9fHyOkgVFtpmbybpGMI2xleNVqMoB
0xfW0NUn/IEQjlDTW6e88vYhVs0riJrmVTo//j3KU9z26igR4Fc2zB74opyT31ZT76PI2C+SOU9m
f/TWYRIojnXnaU+lvEWhLYdHXq6MZO6f9BeyDq3RUw2xDnLAQPFnCsfTXnCE1hrnelbaM0oc9Ilq
rdWCnV1iuKiqQz95A0zM6+5SnOcJFQcXCXC5ylcHkkHPbUshA8Os9T3V/AJIm36Upxn6W7L4iHEa
je6sbxR9WRL026l9Hv6chZh28p49xF1Ntqw3d2Ij8NPcH1IJelbo+vZLDJ9wNRIbFADvw+05/DEL
yAT8Ym4+I38313PBC5qp+vkqlfFrm9pfLGR5Zl9x0VfEG0+GdMvfH4U6nA+lfmpUym433ijMUoyl
vbpIiAYBDb+6dNqzRyeYMOEtrzeSSQpjdSnvq+UtaPFYyx1TOVyYIJpCJKIvs4Fpv5bu5fV+A4l3
r/XnEISCSKOAuKcwROwL8DxSmxkmc7+uQzyIS3USrYyAfJUWWv9EYEdQDsIcgw91IXluGg+Zii89
DVRJJgLQaAL1j34UL4poFIQ98sHVAzklIqJh/kRaa2nP2xS8FcneMJFrnRppMTQJay0iPiLI+52o
yOPOmGwjLrqki14RtWNkF9mh1S6HuWBk0Gt11JBvHI9r9APczFN0ZGODBLUGXd7bOmO9JO18RHge
xvxtkdI8kjtKIxtZ6x0xec29HZJOidZMLP/2TWVGnRzYzhmG7B5IiPGsCh1DkHyaV2fxHgmZ5lLk
Af6l+HoNtKotE8HgYIBcHOBX+oCitp+E4yHxEewjA7Wj6/+b6OhShqFl5/fFD+vgyzsvp2OLp5Qg
1ZBtQRUqGBV2r9KUUojyEEFiPOKBu7HH136JcBIQl6s1PdJC4RESgvDOF3cV2Gu8r4uIpNz8/UEd
dDPy5NlX1WV/37FBO30GUp7/OsAc1el8pBZek5puF7W7g5+4kgDodYCGPUaPKPGZpUIMpzC+AudI
dWpr5xhNVGv8puV6tAI6saS+Z1Dj17GRKAc7Ty6NchgJV4kekrXSa6dBTpeFiJHnop1MCZjZWiac
gnq41719ZfY83VcD4jE1CuzXvQ2pGcQhVHXHs6xnoCVVHZkCU3FVN22NC9WJleCReC9fHav4bxnx
jGTsW4QZhyH4F/pOlJXxuuOcEQagmDZZIrDDIjjpoyWxmyMmkfFBPnkXAeNVXCoSSEDUU/EpS7zK
l2RBo1RoOo8p+Ml9sByXozIpQmTU4tEB9oKIGKYQKFD2lzMPK/zEX6kF3WH+ZX1wejYZVMiXpYCr
f6s/GTjtrx1Oj+MUuSBR+04ATtpyKBQRFs26vhMPcFijh+ER64Da4Cg+ICdxFuk/FZJLPYu/4l7N
cspmflLgPTntUFCYW4XlLAeE0BCSWaWHfJ0SocDm8if5S++/p9JZfTjPDNMMexxoCdODgvgXgszD
eJaKHS03LHuK+s+JNUAjOX/76cy25M4IlJ3XfP3icRKt0rx36K3Zon+rdAFNEfT07WY7TXfg+1Qk
1Izn4jqaUVCwzEqlsS8FUjerPdg101aKxLuw7tH2ik3F0R4kID191e8SR15Qs9Cx2w+W4L/hLmIK
SXC8DWOsOfz7tInbMfQRRDC4JgPSMTXShHgog/xZjECpBxH86yLOn+ZDAPOVYVVn3tSYUdyJpEcs
DdXZ69bTs93daOHfaaqBypje1Sz/tUDphb0NnHxHdU/LCZE0vQquJUEwnHS2ECc16qt25Ro/vIy6
q3vfsPDjJDnIcYFDswxloZcx/wrleZ6p2OvHfPiy6DM6WC/Yr8X6hFoY0uAUFtW0m6e80AFIdgnB
XqAFN45oX8PunlL6S+8LizuBduLImAr/l2OyRA7K4LxnHnwXMsBqTta4LILPURLDnGb6QBOild8/
d7EjhrZ0V4pyJDrlz/cJ6AVnPs4aYFzYj/gccgxKTKvqmTvQQoyNZB/6xs3TBXFzqnFGQ6pLbLLR
/JSUSWqQ29nXz2MXoFzxyuv8JDzrk7ghFJb2MvTkRhdFxRFAcRaE9enVYFxMtW85Z7Cx3Bewk/5w
h+PfDpdxDtvV9SiZFcbx/Q2mX9B5BodjyjxzVk5juqkXbnsg70bzKd3dO7Pds2sJ3+XdRp57FWpP
lDP7kSgmSI/qPmuQFEFIHEZzjs96FrD71Vw6m9MNT/oB0G51b+gtWMc/33tkpA6veGx2qhB/MEM3
/WDm1XsaiXLMSE1EA/w68l+1yqIbs4AbeDgGbAAZpjZHtbYkN9ph8CU5GPvlwGZfdI6LVvNwWabu
bKVHow0S07/JjRZnbUnCip0F9FRSR2/p9e2jjNuf212AOwLF1KLRpqX4aY4Cjfpz3lCe/kMdMzCx
Tmy2X6yUITUPHtgopoGCufOMlfIB4vscvvd08Zfytfd1vnpyheSJ1Wjssbimez2RLrNgk1wSB6OK
i1qN7WkrbELDDZwmiK9eTUT0eJoCGoJ0fZbsjO3zu7Ie0jXlVwtfcuhNAaSBPUGUYv0p7jMP4zPV
w8TyDRgER+eb3HUfhTw3YWXcmu7TtNC92zwcYhKpvuhLgMD1q6l33r8Yp1MlL0ZC/MEcCVmDkJ7U
bDDRleQPBRUhfExXDgxbab27jmwLBu3zdCwQgfUluoVGcxYaEnSWFQgDXD5VMy9gYp56Dr86ZUyg
N4qracWGTcDDWt8RA2v6Sa/4uUXVwu+sYDyNMzRsc4jmKEgJNwJqZ4R8M0a3ts9gHxcyPUO4itqQ
YGk1sbD2BD5ggsp9KTjlTE/x8bY2E+wFg6bK2ORIDFZJ/+NCmy7oh1wKTLabdYCSfqLwyezvWMUJ
yZZPhDC5DJuOFi0UBQc5WHM8l+fHNa4Q5T98iTj00QFLsJXfbq3j64bmT7hkLZIwiBzz1nJJFn57
SX4oiVZ75Q7QfX8cmeTqZO7aePhf28jqaog7p4iNp+ZWZ/nIWvYtTH8deaPEoobrVszkZ0mIsjxW
bl3A5kjMN0KvdgFMNCpWnuVKZ712ZtMdODe3eu04LN7XF0Gww2njNuCygU2UdWr4ixftXaTeK4cm
DrgjzTNya4NiwXCH96R4qR6akD2p+sSpWorJ7hnUxQ7Sok2P0XjLVgTLnUDxN5a77QsIfGle3q1b
rRvHqE1VMP3haGaQYphuQYIQBDBZJ5x9RF6hNz1RKPTl0BuKTl/qFyU/Rl8xHcyPqIHO2XMFdQff
3zzQy8j3+ZnM/cnN0c0FXhbFpGTbM+dl46dJHsg6EZJy2oXs7DSh5i/RfiL9JFJDp+J/rOpGbY9i
M3gfsx22sQ3cBNNfT/qlectmStNGTQojqLuhrT41RKrIqqhVzttu/UG4mDSUx2fcXw2oI8e5E/Ll
O8sNd0ZpeJDKOGLPTs1UrXBLrtWDtNdk4VZ7Qnl4SXe69PA7nTiF/1GIwAz7xl35Jmu5mIBIr/5F
ZPhCsnaMWwkB0uCsW6c9jIbI0yw8ShBqhj0lrHxH2TLK3Rsj/5hEhpnCrWkoHu5NedYh2K+5eyOh
j+sUVNXgNf09AOSCENa8f6KpPkuqcE74o+ol5IEyqZ9jeG9rdOVGhlqsLOa+znq82FMXdanuexUb
/4H+3iZWK3mGGRVS1Y4Q31N0u2pdT+RE9akNQNBML824ewNQNfmypnNHgEN7eB2i9i76LTtTw4BH
UWWpKAiUmE3xCg/trX4nx/nNi9ZKDbUZYoBhWTkaPSyCRsrxiGJqHs1nSQ0CkWBWLN9MIwcTtAjH
9+IA4SbJGXcVxlF1Yd3nfT4qN//AWeHQZBfmxtnflqfMrZAODuUjv1khucdECB7SCyWGqshENVF0
/Q47wMFfY74LauDMo59hAKmnM8MZiUdjFRxVXZGDn1TK1dn8p563pEnAO7e6VtvNjH5h1Wzt/XYL
rBU9MQgPi+REuEM2Yzas5oP23+GhDAVoGHL294zsxhlxnuhS2fNrp7CX+RD9XGAGgDU+Qd93oYHR
K7rYsw+kcjxgwwRKrnSqao1zsQPt1kIvUtddZfdJs6nxPyg/dio3TDf/lCzRB0QuM95EGD11O6lz
K1as/wr0TwnpamhV7XFvboJmnIBRZgCFCgUZwN2qcZJm7lL56ve2DhmxSpM+c+ZNgNaq2zABXqUm
IaevwCrrPLJKp2f4uguVSZB4wYwqUjZhioxYfpr6q6Fn6H41mbRrIPSCmoiqmYd6LypcqycabIFo
B2y1ueDk2EBxzaTW+z1GAI92NStsHHuz57NCMIDqLhu5/TfMwqL3PAm1HhudjypqCkBTx4ebZjkU
ARdllbdJknqwzLM2rKlN7dgXJr9kgV4XojAOs8Ai4fTnrXNOOArH0ETxCQwfwzKGzo3BcoeA8ijJ
/Dfs8ndY6JaYGT+U3TG0gh/qB4VaasF8UrpGpXX+9XcJUm6i7zg7N6gKj5W0fX3HDP69K23DGITD
x38Q1zIpkhOBMapO2kKALvrkm1igkhrG/q7PLRQr033J5whzBsEIG6zE3nD/lIGHHjXehgN+sarY
QT7FzDeTCWa/HGLPUq0vCiqIytJbHtVK1eWkWPzaEkl5GrXl00ykVVIu6KJ805Xr85UcvzegFQwk
5c2EdKfRtbE4M4VQBL+ffXhhHhNN55w/HGBVNZTHUCvQwdAd9M+GfLTHgMoGAS7zWxZFn+ByDQk5
uaMdS0Gp6GmstoiTeo3JpHkD5skskMO0lKDD1kQEjwuJeT66+YJN6WzB0BqHCVvLRd13aSCsoccc
7qq22Wor0FXpkFbe7iwqL5XNjkiNtnvahiWsn/EQ+RzlDVZ1F8gwwsvroQvTz5xumag+13COvFGt
VstlOYqqDcOO+k1ugpQ8oVlAOKRAxLgZhNnzlI70Jw5MmMZdPOolQyErB4a3YoQN/pVP+V4jhcUj
X8nrGFP0Bv5pKo6PR5XmF79uOMuv0QS3Rny+WyjfPS0RObHm7G0t/fVilWUhafZxkwGpoj4rgqq7
jVTbmd5vaUkw4Ye35HUcJrdclu5Bmy2LQs50NLsKMp515OUoG7SOnygs7Pd7khBiJDoxHzgDupiw
DWWVyIx9mX27pFGeJL1Zfc507u1WWI+NFKaFzHR3BHxRtPKmczvQyF1kWp2ujTKuFeT4jVsYH8Vv
N9ODf4jKEax3AUYUWXLzvSPiK31AM21pde5l9b9oFPXYqY+6qq7ePjpwvj0kbFEO0V9HfVnlLSfc
X+/0aJLPQtCJcgALYB747Wu3WHoBwfOgKEuABCl2m3WmmshorwNbYslp/KsiXTfVxgal3d4OnPYV
dke85BjDUJ4N1gXiRIOO+sf47ldRk6LHKttwZqo+acBroCPkteIm0ygbbka9crFWD5Ta7FkW8M0W
luyGD327n1K7xETAP8D4tSfSOD9CzD/f6Vo3le26wqjcc3hR5hmSyiVTqCOKU4ttrXxI9OdZYZXU
iTjWPPXTWKkdaRiPpl7OTF3cV6/FVIxWtxBRj86D3xq8TZKbk8oOlILQhDFJmyVVdjnA0wA2X7fz
ADW8kvXmRigO2MNg9fcTyx4aNU1viHWBhXgL8saieQFgM+FK3JXBShjUrQDzCcMfTMqXCemE6ThW
2djy6tmqCZa7T4+E6/ei1iXhYWKeMxD2lUT7UhvIPrQD8j9kSNInD/6tdTNR8DBuvSGYhKi7xjun
AfW79ktThaXSkW+P+hIBQX1eQ3SoxlGrQADAggkCGHfOikUJnZF+scyHIbIwEhPw9cHSnAww/782
+WB1dM3mQ08w0jjVrJDfzKWRHiDi93hZMn48TcrBRw40ZCkHseEFpOBuGcyROTdRljVHlpc1n8TZ
fxZN8OEsKtj/r2ADfhgroNjb7Fn6hzUZx6Q8oiohlJlKaMFQbIEW0klI8HRrgdtXijz23F4f1yOm
uLTu380tTJq6vP5J2MyRLsitWdOY/NxyLAV72oIx4Mo0vL6YWwwYihFO+zjesaGWUmMyNfWZykiv
bsEV0/qWtHDl3d8MT7almggQWrBb9tkJs3iMBvJlQv9rIrA/sMvyFmmNryBR/fMJxL1YKcNZnbJI
PooORk7a6H2W4reVHdO1Wm7Xz2aYkGzG+v/A+lNViOkN8zKQ9BJ23yDus06KHRIJ58kW/mL6N6bH
gdWhqjXCw6KG/kR4QAC9GLBhImdRwBQcSWlBRE5E7ocx1AstQTDlqFIM0FDP87MBBJ4FAdeQ3K6o
YoDUMI9Q9jcEqk2xa/i2kZ/jU8hZrXEWwuwJc4ph/Hrh2q6Re2rLXRAjr9OZyfK3xw2Bs9abEDiW
9y71VMbKlchAiufgjy0lrrKrQhSYmfkTmhssQJXvD/0DwUP9pxtxLHRO8MfEChUMqFT4ry3SJT3P
QgPqoxhhZe9qdjg7La1Sf+zSJD6uwRQlYBHxtUvWCZWHCqJyCSX+FGgQduVoBfeyTt4D8STtxqyw
W9gcWURL7/5g1OdrSJij9Yhf9CyJRlBoZTyGY03QVO256pbf9UZmpbBxkPURihSmxn5pDChe9WOy
9FndWpVUqugXCLdv5qKmUDWTeW+R2PiFtR7pkclWQfBFjnW+6qKKM3Wf98igVkpfBi7Jmc3y2Hiz
dkHRKMXCvPzEo4F+yz5jCMMv8RArAMMAskFExYYNstUha4rGGIQONoqTCwOpyHxaNowZB+47cjVZ
Q8BWrmWwW5dkUd2K2WLselRt01NTrDaQ1OP87NoKA3Y3BpY+/K1QEi0vHERrwiB0ITJQjgVJA8F/
rsX9JC253HcIuTYlA+g2/cMeWMQMQDqmf0bnkMgGN05vX2eS5+dTBPU+rXkrilHbrgsGd37CrbyY
/ryOv50NoxFzWuQwjUjXkRPpWs4n+h4Dix385CPGXqHDAtoiFv68X39m3TMefAd9Gv7t8rH+tJRp
S1OL4pQ6ak2dMV8rUPfulwCXAGp0TsxeydZ8LIHVF/ohcp72D8r8EZxNdK+5W29gLUEyydD08EuR
x1z/BpGodhupqZqPq0umNTIGXlYVlWCpUx4gL+xKatZu6Zq55PcK81cUTZSzGw2CQJuGH8oE7jRp
l4AN9JfKxalD2m/l5EsDM48sr0xoxiO0VXe5/te1HbNQ/bviRKm0l/0aIXZ52q5M5yAIlqWVd2Ib
PCo5m0coy8XJFKADso7yMEi2O+8ENd4x+BcCZor6SKo5JRm9CH+zhgXmxXL1GHWXhpw116ixyVB1
YCTKxEJY22l+2Wi8NbibrtZnsb+RuDlTVVueDj9STIR72takK3JUgFYSF5sgMr4rZodoSt1oqfxk
F4BuRLqDDdEuqfJ6o0TQVba1Clw8x/5QQwABd/9OCjc1a9PC7+6BjRpetmza28mH5/Vu5bi9d0TG
QrdkApnoKWPdvfox9VHBoe9o4Nbh8EfUPk02oqjvgpMxcEYhSqnWlYTtYHSIFn1kaCBX2vtCKmsH
rfqyBirApD+7cSLXEC+4lfDwPRwdw2FBSZi+JgT5AaVDmY3jPQ29CPCryntdQBBeC3h02mbZ5O7w
N82ZN3ml3rntgSG1TMU+Icf8HajioBDhv9khVy7JF2cqXhBNJiLuVsbXknJwusKDW4+FZD5qm2cd
JqI3Kp4A3UV4cZKZmKimagYcB7OdrP31Hgr/gtDiiG5O0Tv9AaLi3p+RHIfqzG3kriDn8WksojVA
or4hVb20nApor4woKKW/emYve1vb0bm5UbMb3Gsi3jewWW+lTdU8icXyPkoRkCQ1VStkHJm27iCP
zYukdXeV06F+i4VWZ0Lu2RBLeqzq+Uw+zCm7aHE9Smx6uLIsGfDIdB9xS/P33sH+At+/9rtto/m1
dI4avz5DT8F25aaqYthtINAVA8TfwkRlzU3xleag3jaYbJXdbomgLLY9y3sqeBwQKput+pUeT7Ur
GpiCPdyGR3Akzx5BTmNW11RyAFAxXtLOY7tUTG9IcyuSggtUp/ScDYtjahD88Ui50D71liwqv6wc
DeXwDrplSwAqwSTK8glDG+cwiIetDObuZUtha4Ln6W0/qICuaNefP0x6Cq04wRJeRoZ3dlvIxWPJ
9wwNucWt9eNwHuYEnAKhY2y/qLrpeaNwCTBIOr+j/l8OwV1iUqG9FU6F7zBJtR5DHrz7s9ahX7L7
ZON5u+xuy+/qI7gWHEXoFz4rJgtkZTlE+o4EYyE3sW5O6Pn5/p46c32yXWaZERW62jY+sOj6pVa5
okR3rqqgl01D4Gdkk8aicmRV+mHNdosdrK5E3ene0i0VwQ+bhTLOlDFhgfHSXjfDcTrc8n4s3IGZ
s1xtbvRh1euViCTV9qd5A4Rn3GATHWvFyNVrYeXiqSdV9jHhotrQBB+/DWJQL0xS7Ixbrbr0W9US
cs36NRYuljcGPus9Vcd8ZIpPRNCEcghdBH0OHEAP5u9j3GsA99KPqBZaX4TgQ16iWcok8N9xVt8J
6ZObF6/ThLepbgBcvmQBb6HiORDVet9ejbxvgv6ZccrjqVNomqWhAGEd+0gUuLD2pMQuAuxtjQoy
uj1NMavMIXrYdalR+PpjdsRwYu1uVD3M+N4lBjdR7kM4xCL/2SueBuvRcvKFljRvVTNhE+nbHUvY
NdSl3ESL6PGpRGehZkh+dwcHtJ/e+CZuyPspwJgsIYgRNVezfOfu3F+rvSU/zs9wdAixZ3gUvvQD
7oiaiSGVptjtnvdVVKfqjZxWN0beh9+cokueer0+EI5liWKLup80r04CGsel63ao/1ztDaKikG/o
uftwB71ByrIMrcpACDQ23JLg0AHUcqqP3dwl5MMQCfWYPEmh8+ynnM6EJSYIiQrQZE5o0MZbYxvi
MV15WTRqg/bCt78WTNYvmvc9/WUikISWP+eztMaNeVBqQiCn4hWcD7P/oandGWbipBvTZo/Z2E43
8ODE4g8/ZnzggVYQNwPn6BILJDUZX2TO7t/SClTrPJrtEbDUpcntooxgl5rfDetPgVJG7D1V+cMx
nlx7stAInSJoML4yEe17DItuk+3BRyhmPx9gR88bE94DXupKbI9C+VWy7Xdohtby4Sw6S3seOfGZ
VUBJFSay7a76wb+nJrEWNUUxWyalGJL0i6UkrpuGLYy0VG3Iev58HjPEClYqbU+cTvNTZSJ1jg13
eb27SN6BM8AxlZHvCEcnxI3jYM917RA8s9gwqQD5ZHG1W1P9SZizTJwiB11cMnAQS/wP0rTZ35PH
96xY2/BfozNHDguV9B+KFluB8qiTsfJhRKNT/68qsL+gAfk2g2kfUrXGqL5auREq10KErHQJ90/c
5r7+Rf0wt+PoS65gQvW9SXwVk8D4j86fRIw5pmM+XwNwa+QJtfC17yqrpC+l2HOJo4p1ugnRXhj4
awqJXIKvCheeYdCCsAoovG9OO3ZJYfM8kM4Q4XK7jCg+V0sBT0ZI77MKJsNPBcwaqNBr5iLjQdHg
AX61KvpkFJySEYSfEkpi5+8o1mGpPvrdZjT/5uowmriaBnB98DwpT3duk/3qu4B9gaeYZ6pRixcb
L7N1fIqw1LEHECHJy1twIBUCqyuTUH4/idnus+H0qhYmZkNgiMGywRAL/qzeiugufPP2Qq7JRU/O
UHUWHKLqJ21g5hOawPvpS6Cq/Gg2/6lEIkCzt8lQ4OBB5sTPSYqXamYAD1EYKPZLk25QMbqO/BtE
Lvy4wWJwQSmE8nm5EWYa2TRSXVvJ7WrKjSF/zpQSQqj904uryzpVGB3tiBKM1E/v5aH8ZMeZ754x
/r3LO56ixsik5HTPzQ6U1ulZ4M+pSCe+qNjkJToL5snMLx0FY38Vc1/SCH7/AVMDrfDV45bt+PRR
lnwQAyBQ0d0eRSWt9fQUh8POa3o0pEhP/hcYdON4hJa87dvaqrUMsDkFJ4OEp7yG/wovuBMQD6Es
Wib49eDUJDFpcxJjvOl+gYAbzlXgHnlLnIvYksCDCQg78No4G9fRsK/mqSHzsZ0RRDb1Im6qxGjQ
t9ow/xb62DTO+NPwQsUVzpEIqh2LZ6BkHpdAq9TJBojBbv6hYQgf8yVHdiPZ05SAm8pHe72R231P
dV13SjRv9dm8uUmKItMo3NXua1N+uAopHn7gP/q/aKRmiKmxiYd2o2zFkVQ+pi2v2JnB4WWU15ZL
JmI2WL/3E3rZNMEH4e1d+yOC6YFEZCvupIAB33JhJjLK16NrS81FGw07dC67ksX/yXBYt+M0BivL
duEl4cN+726RSDbPDJEhVfx3IfRjZfNlGc2i2teg//ZoM6M4rP/fNl8eBrSm7qo9us3T/xxBqIMW
9Y+FlGFjB03vBTjotK80vY/Ou9GARCblMZrSJUQNrnviOuUlzwUsGMr7TlJoMyzULoAspV3AZXDf
ZwLViTIYPjzQ2oIRVQtGmTSbo+GTFw1bNzbV9pCioOmViI9KILvtpeHDzzSAwLSPknPENFMRc0c8
JZKMULlZtA2eekokdtsmlfGtgxljlIpordiSIferSw8qG2R7KlK+iql/aHBxqKrUkTwUrmNsrZRg
98h5Fw/CGwIx+dVl5Wby7f2xXdYWeUAikmgWlSrAI9guozlw2uGOzZomnd3tBBCZUVuiITRWQXJH
IRNavFO1dJjWpgWSYf3o0robup0hgDnZLqQkO+ej/0E5mZ6eB6KCv200Wiy8OOqO1gKfIzETdQJ4
83PF5GZZZ0sm3ifWq9wSK//VyfKeaiOv/g+0sq4hSv3OpJoH0x9H/IwkGRyNKk6FnXzAun9OI1Xc
tQqrglzpIZbsQGlcKrjdTu1aavZ9kxL91S9vWofRrOl/I7aAZjCtfNyBagsfGYTmEdQDMeiFwneZ
Nh4ES2F6puHlEZ2GUlMvp9p/ETtJcPsAHWAo6BfH/jBSKIwnjV0QkvyZ8MOiyDXY00gWYTeKGXeo
xgfX60ITL+bwjQ4OusIEyM/vwmTXSlAl+jOFaw8NDVN0DCYdlMPP4nMo8GCEUhEckkgCwVCMTcpN
1azjjtJ0Z1KLEXM5Pe04Zf1VTVmOnCarlSPOWNPiM5hQwWaic4Zpeg+NK5Lpz8z77qjF1YcyL5J9
zOe7+FgE7DpYbfTzspPATWBRMqqGCj/x3PK8C9/AuEveY4GTpAP8BoOuyxv5wPGphqOMjLMPWuYM
zCjj3BsqzdKqIjM0koBzFqmvepvyrGff24mXiPZCXEjPTx8gwjO/tTrD1zLElyburKmaP1Q2T7HI
JCW3CBrXvNGYiYa/tZN+FuqgcVzDdzLjdUEJ4nk4weLm3jPQIDjBN95DmreRTNEUACBZmhA7J+yF
2/4vFzt05KQojKkV6l3AnaLGebtzCMrQES9u98GAyiqijPIQE3nucHlQHR03fR4mk8pHv289+Roc
EXcCBEXR/d7MCsftebohsdB2iBajLzHNU5YzhLyqfKNM+fKbCsSNIIXpfQXFD+RDsjB/Z2i/5xOS
6y616zXZ1vsmdBIM1E34XnzoAdbL4fxDp5UxbhnXOe6cN+/gPy4v1CxcR97MXaCONbppjKRaYfyF
KFx5/ocq1XtztGcmLalwmi4D4md7APaQyBfBmvF1pzHbnuxFEHhlxftXAB+8wNtrPOa9WK0OHQay
NY1FLo01/lDQOHMYd2ED5tMfYXJSxC3jr+Ex8O//kU2BoHwBcmzHiqW5WLbCoS8FXe6QaWDUuOJm
CVRkPc9uNocJPADsSfvDYPyApXJVbxkFjMcr1Hb8k60ILmEbqQOTR+y8pU1LorojJ5uUroFzkRDs
fv6IVLe/X2yfqg5DrgqHOVHhp+aHCcwXLiLBRSCbHyDXz35HTRcYIDy/qMOqlEnMOWKBty+JdJIa
+ZeM1JVPUpmOR+dv7s+AaMyPCrjaeo/7nXRheMiWJHTOP2kvle/G9JSfaR+G+buE77eskOqrnWjJ
vyjP1Zce41NQZkRXYNX4PomBt+MjLEgiCOe3tK9ljmLa0y3sTx8U5cOBOSCT38J2XO/I7/R9WDAY
5Sits5CTgYzN/8kqGjtIRNxWeG6Bjk5WVObUuBrTV4Es8R63O1NbeI8wue0JrqFLoQpVVpHj7Bp2
KEa2vgKY0vGOnEytHi2b5gsWU8xmXks4yY/X1BWjKCK5K5RWpAxVdL202e0n2VLIX8nPVFfsDrea
gQg/YvN0W69/wT2fZ879u4Abq6tnXU9PxpzQp9cPWGS77OKwui75Y7MTJRJ5Ch89f7MB+3FUZvzc
sVsHD7Hch8TCTZd740Zms9RFYEL20PxoaimiQsZAifxe5dIt3b7orsfU5DtA9A8VqAF+ptOEnfAb
LkyLzZN/38mqwa1G/CRgm9VS5WfBMe4erIO4A9wsi2AudEg9m+ByH0h8WX8NvZBorvv9c1OUeyFi
MZEek9W4axdgbvoAaEInUUVxBxBwDEGQ0tvNDBzFHNRsy/VhzwioJqOE6eRaeaUq3sF7W6YLUmjr
yUvLUzF9WwVk6NnextdM/ph/qon4QWGnOiuhP2bzyAjUyQrqIQ7ht+RHohh/u1OomqYOoAbq0QQq
Q9ztVjvTfHPmkZTTiSE1YIBr0b30YqyazT8VV1bovY3L5h12CJuySPXACup61TexmmeeGiu2QMdN
/9jlY4fhvbBZm8urcUM4F3JbIqZppTknpNGLSYquYlz834984D25EJDuk/XwB5zjTrcHhilRyd48
PDjqyUOjnJVXCOH2+8j0ENyiT1PAAebAA/BUrbqY/mRDQ0qwoYzWCQAv0J5ZzVv3wGUfbYTwpVG7
azOPOh+s6EDIuFRbqHqdzDyl84wjTUtb83R7k/WWLoUq3zx71S7JdNd73LHCIdkO2dk1I3qTryVC
eW48hNUvJLcjQjQslYcBQhSiHt7rgxeLPm/dsyC1kCQ5FcndYuDci3Vvw5Ki9DA3Xo0bhfHXhrMN
ebdMBq7FK4Ag6bMpk9iQdKJm+QCUN5UBh+JTuVBlacQGxnQG6gmUZ1Wft9bNp0fTRL83yWpYvHOp
YRnNiyp2elVeW/y4neI10rn2A0pO/KlhISN2t3UCUVSEMCfNwlCjqmiKYygoRTYQ2LDDpjbmMwpt
2nWz0ePWHy4YdGWk07FymXB9nu4zC3Ih0yHaBruPebZAO3z8fc0c8YB2DZ/r73WoevbZpM55qbG1
5uIycImiBhMHJaX98fU8uNRLKEtinJkQl/Gcb8zwYEVmdxuRFD26kBhawcdwY7fgArmVOXqmirRf
ZKNwh2sLP8uOvcjU6wGLvC3PaJ/w63NqC8GSHRBEGoyrveMh0JYMLsE9DEF7SnANOzdL68M48trz
cJSLQnjJg7BNAjO/l2oLCKjtvgL7FGO+nsZUHA2xSIrBs/4wL3RFEHjWhU2TVA+KJYmmY22adax6
g7bRP0DgYUb1dZPHJs6aORsNIPTg4r0zpcV6A8lt1MC9PzYlEfA/eqdX9jvOf1HtHz5uu0/1490v
esoyHCYgDwiHhxLXvlAcG39axmAY+WJZsXCzvnHY7Ua2AakK5Zl94oN3e94g9sXwhmntA1J0pG1d
krxkBdJIJBcQcjm2gdjBIkyuQEljc1WcafdNHwmnhC8jegD9HbUS4eEtDxbmFGqVw+gNpBEOoBzV
WbP87Gch1iu2rsQ2bZkRH3Hr4lKJM1l60XxAMKu6n1nQx+JxyFrsPPafJx6+Z2ejWwt/l5gRPHVt
AcwueZbVUHvwq0aShbIV6ba2HlUPg1BthCfBUtZdGcQw+ardTsrxjuTsuc/CpMLZpLfkDMfoT/I7
kwmGH/SIdtqaqT+pM70mkpCn/V8L/Bwhb8vsU+Y9/jUssSy5nesmx9cdA2ehgq1hhbVK3k3DZFiM
hb0AaL+znHNEwbOK06sH4jO4TzOZ59tjDeOTjOU/GtGD3gljP8zTwYHTY01Izz/bsEGPVrgAOC/S
ZakEuIabqxI3aZhShQRPZl/F62np43A/ptvIpJBmuSAjj/1cyEkXAwZzG3Rxs9JPL/2noMP6B9dH
2JC3aBq25J8n/bEIuTRuFUt5qGQYmdDcA+w8wm94aDYHKBsEgoBzJUM8cZ7ItL/ofWkPLrdIUho5
2LBix62uum9EEvqiHPX+g16tIp+D6WmXioDUiEie5NszoD0A4COENwrKqR9CKWij7GfXzEouB247
CJVh+BEWtQ6wQyMyGU0X7spKTm9sfwh3wOyvjtljbcVTGcPFZDzHK/LvpJm61sM07y5oHVoeO8JN
u19McqjDKRfjY5CSr6nO0/6rOMgC3wBrjbLSzmdu6Iz3xlGRdxcICHLO+9C1Ioj9Hzk/FLuGKLoe
0WU/W6rqeXcm/qj0kaEaVSSje2orpKStn6gL/DWtf4HICjISixMNQutuga5IK7+c1ry1bnJPlrMl
szbwJuCIRezllRjdlfSltjqA0xR/hODRcH2h2DaHcs9bB1Xh5KqyydgQvmEIdEU7g4VIkaXz/7Yq
7Q16+TCaHerCiODhOBkWCnQ1NPlYexPd/dxUjLfbD5DhjT1EHMiSyXqbPTaWki5rGdzta+Y6o+tL
iUyMlqveoW2gP68EG/58gjNP3ht94T5fmUL5cl4WIZXJg5xAwQ0kENc+lYVc33eIRAW4VFuWDZ1j
svvr/Gwj5gXZ8+S/jcdahC3N/TfQ4zgTYx8POWrJe9vWJXalwyz3cAk5XWKInuQRpmeu15TakyCS
6liGqWmEs4dVfWyrdZo1RMioaXaC3fB1DsnIZcxoqO+bE1mubMOrD9DaJPvaofVK6JIjDO5S2uSp
gLzzuKtuY+U3pbm1k0JZBFeRuEAseNcQbcTCqn9m28JKyXKbpDEbTZdpKp4UT7TXCi4febL5bifn
RsCad1qo3L9OWxQz/B9Qe0suAlTmAd0d3CTSOPFVcCRzCeHNjwDzA/OiLOZodfBKbdkAZ+rYCVBZ
hwKa4Lhng/7bZdMEGCi3H1hbYKqnn0sM/+TtHIiqF6Ck4tPf8+QftIbhyCWj8CQC8IKWxbllyabX
N1ETIkqUZnqk0LUQroykz6NwJyDoow6QG4woQ17HuOjsmMzkC9qY0HId7QaUVRiO9WWPl4VKn0NZ
0DgrV31H1OWymz7tyxeo1yOEfPniTAWn7fw1flU/oGRqlqz7Z+6+P7iZ8PDIOrVfXgW1VtieN+Uq
LKKHdnLnF+3daE4lKWSc8EeXk75qQzBq8eKswTD/wDnyxXtcJbCGy7gFLBU5bL89GYdSUYd5o8b6
xiugS0ChpCPeYA9MieZZuyho/V74NVNnoqjESQaHJ+qrI3yuTJDo22fGyuzXAX21z6xg9bHdkNpU
uaTZu6UGxXmkltERQpOcoJjRI9/Gskebsn2jFkhIa+R+I5R/TMVVvJPsI6ZGQRHmVG9zVLMDd4rm
3NE4QW41iXF0LAW/EhYNtdPjy/Y5Xl0IGSIu7ukysvKHL/6JXyVLFOeM2Gne5JlWx1flThB9GIPs
s0ZK8bhUv9OGT6rItChjz4v+C7d7XHIzweTmOG7LhK5MHGNVk8992vC4nXGwkfQ2j3ud+s8I1sRJ
4ot8+siNt0baZWAOkno+ijyrgGavevTzppiSu9qnWSxg04ooq2ucIu3e45BKx5be/1UkV3Rsv8mf
CAIQJaInB8ZhP5HWy1Gt9YEuZNVnReiUvNgdOEQU6DYdNVgEq5h5/jeMvD9riUhtpeF/bT0nsVQO
Y61cHBM3csD4Gf6a4Y+0Ja2i8L092kXqWfGUhtc3bToiFwnwXwwN+/kydTvgfCfilCwL8OP8e5KZ
l300sxVFBQH3CDzUL78uqg7uZF0pwGsoisAB2JQMg91EA1GNGlB9jEgtuoyyfAZ1dzwVqwGxkwHE
rt1Vt9ghk1/0S+VcJ3sZuLWFr4rUn0YaG5g0vxd6A1T6keV5fzHCFoqWaXP5ClNTBTAh84p0UGrp
FqS+h4so3vg2XHDm9SMj2pVob1mYtTiZSqDq43hmhn1Z7Po8bJ30CF8Bl8GxoHmw2wpZBMJPG4S/
zHbkIqVGuQB2UUUM1or/4/lq6t/7hAkkelCwB3nh3vebJ7OFIN4XfxuwdAzsnfo8vhB/Jdyopgv+
EoQqaJiEI6Z0nVOcBXRbULokSWQqjAfpFX1GFQyQGJlYrD3PSWU9+GChYkmJPpvNl8zw98NOc8Zk
HO76AfWO8TTLePd3wYfMh55ZuTQL84Rnkf3I5vAeTY5TcdbApgcMI3+mhzktgq8mGKse+QYHJOAH
x/ULhTr20O/1udlHboa/aeMjn2a2Cqe70UhIeOn472yxi6hm5l5oaI8EzZJ0qAcwctrid9cciD7c
YPv0tEDvnGfnHkFjIXmtzDKOTdnMqYyBCz2ijhdTKeR94A+soVpCgFZvsVA+Kc4fXDdAp/+DDe4X
eOxHwG3cMQhqlflyOa90ZWP/fQLye4nvsv4+IiD8wcvwi/xal1VK3qbiOzj0BSdb0nUjSwHhdRdA
iUzagWKH8uMvsrOkDvGCAzBFTnj7gsMj7dLiRZ+ry60T7K4CxwSYCB5WYBB0NwvT2BSxdITTo2cN
9HDeA7J3IaARxbjHxHaadsugYmaJjVHD5p49AybNQ5j/MGUhHQ0XE+KWxQj38S4tzHrw3UJcXoh8
bKi09GPosVEB2UuGk7QeYiKS3V0CZ0rqH0acPoAcRT6DfyrdPrzMXJXiw9Cc/juuErKBJzN24m//
aoafKATI3gbtnm2oCF8XGsYfPzPUn3GwumNVkrY1BXblp9Khz1IXTtE516l/rBsAp2k3Hv0VQjmR
ow4w8o/kv06BLa9/FlPhVrLFuvE188ZWzsrVwHFTOmAfWnIOhhF7x6puu8oAEQkGw6MnSq5wAEJv
0dgK7DcYZtz3TnjwHoKk1P31FJLZj8GX4uaEVap2CMesf5+DlVrreCqQ+7Yi6NE7gGPAOPGAPigT
duaBq6HJydjMlILfAXjXZPe8J3kRvpq6egV0yIUAMQjJ73Bb2lSF5vhXa7XvzECWPOesP4uYLI8y
hCkSpC33pW6qmfmNi9PaTldeRDALkVl+R+bdVmU+1nxAk3pmL9RwtirbkQD0odFYlngMCeZUR7hv
YbOeydMuGGd7T/km1BPf9cJ74gU84h+aF0StXlsEOYIoQYznm9Y7OhRvNS1E+esLJi2GiG1Xed4N
cUYbgpBKAowgq5xcVHkgu3BCSQt/1CHAabmaJU95ndSnIZ9b7nuqk6RD4TtBf8XtuIP5x+8VOgHj
THI/3GqwB/2wRC8SmZ8cjbdzQORP7qZRcwLbDcY+jblJO1a5IaAcUIGsQVaq014St3JAWaalXzNC
ZSWgCdaOA2nqIN1iphtmQfzZ27MhG37qN5V/O/VTzcSnSEdAnGHTOOsPjebBJozbBWaFfkhzYzHM
sHetwuzyCPmLjX4m78uUAXtmbTsrzybwVzZlZiP0Zei3FTS0VwTVsYz8uEty4V2tzDLnSgvdaS0X
S+Fn873aGT9M8IDIIfCG3uTRAYUk1mTGhEAauaSXmqwlmKOOKwe/3D9EeVCbJ/WqGG+n7ocTgWGF
kxD/TNTGggX2qP6cYi/M+iNIJ8jiMapExZoa3O3JsDiHNhnCl+VzC7KpOumpt3Eybz2qisR++lWX
RYWy0N8aejzI1TK7HeKhqfU2ZwYeQx3m+Tr29v4rxUfWNCWAee0yUXmiFiz+pwGmgmq0o1TSq1mM
UDxtzg5+ystLFjmebQmiSZgG4j8GY1gaBEXWf2FdAfSZEtNq1pWoQn0Dgy6XixFg0qCr7Hs0Nffy
C3Tt+D2jbTUWP+h9Xbocm3v6Ondj66wtaIIpiFx9O09Hats+IKZLex80XIpjln0teFb8y5Susjb3
MbG6mtvmTbR2bihr8mOWypbYDtdwTxXz9Jv/vZG8yS9DSSAbYj7tSLNGf8ndFokK3kCxkbumsVrL
DTi9nYHaB8QtA20u2buefWkZLWZzRnaMgWn/mwGo7ICDBgSDvXpQWrOybZYsEp00b/ZzF/VXQYGt
VPoc2zioT7NZxYt5c+zn1LV0KkXpnvHxg3S4Ezj+T61pLBRJsND+Gky2aGOKkBzcbKww5iuXhNqH
xgTe5njFfVfDektOrmi3L2OdlCpYbEKENp8PPOx41yI33LHomoQEejqexG8DMD99aOdWYusRMZeM
GDAbRDU77O2C086P20ouKKYuk4BMP/47N9R9kHOvL745GC4tDg0KhUYzs1cLemEKtnkx5ojF2PKL
F0vz3QzXNxIWRdL8royYhFgxCXW0hWwLMuX7pFeFFw//oGkHFZ2Ryj9hOlTP0TVwQpHK30YVKO7g
51mtnvXb5yGeQ0upP0TRd98gZUvw7cvGYsFx84RYZIEKsN3y/kga9KnLVhqz383ef6c4zi9UfkIV
odcLF8Mls+zsmOP3hJ9BaLEREH3EnCh5VYUyjQh6wRcAPWzRQWvSuvG6SN0YoncBAFHxUA+a25nt
CT4In6di8ghGI6WGoURi4LeWj5btgeDlCcyWeC6deOjCR/7FNBVbMbiImiNJ7GwgHGJ3t/ejwL66
VW37BH676We+d1WEpEfLInYhp3rXrjrzyJzjwix/fROentIEkGbdgdCEOKtzPrr5yKQmHBPnC8aV
LTa/4ZHcZLVFjrBYNOgIsxPuCiAbb6U3RlOfAbeo4VGm8/xMzSaPQfIDWLbp/2dv7gmHFVlNBcrc
01lAHx2yVSG0HGa8AKtPEGUZOJlZHydIjqjWIqfF008pfZ2ayW45KsF6J3dlwNp9DcBsli6k1OaD
qQLp46cV0GQj6OpDLRP/9Pxf9UmNL20N9+nPS9/CfHBknkomwCrcQ02MWliqCWO0lPUy52QNqNWu
c0zP7y2FGwy78QDL9OCIHKwGatA+GV8P9mvkL4zLS/MnqguJKakMWvWmUzGEQbRBOFYBOgPkmiL2
gIU/kUDljs9tDCZq6EzmUkGsuD84n2oZaZ88ZE2mYK+SCV+UpT97Rfdrvb1WWaFzV0bucTFyktw7
RiJW+s8X23c8QQ940te+BpXpmb4O/YPFFFfDC90h2oS6YgP3SVAT08bw10h3ntvzTnx/g+BmKbSh
X++wG0Rot1HmERzTxGjWTzL4jug4JJQmqNZnAuYtLGAqm8If4+p67nGe4bMUAN/YwlUTbymEw+0b
CieYslFX1jSXKlwZNDsmsjGS8GdpXjfM1Vuw8sR/RQ59b+4Z1BuCVZcE+VP8nj6gHRgRlIOYmToG
/HDFJeQ6ZYa2ZEk2u/W8gpThMd3PzjHSwAXU8GyD4Wkm73VSDbW/Uy4iuEiXU1aovnW6zQeEfH47
I4cRTpPOPfvClK10BZ5mk2/og5c7GNKUqUtBZeScO83biTe9A3rfzEZ6lyo/2yBwVc3Y83yVYbHR
VKoXl/VEz37UCZOCVfGFa3q5Mw/V3F+PPDZnvyy7A++lOZ9/fTBQW+IlOeDzXwUCzROk2uMcyzXr
YCntx6vmWHT728Rd+PmysMzbh1ST+kAS9gLUayHUOONGZIoNpcnCfaIqPHmAPcQ9sD1nKS+XOQPe
utAavH0jCYpBNzXhWrlfLZQkXiBtW0uXb753s2+pRZQfvewr2V2ABgC2MIpVHRupS3LjV7LCIGH2
5BOhX1t+BgWkXr4ysc/hP2czYtSv0jI9T0k4kRqK2xVKvqz9ZyqXtAb/TJecXO0v0mlMsOXnUGsK
yJfCUfwKaKIMltkEUYiT7T9+dRip+IvW0OM+Xkpn8PJV3mNcCDa0R2Bee9hDpjs5pbVq9RMCszDk
foT01pEOLgjUkbXh+dj+K3Cdlm4PETC/UyvQ8/j5f0O3YuiTA3kWEXtfZqFIHJDj0ayT3Vr+uv0g
wCAIqdw6IqxKBmpYzDsytSuU2BjoEeerl0BeY+T+P2zGsKcTc9BNBInmHfByj2V4UKZ7cn3uqFSb
AZVkyHsBD8c3VqvaGPH5znEw+g+ZANbOpBDSdzAru/UHJVzXs5bp+vigxTUwlrIegG3CC+9dhEJo
Cd/JlT5W7vggZdrR89mKOeq+oUFx8pOxMuSczBLzD/BTuNOozpuSiNwOpbSbNNTb/icYOrY+W4m9
UTLBmKmpV+AUTclEbxHvT+o+nbcFkKx3nexeiV8P4I5dvFVb+iQkvkSy4A+mU24lLoYbXYwpLXQ6
qhBL6CDTa65zgmNDb+TfDLlGHZ7s/1+bqawFg8cYYWH7wdpGiUCU2uRwdL6eGMaTI87rOmtQjK4j
r6ZGdsMY1mw2JAbBPyf0cMUhVevbm9eleJuPjdZkjgKbNGiy1FuX4pVKEh6SdMS4Wdt/Y7uR2RJI
YBYYuJYhcaAPW0B9mlowiVaZDn+LGwPy9XHPnfC47C5epbYmB1Oq4bZT6p9c3O+ZxeyKiUz9H629
m+LZsctB9SbWSiciveSg/4miPU4liONrrmc56h/lclieRkzInYUhhXLaCdzd70rFw8PQaIYR0x0X
+mhYqPakSBtV9y97AzILYrYS89ItGjG6YS8kUlZnHO4M2gR9E84btZ0FoYQ8xALQNABluI7lhLIO
V0P61ee9pDunTRilJIyEBbBAY1ktTQ3P3OwF2QMqywGs2ImM9LF3XTlSCKjK0imX1LkatXezW6OE
K94T/TPwSvL7lRsTraI1eHi2umltcEOOGDXPDEEhzIjR7ZFky/9fjtJVhlAuquu22h2FaobXAWuu
xwULqqJRqD6ryj2xAaCCXRASbl1YljstRnWKUtmL9pmfr3/hvo+RBdJB2rUFWaarJs7MGr+a4Bpg
YlaUA9Rl9+mFUkzekMGuTarQB5rZYVelvhLMoYbTz99fUb4pXAY7vOLRVMXyFaQBav8kAQaOGixh
LIMRUkBSNitSt6ynz0T+CaxdJ7SutcwbSFs8QMKraXyrtB2FNEFrX136gDIxf4wwLhCcS7fOG7jd
AnqQzKCQeU1y6Iok5S+VOWA7Od44Mtrmw9QumYFeG4SkMuPhs5xt365cNWEtVvFporCyaTNfef7F
lotZkqUSyM/f2xS0lg7neSPF1SeIO8zyaQIMAlR5MKXfVHSPSVof35S+O4MCY0ssSgstia6EFwfT
Jyxo87OYqgEAOYScyNatoeMYlUgTtvvk/X3eQGgBDF3+LG4weF64bB21tcDVcLfOGbHEb8tpqcpg
vlsdAv6+8mLbQIlLZDlP9+SFMIdxh7wWoiX76XQj/dWmkcmjcUJik2hcPA+7wuHZp3BgE/ypCfRw
DofY8XcZCIA70c8y62paWwoLpZ6gTaq/TzETDnHf53P/DgM7VBKU2OuTAkbcdq9aQSyjzm3FD+cl
CM8mKRXEfG16wAg9GCKlfgvy3uukot8xhGp1zcvE85hUBTwWlaeArO4zzdkTVo7tJgUq2OGy3o5t
uMgaruwog56kESy1KxZlKMWYHrEg9DxjopohTuj94Mg1eSY/cat4hwk0C2II+g38WZldSHurzgrK
5Z+Ngm7jeQzxs+1QU+bq//rInPGKgNlpb2mgE53wbRrDzkRbZ6gXQ1wypf+zymTwIk55R47YX6ZC
CHN7iE1EjAkP56teeBDBsz0vDVeRfaRUVZaTpsCou4Wt7iIMs76vM+5hM9vJVGPvcQtatPpp6GbM
J9O3pH42gN3avuVGpJG6prJ3guAL4W1QpELld/hCbOKLGI1Jfc1vwW9TV+atFEiv4ZPGwy63MOmn
IWH+B9NuTrWIbCNA2A9raFd8DPgNTRvEpNfbG6YtzWsFc7Mx+9ThrzPHvCoEQMI1IiElPomk/ei/
zkx0wLv5g/axHDjdqePve8gc6H0aW3EwWsOVs/lOeigeEzL+IeuPs3wkzlWBVd46qbeQgTENtCs8
4MGj7yrc5fb9uTyeCRrfmvYbL0HwVzTizFpvYpSfZE0GzuRt/DTNoUvShng5cUoxp84mkbHDzTtf
8EQUxIe3gzwsG9v1MKKhJK8XA2pNt0N4OFWOOR1XjdWp5HcUhFsnSxSoKVVgU20DrH7aqeyvqtv5
CbmSssJ9fCyWR75QeCHwy+XvZZTh9dzIYO/j9CqweqhHPro+Ok7VRgyIoliFuLSygmAbMpF+8NSV
gv16+gBiMfp7WVCzgRm71iJlUS0i0V1wRwyGpmnHsd8d+hMDnJOXApuiI1+XZbfwyroTLoyfG7M0
o9CFJQzoTB+0qb0EeAaxRS2n4vR+GmX09kM3gLDNHijkI2nVO8NY3cDSDwIi7KGk3wiFzMxsIIcq
1U9NZjdFKKLx09QMzwa+wSjsaQ+O+eNs6Jk64Yw90YMJXt5ZC22gBKzGAXRpwT+y2JKSofCx4zgp
E5rS3Kzk+ehT3DS0wVxRP59DY3wy/oQqM1642iJlFlOtgcU3n98FRT8QJKUMhA3vKBilFXuKXgOw
Tfevvc0n2XfHhXu+CO7zWlXTqXlAXOfAQkRo3JgUyS8tZwZZ7fPJpzsgDTwnq2clod/CaOaZtaAc
oz6vx9nd8GdhDkq/uJO/JdlspP//sXuZQyZBnIGhrf9oTJgDlrFxodkiTMCoBGIhxyvooblxeyy6
S+69jz/dX8RaIk9x2UcUOypbzgknYnpv9rYP9s/s80UMjIzpnSzQIJKjlfml+NOaENgbBRqbXUI3
hUtaSKKTZ/cij6ayxSXpX1L013IyEm0YtjE5YZqQSh1/9NEyZy6E+xLepFkUYD40rhTc7+GXlqZC
wlHgitM5yjWLM+DnwetkobnXz8dA2riMPChPyBKVb6M85sHYZg7+SfAyPNOSQANR4phcd/Ocqw9a
zoJzOVOrltT1zzkShHU+gSl/EW5lCpGFeOijerfK10NCiKg1Jn/ZQkp9kUNEYhJo08C3edz4eGmm
1UY8n8fHTgnHsv7hTvec0HfbPjW583FzffMxPzt5vJycrWxUBuIiEJHEeb/DpE7Nl1hRgdF5F4wh
a+FTTuFmsHYrs6FBNt0TM1PoimfZfdm+wXaDikiOc8zNZZmVhrp3bZyFCdoAQ7lIDcNohjmMl8wa
u+0pbu4rniJb5y1tsrnHSWKPcySlwCCY6WBXGEUciy7RTGJepSSNUbwW1yPpl/nhyBSryj7b7gun
76fi0B3qG12sbiubNlDnrSzD27dGpI8YJcPFb7YHHe42tQ8/OY5kHtv3XJK457mBxYlkhVL43jkJ
CQ1E+QDEa6jMuajw1RGhK/VrCloquy7NSInoJUllSKfS3J2tOpH9osnnOpdHtMBXsI1/RfYk2Dsx
w+9AiUwUsmilBj3JB3Tbuc9GIPEbMM82gM9UqQiXYHfHH+CUHrlA8+RT2J9yTvgQWYdv/5jok0ab
IZqypz7T0IpnoYcpX4uQZweqzKAaQEsaUwgEUUqlEn9FZGOkylq7SroVJo+50G2qKFSq34jX50UJ
IiHBGHYlr5scSXYFixlh6OsMMYsLL3e+bvM160w9iTqBLqrIJ3x20fZWLv7ejNCIPEHPtdQuYL0+
6lJkQHtJxfyUN47vufDpxCcXMI16ogyWHaYz9A+FZw6XTqwqfgEq8aja8sYsolY6JkJ/VVqPOda2
UXqCTY2bXjtrZo1E1bKAZqLsKOg26A/fFw7jlCUMrAkUtIlASkYbbS0jyjt6U3tcKjJg/Yz4pSdp
k6pWG8Lm8l466FDMldz9bD5AB5pNSSe1ITOGVjK2QnZafwbXxwfC1pokta2LSqIcxxus+Gh00zAH
YkeZPgSiOg6K7ETG1g4t7QHBkpGpWucCXF0PeaYAj58GcqcYa3t0dlcMajz66Q4gtQIk+/p7yRH/
CGmCQmCw9Psz2wbqkOAOSH6HRX7yqC4z5PDWlXX6Vke+HX2joArL0Y3c8XYgJY522r/wmAd81vgo
80fMjg57sGEo3gwIGR/1TTMLGUV5T+F1p/wrFEJoOogPKGBV9tFomeIm5vY7u3919OWublFehWrS
dFVoPv3uXtleGGLDTxEvA4NFg2M3Nc+3o56ngx+BpfFuHMgOHDDONGJBnrPtKcu2DPtdm7P2OsUG
P4keZzGXEhUpuEasyB3MXl0Taks1ynI2Z3u8i7ihHF80b/yMudKq0Ubp+nDP0SkVET9Q0sbxxoW7
a2PbsJcqu8YfBC4hCs8s2wJ2SZpzHQ+H87OxAVXBld6mKrgyCzX/i9g1OLkBcFtqZbkskOtuEszh
WQ2DE9E3vpJlvnr16Cac0egWH2GmSsYPrAiazd96lHctWMLkbHFgWOAt7Ws5i4i+nhBqK5AXMTsw
rvc1eqcTRw6XcZum1aT7MuTlrkKG17P/gySF2arnPAuoxTTQUduIspHrr/TcUK2+jFRN2azqt8Wq
QrMUoQAEtSCVYetEFNWUCoCZLbX8wBp0kiqTIQy5U/+QGzlSEW3Wio+2HUzK+uIw9xfmJSQcvNHe
GVZYpxfJlX1+IXPt0OkVw/sXdH3C+G2+i0yovdRxwSTGqMCbUKdD5OUgnm9FS7j37dvftU6v3ucF
4fbRFoD+++zfZ2gZZia9mJBFL9HV5RP3btovfcZ6QAj+hyeSvfUnu0lvNbF8QVOxOtAWmjNjPqal
pl00v3tXixJDvF+Epzk8OR+l1RjQGGrJaTJOepbLOMZZm1LEQY3T2CyDY11nC0+9nmwzXejVAKHB
YO1oszNukqsi9P8CMSSl2zhUx2IrHe/kQ0zo/QZKNVkO4rkxlggXxM3y3QGLw4/wywVJ0KBj61GX
Dwoio0VdeHSdiZ5KUAOyxPRxcC/vBS4XbV7sT4MnZO1Q13BLmUEYGJPzU+sR+b2IV5X9yaDu4+NB
/rtIONnSXx4gDIJCmxZim5Bx3fvRsAThrhIfBG1cnr9God4qjOEytrfQiibDmYG/NjncucyMbRmP
/VP95hUu73I6ghIMcLgkVlD/jchoezwX+kwPsKZopPayOUkMjQRRTQj+1gZ0beDpiFb/83D5q8jH
i+7FO2vJ1waf5neNw0G2kvIkmRZrDVnWs9zn8bKinfzyQl7ELWearTb/Fo4tJvsuDLJQ+r6S5R+7
eQXvpusaYEm3KTuYiXHxvuMDr467kmse9caXoIlKzoMcCaMoBseMNHmGyrA73fpgrMOEhJCqtSE8
mfyOxQIwGKwkJgXyxS/A05jJb/YNgJje85qH+bG9N/ct9n5v60XP6BOVH+93aUraPXh6efIx6l8o
oJJ9wzi7+/kDlaKNSZLIR8WOscHD1oZb6UToX5T2eqq2R5U+RxA59mUvMsxzpFIKERzWy/GZJpkB
J0fZg3P2GI6/r7gzcpqP9ZgjIYUS7rNx6Kk4MvWs+vA3S4WNYDXEFCH9LMEfZuxbyr+2NyBJY4xd
0iDarNl11+J7Fo/tc7azcem1rSf4KHo/5XFXEw2aqJ3DkTP9PROWYvqoCK4Mib1vkDK5n6SNGBim
mzErTLEgQ+1uCm8HDD1V6OOVI0wskIxkt9gTU9jmFICHymY8E0ZDyr4tHk1TPwImkNlW7Qe/Kv+V
D5qr+hf/n6zCFm4AdpZWeYf8C4KYslucd/PVfmq2im6ol94OJtdGipM7X5kTlXSFKPbfeM5Mbgei
SZRDkpKfEyVRY8gGHG+hWmGSLmDJNCkBtvj8WmYVKYuhfBB85h2t0kXkakjUceZ09fSRDtJpPBBc
FfJT6ypMsPubpZydlwVAaVOM9/2hW5FUYjPJ5EnKLNH6ViQwSUtvQNbgkjrDTEsyB4XPFIK62CCr
sexSAFCvM2xp0e2MN8hbylqrtOP5SvYGHrJnVw2QXsH6jHMf+/YEHva3koBiTOVRQsmu9kF5eIa+
j5RuXrXGd1zSoq4BL2hYw1wesBuw7FeXjEo3rJoOsEHWDIF70U6TN0XkbU18gH5n3xqTuhVXRQxA
qSppmJ5rVl90llW7DeEw2LxDTeudsal2w00aVp/2MT7FlK2OWw7nSzT/X6dUHBUrEolmUE8VMWaR
FUcdE8iMbj3h19zWdtvmMl7JyQkH5bdYnVqebQblSt1qvylySNBiR5XFHsavcwIixW+X8UmEOkGs
fCz4ZoKE8rfRBNv6cc2UqtC/RJfzubF5QTWqwhrFhVUjW0EpVOX13kz79zrhqKyXpe3R1enG3l98
MM6RtAhAqexDxij7+TkG9+5FfnBshDgf5zFxJQhOPjrIhXVNBWbChUib+utKGA068ztwoRr20VC7
WyQzye/5TQ52oUYM7BrKbSMcs4aMJM0IGBxCVttRnHDpLhMa0uaDlLd/sDDbk4i7m801oa7Qa3OR
v7AM9V20ckMAOC7Tas/GrGlGuyu9Bm91AyoQIX7xcSJ+MvGh3rzVd8x2t3QvUe2et30bvF2gUKh5
vCp5lflRCgpEEbCo1o3asOG1F7IRxSTRSAYPcWAznvmoWb1v976Wc3n6zGqP3E51VqPkqfrsZzsS
BmnZ7otquU91z99mo/0Ejk+X3HzSdsr892q2jLVoQxpQUGVJLUgoiuO/TndhoQUE2hxekidhicZQ
McF3XZXIFYO4yAgxzdYYsI9tfzbrft6jdcMpiN1elPRZarLX4kseDHk9NoMRTUhKOVobx9rn7FdI
kdWkG3pTm2j/EajY0vROWviiajGwO7DbszYp8or1et+8lF1cuLNFaResehxDGInihI5yQnKxtsof
8HEGk/BWc0E9wVKus1iGlhORqsQpUiViOi8OLm2Zn9HRgY9vQfNzmzMbJOULbQUTnsS+reBawyh/
1o/QyDRn4QQCd2+CCaWcdnznqz4i5OgBDD9uFtaMH3irLcDxh6ysakS1GPKTmMpTuxBnheSAD7ZN
5v+I1949BT7F7aeLjSU3QhPdxjwA7D1XMgttM6WC1ZToMe70zcXVWLlSQ2AONsdjDuy/pKOy6qK1
RjbjXl/aCAQxPTaIF7mm3u0BjxNqOht9jOvzYtcKAn1/Q5EzJgiDx6a6Bj4Lw2SNJOFZIX+WnNOk
FtP1i7Qb+/ued2bcbFjOPwo2nZW0BQuni9M6Sc9seS+v8oqWMW8BYJke+FDQkcrXDCFbHzLYmODN
igKTTR8q0czM4MiOkXMme9u7yvKVq2Ard5nbqGoMu95SfITqBpfSx9RSBFO3RrGAsCgrP4/Qv7SD
GCoMpDrhhVJfUq1B+7J6/vg6Jt4Ap7qqz2DtfnupMELdUoC/fz/PSA8XzRNLMtgcA/5Yjwekw+/3
3Yss/IO/BKekEGtPU8/OuCqvehqQf3NbuPnk1iNJMj06Tu7Ig9FZYIDmXnab9bjbzS1QqKYJiZku
Ea8rni46HOb6jbzf+XW4/eBAQQ5WDYFsX91zzDOkmZAY9U2iLbNkaDenEG/sriTRQAaFxDutSuYr
21ICLuVorm/2mvs9LcQggiqnHmG+0th9H8TmRlwMs8J3bImNtqSSWiNdXXDwIHjCgaN+99pFnwhE
PE/oJ14/7exsIZFjR14UuouaLaEvVZ1pGHLpIUHm1E7Bl3tKZe/G862Ps1X+n0DKHKMWgD2H4Oug
CBSNtZ/2JrxFCh0DbJzNS0I/fyVflPXUXw6iCoA0wVdN1qDedjiT5p48Dy2BJSPIA7wH9LeT73gw
AQE69Q2w5lGjF27iS0+surm1LWmgFbI95hlz/ubRemQES9Ze5rpkn+7BEO+b+uROqnTFZDir2yA7
a+PZ0wGpvI+MhxkDLHPTNJTxqULg0r1IZ7/j6y8duQdlfu+q3Ed4Frv0nPTiRaw4kC7vFa3Im/Rn
4fh4xZ6DUNmYrnqfxedIdIy4uFRagUo1kgDvfhWWsgRN9KtqeaChhPI/zxrfpdRGAoB+pqT9EF6m
ZzL+GZIv08jSy+89Vysce1kv5IxJim1Iwh7+AIo247umlEtlfZ+KKuXlr8T0g6YbMQxDbdRPWxhu
qxvfpP0kZtjfLsZH6w8VvFRRe7SxeZkzJFIXqHWXcx9aT4C9je+gQI0qXC2WmrQr5ZGNH4rZdty1
jynbDsWoCZeJMqty0c7FHW09NN/MykgwHo7xD9BCM/LJ+FaCP/XzFVbOBriq+tbn9MyCkgm0w8Jy
Ef9biPG4dO+7FZ3aq4uCaIZA7PRwI37uZU7xv7T8JmTT5ENK2E4KAEYNHhBCJjdHjLCUTmVxs0el
72vbtqJio/beLB+xTwk+bFWgGAJCRBvldiehIP+pCvqzKb9pI5THdrFBDc9dZ1zkYts9Gi+w7oVM
OZ9p4ygPGEIVANQkgm27Fs2mulJ20JPKhOP/VQLtnViRrRzJ8lXFY1/o/Lhu3FgtnRtY13r7fxbP
h1K3SApXwahRp2Tx+H7/rW7WL6QKZg35wM5/uMUlbkyWhsXGIkUlF00eCNUI01cm/1hHeUue/LRZ
1XYfesx7UmLnre2acDdDW63ZXzx0Ay+SwozVqVMeowl0ccrMiRhWNlO7D/dhW02kXccJ2/lE6LEU
iWA2kRDgNJ78TSvjtR+/DmxvUl8+zdJYw0RJclVSuxrgnIsAEjnijn6uKFnNitnCykAQC4/NEUL/
OeAhwJZjy3H1eVBTMyJDvAHwTuyyT3YNMwgYWITkgSNgYRUOa53zuKdl9mJuyIE7efApB1aJ9N+4
XN1gvZzy0LZLeBvDA7duXYwenKgBeMKjFl0PdTVKIPj6E8F/bAGie4j0P78jT9vOW6t3vafhnvbn
sUNfm6yAOm0GTYlffUCneFMDaahBrXOcMsI+Fms+YPZeaSeaDh1/175JTHotCE+4Y8zfsLwpWEU1
AeCbjidJLJBQuTASsYRTwfJppKbY3kPfuIBntzS1MOU3RgJ0LV7P1ZPNk1tDy2d2fgJD1rqPySyI
T9iSJfbzYsCPhzTErUAGXaip73sCAEDKXcmFTKrPROWf1uuoWJF268dy4gp++gUZgTCrKFYnt1SS
KP3nsJ+BB8TDH2VTl+AvfIFSQgbWZqMANBiEvvIAqJjf7slG4tCNsKXuifRil6rGTmYWAjKuzOeG
cWfjGu7JoDQOBqhC8/GjhmTJKHZrjwkdQJ7NtUrWEGdzEMOwAo3dKUaHlbOYjwfMBHpXwCeJNln1
RZH66qyXDjgzciid0ijjXssXKGNWq4sRgwb6gUP7ZWxJS/qhgzl8Y11+e8w0TmILMeKZQu2DzpxP
etKGSqm31xPQU4LQ8e9bgUOZwtKimYbM1bBODtr3ehBMjlLIbCx1+zgMXbnUhqvqOvPbvL2YdJBa
hdt7zkSrNhG8nrk3t4ugbIXN2DJ83iz6za15/W2MVyOEUIGBKJBLZNlW+DtpVdwnnMzyf1zN5I1W
UDT1D2z9T0k/bUHl/01JlNv12xKznPlU4a9zjwIlGw6ruUr6nPIsyhmU/8H2Uf7fI6BSY8EmiO4U
sqsfjMGpnnMwC2bmTier0yyK7pr3XvU0mIMHm3sstRrFSKVKsz5nVtxts1PPI9xldnu+xhbHH+0H
JVGNtKJqRH+HIo1oScxe8g92y1xelNjK6BUJNajbRPyeS7jPMEXuhR0TgqdJYseJNE9C1woy8Mfh
4rrimlcbeLmMOnBJe/u/mBTXjksA9iLJur/8sn09mX4dSxN6W6oL4REJTnGrfvrJtf53KVsFVQ45
rogQIbaUaBz8cv35Q30MDMfU1Z1qOU3LL/4sGQUYpPkkKxuvDS9f4XIrzQTdsRPQY933NqTqiVr9
GVgDNGfOu3BFbvVHhavUdVfKeIwtvJ/1LSNMK9YBff1hYtA78OncU2OBVW1lQgwo85CBPrzMivNi
/Gde06CKtTlJblWgD+t4RRwy8d09bQd2+s9PJbcJylWO6maDAVThtSbMH+VKwdgzCsJvDd01HC3N
0Ez7okGWSYzEiCTiR2JFj1FwVb5eJ8KFvPoVEJAaXaxfUUkiT4aSkNiAwE8IsLcfYxNAt7qm/0Et
778/Zp7V0GOu+FN0DuKlDkFAJCDC9t8BBGdAbYxVBvtjdxSs/eYucQMm2ALyRIJfwqmajYAwFifC
SANix1iWtKf6KfiLeR/T38FoFVs54Sd2YzAjPQmamm3/JhQran3ULCLUv0iyGCEJ8MW+Mniqba6b
FsQxc60pFWU5RxpPDrkk47AlfUsath4NQuf/JHUJXouaLfNN9HFGDux9nYTJcvs73d2Ve6nd0jgw
C7+n0Gv1Y1ChQ+5zYRKCEymMV9b5erNi9EtUCX5BJjNkAZAcROYlnRkEWz3LrTLKr5mB9XT2AB1d
QhxvC9tT6glBEPfUDx31MISwovKFVVmdODT2AB7K7Eoli/qcMVpHW/1Jg8x0kjEwF/OuxcE0UQIE
gYEtaJUUNOImi8SfAHnExaoYkvCYtZRrr7p9yD2N1YjQm3xczvQj5LjxE/qGeK7+34upJBuPNi6E
X5asPo6QVCU3keLsLE9zMx505sznXSnl370oE9/hgQpB4rQb0l8nJjR2z/s8KlmFMj3Wwg85kRP+
10XSu2MTLQZjqHmaCiHL9XwFbD6SsELKHJZ0sUTNuntAw0V2JXbtOWcAKhMf6AVXKtpXOI/HiYMx
8p4COQFvj/f7RoMoeiPs1F5v9KRSGaVl5f3Hncbk6ukfF50vjEOjoBOasgW1h+SKe+V9Xg+Pok9Q
Fq+0RYcocBDPk6+EjYdo4HHOBmw43rWXrC8/8z8VESeFOgwwSO2vgrQ+mZA8nqimOyxYcNKEjWuO
ApTGF8z6V67RRcGBzqomxhH8CzNq83Yt0r81uy0cHpB9PqhMMhwEX2aHu4OEiuP5FgKt95UdtNhr
dObQYKaiNk28/7cz+7X7xJz/ux2lEE4oLvXLjNl9YSnXfD0IFRKitF/D7eeJ7c+7JzuxOuOYOqrk
tEX5I5rArj/FO9qS/Oo9Ukb79tkhRxOfNs2J2+VxHp3ixBmzoXiSmvi9B6+xZkMU4+9vnjvU5LAv
a7Ipnm4CUd57JA+6l1wMoirxx7f4UFPXgMMCDCBEJl+fRJ49Py03JAEP4AeloMZdPEv9MwnYffdA
FhD9GscIo9vDRRXP+ogYsGHrr4lB2r4T70Zcg1DcEI8e9/t5YNeNwkg4i8khq/Phdhy6QiAQFfMZ
OzNmXFCDKs/20x00+nGgzY+0XYPEUFWeySA1MX18UL4IO8Gtct4Z26ZsZRadFsefKNU99UjRCoEV
mf/P315ftD6pkJGHVMC+0V1RoESUCkmvukrqNHcaw/rlQnHxSfNl7pOP+gWvImouykTpwszHMtbr
JYOiBffPtnt5BgT4k27czuijsz8NuoTtzSYvKBBgg78IreeeYbTTM8tFnsoRaCVj/xfQayFy9rjM
uP58GlNXrI78lxX0pipPM1Fq/xDH0NsrOIBUIvWFklXzYI5wg7eO/dj2u6SObS/71KZVrXy/l4JG
WaNVn7JMJoGEydfdyL4gjiX2C1S2gLHHFj4gLtzdfThb4T1aJ+AOO+6tSzKPYRJy/2n/3Nnz0Cbs
qcqe6MieIxi8Dy84BLY5XhC9HvRCBZ6Oiow661Ed7dcVwFG0yali+qT6TNvhDUczYSA9bNdHQ9Q2
myVR2zU+eQc/fuAneC8zLy19MoWX8o1+ktYocvxujfuu9HrLSS9SblE3xMR9qGpL1PCZgvLivr9j
dpY0SriAudPOQyInqzrdEcYPY59aGIVjYxerc1Lk4t8HDqK3aHwIaKx5nRUKedzo6SLC7r0L5goO
HXz3Dz55YeQaDKu3KWHGWgMvwNYgQkSfvZKJ5epB8p/0ij/GmbCq0/7CFbVA0w9hiLDcMbQATTmX
kzM50eAvZ9nHNZEqGaSfEm0Zk77SA4SyEFqN96Njlvlvk7Id42VKe0OUD+rOcIJT1/Nh4LPQAqhV
fWmdyKO/wdojKkOg+LIeUv3BhFPpokGUjR9qwSwPr7kqCdiZlpvlI94dBHZn+QKzwpsV54+5EpYP
Z9+p8p7YCJD1Oxo3OL34OuxxhHWjBPfrA2dv0vTiYGexWuGFHX7ekTh31cTGMNvzY4IuTqh1Y0nZ
xfELArwuNWSbsTCOA8zJhmGNUc+wVtlz59oXAGQfwCoUoikYNMYdEpRnteKf7pZqh7wNUVXZdO+q
htrErxrGUukpah+IoEXL1TSQBueIg/6SO2sxu2dz/le3Doh8FtojKgJdXBtT7F8HGykYngY/W9Ss
qLI7SjhdBs5cF9aXgAu7yv99+zy9pVs5WVzFQiozrQMvuxrjNPNawYulGZthFelsub/2EWDVK1O/
e7nISAQ2EZCFnrMTOnUF5qRgIpuxxUGrtdcjDwQyoFvcgLmFIMGPfUERtYNjRkfNkpAkqgIRl0x+
6Dc6i60+QowfPF25dMN39CEXV+ALRQtymMq8/caV4nhSc39ZkVWkHAPtDsma3BW+gVJ+3xD19kie
qrT1Bdi7Tw3LlsyGpROqgHP4+QCtZuEz8kdE65fb7T7yaYhW5FQbGkW+G3E6kDSp1rHNoLlyu0sd
H3L76cKqYw4//mwFaltxNA1xaYBO7CSyrxxEXSX3PVsKik51mB8MaeUOuUvjcjGghjA5R0DxBWaO
if0eQIjc9SwaQHEk1NOOWejcBhmO90XkHR9aWx8O3FW5nbXwrz9fZIxzWKf8rQNAoPjTy7dYKYMl
118xrLSSdsIZ7cIsonGQyy3o44qanlpFSePPNEEDYhSG1LFea4q+sshrWdWhJmUV20iyNXp/qbnH
NPWDcjU4Q/GH6HG7wZSsZqodX5jJoe+ux1Xu7DTTIkAESKZyGIGCAISwFr3AckQD0DUBvESnX2Zj
gQMOEtaSCyylT+pka+La26z8i6+Ejq1xqWuZZMAKX2UIDDmYv7GOdCtVPj6tIuRAySqD7iNBy8KE
Fs7k+xsxbugbeqbSq2heNgJEt9UR63rqiZJiK95sMCUxVm3X1U3XVgdRxvY4yDbTKcweqJQys5qi
CF0tT3Ug0MgIBSRd3+FquM3FiHBQr9r7hyczRZJMVxTstvtjDNrwLQvzg/ZObfmG6VUKz6gsq5me
+B/E0ip/I03F4Kdfq8WMnsXlfdnptM14lVOJPcn7yx2QZ8rgw7aWSjzRJzQBUsYZLWtjSC51XsyC
tC1kHE/iWHwCh1o3O6t5SZX/0Cgd/ntWsqd/s0Yfo2q/30T69A98Na9wFLcNmVvsxMkjeMsLKSCp
IxKa0S5Db2GYo+ciKPVWZa5CaH0sGch2YA/FPDN+OTV0kmX0cIqVMQGhr2vT57Jg5hN6lmbnEcTH
mKgMwnsqvJfk2DPg4GOV9U40ReTKoPNYPgPk5uQrVfteec4HV4bLyL16R0nOPBcTeMyRdjaayVlO
UQZHJfGb9MQtB1hDXDZEPFsAgwq5RhC8sWpvFOl0dmzzjww6CFlIon2RS9BqwlNVLmjjraE0LMtf
Ng3e2MLZQppvkTtuMfLx1zJXmKqdMyC2/IZnpO52ArwyJJpUcZGHmXwCv/vmD3TOKgSdoRsYQGT/
46iDabXPYzad8kksPbVuc2GIx8k8hg9RUVMr3PJ/TKJWG0AQLGuLj47AjE6E3ljDg7LbAu1qNctL
GvyiC0Ms0VHTLjHl3F3cIGFXvUIZvLfYRmVZl7iITj31yds6BD0gqIuvEiCi5yb5uzsmXfEpBpJu
7nwbMIuzkAdhZ8BGL4kx1qAAfr8MxjH6lVonPbnbKbhN5qjl3o1Mpk5kuoTSAKc7t7FFtJDLjySA
NYs6qQco1MAWc0ISrtPTFjdFlRq6fIE0KH4k/zC90bwbWecrw4BNnrk496aiwQFTvAeV1l2jP0Dd
TEDGhUkmPiH7T9QL6HialgvZ7gTjMO7GrGBnvq4rDNjTX/5bKiymy/cLHPZb7pdAvTkvIKN6Yxeq
GTYg5SQuTzlNFShXCZOi3GQp+1LMdNglOZHi8dkTMwLXc+xJ+LXKJuD4T0xasOo2uggjBXE+gQq5
Y5yB0AyD72FzFin5WUXZ8Dcr5VQaUhhIEEMnkVrM7yKK4cxWdZ27eafDNGG1RLhct5lxA9bAVW9X
i0pLoq1wtkozrNNk1jqQbWoYzVhX4udsbKHamBgtojPLZtPPVwSu4+cxN0QA2JwJOuia6csoKjcg
8otmRamKcOsF70O+Di7I5VsHI9ArJlelFdJ5piz4nOudm9hYFKUdyQldis0W6bmKZ2PeZFKTvtWt
57SNUApEh4uIjZDzr2BmwLavjKkz2bOLEv8aIIUTZF0B9Cf9z2S5otWfyCoxBgjmfjqohmsMIjcj
C/hKy2+Kvd0uJO2XZh/OSZ42nS4w6jQPnAFvrA3qm6CEzKmXgOgwI4OAgd+mS4DbEubElBDFq2mx
sLh1UcvSrY9642zxkq2N7MSZYTCAHKjuUHIcg5dK5LYm6PQAQUzdzlOn1GiH//gT2URVuiKq7v6i
zrAfdShMBUtlD5zks7rwGrhyyM9oDP0v5F/1D7BOwz8f0LTW0AL40DESaIJyZ6f+pgUYbyZvoZ4a
FuzKjonRzfI26eVpNyXczRZ1KXyR6k5AXhl5n/ssgawCETWWmu20uF2wXan6Irb1BxDbmv28YQ6B
z64G73Sa+iykyjLYWBRNsYgWIY2S2EYoElbuHEVPV5uxtV2qOvdWUxES9P0LKHC2i91sogHlD073
JYT5i8yS25b4kGNLcKSmQ9NhNYsNS/PhoHy2O5MRwy3Gll2s0fDD2NqPUb5GJHbTJ1jQH2c4WXxF
9230xa+shnzNo4f68GVWIWD3KRGFNHIWwmT6JXjhG6Z+crWElZRhsXK3YiVBJMDN76pMInAvZyVp
WINmj6DtbquPwdI1E03mkP2bUOoDmhenPR/cXpi2aVuNQQz2irt/QWCaQbcBaILYQnXfy/eSTJjo
bKqRVmsfD2F0qO7lTf3sMVTXKu37pSMGsCDcuNAuCdscqziuuGO1GdOtH6buFurISjBmp5qFJo5t
rdm1ZrwUE9fGyWushpovotfgLF5yhyf9b4+ESfMfrmQ4iPVZixjSSNxAKwFCcaQfvUHGXQPjMKSN
3dA47KiDnZ53rllzbVeStg3KOMn5Fg0gO/2u2ebvAKzcEamEqiqtCgUgfmCZpBuWQ56L2zHpVxiN
DUWEs+1yJ8dwzTviGO4qIiTCZaC2kCyhcH/0K4Y2yKp6U1JxMGvXNqc22iJ2oKLQxE6DKLKE7/0P
fUql5tdYjID7TLMFMmwGyDoqjHvlta279Yof2kAZTYrWQuch60OvD28QcNcR2vKCgdWWV6jcvFg5
vDK4vU8+CvRQuG51LBoiMG/GP8vtcsPJbHSQAPEI2fWyXCWNgk+Xafl6qOLlt/4WDLLhwxS6gOlt
DjUs4BzL1EjKCZ1jBPHSp7XYh+ZG5YRdKoMF9BjfX3n8f7gl8BizqG7Lbac+MtpQ3zPuvRCqMClz
T/ix6r5cjmyNI64EDfdchEy9xkEP1z5pJtEWH9qYiuS7N43bAyKujJ3UUPogwwVQB6YeQG10xA9y
zJrt1DJ377gCHlItChq71y/lsYmVAp4ytOS1Bd6WGhmWXmVjedmNh1eZVEYJIHiX6L5Es40nx0/L
HXjmlDsxRVIEjeKRltEXm5G9qlp0clXATnA6AJ7sVi5gspw0w80CGzngD7txIeTYJulRHPHWB3C1
rydbCEDzosDiZY6OwQ5bFMgSv3Xk0VX34SioHHfZKPdZvjrasxv+i/vRqd/uLPeddtc5TsjhOh7B
RMQa4+FNp3s+6vedeufHhncJ6aKVIS9yMTSzYrufgCHq9z7hzPFphCzi4XUAiw8jZJa4FQBNcI/i
dXCd38yhqwngBLbNCqqg9lfkNGmsBbi+3KJgWIpQWxI+rusNq0YBvYJmwyQ6wrxzpr4q1l2hTXmh
w7UfEyV+SDYIwV1DDJCqTwbBP1Tpaqg/JnIZ9adRHyzeQZa5hODWjManC+09JvW3Cl3Y0WTosT7v
n7FJTTeciD6YaADB7GLpJFYsaoolNNeLgQ1+pqMCp7/ulEonshORd/M4CPH8bT42tXsctFTW+Yfs
ek6F6BslNvznFO0Vquypjitz6r+zTN9sWDXJmwxTKc8Pq4DH+bkJqvJE1nE8PO0bw3p1jqjAQGkg
SdzNPp7cviqaH9TVWZ/mNhPyt/262LAszFb5Q+LS1TPI4MxpKDFLtLpKg3RKwMngsFUtfNTJr9co
O4zGHBJ3byczemaV26tmMRKR8GsTW3RDt/FB5Jp415mbkU7TjCzEtHZ0PvZhk173YMTOI2MjTkSj
DhVYUUeck4eBpRsII8qu3vhBBs/0cbQfDJm2W65sSgImjXzky2ys6hYbqyskVh+YevCbjkwvYlQE
Y4geS1dcXucC1g9eh6GzcXKv7y2wVBhrI2YYYlPRWqOFYJyIQdxsxZ54yzs+wazf2Bhq4WvX76LS
RTUkTLcJAk+EuVI3Rb0KhjZPdDWuMFXKhXb/bzqhsRLo9WHkP39gaSfdkt+ZC5uBFuDJC6FSBXFm
hJtEUpVaUfCJwt9quG3bmhXkwAKQNy9u6G11nUXZPdHRdb6wHKXFO4k9lPi7nAGr8jkwtCaSX0DJ
kUv64tSxhz1hl5RsQxXCHzrCPLKzBL5iUV+6Ntl/HXsMunkBiWMtHeTU4sOygRvK6U3MI39RrqXV
7MTyLvdr4qa4R3HvexbkF9Pi18O3PtfdsCCRtfARKW9Ep0Xui7fGyxr9rSq2H9d/ENFPZtIco0cK
Sod7cFi8MNtNYXY/Wv+NUDjYIRQCjTogm2XIs6uUdN7fS0TTrrqkGadXXvPEsFY7ZaypKoj+xWrB
UsaDTeC7PNkVyi7ZH77XX+7bnLegMYJkwhgpmHx0bKrVzbS7SLAf7T9GKixWfN382RO/5hg/5cbE
4hml7AJdEt001YRCxnwxqXKSi2hGxlNH059x9yTWqpLu57abZSAxuwSZRHMz6VCKz6px56yvjVfm
v4Qi6pkarxRLwDzr3HSGpRuFZ1E1rFt3LK4ax7DPelu7IAwpOJUfEMSC97YNKi9vdbm+LK5TIlgG
oJeTahF/P2/osm7IyCRuDkfiF5dwN9UsvhiyyZoEgHepku6VYmfnV9ODUXeSAY0IccV+FnBegLZi
h9S1fqVc2aN+CLC/8OLKETs8NH5n0ThqvvPa4dfubTXPSdyiAHgc94U83nbvN3nMdthXW6Tglc38
kw6GlZgKhkOqXE9cmtBqgqTzjmswLF2oMwqcUx4IuwJiyg+JgbcNZjXOr/bQ2b4IMXzm+n8q091Q
DpXQJLSpQuR6XC/6InOymKtBo64xxljkCLafA+Oui/bGsAsjFTy7ns4E6A/Zdijol7TnNlJHLAbj
v7IrWZ6Xo2kDVttyh1NsqsI2s+sn0PoSX2d8wbPNVtTZRD71yF3s59Rgn1MV6z3Y8ckhrnhZfOAQ
MVR1yxFuipcNyy6NVWvV/qIignnEnznsUvp4CgqPwBJul8W1CqTFLnTnRCw/AGF8LqIIhAhZRLY5
du2NZSXebtLz9GHzVn3IUtNYHdMm2tehA258db6ZI6gnlNUxJiIAPIr6s60yFQrM8KcHsHEy1Iov
3c7DHsNNT+xBBqhDJqMzyH6kWe5V25B9hmdd0VDRNwVg0aGyCL6AMtnNX8ik3YJA8RZc3P7ONOo1
PZZEfpp0w0bzzMDbIp2iA/Pg2GhxJ5Z1YoSdyfjWvsQ/RhBr7/KZVko5OZ6BBVWwJwy+rPHl7i6U
MdgdA6BbL1b16wPvNkQnSjPGpitgY9lgKltPWat4kj72D4WPYCVOoLudMjtgaCeyOYkkyFC3M1lf
ymdlkCcvp+FbiD52Q3rVRCnrWwdHa17wqDS2t0dO+VZKGA5YtteVfTMrJfXCHJNbeprfmezcwgAC
GWTjqo33ev0TR86EwkaK/k6aP71Tk0WwpVRc50ufHPt9ZW2DlVLctruAkHC6Eoq8tILvfXiv0Ngr
a3WtL9YZJI+LTDOSJviVA2RLehdzaZuK7GreAM9PH5X33eEdIZc2ajJavLqgzCU/fTuLijn/WlOp
2vxSXa82WTNdWtBLRO1+LbXL9x76UEqFE0kVI0qa7+b9h/hRsuBbqTTAX9Zc3HW+IS+38su5oHWp
sBOBLZBue0fmmbIR/x5C6f33pyfKrflEGVpLydZyeL32LaQG5yFuZIjOuIEH/b1aoMfCYKkYQVlJ
68/wbivhJIgdTQZDfUCw+Ow44q17qiPF8PjOUEMhlWd8s081joUUmNP1Ty3xtF1UkuPrffydH9Sn
qEAgJeBAsm4wy3PPNf4H1FxdpszDjrk+S2Vf/qCVZpcTFVWEDC4oNCHk6rti0jTPqAdsfWqizikj
Zpuvkqa/u/Kfvhdy32oYryv0iA1wbtDtOAnh6l0s+aLW4qhYgbA7O2vbxsf1RLL++UWp8ZTdyLYN
jqJN9wqo+6USFWSkSD27NuPkdVYq8HV+1BFmOW4xpa9m26+eggvttGN8YFgz/VRFsBx5+ntZ7qeQ
xuCS1xWWjxDmnt5vLRYtbIF4rZUEtvzU9ohHE0lXpKdmsVkIgU+qKoduzCW/w2rtYcttfOuX8xA2
VgkyKgH1uIhXe3EmyeXgwZAbRgOYYZ4K68T69goJgzFLelNsyKBoapEn3PLqhtKpmxZ/M7y2FqQG
iIxsv0YYzDuM448NRm2Hei2GmG/1hAdFbUKhsrYRFXajIV19lj4HZkMU60IDz5N1KeqN9kRMnpJR
JvEDT+tvmGESubakc9O+zB24Y2nBGcEE3vYh+BY/qV3U4lc0H41PoELbtRuQiYRbKzjSBxM82+z5
Gq+upKiTH5mI8yffVAhtS5Vs4O10862abPrTJ5ZQOPYwOXcWbzmv2+H6JmkhaYLi3fO6KPvXhQt3
B+mEXm/uVN5xJR2j9/3VHsF63a80//TwPBlfNtOkMTJVda8yPaX5OY3oeIr3HC1+es/QkfcTDeCQ
wz4P3KMpRbyA7z0+Oi7dUPgEmb+TeaNzJSQdqBKQv4U6xm/4SNQH8gtRkp2FemNT6qoqINdtRot8
neZMOgCH3LWR7U1CvFpgMGIj89JeBNSUqUYyfcp2PCacPtTFR4xaftsQyZ9HBiALBh8jIRbK2OmT
hoW1DK8reEnJtVAVGCLiVih12ImBCZyXp3dknI+u7SroyNJjoURp4yOoa+nEEscxCNhqYEePHBHQ
vjVVyDRSbtjQ/vS62Az2gNQTkhlAFg8mymYeT1/0HhZ5+N781U7+40oXYH1ZUJX/FssDZvqQkhLw
UPpBQNWU4H5r0gi/Dhf2JZpOXHoyC1XW8w+XN0j8Vqrt9AcObggwkXdZBqbsdMPyua4CruDVpMdn
CFgFxmNb1leYEW2HDx8xDN/XConYg5mqibKlUisNaxlu1oHSeqNkAjTfR9MTBgyG5I39vJHBCaEZ
vp1mVyqrlkiex3ku0TXktGRGPz9CUFVoLBfqkYGiWYKy6DzKxVLmXdAXy6R3buU2/xWdx10Cxc1O
Dm2RG0gJKRsKeBYGpOLGE7aKE+0ug8F7QjCKTLJL83iWwqQuYi7O0s2ukHOcXQnHbnd94sh0YcL1
ee2fwxc/vR2oLsfUxP4Y62ujtKewRLqukSpqUwZ4EcDN332lp3IB0lfJBQkz4D1hYe34pTzKo/sd
oI28n+pNB1RybOZi50nK8OplzF824nbtHaF+Kk8cHj5SiZDreVA3s7p7lMLQQrSxpUB5Yafeo4Eh
Y4Ycos7rgvrbXJKBZg1dGa9LSX4nYWuYJ0ZJVgHmpXPdL93873AZ0AMJfJy+fN4OvxYxO38TF2Ih
ZiN6sMb57pwIg4FlDhnOlrK27Jg8rRdj7Ce9Y9dcHyuIqy9dvMeUBwHxRD3iDJmWW1s9UbKTd+8q
dzrrJBG21QhCOpoA1XGr1peBix9XS8hnU8IHOX8z/i9mptqqoQLpAqQgJbczqnPc9Mhg0a5eX0QO
muZqLE0oLbIYqZ6pgWi0SOQXjjb3/paiPCEcvDbJXtuh0TG/MTEXMColCnj5zi8JDoWPagRstXmj
NGHjNqUlTworptCUxxGNX2TOx85sBiZgdy0UIE6M6WoAgou9M77vnWK9zltOIJovtAvnWtaWYv5W
dgMUqYQ9JtCLAoRkPyaDG5Szyfd1l1frLPb582yaoQDImLmaAyFkD84vxh8cgxD20wQsruqJcgmJ
sNkC8yJAx2ElUTtIiiDC0vo1o8CPDS7xVwx6T+Qdx2NRohPIZSBA92KGkyl1LQxzKjG+4sB+eVjF
mG7GzS18FD7qMCDPEer9Dt6Lp92Ujp2G1Mi7dEAjroopARhbgmRQr1kfwlr3KhIpllvOEv1p3SVL
N/XV6B2Lp0HFH6nbXmQ9pRQPGEzez+aQ3xPIv09G2AsBGAOaRgDzi/XMLkL7KPNPxBC4PwryBP5f
jvimIjmCtrPxosiXaADgPt4LDiLICufTX44v9b38ns6+6+9T2ByerKu0t2YOK+TVJXnnmVw41Jc1
wnwJ57gvOjjBxGXGyR2s7nDQ7YO0Hxh51HecIB6/pGI1cEBBRAiPGJ4CTDveMXiRWS04V7UmLh05
6BJ3ewzoq95ehvuOTaW5Dh1FrSVGMEwD+3tukwfQQ+iojSLYygFP7qzTdaRNHN/g9vDxpwYhnuKp
afsY+l0bBM2dlmvlgFkF4y9WvJ0aOTi8iXoSFxOFuHYMR0qi+suubZuGmQMaRjeQAdW1OwI3iE6c
SUXIrLIdZWGAu3HjIY17wmhOurn89ZW2aehMEayep7tSOTJrWns5xT7z8Bs0EiOf21pTSCZlB8K2
Ywue/ytslqo+25mz2llHh21c7BFSpTzlZu79w0vGY4nNiMmv5jmZDe4G/IBhSietYTa9mruEfkyW
MMc7J15nA1uXdNdR47ksa33yWn07pqJ3Uaa/r9pJXvI9V5QUQ4siZBexdkPh2kHH/KOsnwLpw54v
1xdTnyuYq0k1MOjwaO27pnvAYMEC7nupN79P3OQPLED7DRpZXkiDgWwNPzDYvSY7fhh55XAq4Lg0
rOJYWZ7DeFGm74VBRqOjAhynd1cDz3krppCltVWglOZA3bqD7tbiWQGJPdUwr8wLp1VurWjgOV2j
Uk1vC1e4KmpKDiD0Rc1ZjDX73DMKTdtmojafCLQwQ1hr6ozlKXSOoRZ+fvFcNgLdbHFes1s3y6h+
NJPz66+Y9evyfFo8WOfKBnwq0z6VUqGasDhKrgxuF5IZ91KGxpHMnHcp5JHzKG/qb4sFr9KZrY9Z
dOE1xs4aWaDWZunvRrqjHbM8fv02vHMOBX1fpK+dMP5VSUd7EVrydw73Nq0+8K/7NiV9fNgJJA0h
P6IcEy8MouMNsebTTdYMIwA5iyBRHp8+LzQQ6Kk99WBVX2yAa6AHcKhTw0dCvxBlvCfg0emArZVE
yk0Dja7QmfUGLVgcZJ8wA0lSjtOozv++8JQBx9IGnocbimcOm1KYWxw4TQhXn1crJS/5oRy48FxK
trhIruoF5fsS6wfhvPoZK4tVwHigIXcXqcL3xrM9m5Hi+JnGKZgrNKRbCVdy6Jzg4GNKUfjecapA
/1I2p64F9WoVOb8OQzoOgDbrx2hwQJRoJ0+3iZ9wkVMFPXmzpMcdiNV16HgVBL11X867QdKJeF4S
vkkUZyvb8H5IqScCuqLr8QnTW0EzFvBdJdTliS8Szre2zqlXLN5k+rgnY8/tCLeLqQR0zvneNM+Z
XoKI7MBMMp6XZNQcUR1Djbe4qiM+BUoZI7dcOMfTKPdFIpIuXAsULOToONgQW27vOf0zwCHK6wLL
sPO8JWzUlxCyCiB2hWZYm3mAV6Cyg0Gqo5IPHEr6AJNJb3HO4LBay0HlXXupZwQyMOqh+uxEaUgF
pys64ipLKkX4x7ul4qsDyFZpkAudCNatgJXHp5691TQyWfIQHkBkLuYSEMhui0ykcxyma6LfBh8C
DUjPNU1Uck8fYf5Vhaqe9GzCVRQuLOTPmeV+so+syg8iElSq1Ko26Xid/j0V8O1SmcOqdWnD0qBi
HlHPMY/mtIz7/dBD1hXOXOpxcDndWPOVTXpQB6/E5yrqZ7+FxjwX/utQCZrbVtzFcWyBH0CYqM4N
Oe9jhO4pEsE+P9F0fdqQPVVb8sj8F4buD56SGcqK/K187EtTqUJvinSg4BhkRaVBrWx8rKxXFcnB
ZoYZIdfFguzEmO4xNH5y2yMA1tM2CJI70YuTEaUQgeaSUkElZ2+PJ1fQeLSBW/hgj6dtz3iZ23i9
cBATeOtxM1J/NAs7hvHSdnIbKVHKoRAicWANRfOAwEM/GPKy1ek55dCUG0wOvQRZV5c2+3i2eJ4P
wsbkoMxWHcGorjWeK3VqLSz5x2lN0sta0xUXQ1QprmCcgDrV8L71BWL2ESoqz4TLkUURKtCEZc0I
YITP/aPLG+XZnwGBBnee4Ta9g3PIgnNxFKTOGA3WVEIqaLJlzVsWMFTI2JkkKLUs5K5oYCPoqywg
FQyBXCfdfFPlYQShsWlo9GmDZt0mxqB1Dc1RRjuWyeDQ0FcANlt8XvhInWPXBaqApOtOUpo8t7Jn
C3VmwFy+jrdUf/+ZpNa0PupxicBwtZov3OWroDHKP3Bd8adJuhSdJ2vop8f0CfduWcXiyMp/9PXd
jb1NtC1+Q/IATKRarandRrIP9i45d6rEFkiyp5t+kVcm6u1eUUk0zmSjmkaMI0XsUn2d9oCXIjv8
K5JavSTdU+dqt5KXjjbYIcjjncbX3l07qOoTGkDLDXGJG8P5CqOnUZaYFxMVl4WOpCohEUSlhD67
ZF/eO+SPbkV8tSDy1ixFqSo0DBTlNEyZj3c58TcXR/U+tF095e0aARxf2pZsItgogPerd5AEcgOP
3zCMlxruC4jL7LkRNzn86az83mVOkFbLkMloP/L84OZQuEuT+VDssLy7CdVPFnVTRKqZ/pGcsvdP
qKhUC9a97PVJAuje/YOGNtA3XrdVl4Z7BeOAF7TMPUTseu9ajlPC6MFrCp3j++x8buX1BPVbejhg
0yR/L9lERTmPT6OVjjF7TFkXIVT/6xNYmUeJpbjnpTfaaT0S7h1oXZ8ZPcZfXI3RGF1UDgTroESe
zXBIrIZX8O9DGwqzZE0e7frHLcyyuxqU0UgwAqtew9aaBDSoz6h7S+Ic8VLDXFtLkE91EEmRxmeP
YTR6faz3lo4jC9gpnKGcO9/6nbhCr8zsFjbur6Z+bGMl9+6WrrHkQ3Ay+JE93qlzvOoZTIMtnQmV
XbeQehB4FiZlHH6tQFr6G5e6LTQfGIMp5WpZEwSvxkaGcQ8DKDVvNNfnhdFKRj5wHN0dBH8Kt6NR
hTu8/9xBcaEfMT3Z2aIr2aBVbBDJAzWrI+5ZYZ6nqI1XfmCiIfzoxqwoh5d4b6N5q3I0kJkBH0lG
Ht9XjTMKEa8LV5JvY+/i9Qhy1Em6sZcsBEZBSDrudamjHVIZG2oEdEPAyubGhd+SVJr96ImlRATW
8E8qZf1XEwOgXaM3oIdd23mq4tdb3qd9L680HTDUHovm6nMsz2xXLpQhiEuWFhcvmhBRQJQx9hDN
YRyN9hl4fybfH7CKBthQexxF8nDKhIpcABWHm327VeRzDLQjnTrs7GYuIOzRuUDQsp6O+InxsPK/
3kHj0ENccmTsx0X7RbMqZ+ct8RfyXBqfQ0fLc63Y/+Wi3AbjBQnDYMZi7RmRMyOPHiPongqSdKK4
5X0EYqC1QWfMm+ebeqEk4iFJZN1AnjhPz0NUIkUI7ju5c1TAaLaUirOf5Np2Aj6HfjzM6jrWGOaw
3yQcSpQrUV6xSk9wqYzHE91BYceSLba4kgRs8nrhS8Q6Yka/nZLg4ZsOL+UkLA/968WAkLx28wHN
ToMoXraXWEgV4TG41lG0bkc/3fC7fAxbkkbope08FpUOJIK9R6m5Waenxi3ZdJF88CGdPzNbjyKo
LEcsUgSWmupDwJznNxjXzjj2XPH8MQmUyHaFBmQ8qD0bTi35vIUjV4oya+7siyAZMPuO9AinqlTH
V0s/hCmCnehscVrenOgfhGUcAan3/8Reev2YkYrVwjQKcVj28pDI00gdCj0fwNryiH9TGJlBPuEj
M/X03GMbupmuLZNdP2nJn+Fviwld3X2ANRReEvUsBPDGGgYOPUFWd6Y2JX8cVlL/U4Q6io/8qyaS
sehdco+6jUpWrgVlOfqOBn82mfAokpQ16ApJokiVfn4CS61uhTt7SlpBsbY80V2oAAbjqJueY7Nu
qdEfuf7JmzdFzv0G9Qk1TSEwNXak4FkOg2aEe4ulHYUKDTQN8RvXvTvCk+3ibsC3cu5+wvwbH6dN
5zUqq2L/U0Va7YZ8sWMsoBwIMRcBXUijKj2V2SPlQwY//jjJwFa3BPjzFjSyg+ws6BN1LWeLqV+/
kNSs2Py7KGGzz4yxUNgMJ0NTcuVzjaCivsdrIYhn0A1v9Wx7V8nBTmLG7uwY442fhcId23nGWB6g
jKYV+6cRL0QzngEIdIcj0tDheghqLL5pJR1J9sjYU/RjmyBUqGSYztS3aEc4xg4VcDNGLQ28BjF/
uHkfGGN1vshW+7tghupoq/+wDqmqEv5AAyR/JegeaAiK0VWa26ji9S6BGhJz0X9ZN0OlWlN1dcjo
7y/FJuozIJFpDqL3VRlONo/NRdcaJv4mXbiKeogjru4OseLUhmYbKtePeERatAKSccam3KkhLJco
DHHU8FODK07kKZvzzloJ1n/stcihMfyMf58PENvoTWrE15Zflm5eizCfvUAYFD0o7cOfzriFcY5x
eFwOaU+kaq+RvjuDjRK8Ig0cIJTM8te33wqx7lW2VydTGsQETf+wkwEMy2xqyyf1mlc3SKBytGbi
tMjjHcO6dAMU3LzZmh8LpmvPFeWXnn8xzt+IPXEIHc44FxNWH8gR8mM8fYUlNZbGCyzAtERPtc2I
nPFH0dQruSKLWAzhwiTVUYM+fjy6IKnf6LL4tv+ZwCDYI2otB71siCw+K6NYzrLOW8hLxbqskS+d
Ylda3C0F9NsNzaD5P/WI6DEN7m50tMpw5Bky66QjufEJBcFO1FA57vDkC8M7rOwaWkHX14eBlA9D
AuSj5zooatP5uJXYXg+UxzNbAyfXAjXNJz3Wn1fHpmp2cMAejhksmWYs8vM6RafPxraQg9JyQ0Qp
PneZ4BumIdcjZPWQLfJnv0VjFYypICO0romoqncCZAi8EcymvnpSJQT+9hWzI+qz4n2FM64iMLBc
eIdLZ0kkJ8p8xhfkEsSHY8FNCTk+GsxGXHR9/KnrSXaO2YRA1OTTVs5ySBgtSMvpZFQNckvVLkIh
76Tco33R+sj5uyOyX+GGlLNrwCcuuLU3g9TOuLd8Rxm+ugvB7RrVJ4Jfa9nJGLrFJheCacp9C2t2
ItsS6zLLJ24J2hBHa3N9SOY4kUqlOI54oo11pI8s8PJYxrzHlxYg/3SAvIMC7xW1s0Jqw02xmkAz
6Zn1rM6DablH2a5c0GllxenbkxOGJMRWQsf0UPkGaRcVdQ5Bw8SwXotzV7Xpg9FnqXAUJQS8Aje1
1835hSErZo3Alb9BmwQdxQFuNNk8/lZZApkgaBRGwMLYwXHnC2yT990xkkjo+I5A8EGZX9fS9/bL
XjY28g03G/uJliIwTip6YWrKCNiFPkxaiaSxws/WzjtLblID1kz1npxyLEf/IU86YotPVJr3gkIW
vLtpCs7y63ZOBRxuddXDpAn4ch1ibPOLnAsv+ZQArWagBmC1NxOVxZy0DOyVr9kKMpdzl2kJC2UF
/tzFY44nzlJx4eKmr/igEYIigkog1o8u26hcKmiGb3cDZFjgrIkBTfuU/e7lFs6DleVVpGv3D3K+
h7i/ROZjAhMeuUv19+SCGNf4C98VIqwVyt1WGdFg1vK6SlIH7hjAjQGKesRuaaOD5shpO5Mb4hhf
AyTs4PXv4TTdoVQvrIgEDVZp8ErHdnhiM127h2Q5CtiszIr1q2VuxSLtCn0ei8VTRAQWxCBX2gRV
ZE/wKxE9+6cNSosUxBXfju1kpXlPgUv9lLu7b2Og/lNGOSJXucCSlPymgvQqjwRTVx7fY5Sk74em
wbPtoNNxHUMr1Tycr08i0yYV1GxqD5h48ODw5qeVxRATJc30CCS/MxGn9cjTx5esFWPX5h3uidvh
gUNVKZOBhupxk+QQWDFJYAI1GKu4b9KT8CWaoelJG3DAs/ZLryRBRidWH+/MYHxVIcnRjgwnM4Bn
/myUKuNy1V5vXEJy2Xpc5EEzlRzYUuMlclLwPSPxtxShli88Ew1umw55GI5DIptO3YlW12w8h2b/
lSIgElqNKRjkt7soOV0a1hM0UjFsJxV9DSNp4LVrR/v/C7d1hHId4+eSDDGpVl8/dR/HUU5vC82f
wzs6FlTow1p9HR67BMBWpxAb8FdGDIIUgdcL2O0euuwymChhzoCGEwIz5k6eiFyU/lcVozVoFMht
ALl4mMHtLf7QDVTHBDzdZ4aY+SBjg9AW1XtV5IcBcyj67mNfMdg5bAyQJAjNbFZ+Ev9qDfpMaPg8
E4VxP0DqFJ/iRPsbAXwoByhaZNKRZFUQXITZ1KGEylk5rZ+JYI9X1BWLMrd64DVEIrCngJHmTr42
I/m67E75ZlTIng7siEF8OPQ+Ud0/ObcYhNiUlEK0dL4a0JVl0r7LQMdq9hYjUkC3WZnuNVLQ3Ip8
msXj5Jxb5pZQ+v//iFJY6s3iivW+TsxuqIjG741Vw6VKbk7PbaekgOCohaaAF6reErx0jbtTI1IH
zFFxzBcxJrEzjxSFpRAEO9OYx00wYvedI8drHesl6RsZCgqXloKRn8nU0hyTczeUMWgQxpmo4V3d
4yzPR/LyKdwbBN7Ba44N8iVnUNXiNvCtgfShmqjqDrlOXDnZ8IZnfbhbDojpZOpcCzd7AVO8E/uE
fFQxcNYGB3k3gwn1WJs5rWeVPDGtXkuaP91ECUmHsZyiwpQxcKJZG0H2TubTA0a0wLZBXROx3lUE
ShLoov/o0+ZlMOkugz8TBTeBXxDEtnOMjD/i1chLicwJHsdCWNO0AEs72Xxow01CNRjTBaKFrYhn
nx0oU4YcOZhBGZoqUD/xdpubHMfhUsZQ/RBMmbeHcpvqs97sMjpNe773ag2ONS0gJNgpGohgArY0
k3eNDkgaQb40E16uvT4L/EsZrlpajEYvSA8/XN8ZRv0sXRLV9CXeHU2B8K+sDgFydiJG1787Sd0H
IHuMbaxNLYUwldD5UmU+a95l9Kyh6ck4b+GUeJakyf2HUEPLhh9nDWqAC8Thya7OHwGVnCl1xd7X
PpkWTRXVSDDBody+soBimrcqHKUIeQga5zmNgGZuBW7GBhS9PPDjAs63KRvFnEFi+1ThNMuYVDBu
02VJWFPkqODzyN9tRx6RuOlKMiiEK9i8RTaM9Dnqp1efIjZI14Ti4NUwjrUT3U8wDG92CzCgX0HQ
/hKIEhaLYkNH+2H9y5z3so6SaJ83a8PyiGxrn8Z8dW/cJDueDEKILe584SmMPDF1qBFbWgDjJ2wy
4Lwccjqw1jQFH24mGXh7ppDo27wwfzPht0y503iit/SAmTQpmsWpRKWmGLgf2sQpt5gkiUegomwe
/pf5+ttbDaE6rajT3T3pNiSZ5Ljfl/B4GlpFEdhXjxLGZfpdrc0r8hY2q+IFk/Ue8SgcoZimR/QU
o+I+8rdSI0mCeq58uPUORN7kSQvGnO+HODbKSdAApBIS7y6WDPPXRNFuEJl21CewtjMEmnXUIoP7
QUPUMY0johKg718Z/ZXSIRno5pXdqLutc6fH7PrOsGxeEswvLkIEBfW6f4X9U59coaY166WF4K0L
gWefR+LFBtfECCSSeADGHGJLc59AjodtWa/UveW1d3UEy5qGPIy7cL/uflQWuHeXTU+h+M6gUYGP
HNLwTNi8Kq+6lHAeCiWNgAbhrLakqJwQcHikf3uvLs8RV3LGac24KIfRoBkNjXXCTH3n4FA+Ghbv
fRxLrnjSMwY9woBcVAfJ/qR23J4irBhw0Jiw4PRxSgwKocbTBhq+WpgTyR/R/2nNutMKfvRJOCMW
UGSWP34QiXGoaiVAmM8CaNGGZYbEH5UbtMEXUGopqyTEEehwfsaGqUiBT+J9fKJZdzTS91vC6Rv+
zae0+OmzeqHXNkoOBiYd5Z+Lk/RhjT3D71mh8vkQYcw8Sb9kPUwN6eeCSVLtpiKeKcLnv+G3ks92
ICYmRbavvuAjTIhkccIVsutLgfLxUfSVeX+5vYD1qNd2w7I6seJXuDkEWRCO8OZVHteLGl1zoSeN
MNbqSzZ07EAR7oGSV3s+slmlFMXyZzZ4RJBdyQvLFzyvkqavJYdPNtTQeDonm5f01b6nXdRcaHU6
CIa2VcnoFxZe/CFN8DdAPtQyw1yeLSma/55neZSTwj7DCmem3+eG2ACwK9fpDIRIK7fmTPaasoD8
UNjn22MGJXHt/JkM/z8ycifhao+eLip+AIcEuoeQyBdTdauencEFPdmBe7amKe2LSHxlLddINdiW
UDWK87ndk7dOgYIFm8bwHxxZLN+7GJew4TOAwpsUG2SdHMwuXSbv/ysNbpP9Eh7tsUMC1vK2d2HI
sKq2zUCvjZmTQOywDAQFOWDku+yFoGzHYtJLEyKauAamXalj0cfdFejQJORO5V/dGSOIBMA2FmXI
/2TKQvsrKjUAwLGQWp/iLjkiQb/yHn35UBx3f0aG/43h/MCaM3S5D3+sjjQJZkKAHG2EAFLlg3HR
T0Hazx7r9pzL3RrQrraliMNv5ar8yfJlYuLE+SSpxtQaTclCNBxKXYCLz7VKHiu2pBsHiUAD1DbI
CRTIs782WSQI23m2QGdQ1UqDcrtkrH2Rt/MTKajsQlBE4zoWnfj7iI1Qh6EScnr84bhZXRgrwZiD
Yw0J3utlsI06mX/WIrSCmrZYGiNHJuSp1N/yiYUE8Eexy1/9BmenPsOFcqfKNI4wrXhbrk0MzSoU
qwTX7hmdDXfgYrPTzyuF7gF+3li2n1k9UJKRUXi4M+tFbaLJjlz4W3wdQa+G89EjEgohmnHFUpMT
q3iEh/rGOR3x0d9u6Yj1RuL7NQgBELs2ppvlsYqiw+BYJlD1OejOJeQTxVzg2jE3tPazgwGMiSnk
wfFBXa0wvR1l2LoAQG/9OpocvS65HI3Z+EqN+qJZL+HXVK9Q1gRoi734c6hOFIlDYMx/s04WFYPp
PyvshlkQGPOpc7HzUSwkxSKeBrXS6HTwZJQwz8IDIIpykYjJNlx4/jUcx+ePYudlxoWcDsmdeqiY
MJdEv4kpsGqtR8M9P9tKl2SDM0mR2dfrVrpUz3dQt9TcRY16+h8FwOXgBBVcJKL6XFg7lvaLFTzn
dqDjLwZYy4tOYN4VozSF+fAKz/KDtdolgi9lLRxHx/LYzCz9IQ+Q0fud+WFMDR+4ZvLjrd+AncGs
blLZQXyYhxU9lZCkIQW+9yHe+0sa5YYaFm1CgLZKjxgaHNHg7zVxTBOw7HDH+6okA8NcLUMQgh69
ewWHt0KFhq2VTyXESEC+fBlRI4rr3go6727+dSJFojtqzaZgVLCT+iOiDjWLzWaeIw4/9Tf4yAxI
286ebB70uM8dfrRcc0OE5JWaCOmhFoCwPjty+GuwxhHanVtwDbu0NRypf/Nme9DIEKPJVWeCtm6V
tZGjzbmeqL3371ndRklvxdffA1HVKQcSurdxVMlnbhbVi8c5ML7Gd54Ksjb90oxsD9zwGGpC9Loh
m9a808gqydGxE1kySBXos0s37wCOqeVKC3/THWU97zOkdxfJh+FJC7NADims2qU3mwhnQn9jPtNU
pTcKgloIUB2N+k/dzu0OF1tKxSVc71JiQVopYo6JVdV4F4o7M1Fhs0iroNbWfch/R2z9OSUEVEzp
Km9Iw9PFdaJVrBsWvdwLQvL6TId4lo3EFGiSrpsMz0JRlas9Mv+LXFxUEuBWHLyb9ODO0frI10/l
2zQet9DwkY7VyENQM1aBym28UeR8Zl1NqLJQ8fgDUpQY/yUxP+X5OEx90AUtfo20NzB9/104vM/a
mffNXLW5Ch+X+kMfXl01vrG8AU/uMprbpDflTh12ZmQb91HMbsx5Ff0mqjTIWXeMNJRFLmZPz8+z
mFSB9sEBZ+zS4ewdmdoHzKjs6zPVJ4rPov5INiPdSpznLYgSSVxc3tPg4q+Wi2OmmFxZk/naK+ST
Ib/lcUDkAN+OMxZVGEJq+EjzPnF82QzyybzihsZhTVkA7YOtxq1dUWRV5mIcNSdf5xMhvT/rKP/5
tjSF9DX//MfNvbKvwFTJBPyLOsDvn9Gi6W/XdzxNbnyfqK/D1zAQrb+y3M5haFwt2/wAmaSBZ++p
60+4Foc10X3nbSe0zbc6uK8lmsCZZkdTQHmgih7/ArastvAnNsi4Gz+SnkPR4C5XgqX9tPMHlodM
U8AcJcIT+7eJEmbN1dOCCZVbVVeY47y3JGan5nTbpOucYHjT63oZvWk40xv6kS5RfYUnKGBywL7d
aB3KqJo3ITQvG3wqCZ87EOtRpWB1XNibX6TBwY9k8185AQ1UjR2YT84SuH2f6dtoF8YjmJZwJl8n
fEWlAWsk9iy4AXR3bS64JLYs2Y9ecoytFjY8vavuThQzcEKU93VfLCj637qEym/MN9gJOjLlxsUi
scK1cbm+ucHTVhCsvv5iu22sGCG5oswzPgQwLJVqITb81BZqLY7BFql8bX8e5LVY2dFKYDNZkVsB
KgjSQ/eoQXcLTOphP7U14QqvopROjqWvE8FpS3G3NLSGBdn3nH98L0g9FLF4KHgdYizR7nLpiQhq
n0RXn2ZZqkOr6zKhKNKtndZcL9DcBDVKvrUaHIG2ICigWGvZs8ys+1d+MhZrqDoWNiGZJyTr/hXE
x6D7G74J8rtS4RWAnKRtnx3y8YK9fguu6CwG4AEqGm9XYANfEeyrUFq/Afwgpy1Hjl4GDxNAQk/l
rLGiZc8292/2XE61RjWneU4uZtJK9jh7Hvr0KIqvcNAXsCyhcFnJKp+TjWnYNyALt0Gkmaz96pGV
cOZYtBQwmOnpG57XkBRDc2A0sH3sUkDzD3RLSKlKZZjcDLeZvQGcOYvTNoGalH5nvjhmb3SSOGco
HY9tHnyDGPmpvFeA7iDdVUhc++6spnIjmCi5x3NbpxpJlFDAfmwMhcloT4SalVbHWFpj6MHxyONP
qszr+ZNp9XI4eZEWCJTyTfOBVyw9YqF4FX9Rqh7QkkZXBs8U3WZODM0LaaayKxN+Kb1mBR5oN2pw
4Z7LitKPd52l42lktSfR/tl2agUCLOy+LlIxlMxe2m9LjPUrF85rS2AqgwdJZT3nELHCuCcfZAGp
mtr0QrNPluK12SoySVFh52MKCW0sJdN0wYkq4GT1kVRVNwHVe2ZMb0PyFuetA+nDSwt7nFSffKS5
jg9EWKkephfxjEKcwaQFizVlHn14rRVfySyNU1pFTIik1f/8weDK/YZPIn//Nsw9UlzzKHzAsnxG
jbBYSdd5aE1DcUzkAcj9kINfrb0gSJM+E/Aec/BoCVuyE3WSj1Z81WsucU34YPe8ZJIo9mj9uw+O
+irS53nmdmBfDt9RLqtvVmPheNBxagF5HkCMu7EorZDz1qB2BbiAVsCFF3CQazJKQ6LmFFRgkqXC
nb9Lze8nVhtdqdcabiIO91ygGoT603OeeoIkYPe1vuIoC3V/5TApMvKgX2GIilWZZaJpH3fpCDuG
lFgQg9BtSTZidTIgDzW8rDyA9wUm6Xvrcb4sQgTKXJL0u5YqGPFjm7zepHy9+925AwU2H3stqPSB
xQwfuFIvAl7U7RjGzUdQbtC2uG9D5Yvk+++RQhDaGAx+XN2icRIlcxyYB13I7vphDeqg39PW7NAw
onY0fe4p78vvgk0XCRnUZwyiBAyERAbY6CuAm54PrkD2GtsyskgOqX7223y+Ku6l1CkBfYUEEFpp
vbS5B7JwQFMxIq9QO1h+oD0rs5IbXV7ZJEOZvPJXkZYF41K6eTNvwv5bSy+UYBgFv5TcUsnoLdzy
S5j7RkIoNkUAq820nKprC2oOaZHEoWTHqGEMVwUg5KJg+WB9aMRLqlSbbeY6d63DgrRZZ17VHopQ
rcJ28S1Bkx08ewVymtguxxKlr22Fc7tH5FHOj8IwUqyjnpx4q86aLzNskRnOkL7MTQr/bc3B47TQ
0veBlPbKPweD+yQySeuCFZ+PYWoRcnpqI9Fi2UEf1Rj7iVp57tNTHQvmNll2W3MF3IauOsJJC0rK
ne8vojSvzfhvlMjEWy2+TQg+2i8Kd6lL1hCh6Xe5bQMWZKKXBcr2MVi4i143yieMjbD56IEWhEZx
XXnz8v3kzfsllph73z5AjCzT9lc83JPE1cOIcy0vj9yYpDldnyU/sS3I8WhDZ2rr5CKl4dFbQ/eR
xyQ9KqSAGUFabxhv3kR7R3kjhJDyFG64XFC3dJNy+tNXXRBtzdtZA9D/LnWMCYnPJn4hHDB0WBoe
Ceoe8Vo+x/BavgcWjaTA9FwB+kgvaFXtGZJs9Jo24KYlscUxvKQfN2KuewbdiVBl0LrN0q2EOJh0
mFqqtzlNd6q3gsOLleT7wUGuNt7mm/kbZzXP5EPqLsbil/dWuvv3NULos0fpeQkQe7rCeWy/99Tc
KCgB8Bfy+cS6q1Y9fpktsoy6LxYEetk6REqzQGS/kgPRZRUJBGl3u8cjfXZJ0HM3PLHHqeikN/Kx
Dt2Hr1LVMU37ff9H8D8PpWb0VjNJsaljAoSoIV0Lb7KQnEe3LaPANX14fin4MtY9CIPAtML0/RS/
YArr1caBtX9GJ2u9af+gBPsN7bAxFAF3dJ/ZvJFZZQ51WRDxkquGN5GLJCiUoH7h+I/NecBOADuY
F/oUCc32ToaT0fXJLTjFsSiLUTgJNEw8PuhplCn5SZYT8UuunT4WQRxn2n7pSqLiFvz8pTEMzlRq
A5uMvlh+iC0xrHbgTYQtPgW1uFndK/2HI5REkI3vEF7YLxt1cstjPDfw5se4V3anKFJKGVohFQEe
4d7uOEVGk7nHuMydHxS4d2Yg4OygYEmN10p5i39kCbW/0zNdvEBa2alGSbhl0XAKFh9l4GH5a0Aj
Vd8VDA5v4yz6hM6+crGD0hqlzzCbpoJG9uwaqqPB6ctn1a4l9PZC/VQR+ZE0UHGD3vhCtj8M+7+j
JVWIXRQGpTL56sD96jyRE+PNTENCgeRsdseu9iTCQJ9O67+F3BVDTd81skYXAIgrRfURGFAiKo/0
pzKpTLzct90LE6ddjCqojeWHKlVqCqq72gxDmQCEjULRUT6yQJikTf0/2RUT/nSDF1ecOjaTRG/p
71xMvBiqIFVhZIO0URSqU5jfyuyC228LbeDJT/i0foOjc1v4q+QJKUt4ssCrtB+AVFS9I/rSF5HE
PegDIwbLiw78vxIvl5JpHSy3qkewNLdF/KTnjyVBrN2Wj2knXH06qUief/jrG2IbDA8jX95HZ7NV
zUbQ9WZvdUYkfYCzC0L9VUGwNOaFKixAUaDFBUZ+5x05+6Wa5eX+fRVorCD6uuTysgqQ/vU5ND68
lieU8ANLhR4Qp+Ah58OZQc5vSclry9i4py6ptDPHKKQnNcRFP16uYIfC0XuWATNBBUYrGY6iVdLa
sDDvCj7OAcGdIEixg7KWtjDNaA23XbVISDZo7HTl40bTMk5EELtOQDuZwvNqaGwH3wiJCHmoIz6v
W3nQKT8LXgmv7GNgCK+9odC2SSDlXcDyr7CEvItzxP0EAm731ozsv5iKUC+v/Zwuqo524odFickR
iGkn9dwPMN/ioZH3qjfT+sgLvpr2g02kBmkcxQRYlLW6ELtyoJP+VBkP05ZDw/ZE+IDODwGNwxR+
R3vMdTZPig8xGUPwVEY7JHqv3WKplErCPQ2rfr6tvT7U1HrUyxcSJoxXghZ8U+4aVlCcNhMjsu+r
jxiY8M1Se21kuc/8BW4IN+j8oYkw7hBn2iigQO/aW9HukGOjcgC0+Z11uChvgcC7lORhkCLovIXl
E8hmkXCa39wd2dIz+wGWR0PNyjf2c7n7JGKKTYSCy111tEEqTeaWDNnoOhGCc2Ek5swtLay+Ai9n
lpnqDM0sQa98x3eELLFD6KjaFjaD0ad3eKX+bPAMcnmZlW14Wp8ut4wO+TFatLTpW4EAcJcFw7dc
Ee54UCqqlHZP49U1pl70QsZyjo14VBN8GcwnGhJUiNNZsawR+3OWeLeh+J5H1MXFcFHyGqhGGiNX
JekBAz+gnJFjORG1gh302O9ptL6mm6cUHtBHIVqCX2WtzJGb1jN8ygvgi9sE3VeC/nxlH0YcvuGn
DwZ4Tb+DyiT3IZz8jikn6cJlmW+RAuCNa8taGBsbfruj3vVIJIISpaM9Bwqe+LExxkVyHfPmvMk0
uZeWzYS7uBzg9wanEcjQSV17yTYw8c48R2SddOizKbdVE/wNWbrQFUgbKxE3urR1kuJL5qus+yqN
peA2GMV5z5+dJuKefQUvR7eX8JFRClb8JfzReb7zQVk+AOA9P+4Q6dQ66cndzbnObfzPoRKJK4Gm
GQRh6jRhrPZaYykPoqUrvr4DDl2WIdtYJRt4bwXL1tNrXWB5xEZeCM/A393WmDpZuE1F9oIkDqJl
tMEJQQOEwRx8721EboKxt2CTr9zFB/rtP71pf5WWhoJLU3XPp/uDV7A8P/E1eB/26gg4NEf61Cat
lgJOf5dLOfH4Dp6bmGRiKggYAN6MGOiGKZUfyyzeA70JhFpcdNGf2TTtmUHOqa/sxb4wASd2cJxR
/YTBHLh4tZHg13vEfZCUWfrIt5J6ujAASOvTNKWV64GVO4FhtHs4Or9Ze+P7+KlOcNESphT3340y
wVgHTkquPuYQjMt1qBmpOrj2c6CRWqhwcY5uhgjcAoyrbAlWrux8BAHdHfR8iilBegy9qnfj3++R
rZi7Knmp/g/fhgHaHDddZt494/1DW3Byj1oGhMXUEU1qF6RgQ16EifD+dOYwhyFa4S9otD4x+zdR
HLbRu4/Gu6kyr00zixga8nsVQnqe8fc1jCkH+N1qLPs1E45IsRZBk8guwlVeoFfuwAenZFiWBMkA
NlqDek2T01n7tReSzQrEUZJOd6kSR5Hscwzlq/pW6xHGVsw5ArLHewDxXL84doVyh0Ud7gEqCIAb
k1BJGEe8KRIPC5ceQdw9h602Vq1eX1OLjcJP5ZGdJtwwntOpGzuiHPvykA0Z3+f0kvCYENpPjkip
Z8uLFX1O5LzJ58kVMTCXzwAj2idSRkVMVwWF2QBMUbUZldJ8nsMd2dX6rOGBa5yeV0dUwE08k8oI
8eNt8I7tyfPXmoBbeAMwNIQdESndfdEQGQIuYAVH2MMxwfEFO06BmwzDqKw9YWCAbzyQmSZzMNqE
rzaWKdeWWjHrB247a6Z3gJlLJOaZ8GlEsZ5cWbSQk+hSJVCoYjlmgJLOhAE+IL2WyDbM/MBu8fgs
9qaTWzUOE7z+fMA2ckj6ahYEo599MLQQ+aGNC4o8/93Qri3XFUEu0JAY46A3q+JDgCSAcOdu5+9H
VN4+7j79A+OKBy3JJYr2bKHDWk1ijKwBVDVJ2cwrawrJzg0CjR1uyPnFME8y//4gqOooHzwUzDeo
j1OybRoAvT2JUB4oPAS+QX5vNYLZHw+s3adpUAnmRuyZSQgLO8ryg+M1Pp4n3f3NUNiqHTBO4bRo
AyD9KgurodAiH8UdirCo0HImM1V8Qz7q4NelUwWtxtaPkT9nwgeiqkLq6SXdu5KOrv4DOu0uD2dH
lm+Z4PMcbEwcnbbCsvrDss/TLwivh7aCiOFVAC67stbxz6j7kTSVIS0B8+QOwHWG5bRO+tZ+OaCT
slC9Q/i3FYZI3iAOrhf58gxjv+XfJ4oqXdH6WZ17DAHlso1zQ221ty0534ZYttRlcFMGRKICoB22
LzBwVaThnlFjC/dti+PE85wkD046CpyO2kt7vri5UDTL98KtHPzSpHYHBrk9HE49gpSrJqSHS9hy
M2Mx/s6Nc0x/WhrOZAFCZLagvvDpjjxi9f7MIlUJ4EvQOxPYPPCak/QoyuofdJqAM9v+uQaoaw8A
NhhtAj19bO96Q4WCHECYpkOEbdpYhomvEVTGnryNmn9pDWjaBx6bvjv9E1DkVZCiENI1XTP33aMg
tiRZFjOIavR8YCqsZt1LzgsHPHXxRuPHDOcdQPDlj46ClbBZH2KxKGcKvtp9F/1gyLAtYpt5TrwQ
PKNUe+TbLKmH16HVp3hacNG/KPAQLVesYffE9JKwxut5uOv4ThD4iU4FVX9F3e+OMBGx1IIZWbXp
iE+YYYw4vcZlLkbJdNe9vYgWiEaHcl2LmxlUHakPF5J7YwUvtbKMcvRudhnTTvUPRfaaV7WtYywd
SFqjpe2NNztpM5c1ztBMrNjme7uiL8ru81fdw+FtymLGNVQqyFO3w/dlTfAOZgWnbtNcC+qYVWL5
k2fnWwpbXMkes3fNQIc9vq0hFDaeZeeu1gYI59ufHjsjEomLVTangoW7n3ysH+7WVjoYMdrDHKa+
mfyjw2gJRyCVM3zCO0qC7Y4WBDXtV9SJOqki9JxtThDNg/q/amY6zhGTP9OUgxsH+tYCRE6o5YnO
Dl/B9zId73aq998Hz/cj6WTglvzm13rM2zkkGc8StH54i5spa0+9ZKfFpAhFn7JMNIYRFwxHjNW/
Azr1kbnqWtmwWnmMpAgPorqzKfYG5nV//fLwBpmL1PNw4UFq+ESofdI4gkubk6+cyfcxi6Xyim7L
4XlSXWYFv0IV5IpoiZiV3BT8RAJMWR/kddkQtMTk5BKXljGjfNMv4ap2iEx11AzIsSe1LHLFzJ20
qdy5si4b18Av2giOscacL++lMw8eoaq5fdSOAUMux5fvurrQEOBH7tpQrELGO8G3c2h1eJTCYuG5
n9kBfgbjKVx+Ck/6ZUF6TjLHNwvhzZHIGl0Z/InRlSeiGKbGgKswtwCRcrrn8i9GA8DQ0jLAuR78
OagRLo4MRPl+QxExxbGrzB5sYJZgaeka1D10pKQmjJ/yNpaCLQ1TLiF62fOXY6IS7DTDP1vQE/pp
xKcH5Y5n6P7YdahRReP5ZgLfln5llizR+4aVepf0X+GxPYUpPxjaaLnDxCXCIpHkaBPeCNDeePM0
ZHqKn5zT6aTOx/enCk5wDTh29DGfgfZvH7yx8B7dFxqMpWojYBha1eBDBsb5hFTu9ig5CS6lvaXz
FkzgOw7CXR3uiMunx1Kb0XZ5B6e6G52zPtVxxH5LKUikWd1liZ4OeTLlE+EZnFwIcecS2Ftjy2x9
8bU/B2PjopOGnVXr1q73TBd/QDe1UB5c5pMYP6iX9H+7dqwYuYXV9CI27bUOJV3U3bV4aj/yYGWf
StBGH0YkgKjKTHQPO7Hj2vFN6TWmrSOOmE/k0r333nRuzdO9y9VLhGmFUXD4f2Ps3LJeALeG+rRK
01F6F7DphzA8JKEdHfFp/NEcQ2Skbbhan4F4mH9yatEUJnR6W/esaqiaBPImJvIseOPWdHkraWFE
JOtgz7izODmrAsklrn+yQV/8ZZ6cqI8cfnzQ4q6y7AtrlSw1PCVEgTZFXUxeSOdp/j2nCSiOJjif
AW0fYr0mBPtgkqcspmL/u1EaNH+hE+Kk/q8kAGNaLrJp+eEj820UZXBGWPTHfJmqgswjnvnE2VaW
8OX3EsgYVtfAGUug+6A3j+gd3ci97qvz4y/d872+1F/wdO/cjRNOxEqlFvShqJmF7O0D3PbokGKc
ax/g5Jms2K5qNgzaFgBM3em8yWlap1fT4bdqaJ9RV4gMG63YpPsYmPZtv4ikqFVBje8u5g2XaSss
4sYrdkAF4JZoibH/memq0X8eQBVuhDL5BCkUgtG0seM2Zw1emaViHkXiBQqOWFv60QSjD0FhexeX
5NHT+mcJd0MB3LPA1NIZvQ813iMoo8jabShTm6Je6Vc4ML/n4uMt4iMU/khBYlIts8XgzuD5N8VA
yk8XEb0nl24apjRUNdj655bba7w6OrN613VTkwWaik3mzn3MfNfk6xbNffcn/4LDnXgcunhYFsod
+5NNv3xgHdBBd4cS1xh9/5etlnMVSX8ZauJENVGVk9PjFnU2/M9c+iNa1XdCZQzb3biPc0bAQBL7
gZS9/MmtyzUOvXbk0fRCcREZiM3nFcMbdJ7hLkwie42cAASPhk+VlmdSDwuxJfIXASIFIwOzHybc
kgKxYFeEHSTrgdylXNTkQ+CtOYT9EWTtCHNEjdm8efDLPIjUXYVh1UoJ5eeJwj0aVihSFhdZ2n5b
/f1zDZPgS/lTDc734lPO/fQZYy9YtggYe+nHNv1zZcbUuIQSgvErAS/U5ickFWp7Orj/fL4qxFwK
pkpKOc7uWLVEwT6fYktx6vcv0PgozR5QOO+Dd1QflIi/9yOK5D1vgqPFLronOuWK1hReeeBXj6+n
Bvx6Nhc/eyHYTPDHCIVIEqAdRV6ceZiDoWLGu+o+0u4WLAHsA80iIehPt1LhZJP06VbYYAYu2PTR
FJfyqYJgfL/DeVRKXPghQ6QqzJSD+7SiP9du319ydMpTcWefowT6xdg/ccF6K6skLh/8hloWpmrm
5aRoLR3M6rNDkdkI4nYTDBOxyBARE++BF5VPqcQnNjc3rGFlY0dl8OzbIWKaaZ6KdaWE9Ac+zQvb
cyMx92Zlv8px3M2OX/X3haPdvHXjcaMC7ciOqr0wZd5QpVntPYgQLXwhK00aUN6jPCQxG5Viwxz2
tW43eHZfgLbYDI2pbD1dZA8gsWthMm/j6RJNAYZBd1sitwMfLtOF7PQQL/O8CbLRGen0p/Df84AU
u7Ddqr0SPTjYRiXMJsNNjBGERbcqZU+e0CipnQIVdVbPp68C7rAXFP4zvHdfwxg6WrcW5nDjpfRl
ULWHNSBDLe8lBIS/0bUrIrJ2JBusXhrvdRdnS7y17DWVmoqq0FGrFw4zKW4wB37qfcPbdQokAMET
GvTDL6opPrMm5nELMdMGX4Ph4OQ5U3NfUWb/tRdINY6FbxRxtmwAQB8/wFvteCQEV03Jt5IKEnxt
V/EsIqXWFMe7qabGYD37PeS+haoounL/sMiirfYtqwf5uHsbb6haNhwj9JuSUU/Ncbgw4FUvYHX0
G+pRIeG2E7EoUmTw/2h6yq9u4APCfPwrApzmNujdHxlWDDlQ96g+2MqYxfY4CesFkHnvAhr9cET1
DnHhvD5mYG1+YKN+tPqbqmLbkK/b+GJMU//cXqsymbICqxz1eQcxZJA03uFIYXMUmMwcBL9MK+Dk
AOwbPoBbEiG5gVaARV8oNh1Hlxsq6jHz6lXZwjsfP71kpxmqkVwwK8BDRUYFGPRH95pEjOwK7b4L
f9tqoTI2gEzE4osTp2b6AApGLgHuNJvjaXohEAZ7VG5ldWXEUHdsAaFhFcSf6NpAAhiXIKrl7O32
MUqemGfGouqvoMn82k1I4cCcyx929DdhB81j/JizoDWOhdoRTbU2ZzCSd8GDUS/kaaqXU09/fo5t
zl3ve5YA5TQQYxnobXhC5T4jxfq2ezWN3yKJKRgElBsNhKuwWQ6anxGtYlEiC5fAyogkOKH9LFy/
x0aCOmnQh10fi19kwbyEzoovMjiB5Jo3kaSOzN7BaxyCOdeeuEb0HboMRznobfd4gSdegLnskPJV
soQFWmjR0uCE9xCoX6bFCZdwwZB/9zdL04M0YqEZBAlJz7xhYHc1dHLpPRkmIIybcW+cF+hnWS1n
lUc+0YoRz6+i693D7Dsb2eoS8qfM1GAEtN7o057bkyrVQ1/5qJn+RI40F17cXp+Bbz6ZR5NolicC
v1wlS10EGzLqqqPVhTfFOi5JNnpaaHT9HtDzHj0iVivk7LsFDxmBTGOJXqzRYAiL4vMi43SAcdh6
B3G5TtKPiwgiJ2x6O4q2OyORpnTFUEOt+K8Wnzw6PUjXHmOgce6J5zCLBLPTPQhhel/9NMVKpA7T
qcO+GSZMuKlp5OQvZ7nlTl2gHgF3bC38TNGqmJX+QjwCeTUY0MGJOGIVqNtBdXIVt+Zt3Su3fndi
Ln23IZBOFegDofvp0AYuubf3xuR6b40KvksjERJCi+uOm6/xJqa3lP3u7X7uAbbN4zfThFa/tWz6
LqLLgzKUlgoEPli24qQJOv/pW3t3DTMFPlgnhVmmDeU/8E8wFMK6a4SIS56OP2b/bGKh0sTVpXE3
2q9gOjUIp615uU+VT2qqg03wp6OdBsQ1rnMvBhFXIJD0GrZ8Qe+sGJYE1meIEzvP91A3zwR7qmZ2
bbhH+aB8ZW8S33fgH9NGZGHz9ZE4E7f6W44DU/7M9AXdRjlfkfPrekKq2s1aJyrylXxYvgcPYT+r
UupIupWqI4hhXww56Ci9PGU/OhAsvNDb9mQXMEJYcho62Fbjm940ACvVkmstbYDZf9pLV9LZbYEQ
amT27umMy4zWYbeGoVoG44556BQN5P9SOUZSGHSfx2W3pB+q0slJ5I75+m3yEX/PgT/Es54GmuIl
Bgeo9u0R3QSg3tBEe+r3e0tyj02cgkiXJQltXIktHlIT2PF3MsYXe7PXdQK8sFVqxAoIK7mTXVFK
CkKNAN8vMIRlSFBbrE2TIY5SuZmdLMfxSHqQaqsqG7H3Kys2X3cA+Xg3lpv64PlK665+SmgdnuS8
eHPs/3MfOZ0OA3uQrUyQNMIHtV51hyutEwVRu2NFCQCwCYRqj0ry4eMA2wshWlE31TMzfFIVdDg7
xCDFyeJCDReZoMZpliguMcLtfruA0zbOvofA+VkNREaQz5T4bS83py4wSIvulbz/SAmT9y5jm7Py
d6r5lt9OQua2Bd3Ix+KEEsuG5Xbux/lGeOXGnCxd36qNnTxNUGqvQ8LePdw05zwlj7hcXHKoINti
5YPxnMo0i7G/6qZb6yiWGNvQhHp/ChHtesMYcYFw+e2aeQAuVaSsbVvzBIcFw2gvHeNJx9cdlDPU
V6CVYXHQk5y3iIU0kGE0aK7wmtfmHqgItHKWL++4iyy0vZGoE0d8XPtOpL6CWx2KabuAO3ppyeUs
JOtte/LM+vNqWzF65mXxk90Ln0AEvET+nIicqBwq2TdnIgBkGYN6B21BzS1cfXj3bpUR79K5MrPu
SDankb2ceyBvnmR/1PjLMAtPI9SbecL+T7eB4gZ7skKz6Jca2ZJ9lNyUrw3V5g8+s6gPqQ738Ck5
ZvgS449x16JRfcIr/oAO9hKkN3i0cPL5Kiqmu34GE//TaryiWiUyEScCsI22YyC/WjScdHGU6/LM
SBvH1lfPVgoraHhDG2mhBhe5VM5mWlYyH0+JMEJxoiCNIo15xxaqSAPwHRPoOeD6SqfjALtOB4DD
1VUwNQBDfQD//f3dw0nXEPFKQ/J1HYrpw/OvOIDTvELIhofQMPsmjmfk1SLlaPfqLiKUsSHf4y/U
HXDhACm4eLq3dUONQaRNAyhxSbSLaQ6mWjIgVQt9OKO+xWSjUfLmZ+wLJOgTXGDc1n7dHzqMkkB5
kFDZflNPEbYRsc6PxkuFh4EvVFKHV3gBmMXYpyE1e9tqmH0mXqBQaiy/hv2Cv55DpNsKh45X44e0
hRHKwttLNv5+ADOl4+QzGZbSCr3dlCGE40hNFp2ZEwuchakca9rSnp1wwaHAPP5r+xWIZATYgshr
DDTYjVWKSZ8kSMmC0OorD9ep39iUmn+Y6JGfB8XAMfxopuztiy10JWXOpWl6yHlHVyEdOm2OWTDz
YhHV39jgDOW5fjCm3kmkyJ3OojPFupFQkqsd5K/rs7LL4665dyGxm0WcFdo2+zgTyWoHPuWMcG02
eRUgiIkDpNBijzddP16/JmfEg9fpo4vPFPDkNKHe36QP9sKmaaoUrvjWgcmQnz6DVWwp2b2ifUZh
xqR6ddYPMEAK28+VRuOHfpdMlRORiBAz3s9udDFKvY1vVlgnHQl/C1UDNSj4oyGBX5YALIUQTld4
iicKJwhNC7iB7brjadlBCDYscdGHdvT/8TUa5yn52r4/h7uCgAxk+QRSZJrmBR7em0K9x3Cne69i
1E4kKS8IBkB0VR53Rg3XVU9eycmMW62ZXCMf9hdwooPkuLi/X9wtLTpNg6T2yNn09XEQPlOWQ5on
YeOjRO09yw8mUySRwKptx/LSham9DAWfQ3/L5sZxOtbp06xtw5WCq0LycgYUzBUmsoLQMWeIaHZB
RbqVDMEWtw9QMEoP8g9CBkAOOw0pIJ5GYfzU4tu2Nnj7EstEDaKk7EbY9B1NZ3w/D89ob9glnZYK
9xfzacmUKXbG9j73om7cVyuQ3fNyg/f0BNslOqHlyF6chfTwSXzkL/WfmpVJT3b21z4rRGn6MoWC
CDGSp2NRd3VsRd+2ggFHFZ45cvxlOcYTgZx2x/DDkWPycpxj+XrlCNe+jlTZg0jTKc5o4h68oVpp
pawFKZK+IhrPhswz7G32tL/ejq5IECDu5pcC1mwVyLc6cqP6lfsSR1HVydbm9k8l/pP13xSLzFGz
J1mQc/qWJgJDguLGmOUh00t9Q1VSWq4q++CgYjCGM9/qri+bDEwaYie7seb3LCpnvUEosQPfkGdA
xKsj8aHhqP2xnb8+4DFY/sdBup3Mbck69TJ85ZGjpR5gOUBcJeDUF0vxGPq938AGDy0Q+8h7ot2V
nI7Js4BCuZ9y4Su2DBZ+DHgSZx2ZJPQ4xJDmBeBxCPkgHWZWVx0VCLCKAXwZHJyndjV+pauqkvdt
q/COqufdZ1IQd/+NJXO5tWdMoFDGc7kEvIvBBjidQT1wc37+faWtt9bx0pMQ/b8jTfzBQ/J87pBw
aFLukUvhBLXhszLwXt5jIIuUAbjs1Zqwiy7q6AwhLMIdAMqHerjLL/BHfAMLSnmkCT2sU+ZAOVdk
1XDYWb+d5PIgGVtGf+w1QPM1f0J4XBNOENmmjijM3seUTuWodNfSWEEKHOMPNDdrgmPRMiL8+A8b
OQ7xaoP8yd+/y3AbSj+zpUIY8nQf2KbiX+PRmPvMIvQMJN5VxLzOJ4wgO+hX/XyH/bLTiEywUQgR
iiigBx9r5zYXlg0MThhuB0LO/o/Z3I1G4Pkwoo/rrkaKQfvlnAhfIuzOxPkOlcAuOttBy1/Parsg
7Jn4Gl2ny/wdEkHfx5afaM9jn6P4boOjTuplDtexyzAtRlNZBfTPLmUwiWGGKIn5T5mf/QVp6GXG
Pq8f9r/ucKJZyn84Mtfeg3AhHL0nYNQgGJGBdVJBPrVW2WTxjNI1T72QQxsqyHfTg58jCSxC3YJD
0oYULF17TlyYFy8ctsfnHlHgrv8eNa7fJqWOmAQTCfqSip/iuQZ+QV7+AMUNOypE/huyAscalw+B
vx7UeLKQ7mTVbJ+41jbEeXtsgh/vsDlYsaqwWEKawXzGXG5ruSl/SrYktiAz16bneWIxNqf1N9r/
Kd4dj9Yn3vffkCc+qathGGXoQ4WDzvLb5JmrQK6qiDAaLc/0NJY5lKpOQC7PpXEAsf4t8BKAYHxN
ojM8++BRXO/5gdBfhsmO3UeVz4jqcE0wKqp/I1de2N4izDN66IOp5jMmYnVJssMhOh6AYVa2Q+TH
XWbJHxVSNWSEEERX9u+Oy0DcmIBQ3VqBSTTWEKpQpLS+JZTtM9kx1PC7a/RCc3eK+mXSmtP0WR41
WZmm5sQwGAAQR8T2EceMLPYMxqRWYt6KudSNLqIhzExId5LHLIMBEAtF8n4QpaMwjh9LYKOW2rhz
P9XifOkC6JVmb7TJIKlpLgTPOnfRUucAJFBhVv5iXq5/VRj/PJuX+QFEPH+xxYFtxGfOhes8lo10
hJ+JA2whUbvjzjGoq3G6aAWMYuPNiizNAQz9HCsJIFNS3aZA9CzB3MbAFyOaaf9PXDF4+RCpUz9h
Jx5sJx9k3JdLjz83G22AMYVqpTvhoJ5CKCWrNPhmB9ogE9kH2+fpe1xL34I8qSxXnI6vfHjWiSzG
8omlYDDgDmgbrJotSaiu9ICszEOWMCc+b//vG1WYw9lTNeZMkHEl5551U+hsWu7UDGSfHRe0B0/7
O8MRWHh3SHlPxaHobfWEFQZY1cbHeXeTjG5yOnFkiwjG0kVTRbOLSUkG1+NAisUUbSQjvgD+Z7VG
C6G1c+AOuFOioF+OnPWkP3BbXOOF2diDERi/3SsP53gtRMb21Gu5/zn6BQNtRD8wnc/hWcMu/j1s
Owtld2NL1m4fD2E5J0nafZCT+rQHl0BZaIa7VhK6Pvil33/MJ+ZvGatJLrwU5bZWIkmJNeLnNWmw
aVQPFst+Iw9XMmJQlA+MRF9XO0k70EBqjtD0FZjrVKTaZneWudPEFHoN8KnF4flMDV3PHfPxRddG
XjVARZGFVjp4Rx8NlKlo/uSXSJbTH5kR0jouAnTVh0gPLq+EWhyVHLX07PjZ3Y2YITuRonMFkVat
Oo5V0AfItw7Cm8s6Tx4WJyVp7y/zpanqZZx4Kcm6DTiHcWTF1ApmODIM3l6g7wtscJK1zucHXZDS
qOqi4p8Cd2zhlH0uGNDTiEN3FBlFWB3XBvIIf01kHxB/sS5MDKRHlUYKouxUVUf8EP+R35AicLOU
7Uj4+GlPkSlDtnvQa8DRWy8H5rbkNYXXreUTIqLMBLlBAM3/G2NFUV8d/YClOdLjBWrcePXdnSrP
XSiI+JhN8iKmRpUUc+I0KIVokt2KIlGmM6S4rGrLHzcPLsTr8z/Fh03zV2p9i06r//egKY0cP5WB
3kItzJSXQXeugjoIFCebQEqijGEEOnnAlBQD/NuL6PhKsfDBTOwDG0W5kaB4KJx5bgQjfreFh/bt
0sj8L//p6mvMMMukBM4gnJulmSiJtb8scFBHbf8X1VAbQnIZ7x2/yiXHv5ydMHhEx+uQT71VFDta
TS741w3ZGIlqhC/zglyV/aV96STWrHlTUZDX0l6dS3nUpbs0YDKJsMqxProhtVcOnCQNwmAaeker
B0MtXdjIHYnrNEQESSysJPT8B1TTnvYqUgPqaJpv2xxqRtgKWEVWEGnlaONA8/1rozYgesqMAMwk
qSr5cUkoFQJYVACNYWHsW6/KpGwT8Ktrc8IU4qu1F1up8TdR7pTbd4WAMsO67Lgy/2T8Gfw6fwne
9pvJGcfAdz2K1cdK4SCXiO8bnkI59noXCCqNG+80UuA5lhaz9o7vQdTvzkeb1zJx/d/O+5RWssya
5M4uCHpwlWXSGPxUsqJYeQ5kW7y+xQ5qMfTxnracf8xDtIuEK/cXo1/OFqDMWRQvfnQHIuFkOk8P
A8yxi44ph5nrhoxNG56AdtKgXtBV6M7g/jVlMFmutZ3pVTQM5IZpHuUcgMOVzG1pKNgdtbAl/pqf
K2czbSk1gdBNH2v+6iBbXW+usty0d9iG2jsZUvpIiS0XQUca2bEL/wYJ62U/5b09mZdGycUWQpub
ubeiZmBHM7kvSDZPhzQPf3oxXP7mXMYTz7L9JQWzeTVQlNVX0TFFcuMPMGQ6TtydjDvM2bJIBWaL
ccpE6nIZh+p5caOvWcqym4fHAva80rVOwehX5PeovSnmMm06RVi33awjnGu5UH1VjEdJuw5oSHuB
kkPFLGCRHyP0xHTUiOZfFjYgA2VLQdUB3XUTdbXcBoOUKNrsH5JK7TQw3+MIVshb82npNJrvtNSZ
pACuQOUBB+tmqift9nwrZTetN2BX4KuaFd1RAgC8lU9oGNf39lgLa8c8aBgcKGzMF/7FqzCazYzG
eGNZwNNKH0HIuptveDDbPjgk7/3Xs2/T5Qpy1wqTnABmMIAliNAobJQQDL6KdsAxHpVCVOY08cIW
VcXDXTBMLKBshYJyUt19EHDG1ODCI84RJWvNgNdotfHy9M4pGhnr9P2EaKQ2xqU8n8DfcmMVOb5U
QiXwPxOLwLBlwJxTRxBqX/9YSEzQIRgMoJkqRH0fgoCR1NrgYWGFvHAauJLwVO/vxRCnFWiUbyVt
A2jL2MWB5yOuvtKWpx/rUGu3sPlsZUoWbYlU+lhYEiOo8WhbDelhHk1jZMFwbBWDBRyBP8xhbwuf
D+33dwhNdxAsk9dPGFCil+8hlvoddMsoJlYIi5qcyf2LAv+Y/EsBpVwc8Gi807tYYa8BN04So9ms
5HUT9Yba/WcBNnZZn0+ZVdWZVhJMvlC4Bt0awtn9A7v6hKO1rUMS2F2fKKpt46FVnU7xkXg2ZuO5
js0Ef1CgLkXD1TbK5i8qUoZLRMeEQSKeo2VL/Ne9qk4gQKrzebFCQwOTichu+dTjyzV/w5hb0Hfy
xxukYHoJ/6UcJ6hDWQz1c+0KOOnBKmtZtnjcswohWkQBW6bcym7ZLPZKf5sz1mldJy8PUwdljuEC
ShOmK26XwyLuy/ruqIurGogdfs5xR30zp8mwF6CuMwBcn05dSoMsWrGVtjm7pBzP4f1HOw6gJhMk
MG832Rb6zCpu/72qIpKv2CUE7DY9uKdJtE3PK1pPaZ0Luvnlv4xW/BGy7j5nKm9mIYKMa5tCHBC4
C/pIY6sw3gpOu7fFHQT6gdD7zeVmywBhadC0neKgmaQPyuxUMT8GPBMXKCuFY6MvTh5qepmQIH2u
1S5vNifV3RdBFWBY1zbyxPHWsCHJqoE2L4zLBk2Is2+n7LmrOTqcbHRV2a+1r0+FZwayauochPCg
YP5FHX4gGJodfD14qPPns5xgvwfkDJodxYRKaYBJYlDjvADamaNCQCPbyKd4ZaPJMlMCNqSLRNIK
ZPjfksFMDIsWUuyXww5EKkjjTwBNRc3tpY74JWM694IZKeak0h+NsSTaJ2AsIxqXlyt3n542V4Ii
XisMNBsTU/sX98N+JeKeg5nQgT+txvFAh16ekMhHmZnrdUOtMwcwt2HvVV588/Q3lG2iqeTpbKqZ
Mhf4cBmQq0TJIiUGnO5AECke6gpRS8Jpu7qSFgde+VRtzonJEzjhemTZi+4MPBagPQfa3qigZMTi
sYN+RKVvfmcpgwbbmxQjNPuvC13JbBEXCb5fticfPqpk0+g9/mKylBIs1ONUE/ebwx/BEq0gHRMC
L1rSr5ZH6Rik4yMU8i/GN8fI03EasX/dsYuMObVnjkaXkcNiiS7Cwp+bRRmeh9ACfsLgWSrm66dA
m2Vx8gc0LDVDtHLMZf941+pHyGXJnTdTRvTyl5zhRJoX5ccEuwywP25rJceHZgLWdv2KGIODsF/D
tLhWlWODORtztIL4aH/fmC7nKWP3u7vWZH/0FcV7ejJ/wi2gd09MaDzMvmWUfVP42dADgBBr9r+y
DSULVNvs8JdSglRAUamNurm5Xj2vN4vtnOZHndlcFcP0apqxOLJpdnYjpfWVWoV26xxAoDyKiOjq
+LnZX4c7ZoEJAAdR211kKGTbiQpCc01Lsu866cKF7iDVre1hWXcZMDq3+ctgHWzDp3Whxl1Lti/y
Yo04x+X39Z69A6kyPoMhn0VVRg0eahmT3GIbaUyanIZnBLCye4Fc5scjzXXiv/KPeMQ0RPNcDQZ+
e9/vH91vqcK8/5QWlRv1TbsK5HrfH9QPxmygvtHRI8nofLMfrP41vcidoOUucfITBydHigcCtOeX
kRn8uWbS1g27lj68DlPMDF8C9ltrAfswi8D0md4IxQHtYF52a9vayQOPZb2hbp/4WgfDolqQkXzE
jiBmWMX602xjvjymsFQ/9Cr++W+gmSQj6uiCMvDvDSUFzRXV8o+mKQEjV5sggwvS3vZNmSB6Z/ni
KRfXao3YA1dGNcG+Ik+a1okAODk1sSnCVg4ZGnojxpxftNkbI/SmVMxUFUznaNhlYPP4xY5Sljbt
ZBPSLJqWX+2lD+jfpWsrV5fl1Zrf5Lh5UIy1LEewG8v5UbdFR8l/yqCjZ+dHpHwgMF/9jFJWRNg6
OfZ6c7WROhklIIzUOc6SBfObkySMr9QI9pruU3G0jOpYhJrnizmhfVhYUlBYbh9w4lKe/iVW2/mM
3NZ97beFpvTRYBSLAnxQg9LXGlMupFgH1KpEBOvCRX/Cbz9NY4ZY1rzPP0f3QE52vxPs7KnPEaDe
f6Eu6m9tm9eEnPaN84QpuwRyFvwoUIch6D097MRfZ74Jx31Gux3Hgqh4cK3fnNAzE4BfTKDxDykP
4TkRdJMavE7sjiN3ObspzsJal0QgA+jR2SdPe+yz085OXLERM0J57WsqJKjSSH9dhd2Vr2huU0z7
TFyKGymqmNxwvrY5p2FdX1ytYEWZJVWMaA9SkZx0hvyggwHpy2RE8xUP5lJ56sffffWvLQx4quSL
O4Vd/Oqr+6plTrfhmlhKSQPYufgNLbiRrPiZ6Waf2vFH62fONH/hlWL/EyfCJ6NcYp8d9vwnmmtP
Sl4W+ASWumEgBkB5WiYN1zntcEC2BJ5pOQlLXvrc0m8d71V1Bh5oYY8ytIhvuJDQ+txeqmUdK5Qd
PA9o2gIqFBOVw+e/zzg56Zylhkre5o73vQ9bXH/BUDqxYw9K55PTbLkPzoZziXcBM7qKPkjYHfJm
7Q6HSmEpp5DKu4OmZkjCBt1CLZx2M2FjwlGbCM9Cn2FfIfD+qzl9JVgZK7vqHXrwIY3tS4QL3EgB
mWzfVsBzUxN6OrUPdpwKXfSs6+T94DRgw0oubPkFmtta2HOuhqETju289VbGVno2mlwBV4skRq1n
2POVI1EObE/wbmp0SxAoG3jYHwwQVEsLH1qP0qpINzLMGl6C4DgEKjaFkOHO4fo3CKmmt3htKl+d
ESJCNAEQIChU+UlUBYXRM53LVGwxF3pMjGwqkT7coqkJZaMcrJlSY0Q07YnN8BbKQ+r08IO+Ckzp
cFWSkOR+rPtyySIS/IAi3omWioGtIwTsqR+Pne94ZojEVP51/Cy2G+9KWKLkiP9WKLluNHnglV3+
KCbPLz7R13ePfbjaNF2IjDUhabj28SMY23Jc9L2nKvXGJ2HD3ikHLR1TgUG92cHBfOCtdhc/AccH
3TVDtbXTgJXQAt1doXlAuk4uPWeildiugpBpGK9K9bjVCuBBhQSismH3CTOh6HPY445jZGF5dJYd
YDcUGwmfbjRnRPEf3yDCYYkjwQJ6omet1NFDGSdL8fPUu77Gpwo+u40cXazn4nYe2wZjxfugd0k2
hdvWHmk6h0PzH77wEF99MiGIwomgomv8VYRhaC3PQWHB/7IslQ6G9wJkEwoCoIiDRgSkXTNk+LON
HxBw//YaWVCEMh1t+f5XOf77m7Qi3161CFwdcnK9Vo02ELU3i5nmvMYGOddtB526zKXqL9HRHCGv
iJeyAL+yA7B1Jhv7LXEDrahXPG95XGf8+XYfiehMg14Y1bgD6ZooCPj65hhdnUF8urEHQWCXzKV9
9HnctPjBA9invTrzYeMQwAVzAc95alU1tdUOCcC2wn+ha6vrep2OaJn/fnH78kh48Np2QCSfrano
gEVs/9V3GFQzVGW0M8LyhsLlclBCOF2/eV5qKkEJ9oWBISlxAaASTnmeyabH+RGHjn3ZrcmyiLiq
0ybrDi4zuocTx9irHdYNvsL3rBo8FcIPPwxvX+hXpQKhTZRTeXyuUyq6Ohr5q0e5I6K5ZCsSUzFl
T6/qj251DLoRH/iGbt9JNWyAi4jBa5A3NbCw7vb3aeZDVwMfIOsmSTo34Td7w5XaKNNtY+KkUsfD
W/ginTqnkXdqDcKrlNQeF3LqUiQtaJQOGuCkWpwKlAWeKZgU3EwoMsgt+LseREAbEkrlzIdUzvhk
+FXBzLiPQiKxnKp/csNHAFzwGKEyORrWrRbmLO7h5XNkQ8inLlcAfLyF1QWIlDY/yVoISBjcLoMT
uoxTlHG1dKr5adY6nTTVUGqwnXG6JBOfj9Qd77uZ3kov4uzps2gRVAi4mS0CVGhDohUGCNj0le7U
Tvc8FEqj3X2+EpSoKF0qScWqTzWGRzhYXOsre2tP7hIeiON+hAzGe1u6dugKOWl51O3mhPoN7/ke
f75i9LUhCPLdODxF/pBv3us5oxCTt29iY7+j/CE5QzvR/fNJj+gQnfZ6aifer/k6eDwcd2k9pXRE
9TDIgixgfk2ZDntxw9DwueHRp5jboJI0dPj9ziH5SXczy8Inq/G+zmMVznALgHJwg3CGz+spNGBI
JJKZnaf58uDsjzKGXk7AN/IPuyBBRfuWsQJNLVmpHZ+1TjegWvgRizJmG3IndNAyw/HiQ3blhCrq
/efxLgwSodVZHCFUSAB16t3KjimJjo/hWqJlrAbGSPKE2U7kJilVHssIWaiPq9psHovdVLYXxz5R
OYZIwG6ZnABhScR2i88RDhwqeE4DqoS63P2bmyJaCNZGVOSJq/AFPNcqQpWmdJoK+iIWaKnic4UV
VHfFBxYMT8hPPVWUPhr4goGt2kPwLggwHyy/TPyHRBcvMgJn2B7Gerd9XJM4nVCalPFzgAcUjWoe
V3tcRKQV0vnHTxycIsWDyOg+yHx3B5QbV5+BJ+OGPuHLJYxmHfJDRynsSIScpN89wNiP35UOmwpd
1uD6QNEudnHdPvfborFKj/QfyIn3Tbt5AIQC7Px9/DL9Q3zW2uhg26G1P0gpbOWD8PqeONejf1LT
rvGfwOJkgS6wf+z56gVGkiom02Feqb+pqALq9JTrbqOq7QKUkXtwEn/oC3QFF4YB9Q8ENlEcNMqp
heu8nI+eIb5DAnS24aByfLXhiJ6IudpNQ4DztR6zQyylV08cV8PAAUwFJMY6H+PhhDL/BTZuQj/k
hB9NolaEyWP1pRVNHxIT27bWvD3gvf4VRt9ffaR6UA2StM5EWmeluz+6yYOeIimmuAYo5y2WfA01
TvnRRaOyQ3A686cXfAJrIBLeygVCdlf8mRi822IIMNVnjV7FSXIJa3lTiIUXe8zax81/j6g2maXg
wtheKYi/YDoxTy5/2r+WTnjoxfxadyTQzKvjcZ36bcZMHHYP3+rpfBFDo2tBwzHh42c1Cpg4smug
oU0Ys4ZaqGeRXSnGMcEJ0/APH4NcTpvvy2hNibc1KOtxGJ4EB4YUqEtqkB1TRcuUqmnPvcXRb2Ss
QZnzQaQE5ALYgK5Mp26Tg/1UXOy2sv7QKLSOCEtX/ok4N/iI6UFoWJdYYFgbCjLpJ/IJSGcV5WKx
KmCfKH3DcvbsWi7nXeCADwgEEtbEqUCIoNAorASolI3pfVj9oP5dphQGntK+4fAc/0cmbbZy8VnA
ChTvoHsEKy6kU8hxKFraG0eGU6ksS007sxBvwbnPeA5gwOzyBhQC/ZTqaWbm3R7Fn0IhFCgFCWSD
75sIq3PCDKWhP8lXkNeXT8qtpEtkS6/3sZMN/F02NAJLwbI2Djo4VHsYuDdafFqd92j38JrGFYFe
BthQKgphq85jLege5mXp3v2Qb2jr3Ean8HEcY37QKHjixiS7N550NT/xeVdgzpRSXjFuePdtdbHm
dI5TJHPjfKhTYQ28xSq+32o1CjIBBNWlZinjm6sD7FhM2NdcYStE71aFFdDDKXPD4JBSfOg+LDdl
8DcV/XIToK3Wa4PBx55PRJlq/jXnvurcAnqrbNl0AS/2uCwngYQB+ss/2qYOTFm4HqFFCMKiOiOp
CtCY3eq7nz2xmcXxb1+X3aXgKD5OcHZzQBKhRsBMOIuwViN6OYsAoG07xVvylSTCqA1xIZsU8k7w
iBGEzaCWHUk9GNPmXWNsgiXgko9+aoHmU74NeXqO6GNfdB1VNq6IVHS94zm8Gj4teUlyz6/N+MCD
ThbWJKHOHHjZggXfWBee4fH44+/wrkwwNGJFfPAkpM1FfgOgGw3ac+4DChmPQ2RWRQDgczBmIUzt
EZqfVmtfYANtuMw2JgG4RM9wX67QUcl2/GnRu58mJWP5iXq4Xg95qNvPNLGppdoqjcHhaqlZ5CVR
wKX+LthNHCN3aBhnivg/Z/PWiZJ2qEqK2KUiDtd+ETWuT0FSUFy1SobtRe8F5ZCEMs6x4/0VlpG5
S4d57sDchD9/YLm4Sgvpup9NQ4kd0xVWRNIkcL1T9+1rMErdWYdPlUO6odXwrvwdCW/9oqifqVew
R6FKbZmC+d0HfLaaJKik5Lnrok22CFp9w2GUVld1BrFQKSx+Tz8LDSOURaZFG4D1SgGA1L7cnyqK
zbEkjpoh2NmUQEJoVifYHYYaWpTwj8xPuM5CYPTVgCfmjsYWLHhHGWZijwwMUkP881ds8tfggWh2
F6UFWEPPYVGd/EGDbg3TqHcTGFUkan84vy5hyA5jLdt0yG9Qw7jqtthlZtIOfHS5RoxngMi9X1rV
OHU8nZWdOxeMDvQvgaaDikQl8eheGIgIs52rRweDX7kAbtskDJXjuJQCroSM+k8MH2XznrxFufbc
Zj2r2F8WD5iFAjCkqFUhdnubPAypmJ1758uGzUJDc6BdSq58XzzE5goKPhEhM+pzpM6qhlm6/g8C
FXJkn/nOOQi4T7qz31Mw0IB4jBNksHm4QapFdRYvBZHVFSWkvRsJurJR0+1igmrJI2UUcDv+h1ma
iKJSUCPbP5DdlkyGIo0vSile90gZhW0OFW1+/4fX9iCwvqdwx2/romxnSmcnOm/19I1+lwNrEP3x
ScBtkgq5d1PLC2tYcxu3DTzULoAym0KthFNXLPiNfNHAB0CSRguR40XkOcmjW8YEblOCxHCYMGrp
qVeBeIxsjJjA6p1Bue1fnILLIy30f8rP/duRPaYUN7iQd8BMyi+RKguIktRgdFFvCBbv2AXneP4b
NR4UwaDPc9Ai4Rxi8bDKxVfUEWLupj0LCOvtgfr+M/zj6Xhy78Gb09q23e4n9QSCzsjMhqfvFJqr
8wQ0d/DilnwaLAOq3Y654beKmscKmKk1lHCn3OKs7XdbVwlS1zBWjJAGkqODcHJYulzAUaIRnXO0
csThv1oDyrpTmwlVKFBgYx8QjMr0hzWQgpZeZT68+NKENwQhqU/IjwNg2nAPCpbwRpMqvuyWGLJr
tdrJ+3S6WqW3RfraU25g/MKces682xhiT/zG3goARxgHykfom6CKLWjIxLp151gbu6BbEosxJbiZ
vocWfrVfU6it7VF4MInCdt9U36cfO9JRNS1e8vFoITcgUMyr78yd6R1VZQ9zr0Xu7lfC24C15GZh
vfDwDhPibYI/yJJMKQdZ8I7H5zJ0hse22GO60rt6F8leSjzq7O3R+XfPp0rS+70j8oJgwj/iOE/P
FBjeb+Fo8/qOihrydW2vjZ15BidKSkAX6hWr1S7FL42RbJcV1lqJyIcBq9pP+9R8TA3il8vw7LJp
sWifu8iGhMsxdYukGMW55OPE0HuEZ0SwWU56BGsR+Ya/F/R9ouJCKYe7hKSqMZuh9E1svK/f3Ew5
2OwK5sgdq78MTxVKLSxAA4cQnATv/zKvkz7AxG5C828rRbg1zNaxIKRqYFEa8u9rV2r/U46XR+yP
C+60jd+Mym9yaZOKdGHM0vv4c2wibS8zgrNvDeza7rv3yTFb/H7VTmK4IKTWfYCklE27SAaS+5y8
tWllxniMpbgZv3E4re8/YbjjuRDrRW+Df4PVlU3QXJ5uHr3UN4irnZ6heUiDR0nUx37IJr+OwEq7
APH1JvDyiyly3ey6q3UG+hAqhSLl2zB36qZRLpSqx3USPkoaowu3dn6xMRTC3mT2YGOXNGOvqkGX
V9LcIwzsSSogkOFq4XNS2KDj4Oc2KB3W9l2DvHpFltDxnwW/1dZ3GvUVjm3I87zGmALI+C4LaJ3S
ZQ07FBEkM/Nsed6zb4cnIKEJcIh6sbRCg3uLNCnuLbSygAyVJj/Yp8Azz78vreL+VzgK1YkiJUdQ
nkjxS9bl75NracPbv1Yqcr4PRXT4l9LsveoK23X1YDmqEdHixv4/h7W/yNtuPCmZ+CcxVeUt4VBQ
aYapUWZOYRWKBcutZFTjStrHI5GmgZ9nYV2oVLxHgfsM66kVkhbJD1WIbSovIfa75GQRRGPfP9vv
0pCnIfs2qHFF88Sk3N1ju4SOBkA0S7u1LjGmVzfl87xmJSih62XWDUnoU4eONxiNpkyYK3P6cZoi
y+f2g5oFL2zA2OL39Fl2vyf12j4ZjYb9arTDZUYCgMV+OhzbfbH7l/R1T7Eht7nam5fO6SXnJqES
jgUSAWgQAiyXb8mdnhlm6VFZivEsY1/ulChfJ34ktO09vc55ap5frmPlmk5mXUdOXEgIKCBNAA6u
FXZQ3Hvq6qnx0ICKAABXHsjRIy/0yjaWjFTmsfN+qpphqmGAZZgtrKQUy2oNoiUPUke1P30rxpxd
JJfffHVVuvJ5XeGO0IuLsbR4NFhqBou34umYqXcK93T1avsglSqf980Oz+WZ2Kym1fbEbHhZEZv8
n6o9BUFQ77To3zC20OH/BLYRANrVD5wT15Srm+f4x1Ch/4rSL+4RVSc5GlWQaBDscd06N7U7VWp9
NT5vGIoYxnJDP6Qqys4PP1txBQhLeRDjRl8fUcJz9CbjOhvJAlJpKv4UbIL2bLDIAAEupvK4bXcw
6FygVW8E+XjwqbdWuT8b1xRjhCzNhFYRcd+5GGaISKp9WPp6BzXHXJjJd61YlZPOjjRuggizwhWo
MIzm6IwFGKlHo4FH2v5HTyc87eEunZmzdFtfpfQKqSzHG8SK4ZVDbf5Jo0zwjrhbQTQ2M5zxslPS
5W0DvhKndbvc+z4NLZH1ZxXcMIR0RSWuNfYBQpX4sh1pyGQXEiioQSeDnUWLdvnNJ164pyohJmbH
kpf4Xc0mGpvOYlkbmMngnuE+lPjuC91xk0vMGesbAVyb5qEnjyBfZxrFwJtreMEU4KWgBPhcrclU
r8GrOYsrQSYYqvt7aycP16Js37kc7X4+regkiLDxAb+LeWdv+99+HrWdiToB3x8WYlLsLyIMadxt
tZ8MKsUwQW8yUFfTx+l/wnb57Sb9MWQy1EJKVvJQMFjtGtq7xPutENWhAUbI7Sk9DQgR9jAfH/US
5WxsyNkQO5fNWL9S2NDSOorE+zFngv26lKHI0xDTkCAC1TzQPiKQab3q55+xDQi92ZBU9gGRWSk+
/FybVFXVzyrvJfvo4Fwg4f5RHTA0B11z6MatDuGniGHWeJm4l30a5kwW5TeDaGkgPALQlbgltcuL
hpV7MhygUneST9I92ilCIgD075RyKno3I4WZmWWx6fupTYcltBrM0MF9HJhF3g4NytlYSHVfG96+
COn/eC3woMsJxNGedQK5zjTr3LaqSGWB6UteMkE1Cm26T0kuN6F3fJVd/WpX+ydIg7VKeZsh9B99
crmouHAHl6faVtY95CAcDDmQAvrm0jt7m3wX4HO7P9DZaT+wEawC7CWXpp8j8dZ97HeYQ8fct+j8
wnKWUejnbsfjkQ7wagJjf+vrviiNj/iSTaxH7JvhWTlRkFWAThLeoxWzH2jKu3IRK7BybELvaPC0
LKU4Ox6XzPqgfwguTTVePg1/TBW3uWWnZ4B1BgTJykLH3/d598A+Zz2xse0ExDFJeuueES1AiGoY
KJ/v2PbTlEjtfgrJDXsW7ZrsyMk8dOZg2cjZ14tOBXGrj0gzlrEjH6+4iQOoDOiuP9G402bDfcLS
4hTIWE9Gz39KyeYCtjGqsCdCFiqhzLlExLhtmOjhVZxqOuZpvlJEusd13I1TGw2OBXUSrL0y7Rcd
CHIeZsGpPYzdvCqrEPLXLZC/yymPwL8anc2oYEDCON7DwPTMlZaWGYI/fc/44D857B7B6cRdBOL7
6AbjY3vcQniwufsVPfhwxiE4DEGZT5aU8nKqr/od61gjj/+LlK+9PWtZFa2DUy8B4jC0p9KPBkxh
zngGdD/iiNYVtnopiusC5pqZYKhyh+KU4exmhN7UxJhJ/dM5+/oLUfJ75H/jELkpuH1kPlnOZZ4b
W0bhlEtq21uPlw75A/JUirTPSckXUdsxCfZ4vKEC8v/zz7aZwY+Te57Bwnijq5PhFoOavEZfHoKa
IjAEA2toV09z99YanPeEA8saV6LeOi7lsJF8X3SBpfrGwW9hM6xf7MXI66fy1aZh6wBxCNYvb5Qi
vaq/bVlTsEmp19ogMt7F68gMlZDDEQAOlvCiu9DRqn90mlL4DkwNcOViEbElsQR4QxMs8hRiTuLz
Vy7cZKDjsrZBOjg3XTJiiB3J5HVDR3+bc6e9HPB4XYY72tn48NsPoT1IvK7KhA8QXv2w8ZZk0CEa
iMpMEGlVpPvcFChvOMRopTpdopKcn1WwSA/31GMr36soIyBlqpTDKGExLxB9m5M+Zg9UVRg+uvx+
vw4Bt057WyGTUDjjvSInmNGU76Eg3j55qwByCVMkN6VuBFiv4Fadw2zNJiUVy/Vy1qf/oL2Q+rpg
ga4gL6zR0Nojm39QVo+wuGuTtqQsRI4LLbVCEZhuNM1mdlhDmmWvyoOQ3oa8HOBjeEYh8um6MICu
uCMmUaA1tTLyFPAyDVWIxvFiREXQMI86MZMzJqWFMxiwFHODIcQMnjh0WiOFGeafXXm4ypmIDT8b
+8qqNk2HppaXUcS89EVveK3a8jy8gqpdHbMdpUQYwr0wijhureGs3qhKDaFDWtwqblcH+cem3/YT
icb1BX6afLMOTLu2AbU5Rn71Oxm+8FFWckGR10sM/TwH/ozmPfzmPLOiefNXffAb/EQD3x7GDh0A
fT0wFXSklNrngvhwi62HzlV1RDmkjs1bZDmxeHAWj+M2B4lIftuk+dhR8Ct/CnvP5mNIBXv8j72b
RnMhzpiZWoVnyZHgvCrirPm57ZusaMfz08p6Ncw6vglOjPIalODmOi4f1V+MpHWrMn651QUEWjRb
g2n1lrUsA/o5OFhuUxFvZy6Pvosus9qxnS89jrcZv3aWXNPYN/BhyFwssy+A6vBq63by6w9Hny7R
ckyakSqSkh3WumzXzNnPPDM36h2o5yj6J25dztXIUzTCZA27bNC1B/uMrYb0llNVi/n3Oj+D9JHu
4FQMH9NjExNaDWn0Zp8w6bWGVY8FeXe+fJARk9cNAQXE6RkrZ1WOuIWqqyRwVTzSsxvlbGHf+lTo
k0+OxOvuuHPVV/ThKVs6/PO80W+vtDbIIH29N12R8i5lg42ypo/20ZLJCS9i7/Au/9wJi+ptMllh
XuFnWgBcQ1+F2wWqHo96Ot3VLWF/4AFbly7UJhE2Wxy4ZGPPKQe1y2AMcUQHB41aG2mXpThHch5b
jRzwcGMQbIsWZjhynE9rNa7PvK7Cl8idkX3e16yEGGmbpV3LISlkgCxakd3arA68fEodzkb8CmOT
A58udztGlo4Lbtzq+zG6uZ10Rq8MNiBbqnaQJlMAAZgj766TXdobcYboQVvOzBTOcGMU4o9mX9IB
jPcAMpYcfmE+vwFHR6+T07CcL5t5c5IDH0BBajaPCWttEdsQD6JYIi+KG+HbDMtuR86aWHZxBWSJ
rk7AiXPxcU1Cy8Jgphei3K7Nfj/zT7agUQ8uczsagFxf7XxGuHSWeEsZs2rIPNErrlvjv0he0lbx
53thwaXxv9mJNxD4Q1K2QKosTI8lN4tx29cH4XSHRaeV5yzHOOfCcLVEEFQyhnn9uZ3C/u4pi+Oo
XULqb8pVNRsW5VOCaEF+gESe2MphnkauwCWaJo9SgLeJYDM+hUcBDtXqplZvuvrRAWrx/fteSZ5M
aZ9NsU2ctshBu9W+V1dTPtvLBPVPawEMLXAkGCwrHNxdz3vXEZOqKv5jpFSMu3ZHOFG/xoPgmCKZ
IhCq04vF529WaycyaPNBv3KfWQoPGETIlo/Rr2UHkbZsCEN3icrVdIyIdl/7TfhPaNOTO12g3Fsa
Gu0tBUzZ4RAxDIkmshqzkqlEJUYn6yiYQh354SeWhYgpsCjwoS4Yv9JhvMvbXMcckKQrdJkZ2eP8
QmVZr0JktibQ3kQABKzq/jGVgTEVNTXrLOeT/lfy3lOnqDEM7ltTDhG45aM1ls7Hriww5zu3vY/5
Msc2AEmpJmPbzaIuhCcNu+pofjhu8qqK7ZFA0u+S6DWFn4128DqAiumqUifGtYXWUrIcXbdv/hDy
UCIaUIm7XEV8diwqdiuXc3vBvGlTkuTFmUpc906TVlpTu02MlBHG8Ckc4sP7BsXtkvJhkhQ2Jekl
YqdSkJOhY7NL1RQKab9UDveOtrPAl9H8BU5pTvmqbDHjSig8oDaaECcgapYHMFzR8MJgKjhm+WwT
mXkXKIdMjBsYdpG/6gZ91Kp4HF1KdKDIoANA6BMWrbOWeg9n136WJ1EcM8gAWGU7joFmZF80Zjea
+ELXvWAnH3Oa9Zgctc+gpHpU64MLW7w/3AOWyjtKvVkNJrWgBg6EqXpkjOzzpaB7f4eCt+qGfoRq
Imbu1CRcUQV0AQNu/fQTP2VlYxexAidZwYtMdR2XcBXiiw8A24V6Re+HB/NU0H2bmGRsHke8f2Zo
JFvSAqvsan3AqsD+NCCVSOQCVn1UzV2WrJZkt0GWY6F2nCHPIthjnFQghoB1wwuwWkjd4yreCm0n
hSNLnwLOzMR0GZO/JMMk5poVLKT25D/I2n5y5ZMsnwSANH8dgH6SFduKhdvlhX9DdOWVu8NGvvIS
x8qrcnFO31kRBYHauYRAll9OgNr25m3l62Fx+jwL6JSDvjq1js7G/HHoys9AtVd5NKFHR8hb3HLZ
7VkbGw9gD2QtPCgk4DCjtQzJHzHD9VAIYovmHSZSMOSZ72FBBNgQ8iCXC9bMLlfeqcwqS6KRSQRA
cH1AgklVOim8OxVWUMcH8yOfqukSSe+lpFRwAxY7jcKJFStLAHxU0Igf3e8ZPtw70Rp35zOwiLDW
HLEBVTHwXlGK4VDGVCf84VmNyhEzIYU5nlWCcCzyJSM9x++dpFOXJcoK8c601Vy33CGGeTnKT6l5
B2uDgcvkBlpkRuPSLy3RBOAaGR7STNniF3ma6D0JY5dEWQbkcKnnpZ1DtHnrRvWlqejdPJ4yOCIu
tCm5nX4cafs6VXCvneL431kUk6TbY4uY1+OLOQQ+YP008dAyg+omd1bCeOVqKWMiBAbOE81hDEBN
801j+D6ASHFyXmbrKF3UYgGa+39RNHbsqaUzMpIPMF1/sicXuBwZBNK4KJAqfy4xPX+I1HdhcymS
wURYrr8hZmY0sWl8Ywy8A2e0G7X5B5cTOXLQyeb0g+yVlsujet+2C9io+xnCLzQ/VM3CErKihAKx
RbNb5mVQtI3qquvLZ0fh+2bkWj5ACHjJXDLr/rPOQi4sp5bebx3OSZvW1a5Lssq1nfSbqWg5t5K1
Cs8IGGAvhIlnKfCMny0fl8OMJHokTCH6493ibcBgRR6V0LRQzyyf7uGUHd1YLjEj+36kEy+i8wuc
d8g4+wbfbqQeebhGCT02pH4UI/4lc+sMxnwdajYZSCMlJPBaSTVztVIZl/h9L1RvX1uk9RV6g1SZ
P4d2YdA4OrpLFZ/eMeKnoIOWhp2kKSYkpChsz00ivkxsdYP7gn+pRsaxvS9iObfTHni8pETubI9T
FMcrNgBccBXiX8QisrV021iOTsK69gZbgtPNNncXhgOHkey6dWaA0Mp6eCrseV2NcA1cWyB2h9qO
Dyj+Zch5gtb6tf0oY+WU6wKYAtfVAszbgowx5/9wHhss315xoaNKHUHqfns17iXAqOXr9vXx736m
TlFx0FwYHTx8y0AIgiY3GHd2+Tv9QUZkMjQ5235NDb377QeBPkkNdgCS6tlNphUBTsE1UlOMHDz5
1DmQWddKv8mHXxHxCJlGv+xHt6YUgxnZOCpkc+5dORnt3Y80GvtEV5ECIBMoGbB3Z2b8FPE4pC36
RxsZ9SgelDw9ce3qdE4j5lRo4RP7FHpp/jVyLII2vqdGh/OUujWUfELttKB4o8DmzoFtKMo2cAwH
yMFmwo9JbWYLzixCNP3DiHALH1miyb/qCscaXaLa+aYhwGYoJhUETicR+w86v7+dvFAwmKOxKFm9
csSeGZtcyjwNFZikvMM+hmuyv3dRB1d5ANX/5scjWSg2oHWcvyagqG4C0wM8VIhzQ5hy+hiiH8sQ
qqEUTrfs5udNYVeB6kCXTNXP6zVZ8OGkExb813jA8H9NCQwedr9nC1j3a1hqrDX82jKLoXM6El3U
Dlc9FqRMOP64NkYFCcTbCJ0Qs+olUI37BDLdHRGfZ++ozPqqss3/n/AmtiR35/0V1LS6bc2Uuhsm
w3LXa4z0uQY/3kiIrJWduCZ6m6fUspjhGwMpUx8oT7ONiasIOzmIU9UYMJO3qZkYOFM+8DMyEq1x
Tvy5kx0irpnx2QM42dbbrMIYlHOuSjotsRz1S+7POdpOy85eBz7xdkmnmIwLXJ0nAhMsnNIb24Va
oOZgnwgK88B265McYLhMKSLNZIzs16otNAJrw19C045/Az59HXc4p+69MasjCntk+RXj6SuL52SK
qlEFeeZJ/84nJE+XMigJcId/Wvj+bDL6Ef4J/ST7LpYmTvC62tLGD1ingsPNP/XGeAKvH437bnu6
w/rVnlSCNAeykLMu43FaSBfrneDWzFstNp3ps15YrvJszPxSnLeuaCtJFrB9SeDugKP6RV7oiKDu
eK+tkraIOeBiQb2DNIO/uz5HGIfgVFFfUkP/KKCmt3PUd87gRMpJUo80/KkfzmObtSxyxGkoAvUx
BjeD4wvTN09GFXyc37hmgj+rkVNYYp0SOJdKlLXPVzX/6gJ17Bu3w2nohq00Rx3DlwLal9NwSIuh
c7sXnTdQpdumGCeymeHDWwHCnWOcdHv+4dvurQO6pkmYke53wyaAqjygl5Ev3xf/V4oN4EAMflno
apk1qFV5iw7KiCZkdjgAUMFEvY1ey+KwJ79rSLUMDehDVm5mvqRHqCm61lww+Yrtt9A5twRRJXAK
36MWLnsiLuF+AONtEPxdePyGQ6E0iwcjtQrFPhVL6cW0BTL/7xGUPD4cgFBdgvGcZ1vpLSlVcL+l
OuCFhjj3qOWR2r0QUY9QuMKwksqAav65wgI0UEGFnaInamtHVor2geusCJ8PPRQXzX1PZDAZp6K7
pxSgV2Wp59Hu76y+ny0NzfpbpLsdJ6Id+5v0i5d8LRGJJwJ/nDFvnJl5zY4grG321qkB6ttjgXok
S+jb/qxJKYBYZ0Wll0DvkfgdM7OVyvAmQQW4/iWNa7KgCQmmP8AKqRiFmJEvSihtIDdqT5YaELOH
sghZCE8lqmCHfgKWMxffdR+YvpPRmgJx3Fa5xQd3INICbQ+TlqPhdE8KbOr94u3a+eTYQfgMgVBf
DyMTAplbwid1h7iuUqNDZbcedy3nvwHfFp6ZcEJ37zDECzZgwZfomCXjOAlAC4WGpVrk5gzCo8hI
Zc3sAcZ1FSKAyjXvlDkKpbIFelzf/B+mjRV7zprpAKN8AMCRp01KzIxchMLt2lqaeiZVIQ9ndUrd
ICbaySzsL/E2JYlE6IXKN9gc/FJ/e2GIGXqpB3lOrcvr3Dfsb1SvmiGpPirNmR0dOPeuvN0RkA9f
WI8PJp+YEE6V+dKApyZvlcGPoOsItf+QOUcBmWr+HPYjavVOJOmQCnuXmNBPOYEQ01j+aJ2L/6uA
6MB4HqEdzbKdmEgNkfb9FpZxpZcZ5dGNJgHevuArv/axmLO+c4OWZcFkaXDA5xiEYV4F3uH/PIVu
0z97kGC7MOHikkHBedI+H6o7bLzml2OM7rTTKgz4UAaajcduLg8CsuOB7/AQvPiS/U5H2j0qHOwR
FGZ3WHsztJkvUFI0zMmi0WrloB9T8SEmokT3v3kng3+d4MJVLU/TDqNhZag9mNcV1ej2Mc95AthP
3tjcl+v0Y6KZ/q3Sr6wGB+6Hx/ovD3THkCXV2ST5BnkvbVnVZRzNvYL1r4OsS+ixGVojBextviMl
puJkEZO2MY8imd809Cd80K9Pcr2IhVIEBEBJBxVmiQV7cF55laFpf5tyAE1Yj1ORMVt2aNSXq+vx
5MxdTd8fp4KSFuWlccnSkVIOlvotbVJhebmPH9VIAGP3nq+Xgyv8jt8ctYh8aJGUXRXoHp+qjLwQ
5QCxLsyQ+keZLNo8EA7p0T62sgjT/rBVlXJON+dS1r3vmoeVtiU8F573mL0R+rDKT3u8lLse8rjv
txTBzFYjF3vJkuCLzGLW3TQi/IgMiwrNPo9vgZh8Y/urrWWm0e35F+/kkYN5cZuKcUo0Sc6y5mob
NQou8QL19u6lKif4MTLfLtJYWvi3OnfR2Ew6DgRytCXlPxBBOeBmKWCHMafqAY/I/iu6JohwfkdG
BZnOfjQFIEA56/2agvkiuCLJqDl9eeW20vhpQLakpLFOtk9NXW3XxaEhw+5d0lQSYBhukrfzsOAs
3TGSOaXV/5BubovjYzq8odtkj1rEZRjLUg8Ql2rnk1+/uVmDXi4E8yDlw44EMUQ6l/ngiqJviRpj
VmH8z5yrigqIdLpI4gYolCPh3mWdDiF+vNnZs7Wp5iedZ0fnXCT6ZLLIZvsESbfiIHuN9aU2XqQr
Br3dvKeIVvK5Bq2T1JlgarSax4qkeWa8tA6lACKzLeZu20kJIVAOSdRW6YgBk3Sqbnnh1gxhHYFv
wvXPZCdb8heQWzPJMywgfvdUbnXyEpkxXZdsaKqTDbUaxky4FzyHJev6tXajQsYsZdT3UhSGIAwF
WWWmlWTLX4TtejEB5sOddKkci+KvelcTwPqd9A/5qBGPBpN8OcB/em1Vyk5pJhIYJelkXykqWn7w
Qr1Hy9vDJJvCFiLlzkU8JTGzE1s90wIRX0RR/Kc5nfyoM8rsIOcIwy+nH1bHT6gNyjoN3lNmG1SK
5KcvntFVuN1g2v7mIaBnMNwFqYdEGd1g8IzeEFMztDwAX8RWF8ulaW+n+Xx6e7WbEIJ7ZPaXMwBD
LnoB1Mz2akjfLm+yxwnDlSGccJ4xI9eapbygXZX1QdZ+p2ZrDE6jFvIHvS93i2XOIEmcZYZcjhCl
1uW2fQ7kxgmN1PBslHQ4B366u+m4yqe6dVo/GqNcfbo2J78q+kMcmia+tm6jULRjUfRuJPaJfmVb
uMj6XqFYRF+tZSDlEWWmN9iVbKzWP62+/IDiqAKL4c0SchozNFXHO/FtnsSmibyKykCRAYhJm9lz
xfj88BETUHay1G+JaFYIIAH7/ehdDMs6v+57mnzXlCtYhAzlfj1DSEL1oprvEkcp8r6waE4A1hpQ
0ZIL6L9HoRhzy9Ng7DxQHP2HQPnCkT3TAQrS3Qh+yMjGoMxWFLGIyc49151bsADTUy8Uyo+1Grp8
WwcfvPRkmWrnh4Z6zf4rmS2AMGinoGsYQhbEEs4xaBOUCFe5dLB0+Dxr9EC8spGjsHkYOqrEUTNU
5zHtfjsUVf1TdGpFJ+TIq3Wjl7fi+Rbn0eka9NfBvfB3ztyAPeta6rKwZS8AXz2/7ssfugTqbr9m
87Ovc23H7K4xJ1NNAHgXN8/6G6OGRCV2CiWORsgq/yrtXR4YBqOcjPuwo6vgD4GeWWgX3ZOYBXYF
voc6moI9MARquO4DnhibiiVncdLHMjitlU69/zZWNTTmCjcGe3IFBYwxWTtl8FdILa7MT0CrQqFG
avzHKGtVvA2unSEK9o4cHrhn3zkdbhAs4+LOcQc8CBwO2EJy8oZ38wahyU2ZKQgTj+F6MWLacI9G
Qa3jjZCnF6+wRHlsNILIGJZ9EGrBbiQefUvdOtcaFD72TJE7j2IQtX39BkTqEVPLm85UhN0trLJD
pAgcdNZczg/FJO1GKlTG5iVU91P84tbL3yKxq3BU8Fx1FNioKdxGK4l3eFCDtn5FLHisRFAyZUeH
CsPI8+n4TYbuWAK4wOVJ7ncANrQu9j1TlVL56zzWkRvKq7uCCA9zggCGhgQl7OOJBSelXh/M9W2b
81u5pb5GXan2jvoSZ/lEzDCcDZqYPmv7PV0JmOe/Uk7OX+fO8HFYJ5wt1qW/xRbVaff1u3duRmsx
XweHPjUydTKI0MH/0IfebGBQZQ/4QMzjrctwGCmipsnPM0N4pyUL9lgmv4c4SAeLfwzSWct1+gAt
wBNk+O9RhB2Jk/j+A6v3KZBK+CNLyi2hDJ2Ltb8SuRkysRpOywZounHTu4OmmkjI1dbNc4dCpurv
0N0rGs5RaRe5hK3bULwX9QF3EbfpYWBAWErKEoClLTZnIfBQv31b8K4GURAkNmfLnHDk5Qbji27F
nkFm212acyklOXCRUXYvqJMKL5dW+6lykRoqBXmi0uGzsk1jSZJkUdT8uH0ChdcJI0FXdEQdFbVW
/A2nhuoun9HXDIKTywBxJbUAVJBQtgtxPFtVtFX3DyeV2U231lNlcTK1b6kYKE8ZLL3Md7+Nd5SG
+nPBIffSY2zV7ruyr7IZW5QXnE9KBDRTbQ1pqlMG/ON99KVljX9mMQ+YGJ3SzkNp+sjUiJbdEZZ4
l984YD1pJSToQvotar3jHQ7Sbm2BuHywHFcszD1WVbmOr3gXPNdwnhe+d1uheEA4cy1MGD/z7eFV
VUgVJ0dtgTj643UpEXj99VJSYk4gz1oJIZHIPVMX6JlhoR5xdMRsg9hxceMOyxp3NhIEkE7njiwY
2TqE1UbXZb4McVxxuQdHPkwf0s1FcAaWU191SLD7mqrrayTkL3YZoDfd91jCE7RBnpil99LS0YB7
O88rCzcCUEIesHGIsgpSEyJkhtTolmhoFY4crd4AjfIB562d9IuBZnawBzKOYny8+slP5OMCum1X
T6dbwD9qBVFZ9kzisEwLdua5Wqi8DRI8DO7OXn1vXaX9OoTJ67yLduFzGacVPjTmNPsVpkobETv2
awL07UoqU7DlqFsXFQKLlBAvZrNrKnl9xQOjC5eYRXC3IQJbwr68+1gx1ltIOaPx/s9xnCC35FqE
n7VDmoDvaKRuQuvLtRcLSe2eXLY95xqORfATKzGwHepOgK6bMvQA5bdYCc6bVHVQr5d4WP80eRh/
+kppNTNcrJXFWLh3jJv1+/+Med2oXNycw0dSsSL/vVDf3luJxRyBxwPPU3L9AvN0TawlWKX5N9UQ
LyJ7Eqcj/WtM7bVpgQJlqUL4++RwVicSBiKt2XDSE9NReNfxhF6nzmrlmRHA5JMbcsCktdmQOmim
peAeH86xb4tpvsmO7nK1A44POzkb3yemSt0dHZVtFQC+IqsX9WoENgDLo+CvM6TAhFDZwHPeGPuX
Ioi8oqapePGhuto6Ce1bA0pYQMQzM9wuMYzPZdt6w69ixgP/VJGFZHe2wPalYsyeRkgJo3UdVemW
lEOwD4CcOZQNBrtL5aehQNnWkHgPEyVpxXd2y3ND2ASbHT5IVYibBTHrfoREDd2Q4UFr3UQaA9Ua
nOk8rW9wOeX9hbV8OVPI6yGTitK5WtFPQY0gcrX33io0aBv3Pz5AdwNOW0Dh8VRtqH2ymvQyp7ll
L30siqmncAtUjIBPAv74AMdtYf12hRLJkfiq1LtPEKhzrBQE7dwyUxdOGf2nvg1jZ9I9rgDUOZs3
RBEG8QsDlZDS1qVz6pD4Gd5VMuXEjenEjnp7DTG/ekl7cmWDi3ytBxJDBvD1hUNdoZv5/qaWknu9
bfH2/aJcA3cT2sm1kC1q1Hj4A1vObP/UHTtwrSYfAeayit3adDlmUGsxrn8C8H/vqWFrG7OKw2Dc
rZH6h2uIn9MDtRGLjx3HhKB/SW6hbN0d4oM7sFVfNzxK4YSmBjpFCVjJzAsN62RYWBklHfj+iHXi
TKJ26+mNO3Qj/L+u3SYxqesInc5UOebw6NjhjWrOMUSXkoqBWmCcb+1DRFjYvN3GFo0iAnXrcx6v
AONynBFEvTmHO4PaZM8t1jEXf6/DMTGKxDQJSa9rs/predU4G/jLAZxPnU5rzg/u5H0akeHPUypE
x5yhmymQXbfDig+oGHnFHWpheiXRg2eUROD+FtbJQqmvehkxPCmzkE+d4iE7X95CX6/p335vAumE
hwhYyEo85JUKSSYxJPadrFBAuQe5iXdcDEIhp0t2gBgDGbQeuIAKlS3ZtgopCs6Yf9QW/HNs72h8
QJxh05YyL2eLZqwzJI31dlXxDWJ3zNxbuib8V0Zh0BYsiD8i606BAi3NFYheXdYl0hv8gi5snl5/
pmaqYRACqzyuP206A4MEuCUYsn+oA9N5Psw5AxVkE6wQuQND+/5FTSCtjpqKS1ev1hkJrPcyg95F
l6JOaQ4lGdObVTjBvsSlm+f3p+hf6idJTo03VJ6hYMRWFIVmju9yakEk2KQ6/j4E0ZcY1KQ/e6Cr
iun/BQRYnD5qu2l/vCztS2ux6MNsvk+gHP3W47tFAtnNK/zmVEzhmhJU5ak6SAQpwN/F+NyC4byG
7CGoqd8RXwO2KycDpISeB8h3KhTjAjYo14rhzr4ZrhNAA7llK06PZcaoTBn9p0cTyZUEqOc8Q19R
nithz39lXgbbirqSuc/S1VmeEBejKc8HvLPazilg0dVLSnMoium4oYn40xY8Mrb/BRCk/8+5rcFy
1pUqRAX1y/GhmdIbey/4SS22Y8FYpcIILvRmYKVuiLyv6Z29qP+xnUwLpLIT4GDI2ywEA5jCkXDs
Q8ypCEpjg4QTbXcGnJXJeVETvRo/fxfeMRDuOCii66dM3mx++RlRW3st5mlWwdfsyKjRbWOyGJ3F
Q+G4BoYSIGb5G3Tg7kTk82AXz4SmC1bcQXIXPqKSIybrTHCjC2pbwq9R2z3MsJPFHEGFD3NXhU6m
cO5MrHK4eJB+u/kVSIu8jj3wv0d64e0NgV1XRLK08WohEErPwwDKmW+DqFhd7SNmMpetHdvwnmNt
IBvJxbWUMKp/wGkWCN+YwiWPjJv4m+r6uOOjE722IUkDn80i4fto8r6UmFTWmCilKNxXKD9ai8fY
+tYMTr9KGoCdar7Ao56yKN7tftl2QkQJxZJqUMMW7uMfZ/DoyRzYFAvClL284DSdG5iNtdtXrhkK
fOt5MD+pfophkW9m3XG1C7eC423dQijOwz9igjxEgPyjLQN7jzFSq25BHabRN10sQSJA5e3NKTac
cDfZtahg+7SwPxbCTjpwhkYHC0K3PH0yb6lVRxsksemhHnd6qAqc/QPTooUjTCaKihpV8e6cuUsn
VrQPJXiXFVTU00QPSdUHj0Xy1xDoFGVTBCR8ukGXktrslWeoKIFl5cODpVfBp+hhz/3IPH7ZcUST
GsRUgNPlooKp5iZ9GAzoL7ossWwzCqHDrXBFePN2YFJ4TkabTaQRc6yoz/KrNMQ/kalamCPO+BhZ
7NG4e1VWXR9EJw8ZCCIQ9qRM6PHTPYvdk/QlPFeLbcU9Jxpp/zROAuK96KowfUoLsBmysx10cD8+
OnvsQx9y4VEyOcUx0Jo6vkfUUroEIoOVnJmBVDPRDi1KiVdBi9sFX4MYQZgHaRSayWrFUWvT8hDC
rEiAOf4suSS++S/f812VXgcfjaK6UqDvQcejcGDEIRWICieiyoN3xNA6AATrYJxLF6b6E0T8rXrn
hQ+4waHw7+C+nBEPF2+ts6Y9aJU6HR608opOEc6VNe8omfSURuAgLWWaHnoN8ttGhgepfThuk3z3
Q7iCJceUBLgTvoFZWcx5KLlaHDx3jcpOVCzG284pHWba0FtOQCxnixRtUNAHoI8PiDvpUgJng3bH
uEtgYOiEkyZs9uzT/BRxYLHMtFX2HhqgAztuLk1oYqj23zeLz/nU6C4q0pWywXHxmJ3mff4QTP9K
WSDX8GgbVir2IhHAQKRudJydBgDrsViA+xRYAdeOa9XKvgUk0/qMk3fRMqBlWjLO3+M84ImD8rQD
mA370uNfShTD9rDh4da0o4aRc2Ekt02oCAQaN9YDUxhac7ZL8ux+NbpSf0lHuUvr48y3okvnNOWT
t5VeK2oAcfVGNTKRKsho+A3vAH68h8xDxDX3hNRHOJ3Hsf9+pHnOuNBkIyjt2n0Tl4XPMDkCRiWs
peIG36EANdmDXPqr69CWrQ3kdhSFXR9ItovjD/SYH2aWcyflGG9yDSJO/M+kUn9CJeA/A7iUUpif
7f+vBOTpGan74ZNVmfHgXI5nX/4b62x+gtJW5E3USZzt9MH4DQZY5ioHRsK4SzRgPucxH54WYone
KuJNhvS6gGeXrD+lIhZtp+k02Oj3DnCIsDXqJhHSQevz94SK2BqZAFqA0Yv5nnPIfJrprvGYfZ4r
z2oYkDHfYlUcJOOXIV8sk2404H+ovEY5D7V4yYlOgurOLG+ljWn5aINsEoymqO1Gvj3o2u3VmxUG
9lShT/TUjGqzQm8Njz7ciUaEYTIQ2vBV6debDm32zkdBIGfFDVabkvieUC3dstByOrzERhAM2DMc
LiXp6DsbnUilCOoz76a8IGi+eFYR+uyTv3p6PqD3/sJMLmRrpbVBtvaYOTyPTIjq4q/jDJAZRl02
2odAOyyDKdIuQxbM9P52woBxfaPVpH5THBotOvSy+Taj7SI5xVoO2qHblZwTQRA9lScfwStnHSiy
pLv989gc1gpCMT/eFv6BnVh6vXs/jb7M/4uVlUrOWUxWgRDVowY96JvDy31Pl7+gLsIKsR/8vXJy
H1HTHZ44n4rLMPdu22hLSnDkuemioMFNoJRm9386q38D3JDvKsSVghMW/Y9RUTKD3HYjyw9Yg8gd
3iET8K5rS6czcOQinlmmr7WRy3JBul1clByMBKAwGI3bnFt40DJfPCqBUKddD/XYeomeF8npSp0H
cbCQbwa/k3LcNthRLCSZSPDeJbFT5P35oThe3C2qr6/KsZFQtyqiaS/rbn/Q/9N/RZQIIJlqn+b1
5hONMHwzGyN/V94xydJTz6b9Jixb7KVd3d+yUuTbPjwKQXsk11kGozivgST9ELIdxviJYi06Kwd/
IuABy5bt8c8wVd2+oRGHldNsm0LOj3qY/69NUOX15Gr1RYX/dR0CLIYgY/uFL1P1LAU9wG/1z+cn
VnPYV/RXNyy8KbcCN3Aa/t7gutQ+3u3fl18DY6iDNJD9eH6KmKyTri81kfdfyoIyC7kdFLS5vgIW
KUDFE/oFmSHih5Cfcmd5r2zRgTsq/CbL+8kbltQNrKSI9Yf9JB2GhzxdtVl2gCgvrgJHF1ejfvPo
L57Tpst49ihOeLXzi38y6VQWYEoMETIp/IRKGL7YouTAesbyaac8qAB69Iiu/KKCp8JuMQHrrUJo
Y2k1y2GjYLmRDEE+mypUI4fljHt9sZB/RHPm/KCtfBJUvt39dkB6TcedAsRcUnIUZ4/udV864BL6
D4cIns4X0hT8z21RkN02QSGeFcD4MsMYT8gnWAydgjVs+PPtLtNnCXWyYkEiqlpfxYCL8Py5QKqo
QV8yoMiKJVv2Z67VkIlKIU79SeDrQRAEHuDbY/QQwZ48b4oxnHxcZ3D2Y4clK9NTZ3GsPAFY3Fuf
F3wyk6q4znXySySz1iBCN9empwmlgu2+U1p3yVh05uGhM0PliEq68mgmvSxOUj1L5GiFDWWxI95W
Aa0tWg6R68i+hHkZ/vNu2hRDgsjjL410QX4/MPKZHe4ZrTrIxgjv0lfJyKsd9IQTl7nPa9sHSrOV
7wdxxdJCte7fZz5OLjWfBh292FRBgThFCNgMG9weMllbzBYrzQ2fhNqOeMjprRjsLx8DQdyUXi53
KV9kNIUmBzl5qih7n9+XQ87m9mfXFUDLWAyGH52vysbdZ55GbVtrGHmclYTcBBBz1CV3WZCCaUHh
/nD9I1rxy36KO3eUOiyb8ltpBIjYgim9B+wUy8HcQx9AjqOZ3ktuPAFoAYNkc8Xp73uV5iWDTfyh
sE8d+64NMp752fDfxuzF+Ce2CLW5TPNQISIqMjxAsaSNojPfZ2+wfQmK1+m9H8jwji2PtA3o6Cnu
8L3dqBgWeUgs8YPLytEN+O5WUajIKrLxqKC1oxrzNU1rr519mjSwFxmmFOEuIWGqcpVNJlm8uaYH
j1WFlp/U47c8L8thgpXO073cv0lawAogWYaBXwJvmKobiXVRKjD3Vpu7sk8NQkzX6u/hHx5oag+T
orCMtAPb9wFcImbO7ueAxYX6YX2HdPNUqDPT20n9FNL5PN+uKMmbIlfswRSrVPT18O/wkCypJ55w
kAVIc134inCNu4poD1UPrRTd2M65tkN20tpm44tKo9avoHD16mlnbwGv3QlKTyY4Ar37Q/eW/C9L
nwTkOS68EGS2LMCXcs9ltao032S8Jy+vbQOiQPV16ZC0uF6DnBnh7IZradmrhyIsUCXCTS1SaWs2
CDQZCRAh5ArI36NFv4S/rK6sZoCU1PczY5UfCI73aObYanSRftSlk+8bW91AUSNB264bNZa5uwul
0zt4z9vKVM6z2X+0D8G00g9FJaOk3kiL9nDmo9FFCTuIF4socDvzjZ97WKlUyv1yo11eH6L1F2xU
MvJ3n05AxfgW05oV8noOQ5h56JfIhT8ZmZCej1R+rR+hPD+Ya3YFjzoLTSRvY55XzS9xGOGrJmxR
0F0TbcZXzEH5a0UUhc4srJuMA5BGEvNak706BOkavBqWMwd54jJge5J43Jq8Uo9vBKTKxuwS3n8Z
QfvkEmuXdEDjy48ArRLHoksqkAl1IPfEKi033cR7mMu+TJH2Q+9sL0RdUtE3s4KXMH6dTg+Vy0Ea
0skWVL9BaKZRHnez+sGFV4E6MBvOeH7h/jC3SdSJznME/E05HRus58E0BYnIItdLLBXHdlXM7fo/
91OLcztnyaIE+O1PJUdVIdo7EK5J+4vo2/TQydJjmsmhYCw7hd4J37mMahY9QN0EFVFpD9FAnpkc
R9ISKUILKXlO0uz/PLqPM88JM7xgyhmCkDlT4rkyTLOJ1PrioM4zaWoizenBSyZT5PmlJZiQW6Rw
Rj7XhEstxNJ81sMNGrbumDrUUkJ1BibnsuW3LgBJ7MAfr/aUsaPHM5lE6qZOxWLy5tVDL3ynPMcV
WeFhQVn8oHr+jdzWRM46dgmF60z5Il7T703j2zITOR4OpHnd/vQqU4l6fj/S6ksjB7IFdsJFuyQM
CjK1bQeZ8cCUr0PnDYHcnXlX58CQPqhs5KWCtFbJYja+tfuqf2PomNVMzY3Gi90YKzBlI/sMt5xP
iMUWgAFEZl6UcQGYucI9MTcU85nYfjjbdFSb9/UXi+l8arjzUVR+WP1uzXmVYLCqJzLWC3AcwghL
k5gmIFi1Jg/XU3FZ6nkIj75Vu0pULlsdAsmuqj10X4v3mQO7UmswcaLI4UZFLGlQywH9g3eFLhwT
XWzX/u7pzhOZUS5QhslnxDukuFijDLvhK6h/Ja+QB5hs/uMS1mRx0RPhgcXSBLUgFk5hPZVJiA5A
obObq2whvYpb5jHV+u2oHfLZm6yJURvegR4b8lOl2SbW/PjLspemaZKIvImsg4pbW3F+DoeNGU6S
/aAVWwKaC2+G3IfxbB0NQdK24S2VR6hJDwticTSNS3ALPdS39ykAxsW5Wmk0SJ4GpAyCt2YJnK76
ZD/KqXu3CK2sGPVh1npOQ3ACQSJjU/ORrtXLVq2FhTGMHwiDI8WOGID1aaF49y2b/PubW1G/kM5/
NPUIbcgDaEbPjW6QzMfMBsXlnRYCjB8Za4YMGQEk9uK7OlMgTVzK8ATYZkGYBjpadPkJMJ1JiEOA
Ysuw5JzW8zdpLSYwhFWRZGHLbhVAd4sSesYXw6ysPd83QexQsp2FtTNeh1lvIId8jz8f0IOi8bOf
Q5xsv/LbTYdYZBbsc2Ss6v58AJK88YHGYXVh3RmaONiUm4pnPoado+zS8ISNlfaWrmYI+ceuznCh
mkmbsGENSN99BMWTQgLXEgujXFMV81fjycHbe79r7haP+KgeuG5/SdWVhtyu4nEqy+9y4tyJoxIW
tUvElRDJwVt9zWGBOopw5sdNh9KlhUThE1h198wuntykLV5ZL7v57Mst4EmwlecjKz81wN+UGqHC
M5rxdWOLeeUhF+LOTpUhNAbTph4uRkAeBueBzOHd1rKkUbjFpaYNXEVEbYN5rSYC4tAAbghJXDLx
+k8+FuDQoP74m1KjnM6RYDT/meLPD0RcA1lw4WaXgJ6q3SrdAY3i0zWtLuWdk8TtTi87ljvO8Q9z
zo4kzwTRBCh9v5hPU2rRc0sciJDg7eDa9LBsx/ZNYb7d6/fdKBn+YzfQ9IldabpGoMeshYsP74zH
9kPFAsE7Bg2kqFTxX+fABdxFXG5qXFePPe3cRCe9V/Z/JAzaSjSEDYgKgTetS90HGCI6beaotMm+
NRNBBJSj4igjrTdI4UUc3r2WwIDzV/6YpNhUxR6orRgqbUlGEWvMlAuONavauNLi7Qi1ZYes64rI
PAMgEa+dWAfUUIN6JzrwQ1MAxNyImhyRflqaVUyd/p2Qo1iQ6intkQkMJZ/BbaaXdAGtMM5WB/4Z
x3yhRLaNVZKWnOBaq021/UTXjZGdX5SYCAbmS7e6NWXM6GjYhMnr/FDc1ap886iDBXn0I8cfR4xy
FKJtbfz9m5g0ZIZXp50fIB0MbQTN/ytbhyPKMrhDdCQmVQZBeH2VSmGzmoXhm5AQGRfBmdEJHtJA
elAHs7pA/mdaxtD+KolQviAAi5AgUuJvcjGvMGs1098rpWa1KjYIoMaHNQaBbg4QOMrTMhE+GONo
Aa/oln5WQJz/BabVGpfqVvijrZ9kQwWEs9K9r+UGR9Or5+UX/OVX87qmkQIIexmQf+0NbrqFmaRC
OkhdI95yG2ENk3Kqz+LCa0AYbJRzbaGkOVH0xrBWiUS30iSKcUaLIrNdwh/mmWDiF5f2I8eciR1X
+sY8ieAX82yOt0735V8tijlNvoqJQs2Tf1+fKYr5XQEZgTIunqT3fnblEWxPZ8kHwRMU+IwPfCsu
fDqZ20pU7a2ZFsBpEfZOCiin7THpaxGpbSDIleUTdvrICBaCaYbvQLypRMn0AAdsFm1IZCesM4zv
Tw7poLcergbpdk3jo9xfwyzSPuwdm5NkktGO1EDpDiWQTOZblEbskIInS1wtvOotwyB7sOSXRGKE
M9DqwTSzeAMRhTo3K25UjF2f4OQYHbJ5xSLERaXAvXyjUBJkxH2kjiGT41Sl2dtm0Vh3XfcWIVNz
dU9wOijNpbT31AK9j2S0HYC6Vm+YucN2pAzURYDOMY8L4cWx9zpQgmaejM86aJCxnsdc65k0ef+R
S2yAtqRFJB3cQ95WpPTNvl9koI4vn/AN9HCeRt1wVxETJmj5F4QQrWHZay3sqn6G+dGTcv1A9aYt
lBfU659wciciqU9AOFX2NZzy+4dSMewBgWsB8cJVdOycPPA9QL/KaNC3xEoobDFzdSTn1XyKZ8Un
uVRoOzXFdEnFCrW2HktKoQAaaek6wBJIoL3Zf9AHu7riI0dorODNI86yDc8OixwVsGp3aUwg2q7r
BjK+ZcQm8We7ovqx6JWPqQJAySZsbiOOdjd1ERaychIS1rk0o71qgBIAnI9y773GyDxGIRTisNxe
5WcLZoHUYRugL2hd+uMj3w4/Eg9ipXCK8pIu9x102bw80xWKDi3cDeOqXIp2M4GCu9NTWY/IujJm
1G7oTCNRy7wPAOef5ny7C7qImkZXaDmeksXOI2F68NfQRy29jTeRse+kWiNvUwxkjHUNKUVnAdrT
iq7P4Bu4MSkBPmPo2nlF2stECMo58TjlDp8d36oyQVk7LOdLbzwULjCbW0ZdVtDFVZF4l3Q+F/ot
PF8ApI8loe+Dl0o5jZuoPFqXcED6J7y9sfbIEo3Sg0hFDqJ9usYOsrAAJEbX/LwtV5Ur2iRRAFIH
22dMhlNUn/lFX6nvN4RzHAxB+cvKXSUPqRz5tZALLR6X5dLVf0ito+2dVMtYTWAKcKNDmPtqnIhu
bajj5kBdbLKopmxGpjAomGHsuT8YmeY/N6cWT1QDGfzaZFxBejjUJ8B0thZj9gBDrdAA9xUzVXS0
WJEAUkikqzKHvpMdl0N3DnocOkdj95Ebg0NC1Zf4e+AngXK4fJKbmfRBK9Q9u+7RqI6JGkgbe5f+
NXIYaPLgekgOQKAwaW4FyxPaoGr2Niig24GouTFfc22fJMwN+Cmmipb/VhT1K+g/EvF04fea9o8k
wRpMjRZ+RaTEJLkfzxR3qJMTzByX2xSwMu7EML5O45VmkE0IdRUFZCnaz3c1dk1y5R8IumUDOXX8
Ia8fEQU48nEftf8ImVXFiQ2hlbMKIsDeEPleLcI4PjoPDJdYiZjUt9Y43lkIRcMDS5dy5YWyhF6L
XlZmHVs1BTKdI+pKOojyx0QPzEgvk9snR4NTeTZwzjcreQgy5qYC31N1H4b7D3r7urDp419Tw2ch
gEsnxY3SEx3LD3yJKo4Lw/ka76Ln67UR9AzWCZJG8wXvp6ltlsbCYUodAcsdz55IqYRClHgpPb7l
MMkq3aG4DFO2S6ca6sTp5KQ2fIF0bSjxvnORizYSUEEJ7qAXNgFf95t39gwM8YB+2DUSXQX7UOOp
P7FkESOf/h8nb+8KQvVus//51eFgz9+Hv+sayKjKYYGfi2pias/8gKqkucdMVjAFJ6mBwjf4szvA
fKqyFTlbUfqAntKQMLIiICJcPQS26tQLugQjcammIN3CAXlwhjXspFavpp8Sg9dwteGsD8GrSsWK
V2SGJGEhNizG1UnJUxyncgGkziuNdjC0xFR8BrSz6TMtbAyNxzdE81SN8Z4eN/bMduIyodV/rAhH
wtuAokXmSb7ryDaac08FXQCp+/of+XIq0h96U7ChqeEWoGV7ocg7Cb8ofvFglcdrDgfAvCXbKiEo
10rwcUsCg8xD3b3lolO69A5Zd8mEs3dXFv5EUieAP7aA76dLlduwRpIdRAy8TMpPSSMG2y2Q5BFt
m4akJduij2mOMq96eRsYiKapnv68R8UMGCcSv54uTW2EPwYNSWmXbRQA89VLXKVimglxWi871d7z
2pb+ImMSNVPCILPADHkgjoTu+m+Ph6bCK9hNaxCbBVGkKUaQ7twYAKwT6TdgTUiyv62kg7IVS+73
lcTUJBpbHEiFxBSq2X5gucEqs2nDATGWHO2SSuT26DSS3ZEXHjjryXgSLF8tOHOXO94aCleWg9Rz
d0bHGsCJWHATKRz/yEKU/FuxBlABo93HJpJOQjUpJForAQOk9nPatifS5DP0nJpSWXM9scgipn3o
2ZUHuEdX1B7QskHYSZTBvDRS5zSlHpgnMuhVg3kQaRZX7u5Epl1u8AfCzEoLaZ5p/6S5NQBXRhRe
mm8nb3MwZk7r2yFD0g4v8D4kLOgvHhnB+C7rr5xZxglQ7NumCZSmEHKIzLlOmkhAh68xNt3AGrkL
edyNHF2mBIYWNUyG7mOJDgFvavIcxn8fgCFPJtRLVISHYSnRTNbK2JEMwjyHJxaXOH0AYBxVqzPx
SrTkxS9l6V4SOO7WFQigOtvLAcETK5mRHWOxMpEELG3NIIdLMhcvod6LO87fv067uP0y438d/CyV
bnGRAzeL5aU177HTBGg8YBaYZYjQ1YUAyw+hezWmk0x+CMMA1zDMqB3K/CggyxuJyYkbbXdsU84C
h16KqaTqXfw1qFKKNARWiQN0fSc83RbtAZEO5nUzd1KsJLu9JlkKpg0ZhHod0wIisVvqgyX4auYu
fstkFdiYMeTBxzaQcSr/aNnwK+RHTCyiM6iEOEPVjtRF8fk5+yqAq5hGT8wxnvcaWxpo5/hoagO8
BssaRD8hprdxSV+zOc1v4dX57jEL+rZr9TskOpLgzfvZwswzdpCMz9pbceZuq5PNe04FvvNk9F54
oSyjwjgloT1QUKhlP4JENCp5hg3g5aBppjj89ft3K7n6crA+83Ln8nnwiS6Je8oHNph9eeTWS7wv
vH5j7F0wvcwZ2OKesVsVBzL5r3VjPQpuERPemrHFaSttLTIeQYfUtAhFfu6SBQkny6c/mNiPiuxB
yNEttXAIIeBHmkJqjGYh6H3laHDlCJxMlUQNtE/zX27Y8dlChIkd1x72/igl+cUstd6WW1qjCACf
BxUCm3N9KyYO1xps5akPhRjArNm7iT9gf9g+nacEzqnyzMoVDR8+wmcIMAXAIwL6rQVG9xgDo1Ip
CxVzuEIL7z2o+lLd2/ylvStpT41P5zaNvjzsqWZw77ZyPBSDKpBVpjoHcXYpz39It2JTLaDKkJtg
7Py3hFTZ+LjCtC57iBUOgoxH0AmQNaKUU4j437JTqTOEJLyA3vwF3BjAbZ7msvzl95vebwfNOYtl
G118klRKMvw5k+EskHfMCWvpHBGTfqxi4Oh/Mld5dH9btlXIMoIn5h9uyTEMRVjHKFdk9so6J3xs
cFJwPGPvqcH8qK/Q3Wc7jLAOzi27tkRLWGL2b/cphI0DHZHpnLFYdGUAljPIEUb3BXZuL0HWGWAP
//5pOREmkz9VcQPj7SloX5M+2XvUukWkmA+vvi9t7FS+Z38kiiaeLamlEfamgYi8eWx9x1lByIAc
rS31omfanee17iStf2FlRx3XtuCZyZDt7lMf6yiDsNfNjORYFjfwXi3CmZDo4czPjGGI3F88QgA2
6uF45l7SMuK9lWb899iUQhyTCKaSRdXO01j6KZg7dWUjKCZKU/7vv4wmhvO+XddWcr6Y6Bcj5tqz
vYwgkwXzj1jXeifPMk9XDAlzpRUx1OwdxmvwkVhznuk9gow/81e+C77yaHnR+bsZCg8ucUF/k4yD
cRBgi1b7QImNeCiGVEi1uWLYPdVXifuaVcbfQFSJPE0cphMUEYDSGkSX2bGsDWmXKgI6Ufk9k56v
PFpj6ZtBLL3s2zEvCGEIJeD0Ntr1AhYK247/WFx7DlGiPvVNmpG4/trJDe8AE32kjXicdCK5SUrN
SiaLI9WP0L0jMkG1UjJdqzuQat8VbKFOB2YkKiEq16gwpO8DPhCvHxJDHjAHjuKhi6GVdyhlv1aG
4TBkeoZjXhrdFvRG6/1lj3tvBrgKM3832EKVvtR8rPGR5cyfT5/e4j+4sHarY9vYfhuTLr+2oeOL
VGbMfRgs8IOQBi7hdvcfjZvS1hjQ4ycvduXDky8ldReXPB7ELMeBPWj2HenKOzHJWxgozZfmCNWq
mUUn8LN3VfFJ4vDiwKKyvkmL0+ZwbXmc5g1zZk/KDSsoBhpXCiEmO1Q4joqnupzIDiAnHb7wZ7/N
/EKtzlkRZJ7oVzCeHrwoKPC4sErkT3LtLCbs/oaqhAYCZSK59r7qW9fP8oDpf4384Z3fWqy5edga
5DNbXTO9vXfgRv9FTerILTc6a4Ax+wRYMIWxK90mp81tjnzREHXIy0ocSJXH2bgsxySG5Xux7nf3
R7dX3pmUkrZcQ8SFxYDkBlNZ3lHbAROSJQOdF1xQi+PA26LCsykVL0DUHlV+RoN7Qtla0RDD7E2E
/fEPUXYdakTPq74q0Zg9w1fw0P57WWKNpL/XWM6yprzau6B4pxAV/jPk60AahKuKQgcjqO4QQHQS
U0qFiB2nFmx0bWkekVSXJvFTpuu2Qr1RmCezdnkOJIvu5dG3IuB/arMHOojQuENcXBF2hKhwOCjJ
NFudWOW7VEfr5orQq5IJzlCth6s7PEE+u9rtxNBFsRUEIBR92v6pS3+0V4xNTBobFMXi5vqWg9RG
kS8TrKCQXdHLNfTQJ6vHp8Tz+xHHiEA1noB/rQfUiUp33AABTjJgGeC8yPWapNtN4Y82BN0/afdu
PdbjLd3CksLw75EhB3bKLyqurL/6llBWk9gP8r9LWxj8y6eFOtrd9i2YNABcTYke7Sg9cUWjguFo
T7uhOTyo/8P9LF6V++vqs/16k/CD8tX+kEGfqOEWwnFhh+r8wmlqjxjHQ727HzGNd7wAGLeQjzX3
5+jugjUr8aJnb1nNJ0mv5UvprmfJ/lYJ0u8aq+IPxQFq2akf5jamme/nxdH65nhGsbh4hdebbvFL
x6077nx8KQpKlAxHWdtWjqiFGT+b01xrzU0vNcFXMuAhl+AXZhxYXN6QtloHwS+HWXKw+iCQGYNW
/rFqZ39WcdgeP4m293MdfzbRcmMkkival4ZhxQ6ri66+IaB7MXH8+YFMvdX23MSQ1xTRI8J/u2IY
T6d44WngnYnReeqvD8KSkNpyGFTbWFuVZYygYCiTlgrlqcYdkXpBrPoPfVhMIsq4h2VUxBRS+jGs
dWs+VZiPQQiUFzLnagLnieuCA2jwCrnI898sWikPSXcVZtpyjWcZjTAJFTQ/uMtu6JJ+F0OtjZIf
LohLDWlg48lSvTGO13JMlfe7p/qsv5N0a1j/YbglQ5JFyeh7Ka+ONYFiPOaOUlVkgvqIFTE78a1r
1EucX6x7uPi/y5L4k7H5rt8cJTf15uI+Kcu3Yy4XyQX0cJ6lXiEXGgsJ0kceDbu/tKrOiyn/JZWt
2rPk8dXrTRBhPDK1tG6cNFPaQ74TzMUHXwThcYUZ3vvJHZLRYKC1wA6S2BDKcOCj1FTZfGwC+qkp
xERrwGQ+bchMAsAGVY5HpOnpi2bVWj/4hiTVK/nkO9tRFaDCWDsoUMMA5oLIT5WvcitdsLuvgCI7
XGWJKRBqDecvvoLanN15S9fdnbLXICkkBU5GcgYTL9ZrdWlgv497LqGL1KVlvQBrXZGvg72czO/R
Sz5mAbRtk931OBJNeMx7kifOWJrBwpi+5P3oXwnsIlDL6SHoI+y/b272bx3IIGmwPu1NWIt3o1bh
9Qtj5msaCrYS8LZf/kgh/5b3eojxMybv/dXoJ16/xnX8+aCFPd949G5jhFCAqhUYWF8IRYb76qbb
sIwliakW+Kx5iUK6CJlwpxmW+zRvmruop8nwtkoFXrSoDDQRMOtdmOgMTzk94pbqFlvPP0Hf+s+h
ttjPpJ2Jz/WVbbIsCBKeqdQ+qIBBqu1Rg9fBPWtcpJDZ1VIqf4PB5t9QdW4M1gnbhQdF2J0nfCHJ
8poLQ/yxX282Xms6uT5YsaDkvR2zZnNAVtzJqmWdV1/R2/5elgrriXEAM/4aBkTNN9TuEcqVvpRl
kN5Ici+f4fhovn5er91sarlpvIk5R4Cg52Szalfi6A2J5Fo5fCVtf9dVACjxszWyIuLeIxpLYSyg
0P4IJ4tvomGmLL7IlYB0LhjneGtvZjlqpv6cCyr4f4BvtOhA99AUWzvtmPBoXVlXhejaoaCf4tsf
8feGSU1SUWHAOSiNs+mefJXTotfJzsTpmTBAHNG9MTeito0QLDtSpz05xS85irCgyodeDjvcgF3C
c6Vf+BuoThr7t+kkew98wmGKFjRREdi5tKHEWKTlyrh9EmmTmEJZNabpi/Ca2RE3Wlq+vjxavNRv
XJfH+BLGgE2zYBPdu1mFm866OFzI5yxqquQ4trqgcpqHXrpTO0D/PU21MYGjLzcKdJZR6fxTd+Hg
0PiqJaFEaRk8iJdE66S9hpwiINX8BHm9Uhvc18/aiis4gr6sTVXuKLcg1OznH9jdkTL0iJhBk5kj
GWlt73dP7/RPmfWhXG6i+zSC2bLgNxptHJjLQygzvHCWtdupgR5iFZdzPWv3E11QOWrWRjlbsW43
ZU52TD9U8jSgbu7BZuVkXefUF0r1oQkj2/NuD+Y+9/M7gGWmehq0yBchm10loq2ewM1wB0iPNkrz
4F4IBwB7YERTLsXNBR1tf94kJUhIzJChoS6+hmOddJwfgyLvikFUJSsDnvSHyHxUwA6wJlwo1Doi
xsNNwP/5Ns+d1yUpuClhlDZCArEZOgZEIySSaMAGCbXQxqTFfEjZM4brrIxZv4MiDdzVVaOfvxcm
vQP8MFLxL/C6kYxBnFgVDH5WRdmRA5lXeBqfZOLtZwA8/gZFmKR3eiA3odnMbqfIjMQvVBKB9/X/
eLr/ofVqcNiE6HCsZC2eDzQB+xRwi5zECJyIeyaCm/AtsyavFzrm2vARvLsmbmtKtlBrMEGjCZTD
sxM5O5W6AA9odymTuROHZXLjXErixzHLN6WW58swrxdFYglEIEvF5RkGj+kcEwUBq5p4VjfChvxg
yA9SPGvJ4gvNFXEdlTGcl6VuJTyNVIfJQ264oOILzjnyGY09WZXrcpvjlrIVyL9pslePEzRsz35w
MxfBQwElOMyJovUVWojJAmsMRbNJ5+06u9Kwal6wL3b3dHip94vucXdN2rRbEm14Lf8HuCLViOIf
IunYPOMLTGrv3qvK10o/m2HPG0TODzU8amkz7OBax6OPemnl8ZA0cjYtvtl1zphSoNI0eBel0w/O
ON3hwD8qwbggWeU+bGMNmdU1kkKcGGwXp5eXgtYy3Ll/0ek/7kNU1ZdJTBgGA2HrUg3uBtVdITqi
7Iaey4tOdUiZHmirrOcZlPRnQNZFggz4z+uLenFsbKo4B6qbC2+rksG4hEAYdFn9TNV78g64Vour
b4Xf0LxtG9CuWGP3VHkOaqsZkDAWE7sYf1iVS7LuH2fta1oIfz2JbUHeXRIlGNlMsuFK+WENSSKn
Yy/CweZpQ+8gfY8SinmwnnK8ouDGInvEvIhgyrvgpDZ+BwMpUwSK2MHB76FKkQ+9p6GOP4XK7GQr
H0uRt+ksmsQG8KINh1N7vdigzibyJFvdbjHPqq5qC5Vr8gDB8/3dvGPH01cKzw59ugWn4P08d5SS
Yxn2hOuerZSoj7MRpvdK9RMhwzYRD7VRRYGE/14KOcAWESqd3IzMdQhCOweNXmkTqL4lcT0V/b+r
XM+qLHc9UhmqNz7MOjNs3G/LBX2M7w3ADik1qBqOZe4t/ZKRFaB6Nl1z5WTT5/dR4Tsa7Tr78OjZ
UgQTIJQJwQo7I3qI70l9hEMpwmWZbIEayy27gI6vGbd7515ReiWRaskJoRbGsO6dvGXaV99B7YNh
m5I3ZePJh6COKsF7kaPl7xcrEj+PZrYl+qlgDvCl4EhYeiJgxUEFx/gBUhjZSIs75fksshKcUB06
s7ZoBi6w/2AHfL4DXAK+HXr/fhScViCh3aEHdm3Tv+Jsd8UeWvqSDtR0ZOuZDC04JdWPTfIK2qLw
ZmbxN2oQKVnsaI5/VwziTwWG/v/6tIKX8Ze+/bpaESwZd4QnRF4AIWb/fgx0VHvqs3Zd8n3HQMrM
BcAJhri3QO0IaTuZkfcOwD5f1KAtb/U6vlpHi+AfIoQU3Vh93t/kPFhlMPrtxQcw2H5g4pGy4hLY
hSiuVPjdmNiGvZKAH6lh87iFNjeyBPB4dh/KeHj7bZM6bY+hQp7472cI2YsyMXLQ8QFBsnqxCfHR
O34ukvMzlIaGunO6u0sOfJP0qsKqJETq+b2LPqjV3SQDNq4dzCHspQcRf3lxMm31vj+/H/K1sVyu
DOSdzs9JIxVrXodA+XrmZF+MqH5lqb8bmonIfFf1Yf0eA4QB2zZAupMkDfdNcckQGgKAm+YnKcJM
j9OG33nS4WDIl1isVNwcxXQeAqS7F2kQdv3tC9XsKaFZFz47L3FBg6qK9LGmr7FDlz2eJPt7DQDP
MCH7z205gu9XRS5jUR6XcPgHPSYXzjXFgJDkgAKk09gmVFOA0CrPlaiTmqDlQR+uA4gmQ8+O8WzF
e8r8aOeE0F2ECWEMalHWBMO4Z2zKMuVEpvxIJIxob6RLo94/2AMTf0rWbkBIjfP1BUMTm05wRllb
TtuTSkzuXvVRs5+GJ3sOgLmwcLE7cS16eOrn+kQ3GeoGG0YxuoH2R9YJ1/iosvL0BaxDSzjEkJv5
ietW6BE6e7aCFQl2LMn46DZfEIaxUCdYnlwhtH58iZAEQ4HG9X6q9hazhIp97eZCRIDPQM7zCQMb
t9vaQCzzkz4ObGB8yGHcESbN6+ch1DN0rv8ajgfnMc3AYpowUDVlVbh27r4d0a3dtIzfL9LebuH5
lp2HpMir+vodXXOkcX110ApDzZUvNnIS0u0MY4aRvkNzGftqRzfxmImB25OjDe/Yh3cMp77yLQYI
yfqF22u2sM4rmmZF6lFe8qad0OHDk9fH+lvLgXPcaPr0mNnfyVw/obyU9UWOHttNYf9v55ZL4LBj
O/LXeesGj1EnLg86E+/hesL5Wkg/53pp70TvUC+gz2Tu/r+ELEbGYjWwuZZOmFKdcr1lodzhLLhT
1ih0KnyXg26fXVp6467PHFxi5qVc9FD/rJ2d3ajWqCefiIc3eVHyf4erOAgWpTpuZ1mEYdP7T+1Z
bt3ez+UsjRsQGea2X7e3l8pCo3uPWcf7VGt0ekuk/j/wIhrWVcAo1c+UjvrQiiXTE4wGd/zT8aFv
oyhB6fzWWjghRdQEtTD4BMyY0V988F6J5zpzT15pOCVVRrAdwBBLMfDXwPlapeUj/hNeQBJ8zIhK
JGKK8GgsSIJSr9jnTtKPRgF945l1R2VyVYOX3FuXyjQ5+5KrzkDQ1Qg/Idb0Y3hSwnoZOeyNosFD
NJhrOCEI3/jRWffkj5Dm8ANkcLz8IDiL+LCzwtjiqVA8DtzTPZV+ugp4GvvxsReZadpWKi/dvREh
Qa4yikJDFQ7jZNYZ9D7rnA9aFyMGbJDzo1Gbh3OjJGnF9tz3fQF6+o+GKbRU9PftTQg2DvIDsYME
Hj5aJY8Jg6MVnndYSxQHkKzAAYRHQtLUD+JYyiQr66B9DlNMwIvzi2rEPvBeMnqN75zYZdCrd4ee
mOhLc+hMVQEFbvm58vWijVxw2yok2t+xGfQTe4Dis+WTmD1orAejlwU+Ps1cxlniwV/IlMJtua+d
gKhFdDv8H+By+fsqRRiXjpCOtF4IZVyrOXlazoW0Y8xM0HQbDaO9G/zuiLLpZs0B/fJVyeRpWAGB
BIsbolf52WVIJAmkw/X3qVguBbmgOD4elnB8uPn2E3aKPzhOPvD+vRhi35ot6nhNGOpQ8VXsb3WJ
r/aOSkMB771F166T8oinCSqxZdC8qwnsZhGhWAaIUO2FXJj75RrtgzgRW+ethh8OiXFbRYKO+TSf
2/ySIQyQTUGmi9GeOJfBK4Yw77U8o3smwWnhfxXils740i4bIERmWe2jl5VQLCJOXrnEFgU9LLmn
2tGvqI1PtMQWYpjHsPUjUCrpbTjvgsF202B6PVeci0GPe1YCluOOheWrtvr1Z2OwT3vG1w+di+IS
6RWvwwq8VUiC6qvaa5Sp12VyusTmZv1lTffefCVXM9KDYiQCNTofFq+3Bz0Q4VaEjRRPIi3stdkg
UvpP0l9pukE3JDzEwZYZThcXcyvWYOW7iLO0VHXZaInuZYqDYawE2BCFMdCC9P86QV7bNdT1TL5W
sK1mHm1gOyo344+PGFlRA9cexAHx5jY3IVu3sKOk3S6WUSurTaJkfcq6w5Rx1L3nNtCW0oFGpgCC
BZk0LavdXJTXY6GlXUYxALFtvRxE5FE2e6nuZNbTUbrvmkYqjXDkAeFcsyaEWMng+hfUnBADF1Gi
czNpC4ejW50towmj0SqRsmYFfCHWRn9Qk02Snk9pP2TmifzDZ4AdOFl7F7qO3QEp5fJsmjCnp/4/
BXmegTjE71Lu9W2JxWoTfnNPVRL+wRZo/vSlatD061+DoKk8uFWUjZbV6kKmC2Az2HYtw1l2rJCe
lW1blmeX3SWgw+TRHy3m71EE+Sk7wkVWCry+jF6K071hnIWu0cG6hjwCRGQiGlrXsF3uTJxlkfVO
Gu5xDztSo+6aQdbe2ovnABP1tFJmYtglmf/vbouVEe8ltLINNT3elYDLXqM6laf06/3+QyUyqqUY
YZehO1xCw0tMVSEx3RTHKLpiUUfz0yBB/ig0bEvqvBlztBc0gPIaP6McG5ebSgtJldoSf/E/hJs9
TqZK/e03qx1bqjaCc/PWcqS+oil5LKjr2I4VbW2J89HOuXHKZX3tAt8j0Hl0ZkKAVfo1bPfwsi5C
PTcx9EbZ8X6iINiXkzKJsmq3+T9hXmqBr4+m6HOCh4odSke2YF2WGRq4ajVN0pmgxCgSeDNaJZHS
OYF7dAoHc/R3jCusOUDyuAJ/5eGbkgvzTGxRNBJTqDING1hn2RN0fcYnw+DuPKQPKuUnzME7OpL0
koiY8ek9IaAyVYFvCTEo/7KFQIo77MKuBlvdPYcAg5+XguX3axrspv4Cy51NCWLDDibUa/Fr4XcO
ltOdwOB5o+TFnyoEXFpLv11CBI2QW4poUqhdq/qiN7hqhRBysF0fCC6C/cfypG8aAe7usrrJaOuP
o+4A5hjmB5wHF4siCUpQ5djgrldoFGK9w0nDubv2n53AWWFoC4H0llpaeDgdkWO7TYRXCCm+jJU4
EJ+PL35LtJd7Vez7TWlcC9yKaNR/x5aIfouelp6zzLEBs3jNyS6FxalN3fT1bo607xMeO/2debiB
FR07pJ0HZdeWq3lUgUOzOwojwMM3nxdZlpAD7yd/pslkOJA3OEF/6qCS8T7xR52rXqK3bjssF1AT
lsD+LkRGFfc9IY+93wY9xH+hjAjTLhECRKDqbfYQPr2y6+b1UXmj/ZNSElzOGj3O1qsygh51Hy1j
cxcgt7bw2v/7JD/WiN2PQ9G81Tx4E0+5Ruyd1Sh7PuSywcn7NibmtYha+1DTvEmws+o5oc/ciPxu
kQzMPw3XMZwXPTa1P59S8SSGtC3Z/LmwAxwTEVIaJWM1EfTcg8m5K56sq+BFcjxOrXseDKrIIwV0
ZZhv1SWmN1Csnwj61zxcx7r3ButrFC0ujYA4BCTF2aQAk3ELPR2rj5zFP5pBBing3fNlkcbU7Mzt
Dewb37icsVcDoY97k53vzQ7GtuPJy/bnxAblAoJpoEhUtFf9qDrYo2kGx8P+3meSr622/ltFaqC+
mfPHMpg9ZuooKnb1M8StIgScL9qeZW3aAoLwk+z7K+gAp1ZAltEEMXGpLR+HGNhNISUo6PjDq67v
Px8UTL2NjKZMsONX2qHO87/1G5XdmOdflV7tdn26lr+E7g9jgBzRoFYS1728pRqy7/+kl+Se338R
RXCjV3TRp+OLTwZt5fVtoSB6G26PVDX+tCM6w2wNwgD0kCj2KJENljWqHWS4/NPlDFD6SIu9PGZz
iYSMzenJ+MX6wWSRgbGrHl8ieGxJwGkAuZiNiQ4MVDuEqDnX7y1gtJ9psrA3wwiU2KCMPhNR710w
wCfXfMxUiCnEgf5VEmAoKm8nQ9vNcM+xW5aGRtKj9teaZQ/dFxQ1uZu85Wh8uVhBbRQwRVXk10+m
H+q+WJ7y/mlUOUqirsn7LFFnh40OUE/emMRPdd6iRqYFdblQYEAu4ri0vkfycVoCCsSfskyM9JUE
Q8JDErIFvnEHsUXW9C8wZ6hmZqFGJKgZPDPNBLHh4QIxki0ghkpmJlYn3FqGltMdIX6lhaDBmdRi
ou6/E/GXrLJwVrrttP4X+mcH/mf7GQs7MGgEz6s7bJLgUa1Nr52IMxsdmcTE0ZfEhp5WbfA+PwZv
dxFu2mMXRWDSyzCLnxNhf9tlZW5YDCu9iJHuCKrr7pmI6CxebgvNaoeurCS96zkVFmb5YVl20lpY
4KLA29LgaJhAyU1C+RYUXpuSIOJs/JACXukwnh/0XgaLN6EaH4oHq5eKxsZNQDGM1OI/Hmszmu+O
obxwZtIcQyNvCCleo85DiiIx5Z6Ot3OLHUUPYB5LEeR6BmBBLvtXTPmhmmpnpnPylTVpBaMTtZkO
LHmNSBjivbOs9wZdQPPVy/CCMDEQ6EnlbjFWXEsFKTsWiByYwbvIBPtrFitkFoUytEFyCeaaTrJN
RWZFU8zsxed6Ewk63SruLjSDh4ZY37VkHBEnCrdvUNz24wxyUJmf1H7u3T5xq9itivBgIJ9bCR55
4jv6YJttE4Ny+iimvnT5/6XSQ2/rfOxz0X5+gyu3Vek5fHKN0BCJhWqke255TW6RuJlr5h7JBQW3
j9xdXhOV+6VbYpsmfEWHGQ2FI3AJFLs+gLMDT9fVj8ZrQo1IC7Ar+lnitKaP6TS5eaBY6rdWUsMp
e7Tlr4o7vHkPlP3KkfUNwJjcdccmuwt4/lQJ1uXwTQUKdrtN7Se+yYM0p8KmLRgbYJwhJcekwG71
vj0lGd7/yApcVVHen4adBty2ozD532tBxF1+ybczOzaRRhLqPkdf4MCajS/FaHKVPBUHbr7sNqKt
91zQphBjqalhOscjVVxj+wu6yLanWlR8hJzlVqJgpUpQmeULgZfORmwITEbuVOd3f3lBUOd2+zW1
0+0qo+CXAyqEzJdDQ9O6ndIqIktQ9P5IiVOMm9feQQMykEixHt0a3T6spej3jAvlfIhxE3pMsfIr
7wAaU+sf4R/5rGhub7efXcbQA1S7k6rBNrZB+XFPLHou5GMR3ss7q7ubEniHMQwYc6WSFVXEpL8B
U1WT9KDngr1I+dQhwMnHW0cbi6KYPAa1AFShCvTFT95cjm4M4DiHDVLkz24FUr25gLB45C3gGshU
jX1aJ/wZlGq9DePp6AcqHk9JJ6eJcPoYso0wRI38Mtekm3L/ukcOohdFU6bk3Ozzheb7oSCL39z/
r0zccnLsGxEzunVzsiVNWaxMDf0oMsAaCoEhE/Y7OyqSk3e31Ghzwep9BvvradhxCznX++Xd20Nh
KIshjjN1j0satzGUURquGX4VwbZlI0epHVyPzUvicMN4n5/kbeLLjbHyPTrRDLnnXzLytL2GoUhf
k+nXylHgrigLRiMfDiBBP60jwbEG1iUVXeZKEPtborln7rZPwLiLz7ZAwE8+XkvJ6rkCYIrysITU
BUd/kTJl0HAcVBv6kH9SWEOoWDKxnsVh5b8Exg4L/3ORbgCAR3vEeN1c+1FEWW7vGzaSgDN/5ifD
mk/wUKBN8Vl7WRHwyQCfrRZZXXPHoQ5/vAFf31recLvEIFig63t8ho7Qj0C2+bsyPjQfe+eE5sF/
xnQsON9gkNipSR1aXYrCklRMfSEZFo9f8dmXA3REq5oCBl+OjrkUpsPxH5o/7MvvaQoF9zlOt4ow
nvlJjeQ11dOFu8wYPZQvVwkV8Ma5SHRxdwspTN7oQZyO3UI+ADDyqWTeSl0/cAScMUA/obc1eNv5
YzbcHccQg9lkLf4JW6v5fWurQO4XCdyG3hSefVHVGopJKHnNitMPBxd3lEcQx+Nl3iCi8PNBDQ4S
YwV0jmGTzWeRn8rmIZvvt+8FLQA02MIhLf2MUGt7lSsxq64W5e3aL7pItBCyoQBk42pjSkSh+IKz
ot4JrqxVN6lwCVBXVnuJGnCG3l8CI0B1ZBzvezHhjbwy6ZyxoNpRjKm1ud0QDJPY+/hyYjZo5M0V
bPmDfeEfX8K//0H+T6lAp72KyGkazsnkC0J4Bbtx8RxkytSkVFZeoFqbBgv02pFa8Vy5ezkwQjCI
qHEcznDZLJ3WPUQs/JcChiHAMadjQt+c07ITXdDn0FtSNTFtTBhRgyRo4TNMnkbCO4/5xv7rxF5O
2rjh9kjlOlxjJAU6W9EbiJNmB/8ec+MXv5b+4vGW20lmyjsyNg0TZt9PikX/QLCpQp/N61rCfw5C
H2m9Kaw5/4BrC3leHE0WdWRXAnNYHfxtFclK2OHmK0YcWgrODbyoDzs4Z/VCnFeX6UDgSfJrrxZW
FzXhb3z8CAD/w4nOEmA1AGanVsk+d+BLANSHz0By+47cPelag0SqNjHye2YQ5FAo3b6cX3G/hgbZ
NGRUnZeHzTdXRyuaDast/omgOJaPO54bJWUeaS2Qh18IERRRBLi/l/evoJJNduqnxldk/6a6wQ3I
9GJgSnyT7uMs/MNQfRK2P0Wc8QAU4Ap6e5Otd8vobXReU90VpGFBWD3sj322aKpkk7eVzoq7vTAD
T4ngDTvuClL6gwVFAOOMjcnIjsItf649UxrJF7R/4EGHMBk+JwwyhCZjtScPcNHzbHTE2rK5E3pQ
CK1QNgVb9OoucC0BhXruwVJfxBjbFpxbm0yEDQNKD1uz7Pjk3FbzQ1PdEq2t2X7fOyNQpcyMsi1R
QIbExNzsp42wvsjrE0x/YO+lw7H7mMjibwfulEa6SJd+6wNH6Ue1pgQKn218gaWpeYoo5M9cAOVg
bIQIzvLmBmzrSzlXnGBfAMTMCnyOw4IGA5hUuCnhmooGOW07722Cx/KlTMHoFk6+2e319CfXNqhw
rxxtP/e7806QGtOCCx+TGEL3gPNSkYH7l/M0+81Udzyu1eeN6NdCCyuuuLbv5hl3WwLAnTNzs/VN
BEaZ40w6O91I+UxtUx+sjVf3Gj8MufRwWA9Exxreg2H3xKWwTg4jSeUEELncJ39ksPzHr1/sKP4o
IJ31vqp46PdDJe1GBwMeh8/v7ZUVIZP2gsaPbATIhQonKazOvND5qm39mpIbi1vPrzmCYF6SPjcf
0WfW3JymKws5wggQjr2F9/cHOPXrc5Cnu3tc3ZTuU9puG4zKWBOjPuBzpioA+cfSLEuje6tLgQ6R
h4evMzW/q6YPt2SfwiK/Q48YIHeGcROZ3mGmHDlvyHXGExaKiKQy7rSkdx6adeslyiyOjfguM312
vXAk3imeA6qDAkFFISo9Fzem5sYYGZa36V4eEs0Jc6dtQzW/hoxd6vvPtnIm1Wy/yssC7UPJFEG8
1FUT9P29khuANZLTdc12kYnSTi9hj/JUzG5HonCY1aDp2UPcOsQC37eEEcrNqHHnH/OQRZTO53Op
nw9HgkYC9ER/9uZ0YhnItpKiNknw++Ie8yJXLvifBCaYB+t2l8gU0VNT6aY7VbQaM1OUmuU9INOY
XyS1ag+KQOWhCDSeFi8ILe+Kh5vlJtl6ojApiBpWfLG96cZjF3JNn7DBSrvd0Tv4bQD4ru5+kIyL
pASb+8kQsAcUZVzJvsbMDozcDqxtPQqVk2pelbgcd+FFYx1jUzq7g7Ue1yDNi+zANzDwNVKcGBd5
ImoHVnzs14y/Hs+x4sIeSsBhS0sRlXlyLMOFOcoJwx+mQss0nrvB3ZIhCGFAD08BHTk1qIch4a3I
gVgo8aHkicGybxa41fRg8/fZ5uZnPRcOJ17xPRnQRjHQTXvSjr7tGPCSLaQqf6sLuICc4XRKG99P
DcMb2sJiw1ZA7cSCNYAevqxV2AOJylq9mVLPPUWxt+wvcwcrmhEbG1M9E9y1aLBY1rJLxOSt3QPA
MxyUOKVO8HLIhSWN2znK2Y8z5d46eT6Kl7uBSsl4jupREKYZ4lo2OPRymMQukcgOQVodr/oEs+lI
YVpUMfR2OLIRUv+1X45CF3ULtGKBvkkhuEs5Sw24rkvFiGXDorsOf4tSjoZqqsujUtWcm1xsVj/N
vAOQm2+ezweMaHdpJcrSQNrZVFgWZj6mJxRDFLmqlVxaDZ8afduSvOzsL5hAurG+ZkIrWmMsBCfx
mI6yEoFfnUfSQWVFYW0yzwPfQ5d+dYM0iUGwVa4/sS49LLedWDrGswzVjk+CC5Oq0SInHNZ4ibDy
+CPRPUQA5WGh/aFdK+L86Cz3jitDzgVFoL/KP+LBf5/2V73uIbcD6Xs3OPk/skJ3P67S724JdNcE
gc3mupgfQmFzOQLIAWPi4rO1dXuFeiUTXrDxHhear7wAQBJbDiPo6bAsEIdOgZkF+icNOjoxXlWy
UH4unaw1hCDOJl/LKwzaD9dQkQjmJPo5zJDqUuft3xz7x7zODxk+pA8ZK7Z8yfd6M3LUcWmTTvMZ
/FWrW5RfhmzUoZlG3e5naSvzKWF6xVzaMV5ALgqYA8/ilAxbWH9dwpwk2rb95GWAR6QeE2xYiGA5
4B36WU0HbAny1axP8J/ePjvhPbYfaq772VuohA3kifUN9WcAeFyZhdo0Y9FNLjfrGRQCVNexAaXm
9yqFUWSU5b//+TQZj0LZRsaNxyBaLTh6S/dMTcsfzxM3FhdUv6pWMW8epEot3eSzFaRuXB7pj4Rh
nzcK+MvKPeXriHW1X1qFjRNlbwmh5mYjmyJh/oR+sXbaonutOUvLoSX4VnIw6STLoZ7pBl5/cmV9
B2br/4X6uhNPVb662+EqfcF7VnPWWAVZh+Xvd4U5K81u5PQk+gGoyk7pzmpn4jXShGJ6ansVaOCy
nwhq1ch6ZEjvgEANUw+hdBgaI4Z7P5MPVFY+JRjZ8fCEqkiXIU4BjU5gt5kYfqP0BsQ+ntWWYMYM
xNAgx0dbLdSNm9aElrURVcL+VIcODTq0/2O0JiCwIcSSkhi++RnILEZ9n3hrUJ2OXZpJwnZNJ03C
NgsC19nicg60VCzwa/b3MxCNa1ZhSrRIZtSmSLVszMy+HLkX85wU/udLD/KXd8bK9nYHbxWnCdkY
d1mJnfclIwxASCjHbVhRptvW5Lunf+J5mv+acfnziWdD/TZPXGTysiJxwC9Zy1P++daEyoCTsV1R
6viHyLWfLVBYwGMjNik1SmOE9idMMJs7ADHmMKWNDp1wp3Vx8qIBlqoa7RW/3v01BqcUQfAB6dDE
kjNb7fC9jawYxUpppawjC1Duok7icXFlELVGDGlOQ/VPbIpN0kIVAmD2+XnTvlshkZoHYCFE6q5p
N83S+fDabQ/yW+CUTZfKXkrofHx4s9nkecMvSS3vLNDRXuq5xgES/+61QpChKD87h4aSrhuhXRbK
TrmYYkOJU7+3EmmO+9B4vy4tccJSd79iy7UOWawZCUOWrwTKXTX0iB9q7Y+KTZilSW0M8N9Ft7av
gdC86f3ioIbw65550SIPNIqz8i2W6pobRJ7Czkd77j7k2jTRBssEg2l5VP6468pEyah6QitSCo66
PyB3+J1wq3uEgAZICaIyiMQy8QkcNIzzDuFqVCCG+1WctC3DdeKI8LcKGnWmf1jm8K+FA3Ul9MQx
xW/kqSO+9rh8fqFFGhBSiCtvrg2UiOAvn4sKLbF0UynM8ZaPdtvXzswZs4R8q5/Ncp2ZlOMofpuA
jhQhWkJQdz6BYKaz1WOMFK/t9XP5IpAmjtL7CcuSAJEOsHqVN2B6grPA8sMVark4/h46hl9wdfUU
Uqb60XU1pgqznLcV6PibPiz8o0zWS1Awm/3At5ReMmeu9eRotPt5SiuhWDAlZqHe1AH4I+U5ztXU
wiXZOD5rq4GgbeLyTbCZX980semPcRbX5/X8KH5ZWBv70qTG2zz1LiH3ZGRiuY6SRi7tOWLe+qbC
Dtl+cfn8drDrID088EasZYSculZRrErFirSC03bsUYC+cItHlZUzdgVbsE3FJ3LQOewuWMOvH+aI
Hgu4wHMheIzbV9TCjqgT94SUF5/+w3mUeeKv3LnrDu1rj+qKx57ikxIAN7qyNbcbQr7AxqtsuZSJ
ni6AqXn3A3XLmCzRzWaU2zagHUkneSoNNAWk2lL2U7ZVWnpD4S2gA6t8xTVztXYN8CrE3d/XZ6Wc
/JTPK5cuTSfFzwxg66Y/r0geM/6MOUnRbmrBiCf1O8vQgluNG+J6Z88FsD1orLKGuY1sevUurrNW
KvY/CEKQBu5XrbJUc336rJ/fUFPE2Ci2Odrp3Hv78+6e5zgja/mQrbXAVfiSOh+xR1AluA5eA4r1
jrXT1/CZa7cJthgA7QyNnV6JOk6jpGZ1Ht0pLfp/YBb/GljHvteLfRf9cFw7iFsQY0oBbL/vYJHz
CbFxEDayZ+ogBigeROCTZd5M20uKBLOqyypzSHvBrEjFQqMHLUPw72OxMnN0t7ml/j3KYWXxYr1/
I3ex6xEILnqS1hoZ70hPQZPSZ26+uKaH8GnL2lvPJCUUz1l+9mZJpurKp6a4IvIx4dVdD+B5waOe
+z28SjHZHFzVoKTugA1Oke3D0zi0rvStycOJvpdPvJeZHysH2d9OX9IuPZzVgtkpfkf0l68WVMi7
sLeD6G94ENLi/fsN0U0WPAZKl6VfFEjpdxryVI269EHE+GGgqsLC55+6tfdxz2M9zmQi8EMg8iZ0
4jRDlWW03N+yfSDnThMut3vg7ebl3J9kOAl+5ZVukhZ7kZUc3loUf7QpYglxzCL725hIlIDfMXNn
C2wqdzNSa977dgXwcww2S8wr3EZObIH1VBV/tZM+2+lg/uJJ/+rWN7zCXdve/d2PnsB2UoDQwQdY
ulKmJtj88IG3ifltTU5fadaEfwaHkIYCeQ7lHTPE/5iEzBw6X4Iw5n1/gi5ktu28WYLIUn+7k7ya
qy/9ZYeoXATksH7dPNHlTt/nfYZLTdhe0IINZvFe0MFsPhjl7pJMdCTtlP0vCWZJ0+no0Ydh2RmM
EsrSpk21LkCWVsscTX7efiExOKzTyEpxZccvGyNM+J88jPJNAvpch+SHh9+gGWsDxWC3ee0Vd8Lv
UUBIIi47/+ZpvKDeNwlWUhE7zZxGLxl+adM5y2K9UtkYdOe4O3f89t3o40ZyRzlF7Nu1yENbMn+M
MeHMOKKE5XFegD26r9XY6j1ZLECDgJ542BuOenNccYf2mvtLzdcIMYteCcYQ6IFtDcJDtkWs/7nY
DnIQj2sMnVSJJaHxH+IorJvy8XbO5RPfKU6aoPGz/R2eAbEjRksM8ZH3bJ4R86MFGYheD72UA0yA
Jj4GogmqSYl1OR84gR9MC5Ch8thYgNS/Awmd93hEJlGR/xk/KDZ2wXYnbwKDe4j4JNzGEfxJisF7
F/TTJp62AchAz6RvViJzbMg8GsMrrOD/YnIuUpoYynIJ1poFqmVzgZKrxeuzH+zYBkCBG974xUnw
A3H9HUa76UZPMuvZvTjoZhnRZoma6+PiQVPDvCmNChWZt8DFL3KsMbedQdmiO5zQcmeEPznrYwZ4
VUoDLzzotK3hZYYNqg1QSFpHyvyVPvbqLn6enibqhlXUov7VZC556GIeyXsLm4DN9i4do0NO+eNz
KQEIGJ4YCS4LhBCealF61JOYEnAiayAt5G4ziwzmPT0uzZh8rFILU1tyvbzQJmQpZ3Eug2H+VeNX
+eS+JWeEJfUSG5j0gHSRwtUrBS5t6fKySVgpDRRHr8Lw0FtHb5nBT6Q5yNCDjANHwakWoZHPJaL7
6yaZhRrvFL7E1jfJpUYdIiDu6ji9+G9lzqud7C077Ef7Gm2SX1Hoj7dUI5/TPojJgRt7/pdkBkTK
EDfB00NSBH+e2wmMpwL+AcIpUoFJT/YlNR5FKrEH6+u9N5dpAMZLD19/A6f29B/Oy7iYIJkBdeu3
b/Cf9y5FSzI3tKez+ptFHzr3zK02ao4SGONDE/VilcU2HOL32qMJ2pXEygsn1TvTm+awokSExdQj
BZ+4/XUyrP/uw1ht3bWMigxUDQI/NwWiXlxVfgKKnAOoPm+ZwAa97jzvvbJqeA916UIcgh2YzE9V
aq3+G1wfQT+gYQIbycXJJRqbc1WHBu9WI5Y6QL3flSuln0yzUuNT+HqIb6NsUo/cYt/b6jqstfas
8mgis/hcdhr8vQV94lQrXRNnf2GzSKZNUK8e4n34xUli6LHcSTochQlP8rMEEZtaCx0ODZUzeUNH
XOQnfdQa0B0BaYdYO+AGJnjy/R5TxZhmR3XAYzvraaxT0ByYrYptkXrcPVnyzOQ+Xgm4BI9iG/F9
fTBk1zE8s1XTTnl52b9WCOWORzFLLlC6+i7DNNQJ//+fFlzfj4X9EDxtHhzThtZDhDjXfk1euzdt
6b4YVtzoALgc/iIgj/iXkK4M+Pq8NkwOwAkRRAkZJ9cS/Ow9FwkeCReR1gw+ndV8Wz3mEO0+dJtk
I1sKb4L8yfvvdxjUD6XLP2A18jADjSlfOQmq/FLcKTyykchqoiwAq10WifF1y2NlWriM7TWtDgXv
4IV9YpaD+HbwTokvGHlpZ645MvjjUHqDhUq9yX6jQyGiEDaPQX3NinWQgpZxJZQhRS4luMI2WXcr
V5BHHaa48aWTTygAD4xZ8hXgaqzzRbwL/EJfDOvo5O3nGc1o/iWPh6dd6h2kKaBh22ONykWT7Ekd
fbf8Nk00aIZp4IDy44NzcsVEgweIkoVS7zZBQNC1SkRDWMrx0LLjTCGaKs3p4QZVexpiKYLziWjR
62azdfTbca3cs+DROLiCzGHq/uk3oVWH3gbxe6qvDiPa/nr2vvX5BdItl/nmNFG4E5CDpkRaRq3q
vNfkMsFi6+UVxmYL14yHoXbJ4JzSzE1orBc63UKp+sDgmUontbu22opRVFqwOe09bYoxrd7FUu5a
4BoSp+GHVjhAyXzh1DKZxgDpCl2q9JItk0WL5eaiXWtXG0S7ueoGQz1YNmzsnrSQKcmxfE0nGrEg
BDHWBK9wTt/VEzCbDxhSzbwZzhPDQOm3XMGSN6d1T3qhgq4XZw3+mn0P4WcKzTgdVwmlaw2zGZm0
ZEnSTMdl7H4E6RbjnE8xRoNrbrrM+GOF4AKt2HuQPd2uLLusUZpWzImnFhSlhCJ7L5MjpDAppW1p
soCU2MhOn3p8UWOfPSPaG90YZyEZFL8ij4AmANi1pVHNPSg8Jj6+DquRHqfVcWJ0airpfoGyKVP3
9MahorSGIerdyILuLpDKuzewCuxX0l468p9+88PUAkjIyG4lt2iaTGWzZE5rtgXPLXn1ojpkwRpS
kv3VVgelZIJi/nvs3OJS3hSzWW8NEFD9G6lMNS5BcFRPSThJY/IIQWghbUlQ/XySyjSPFwqxQjXM
P1rRrx1t5xHXEel0b6kYWPNDQz9uT3ga2RDCUlVeUc7VhrnFzEmGF9E8wAxqnhZqfvKd94ne2dXs
a7ZrFBJ4YmTMPNEB8oce+R/n7uo01W2VFU+qdsOsImYBc2GiJWHfbMgJ3Ja76qAbE3tu1rCxWTHC
RtZSKNM2MX6ccXCqAOlNxSsKzs/kUTbAHLj3dLV3AYio+EavV9fvW5wG60fmZ105ct6NBokRXW4W
tbHtRTEbJG8vASoXGcrp/BRcUIQ+TST2YcE/m5mJBGBAY1gN91/TNSHv5YRsoZ7VkVwrSypOyuv6
t86GuYc/5GKI6xv8w0FKt2EZabVbAtK8bdy1xPM6tG5YcIlvzIfiRzQ/yumMBVpCygL2lZSDYHP+
la9vE1n/Ki0YU0SNkBH+SmE+kA5/ENqLxI22OOxbV5naGp2OXEiYpxNW5RZcEB2+B8mGbYXQdtqq
6vltf93ONS5YCeKZH9ZymNUEDMq/TER8cIzuEOyzzZ/iAFmSdNCfyrSYAUMlT87Vt9UirKnIUXOw
q5SIrkE9ZvhM4K788O4U+dXsMo+IY2noMXB8f9CFrcP2KmnPAeDlO1F4LPXmJ8fz/i+60BlQuh4g
xwsxtAEjzJ8LfvdehYiY7b5bHL8lM3AZ2u1x4pKasx2GVwWkpQS9hrDygvRB+G5sJpH382kGzQvB
ONayElIEQh0Tbsf6vfWH6mn8Zc4m8yFiNYxY7LijsIfERkdWfsQl7FyEgD6xxSa3RsMnEe/OjQ4/
Dku84cRzzjwiNwHdfCzNBFtdH0VWEzxoRyHz4joVQllyZWP3DXMCy5jArrfTRZbEiixyn5Tn/oak
d8xQMNjMblXaAqhTBHvSaDoz5i0VR1G9AQyKh2h5/BW8OUyoJW4R1pTIsPUSlQAu02sNdkF2B1vt
Bof5JThUVlvg/w/cb2GX1Wb2Z2AW7ZldQfuSOm1nAM4ZJoN224wAqmU/GwWMpW1ziteZlncD8IUE
glfsweZdlVHFHR2aCRv19jz9EDVdsu1uYFU7N8VGO+SR/vYXN5zp/x1b1fn5UYyvQW37A6Kp2ItZ
PSv9QbnKe0SPN+or951FvO4MnIvstYPn0+Uv4os9afsuT55NYqXqDDcJFEgMjooF8LP9aG5vLo7o
ZS8Q6nXA9c6fiEt/Pkkm1VIHyKS/41SX6JHRqC5bd9mLg0KCjFGCmI1XRgUupL63TiPWlHDuM4W2
LetGK40GHXYtKYGBCxPd1lyMpYGoJWpa6UGcLcPy/w7mYbVtY6APZGYXcKalXTtZzZUr9M5W04GP
CjT66Y4vSzkpXaz2bJxIcNfHK9PzoZ7293XkvB41vLvZ80E6iiDgJFbBR6z36HZaGvAwCpBE4RMh
9RBujx82m5lWNxx6GmhSbgvdhXd88Wq6zNFTZBBmCfgjOULqa6TOSWH3sm8k5dbykD7xSriLX2y1
X2MfcaB1j5q7EwupeGVjY/oTQEXY4xI+nwz7BGfVmHZi/B8YPWF2ni1eyr+8iQMsTqaVpjhh/hjE
d0VB26W8I476G2aMxsrNexlYrkvnkSIpkMPeLv5sUGQhPnkgZancsMRG+gcixy36HkmLFvN5x/vZ
of3nTBCpR9fFvMe6Q6J6eyVggexpD68HVnT2fEnv1GaVot/02AgpVuWKjW8oKBfqjCV88uP01HP5
6aVOcbrvqmXJdVePeFWywdg4XM5XhdidezTgNt4g0NErYXzAN14S0i1GBN5fYlRPw9iKyteDG3fe
NZcj4s3mYAGOLT4RMMt1vlRUDVVTe4bqBo+XbvmDsp/UOQxTkNw9Gw2WWNXlSKe3FIHZK5wyJBcB
2+6WviQ0wbAn6gUDihs3hhgpcRfxL46+W7rjGXMX2s1jvYvNxLKNKfNaKpcv+ykOD2KFzJ2M9qbe
DZ9UapSXFGJ6HelcsshMVkXWO+xgQ9AJawMjANLBEgd8P/RYhYqsWM1liFQIio94ujKbl2WF6/vI
63fL9sX7XaTWeG/U6I7gR5HA4auxV/RA0AIcGSJljsEqu8MuLXSeh9mek8gaS6vPD26U45pYDRHs
DFwLId/b1wr26DCVqqdVoeuLfGwi9CDp/QeN+8LQHpddd4xEpELP9kYhGDDqiwK2a2AX6QL/G9/J
TlAhrXIUQd3WOaeeYLvcK3KGfHLQuMqKbEhc1mSejdxf5wreuTI/8y/GqC1aX3Q79x0QUeX7xr6w
maRj0eBy1B3vnVzVO1ESkOhQAXJ9O/wmm+LBW5qqZSCeyIsGXW6oR1DCDj6oIgalKco7ldscommy
ObvFFGMmHHjdZ7a6zVfoi4eIVNfEEMT/OechY0rudwjwTo1WwBB+i60tFmnL5q+aMXIRvUh0LOt9
3Xy0Nfkc+W11HRcauuQZ9TQu7/TH2fWmj8Q/0f5hIINq1Ln+0VLXBz2Mq6mDhgDC2cnGKrOe17/B
ay3wMCappKMlMKO27I4svXM3P9MMQqCtqGGJwSonkfD7dszzmf6+E7mFIi7TDljJOene8k22zL9j
v6ciUgFMViJa6N/i+Bwp0FyD4pjuEemiPHzJK6q8ciOZjNBCpiyvmXyOqtKcAK1g82u92dhB3pyy
qd4H4ApM8OjgikC/J0fkqmA2kZiLawzp3V/YiKCzsveH16U/eCfbydOMRtHTavg+v2siNUwQYS3b
yUCPaioLOpfL/DpzujX71gz1YShbQNcAhSYjEsVRuCjBALiOxNsNoy4KE1qapm0XOEHRPL7T747S
1xhV+ZGICprSPkuDtjOZ02nEdtNzrS14IsmKW/n2xrnF689XYx8gCt6yD6A1V1/DVLfXzYPXP7Ii
Lm3936t6Sa0fybaT3z5Nr4iiqD51OYbrTzryR2JqVlxKocHqNv7fkhAUkNn5eQ29UZ7HEIkrTXZZ
P4kWjl52fFeShs5bzRQ0HVGAY9OBHLoQB4RNPiA2d/477a/cQ02hwqN3XTT5Z65I00R6OHAO9yoD
gbi4zTgGB7EZKH2sbLI6FZ3JCNQ3mqykqX3f/m0lrET1A5sqbib/Gj8Oaoaa2KucHw16uJAq7exL
kQPHeNiG2eLZJxbon2bLc/F0Kkfi9ELf3uHuY21dEIlBgiagG9dD213TNeZV++K1RVNcWJvcrhz3
XaHkjyIH5inAsRnR7R9/M2BB3ERdhEF18aC5aU/24GYpDjej/GYxQs5g06PQwncVZf6ldHk/4ima
y6ASKd3RHlLjtdHsv7O/rzyWhoEydv9A9JlLRCGuMMXkPharCSXpel/h2GIBFW/O4KegWaMCbhR5
yzX4gCq+GqbyJeJOLDnbLvnGVz+OZx8kAwSxzcBjJbibfGhTy80BsbBKqJ3gfUJY35d7hxcOHC+X
gPrb10cISPC9Gf9qE0zmDGecXFfXyT2WMisgn1u0L0IqI8Jf9HlaxUtIrM0lWJF6HO61lJV9i4iB
4S4FcZPxFafPrC7+avxYZHI8NGFksbboTOWFM4cql5qAoQNaFLbwTSAncsgkyAdk5W+64snuhDPg
9NSKAUKqwBWHLjZbbFaFCxl78SG3fbBCy8oJe0fpzj9Hr5Ty7h+kRHRM0SdsLOYGtOtkSO5VCJnR
m8XzuZNzv/xmMYpNMaKEn6hQrzglH2rCH1+gj8FpHq78HxWGKi7pn8IwZAo7/8m+2a1dTFAIbnYB
mTcwTrzxGFrioL30dv36bT/Sodo3evmQPF5G4p9S8pqAWgqcetvmcFNswzSyVYZricn6KTC1Ku1y
K6uJNR6zL6rcxJ3OmHLIRwlQbDbzYYfDVbZJoyPocXAW9GaYr1WnnvYunOImLDVQQgAcpBIB+UAw
5isIPojVDQUt2UQLh4TQpySnJrEDLt3Rh9GFzJgR6RWnG1nRZcA/9S/McH7N3NBqOYNR5FR1W5KU
4Ovx29dAgI5g60AQWFsmTiMs9GSN9SJQ4Yb+0vUDxY0cpedFEqqBP0YqrZYPcYys7sME9yOEVvlQ
3kkuNodY4FL+5Qb8ulhvEQW+ivV0URcBiNRSNRTnJBiulzEW7bY8mLsMyOdL2Jh3k3+1VF2zK73c
Yi+CtREf3vCu9saM2S3k9fhLxo7640r8GTFtQ90r8Lob+IomDjSOfh002+68XeEQxXKOD8UIPWdi
jZo8kzRYagwnwIxmO76Ij91mCJi5GbVHOULNj2H5YcyGDZG7/8MtaVJzWNuQJrUkBNV9LEbSkmEI
1Dg+g/ExPE/vMbKDVckjlY3pLOPu9CZMnTgjySUxrbK917j9KtiEz1l48cxaDOeJfz+CW9tvI70w
0matol4g6xuck6q8zhBVYK8aMGmCObP63woPC11n5bKg76Q9D1ymHnFdaqdxKWHClGsDeGpAEtEo
tt4AOz0ZeFJ0x/tDeODDBkNUnVmaJMbww+hKisreJ/ngzmhDcILojLrCBKHGoNMnHdiyAFY0FlKo
i9QgHmO1zzC3egwkAzB9oxBA5X/B8123HQ6XlGvQNiPy5a8lEbWOR+a6LsfCr7NS/Jp2qagcQpkT
2OTfePIEgD+PEb+iNj8ahbfaMJb3R40Kyet9JpGbHdc8XBYWQM4w7aXdLhPeZfSL3/cep/oecNLa
9hIfezgtyFCXra/5PWwAEm/btV+M2B5A2M7Bi4Bsc7tk2kMvjJRZ5ULsCPOz4EoTCqBiMXmQjFAd
0c9Iswkw9O7f1E88ptdBvdnOCKI7O0x2jsexpBrm/N6rQ5TvawrK+ttORImBXOlKefuMWLnD16PO
uyY/Tgo+sySOm01upyGK0bVBfHCdBD96TEWdwITIJ4VrPjM0Ndy2QAUO4ldpZhfpiQqKQvr4eg3p
RtJrCTd772S6v2blaV/DPm03UKaNEmlH1c9RdxOasb01IWK7UD+2Ak2sN1jAYuqWi8UEIO4UN+Wt
AsHHlgw0nhTwBXY8FqiyrMLfmyhfFj4nGpOr9bxjokYl5+HbvJDrxw0NKgAPFFDBPSviguWIPJS0
zLLSFYlanC1AuIaR7ziQMrqutt8Nklg4I4hs16JwF7Qj/nwnQiVbheowBxTDpC/JEGoQ4pfTwYma
F02tJ4mV0EnMHp/lDBkCVlhqPUY7SzhDZkqEBi01F9JKjJppVBW83KmcOuRh6F0kACJgAMDL90dX
YjATLBdEAmmADBdiSmgSYPLBQV6HcgQYuV9sTAOfoGgKIU9DSVdLYiD3m3TKGd/02I/4sgQKvyC4
srTzE5fM5T7Ub1X8p7x9yxCLg7dUKqUif7U4q7VC/9zMShdOSU00nogogkkbThGE70mI7xBv2pca
6U4ODvTQm7jG/MCG7mZdN12IDHll7g631tAAdPQwoSoIkDKcoHywHG6oQtxfKwJDWOGYItIUEqAi
133Ff6Qz7m6a5FCOkInSioe4HHI/qfJ0dD83uiIiKipQgCxK8cncHchLGEDJAD29SLmA2Hh0K9s3
aT3ecHqJhjZFdmWVgz2HJGzYDcowVW4BAINa7kayRG2p1J1ok1MEP3LJ316W4/4brR6WMAE+iHE9
XhezoEHasMY7/t0aFl4AlZNmfgo9lv+WlHJSIAqNxTWCx64G8oOD2EZ22P06W9PfmVlryOCVXcE+
MY6Y9iarolv0kfqIUpxfzg7dDaiB9mV1Mdw/V2pnu7NHzn3kdHHRLnvMTISTu7jlJJcDRahN7Jvc
1oInkPYApMY4Rq3x0VrWdBxI6lnH39/mNsdRoUGEcrZlIZUrSG9td5jWrE4ZUE5TFuQUGJCE+9Hl
4lBe3BellCDhxeX5URSZdXqukup0trsvjkZt0FNOliWclcb0k05Xh/8QekAH0dJeGC1bD9RvHYAt
e1ThZ9bbTjyPeoZazGs3SZxkTw/Jflsf99lW/r9xhI4aOHWL9A9YJ76YCDFfRIRXKjvIepYaYPeA
iRKBvLrdGSWPT0333jjB8+hG24S2A8hWJqbGRKbWK5DlUrB7vXTWm92ppP8ujlvtcSRYiVAGZe9E
I8RkDk7BTdXNeqoOPcNW7sRKeWex6pL5Rjjzy1K8AYNHtGTD0qbpTENLsQQspdoBfzv83gmMvgbx
boje2DptKZYsJuXmnyTxSTs3ofmtbYpHE+APVyVdZBQkDKxT5wSNpwAxz5hq8fouLFZXvqBvOuEG
hdRxw3msH7dmblyCqGyFUoUWkTBg6js9cFYFG4uxM5ZVt3qhT56ekBCQGluV5QmhxlQFbH3LjspH
eEcITQnHhN2Ortzv00TMNcwIvFmnKnFEw/41bhOrCqSz2KM2IzeViofB7urTAiEAbPrKX9tocPj4
8rEjpf9pyQVT8PDFZnQnc8hjTeRML18+3f6s9YS7virfluazNnBUkFZozZh7z+a9yMKzryTWq+s7
yLvnuwi7h0jNKxWyTs2QoELiaEdUcIqk0AhHuTJUEjiKnlT3ahohYfVjn8w9ZuP0DepINQrvrVmn
SnWJ1Mevs4FiLHn8LqYi8ODNwrE2VOy0ocRnhNTy9F6LBf124br+h82jNGFz2IZYbCx4W6nxC3YD
hZw3c+Fq+awntQItmhT0PRCvt98Fdq+2VpSzC39pEBlO9hnRVzFaCs2euwS62h2ti1RqFHUFrG0I
l7kcKSQZtszj98Nmel2CV8TklyMoK1ZhgF9TwBOKt54PN3Ztdxpi8laFEPXcOY600edUO1ewc5iz
na1Zpin5u4N5DzzVi2L33Q2/En5JV6vpFjkP+bWYlp2qZuqHRRpV740GkB5hF9NVMGqNBzT6w8B9
6esB2BuvUzeJMGxYoQ7f7HrgwO0LOrTjvBoT1m5YZ1Cnd8Wo3n2rOSn38grNOfnhMWiiNtEESWAa
Y7R7uHQQ9V5B2K0d0gZ3decv10uRUx5Imd1d9HzBi7mvubAjlrzMsQottxr4iYpVtKbfWPmgINvq
7vgUy2dm6w74kPFxROUnqqfnk4KCmGV1JTzI1FwFvIrRvguHo3Nyrl60Q5GSFCP8HT/8X4QqF/Ho
NCLKsXHHMMcmPdnwM8u8D+GITQjQI7MZR2UcD+PUjh8HrQ2RtyY25LA6Ld9Ig0Nb3zSol/3KYRCH
Y1i7Jr4h0j/+RWQdM0ryyouasydyCO3rD5fYoqAvcpVKgO4vz1Tl8iYlUcLpeD55sh3n+jHjjykK
XlnNxrRt5IZNRKMChsA10yyBWgbwnzJu7lOWnbkpM0MA9EaEAx9y9breFI6ZGAdt6aA4/ar466W3
2RrF4vvozpEGHtF+N6J/IDmRasvl7FpHNu0aph+s8OuHR3n/PBTzaydSrvOdQpu9+JX3jVENNO6U
698mIn5KlLqQDH9R3XTjkx7zWYUMXuGCgWJmNASwsDBMxLCi1jZwMwF1L5ZBJ1BiNn0QVFlDybhC
WmPOCHQ9lKCZrTqb76d9B7L7VNGBjHGZqgR29XQ/1VKT9dwcJZwlrE30AxW5iBXdtCovrhhfZImp
8FPwNkvVoKoGiTIVFNIwTxTa1Xlsck9LmmBmIJnBankpBiYtZpt651HUkG/V3/xZstXnkriYbNVy
D6YSOSCXQ34sNPhqPSq4tJcE/YlhmqRdPKtYdA7j1Xy2uZz9r37WbgmyfAgpnxcfmw620FBUb0Od
aSCAODoKDjUKbvstQQyNOoNgssWvSYOadA7wPNl4Q58Hs1T3E1yK2endCteOFbCb3HrGYnItzxJu
/Ub0FJcqkt0k1a+8MW93H9U/UrBMOLQ/Xlc8zgwLFbqadrX5ZobbtK9ul1ujNU+IwZnSikp3NenD
u4wzVVffc3nAgOm31g4g7tgTPpMy/n7ewn86l6jp3T0BzxXHEiTC58CZ8/Ym5uoLOuLWGZimHCZ/
rHox1SxLfL0lVXwkXwBmoO3+Jr7uJ98uqBmaRftShQ7DXuF1UHGbUGHRzfMsbqyzgalJ6/9CRnEj
inr7Rl/ComJb4i1xL5SS8uzhZHyQWiMQR+WzVy9t4msdGF+1LIUxpEdDhngJgkls6csqVPTnF6Fi
VqwwFGXo7Mo22ggvNDXB4SpYz0IJ4qOzLjNGywi2vOTSUVPOQU63Yszvj6zQHDBmiU+opqLuc6nM
+XQVHWxEGV0uxHTdFYJLyl3U4VPS6Id7afcxp7UV5iDeXFzcGD2S1DNklrn/m5zTfG0PoFTo6g8Q
8HyCPffIzWYez6ozuTMMa2bYOkYFqIa4hctuRV0aOe2LJ3uQb5NYIoJEARVzoMf5RWSI9nbWP6mf
upMnQIW0KNzRR0fgZe2VDAu7OUthQN7lsOwogV/k/repP+lgkiY6NWMEm4VGoukOvmOl+W3+JXJY
V29PeGvoX2jMltL3AsndvtJO/r4LXiO4O0RHtL/HkxKUvamPOM+7mvaYOIDrO4wXCACpAeGzh7Zl
Ye1DLZhP/35OGF//Z89K5bt6iEO6r5hH1HFlWCyzIr4bBzdr1wPCa6Nm1BHV1xOi9UISsZ9I3GfW
/8VuS+Y0isVxpoJEm3okILyo7Geo/R/GrNUDOCAA3mBN3wdyO7PqUXZrXjmYBqvzGWeiSN0zD0iy
Go3UhWXCQmDc3nm83AQqEQvXZdkYIJX4YHnpoQxCW5hR0LvNRkqs8jsT9xWptWbzH317U+PmKW5J
0LdWeHxifCSogUbum+nAE/zTd+OXtj4UXRSNpv9H7T1+is8oj3nG/u6hRrJoxPDXPHTxpvnps+vV
CiLVm0L0u03frYVb5ZrbD6qlD8wZJQISUaZytYjGQm0+WTJzfAfZO6lXVfLojLs4BmIFfKlKsd9d
Y+KzxdIiOqTwUWlE/gW5yO4NA8odSatkBd+l9vrRL+I8cBTs6f0Dul4QILnvKPbT9kzPOzLrb98o
xxJxgX1yE0QQqGsVfHYR7iudD+QZu82JS2MZlGwqpTwQ2TmmJBVyAQbooAvKukwowY/VvhZ3NC5z
OC8+z0s4YZM3lUsqg9A6Juzmt+mM9Ql71UWIgJ2lMPL8GoWDw1k1KNfPNAV6MOWXYPO+clq9Y0Qb
UniOXpvXaXNVPNdr53QlEkrzuM3qKTEHofTz7s6+7ydErvKsek9K9UAZlD+7QzvWHZBvg/KM1fE5
0J6dUq+nvEvWj1tewh+F7GUcnyJ5Egl9ZDh+mJt15kOeEisBxw7hLmdUu7lt7Hrvq9JEbJsonQVE
QbGxxkqZ38/b94f1fTS2lUbvZIf77nYAZ91YFg8tlor837YtVlu/1X7/p9Sf5YUdh943uDITrK4O
If05oQpR33LgWJnLPref9tgHxhMhQduqvd2xV1fIgGwAkeAbrhwOWQuerdNrtXYKyn6QuIf+L2QS
7JjIGHE6MWBDMqWJ0KCZpOSfpcUNtmAeXzo2ASkkpi3TxZzGGy0B/9OnC7/KAfx4nw0PbnhfXli5
R/O940kdll/p6Veax/DvpRd/Obbt7TQkpR6WwD2nFMCxQsaUjab+8363tl5Y1Xt7u7/kk0/o32k2
CacnITNNaVc7nnmkYhdW33Cb7UwzW1aIWnTETU6rPG7QkTMNg51EQJNyjOkuCZcS+x1A5Ww4MXX7
wb45PBZyT2x0u1kGKmLKob3tObWHia8v6xjS3E37Xko0d9l02AMdEy77SmyBru0EXhDpI4cJxN0s
Wkbk5p0r3FZjZLWE7Ed927xGxp/TSVjwRVwjzjt/nQin0tYjHPbsPqvzxc6Hs21fIoC9633NfXgs
WaTgAWc/IHnThYYAEuS4ko3/HASArovLGOChTNKLm5JioC5CKGJFpfxhayyx+HQqGUSHlReqHZxL
lh50ilf3AJoHpUm0X73tfcoHn09A8SQORPNp1JXxp2hRmUorLAFNJD20iTZJI4I7ya6LouYfHqMG
XNvkFQ18OOUEUV4U5WhGehczw4GdeNbDYStKz1SRO+Z+x9k7yXkt3kehTR3hlqUBnmGIDN8OQNO2
woBEcuYHC6fHZsZivQ5ioHJe4xIDOMc8TAEbT7VCfamtDlbvqa5webPgcKdJcNWv3p0Sz1BrmYTf
xqEcD64gQ3kjE7mTRpz/AYAhtbfqQkTVn0MfLZElve5/1rPoQA52FDFJjDBubWgr7SBho8FSPo6C
twMGWTg8RcdNionMeSI+PbDVBZ9W7r+1FTZsjV1RJ7wc3rZnTOJjdlpLaZdVoeaqD4zaLCaaQ+qh
op88cC6D272001JnxiaMtml8ooMGe+565w0Me90ky4Ci/ycq0uK6yLHop2ccJHKWkWKJwQNOHDC5
lpPPivQ7tmaQr8VuDfZWEoqFkqVWrsEbokOG/ypMUAYiVNyzoD24VTT+dbqJDWvIScri9H3sHwZM
lCZ8687/gIiDe6Syf0PaPEwQGNT7kbbqbYN8AxgEMK25Qgs+WP/TVW3GSxC3qzcpSy0RRM7JYsdu
MfdEaKF2onRDDBWgWDGibltv5j7ohuwGebICSwvTbmKIAEikCOmV1k6sLjLoDnc/Wla0BOexZ/22
5UNJVZ0u+yGyP/jKfHyohNVyDpMhkJMAFWXoB6Bp8Ey2yiopdIUIvl9FDzTJFbOKVwE57QrVb08e
OR7juHHtSdGUpzuUD8DXbyupmS4QQRmvjABf7tYuCKUlCwL11fgjRGVMLQeE5nVVag7gFrrVxSAK
119wt0rNjF/8FJVg3ShS9LwriDpGERr5Y14fMvC0KYV5qoBTfMK/YIrespfbGEH8RY/lW5RCsDEN
7oNuvSaqni2KxaolNlXqD7mfqRtHAWaFvrLBEeXzjbjPWrKhrg8/3/6dQlGIJ/AiUIHAvzU4jSuo
XYoQSAAJ5OfwP3NgbJuXbBw85mlWaQB+atI0j4ow1Xnx3UirGhxPE6OqsG/3CeVq+xzSSZ4Hx5RK
jjh0DzoQFEqS1bZuI55oak+tkH6BnXL2Ut+DIf3TgV/8ljkiOJlzWIpQ34ovLBjFS6NgcGkwqBCz
5mEV+D3VHOyIn4nENiP/AXPapu1vYYpLxHod1xhKMsxkdxIi6hNYwlxPpyHT76m5bXM0sQGrC1dF
X3nUvXRT1pEYVHo6p2vSu2LXQkzyQNkFDLtYRwUdqiPYndmowRaLe9gJbEmlqHnaVaT58AAtJ0l8
wwZUBIsF2nuntCOgpbtYyzl3ERH3srA/eVoo6vr3ZSusg6rTus7xMYKcEAAZ5vsX/PtEaRGLhq1p
d8Kk8yR2VivJRXMUc6wYTbtBerpFf5fUSBpZInNLmT5Irrg9qBrblxT+kCXYp+PThij6ZvLMp4Nj
T/JFtJos+mIP4Wr8z/HeV7twF3aXTt9x0u5+5nFh8HL9UV7TOMIsGtqeGGUoPd9xUg2CNecirhMn
MC8fVf6S5wH5nMSyMGZkRufKV8qTPn6Ah3M2koCdRQAP0gAGT4VkFkHwVwluTThWFv3opgGwe3wx
BAicJjnSn2OYCMcdcfHho9gOAvwOVMjRgQ2dWI8e4IppJ/U9qh7cc80LA6IWv2HuimvP11C0qNfP
1asljwoPgq3G/7i23XY7lE9Bglytpn3iWXW1qLqcnz2ri/i/ewgnozHsNXU4druuYU1n8Q1R6fEU
5AWdkqbPt1xXJOmBsc0vkexZ0nNF8GYWGVBAbrfYmVOgGzPyHG0HSjU9nXKsnEGf24cuqYRiyJ4t
gj8Ho0iqBMFvhMaRnGvPXGYp7rYFuNTWkAVnUa1JelsVd40A7DAE9+oNMLiIR56uFaNeAogG3yKJ
Yr00AiMSS8nTniiGacjD4duHjSHNm+V1xkjNG8N2jwNXLH+ZswNj2QbIxX81OIrS4y5LkU3DYDjv
FI6IDyD6xvSC8iLCYfE26bhk9yBMJRdnYPwa8uKMuUShhj91VqaRZvqCm5G9+jM1i6ooJItDUSRn
yxTKE1i8L2JZ7371isrOi9arGxhE+vyOIjlVvjIzC4SjXirC6GWunJ4JIqp6EdREX/yyQzt46Frl
F8sMNAZA6MlP+aUmnr7QIM7FoKfFup2BeHw5uAHxvRZd9yWDK4dijDHwkZ/ZW/E3mUQU37KYfyiE
hwUqKO7/Vyf9NPcyuSQ3kgqtghaz3H/+G/UU30QNX9TZpkA4v2AcoopyFniqIroAGfKpm0AnF3PW
BxlmzhPPjw3B/aGhy0+DvIlj71IuKjQJVUXoKXY2Y+0XjD9rN4IN4xK4zDpJLCi7/64ViysiwToN
WpIFB2A7kdrL35da+hdctaxvWp5cJMRWqsy8NMKX1GgeBDQ7YrAPe5FnOeDNHQkmxA96WsY31CU5
egr3DzEXaoRX68EccZiwPDu0wlCQ0lmPZZK3NTfvZj8nyV95fYgA936ylq6rjtM0te5qRMrhYlYB
lmyvjQNr1+QcimqyGU05ToIsTH1wUkjglfowPT58YFzabn/5blbPltu4G08eIL0kVbwphyMA9+lQ
B9k/xbv63ypKFjYqFl3/kne08+T07XvXjXl2KZ/35dADHlLnxxDiE85OPUNt99UJgCsZrm2tTvZa
2pzzSTilt/BN5A8X3NaFRR1n/aH3Dk8aQEG65vJLFyOu9CwEuTas5VVdYXdJk2q/2Hg+X7RYFREy
6dN2zAaZD4DSIpDKYgyk8cc3MVjLAatxLXZ8SnfHrTtqsm/4FTjrMil/Z42DEPOXnedCXguWI6W7
Tte851SibeOUEaDSrn4Y7kcUYQf6nfpujuyKoO8CEmdHrb39Xwk62g6FS2Lx4qn5AYtFIYHCQNxt
yiZip7FWB/nJRHDFirm9y7x7wrPmGVmvXt+jzEILqDwJrUC27zfBD+vpzxqwVnRPETCDxUEn6jay
29yHgqNsefkoZgQFO0TOjkdiz+BEFOPl2TXywmSKaJyteqgf0I8A6dy1M14USFQbCr2YuGlkniCT
37V2Rh0lQNN+JE8SOTKfmLCiK1xZfIpBo50ysd67mEOaOyvLArDAOeRwDU5SYhTStjLIf0eLROqe
jh73FdZ23jWmWYVHxFwcpE5HdJ7xVcXwucD6l4OQvq0BDs8rT0HE8W+7zJEpEbyAZqzd7xHNRBQl
FwJcfl6iA+W3gNziBCHdLA8x/yqsnnrHQD+jE+lMyeZB2Z6mYqu7dBCrd84vu5GYMMxvDt0zoU7f
dO14dqBaqKW2dAsEGQEZ1Fv/HN1bM1P+EN8BTJAi4NjgQUEOGoXLsnLe7CptCb87eC1gLoJF9jbE
0DC5eF0va5w5zXAkYwNje5ZB373jtTiSgfRWuwd/NmzgOG5fvoYKWD19OHX9QylLO5nVSPtGwlNX
5o0JWPQ75o2PIzTWmImg2a84XSgGJRsfUu/ajVxeA8lWAd2Zm/StMCoFiT8qlyVV2hZlEM++XLAN
wiz4ES1lUns9VOhr9Anpo3DNK/rQjU39Qf0v7xlAgGvmtXcyOVD/GL8nnls5jsz19Yi9G5nS0+F+
AxyDBGYqCbuU5xxHPJ4h3Cv5FdhwCyGX+dfd4dn89GaYDAzs1+nOLCGmqqj0qqcHx5bnQILMN/1Z
lskx9FgjpFFkmyUNJB69KINRf6H8JCGln/fLXC4+NBZ/aVow2DnL5r4KJipf1AXVoYYD4f7U0KOf
U3c3UeDtP7/auxiLLRM7jlO1fpTfr7Pc4rD6ige+lGC0d1DESs+1fekZzo34bYcXMut6FpZY/V7H
C7/UWZ0n3VBzEkj/8/Q1YBiIRgFTQo9T4VrPkTDX9HyjJACSu8x6Tpytnl7TKDHijFudklmgm4Zg
Gevl24U70BPcmNMAP/1NM9L89Rbow83Hs5to6zYXe6sfo/bhoh4sZLyXsBVeqX6/HkiHTNYCNa7v
Ip8bUMMsaJyl3oY1styBrSDCFV2n1/muPCMx6nt2WiF54PEfqFJQpVuQzdUGK/Pcz2roOapymLpr
SbR82HzajNzm3uCQQmjId+E/qKLYGdX3yoT8rnkIlyXMeafCrVFck6UKPmfvznb8T8pmsycRw26Z
F7fFVXLpTi1roOGTOec4ZDjj/KEhUquzpFbZ6JkFYD7gJB/X3Zvw6qbU0u3THJV4qmuCqYyYwHMj
4YwJX+Nr7fwCTS2LpFNgkLnBiU/KzZ0GBke6MqOKJ60/rf9mVmA33tulJi9Lh9R8xKyLv7xIE54g
m9dH8+NloH8KIwx7eiIS7LXo0XWewRC3AwbxThlt8Ac7+rApmaza+pQMI6mNA5I1Qi+IbbBW/6CK
d/Yrgt49FzyGdx6omd4mSC0N3uWGnQ4T+vuYdUd1lQmfUwsHYW6jhdoUsma54r6gPRcWik+DfZ24
ZZw95Zv9xFQ62099EH7Cwm5qOIGxxGwe9E6Iyuh+j3kELcwzNAvCOpdAR4tgrYB08fFSA5dJH6cJ
8mJUmKgVDxh+DEBU2RDCmpH98a4zv+Bf2oy4xXEie5MarekjjQkEkzdc0RgvRtpSqs7Q9sVa+4u6
9OhYqg6K03xHHRtL55Yn46+BYMDBdtOJHaSfcuv4fcifwQNuctMoSo6Rz/VxSMXoc0tN3bQqPzLh
mgfj0rm7D+ndUS24HEvzFoU5srREo5Zy0XjcnR6Y0+UiHFHrr+NcVsvtSB81SAxBR7KEvTZR1dHw
nvfu2OCTAse8Ean9M8tEkkkPf53ddeybccrGaqKyZe1Wn4rKXLrAS1OammX8GuZFokLaYI/STRlG
jQjjnBnzZvi+mFiXmzlIK83VyqF1FN98QjAy+QbJ4tdoVg7RY66IfeAarRUdrT1xr4fQH6PgTbmO
C6Wm2GjBvh9z01/97Vcg+xZajxBD7fN0XotWBMbkg+L7EYeMOmriM5vjWdixolkVfanTNUtbrZh8
UynTTqthqqeLuG62nxkSTHEQpwJrkxI7KXVL674ij7HdRrRzr6Zl0ZzOJ9kTR7oD/QWszWFhBlwU
ZwFY2fqaY/B3h2zPula1HvQkLOTPUej3EjtneOtFZzqYuZFZSdKVP9dTKe9txpF+tQKkpqLNjmMZ
992Yt96bfUNQAAYGqBOK+kDNozMPKyliE9PD3pOMstt0OQYGuDoVM8uhUhdB1NGXyitqNTr+IMcC
bGvvT/2I+gD7LpVfnPD8wOUWhIjuISRcGbD2vfSB9ztuOwPqOyNLBV3BAD54P2Jsgpt6N4dQXCKv
88Ke8N5N288wTf4ap51fxCJF2APB5o1zG3/jnF+IEQlropA5qvtQTBOGUJXY1D5X8eUoSVCYKwml
+12Hv0/ib/eCtSKq2u0yMf82dNEBME3o2d0gPFzyqDeL2DW7yLnhjduZaAUc5V7mI+FZ9rkG7qEA
sVDB5mmxmbvGIPz2dqCosQK+6jo0YkG1ByQuBS2WGN2efaxu2XMW4UJznEJFqre4ALrie0eNPeKW
WHe0TErSzmb3hGDE3qg1mLYYGr0cmq3vc+CtDockxK2CLimy5CmX/kkN4UVPmWQgCX99SUG2Bx+R
PyGjjXOsb0e5jyk2pKiKWcEpYvID6f+EmB9kFeI6+qxINQzmZoidMDXoMohAQnJ7KRbMy5PVEb4d
j/47g8NBvm2EVjknTu9M2A8Bs7ezoc+UYVMl2RuaSOKrHcP8de7Brs/EV1KUcaJ0ueWvEV5G7Lvj
bdc1PArxmq0q5fccW0H7u6QGgNJh84Tldwy77fMn7eCbRrOwaT6rUCxzKKyiene0EAq49iuQoa4N
JqcENppigGN72QQTH5hM0ru2fKDeKPVhhKb1Kh8udb/S7Rpzb/IfUBhnyw0cjkUVfmFPWjZMqbxZ
up9HvxyPtjPmeNSzF8vO1bCOzTZcZzADlDEzuzz9UUi6ifuQ+eWR9Af+qqgC5CZcsCmxl3JYOOoU
8/G7zaCb/7GrYc93jXOzTKO7zPi6mqV0bvxO6CIaFp2f3/ufplRzov1oCnPBNktoB9z3lzQv+DiZ
DCm1bLAYJmk3k8swpQADx7OCg+CxYdgvAbIhZNBz1vp97BswJOOy5XrQIvTcbir5SsiULmel/80G
X7wwek/qyUvEPr0JMn97EYf4MkMDcEtnm/eQ07zdQAburt8NvPHIpnDKbGE+21jY9aZcVk2MzRAh
/GJlgG1u3//ROaxNkqYfo+hBoy6TcGvGhKXAMeBk04B+Mjq58lbYIZh9NeZ8IsykcGXC/6Fe10Dx
It9UDQGEZZDopXqGqlCezJKydU7Hs/GKhLn2b2UFfH/WBsgkc1tlF6mVt1vY8mbQrDbhs4hxK3L5
4qej90QL4HA+7odBX9DcvnRl0ciEDCBWLHOgCUZP2PRq45ZwPHXm8CUvl/4TWxiEPTy/QYZCQ/P7
rnCRoSsnAGSdBh/YAZohVKRWISRqJojz/Wgn8muNg60jsLapixOs10B/dg28xPAWNo1euihaGPpX
spAIxExV19KIu1mOwPa24MtNNOPsjTuRPqDanACQH8DbBZtMTF/iRbLtWHUxkrz+I0/ag+ThP5dk
9bkyv8oSK1UeniT99fbaaOgeFQLXzhS6ODNJiTtRVctXZDBCHvCj+fK7N4r5mjoX/pH1rl4UR7in
lAmNCrEqkqSWTciuswUthxopMR+NaG2RmKByelGXX6/BhHwtAl80/IRb2xrXq9UEg2wmkE3cpPja
vI76evzyGYpdhAtnzcMbX1U/BncIuW4o2TGNnJMPh0Wz18YVRxil5pxG/HeLK6N8CKBTlI5rFpAk
hE2zI+VpU5FG7hRv2AiiYr60HXMSefRWd+aY6OOREAQTsmzriKUfGM4OqheVgVMZ69Gt+rhg2TNv
DmeZIYT6T6pJa98Gc9XZlVMhpFBKWMrd8pnkYWqewuZjbSh1RAhfo+INFHEv6bhjuAdh5U6cE3vl
lOIhiyJSPjDlNO8UxviBLHFy9Qa/xl8vczfFZlvSHyap+t6SBTLZQM4+WPDCNoTQqHaGVoBmPQHC
P8FyO6DTfYO9b3/Wh+37qRaxzqg19N6Jk4qJVjJmHenkiz5wM1+ewwQJfER6du2bAPDnqU574IZA
Qw2i+LmVHGEkhmJ3PwcSk0W0flnCg2wqjHlsaH+nP78638PF7FsEQr60akIRw76ESjrhwq1+FUNE
pWvGV3V7Co8S5QgLhr6uEcpsBpiU4qZe8ehzlg+/ySpyZiNB1wb89B2Hzk2lNpAYHv5DcnUhE7gz
JF+oPt9SLSMvAlR007Ol+ip/EzJpAgkFqVvTewR4JLerz4Wrr4Mk2AA+COVEw47P+uoMOA2NyPHw
+84LA6dmsClbVC2Y7tJ6wVLr/jiKLoFy+vQztjaQdZzpOxOBASyjnOuc71Dcbh0lIbOuumB8H4Pe
zT3YU/togm6rzvzxC1HTTgC44ZXvl9BrAk6g6oUzI3I13xGwPydrmjdAjKCDgjqF+QEW3rVdeEBA
/Re4RaY7nFGQgePrOLMm/C+lNL8py3fzJM/ccsA8LfrCERUd51Tl8jNkKmOBh8mp/OOD1215XTGN
xD3jfXpxyeCHQsLIwzSLYYnhKl3RcUQa7sHpz43q8fGbtfc2DfqAGp9dxYwTss5+QQspwVF4WYDo
GUuf7q4CSwXqyG+FYkdwoMtfaLJPEmPAZ2zAnqhAXoNFmIpmRy+zocMdUUwxvRomKTLFDGQYLDym
unPeDEwNZNH7shFaVwGyhhjrNU7PeU4bTEivRONDBIy3LxWdRx5pad0t7MI4m4G4CPnCqXmIxZg/
oVzNKm+WmntqwOnXrPDrYgUPOPE8tTMcJkKBJSn5Ih3dWuiYbWGf830vzaAPDdSjC0FSUXP/3tkl
Z37wSXS9hfg3K8gGuvLZISpdG8OrkVDOudN7uax7kqR7xs6g7kfwZ/hiUBv/KmDx3EfWG1UKOWYH
VpXDZtT9XFcOPF07k/4G3br82wVo3mspVzGW5zqkcbuHZgfddKaKLnO48yXl8dTWOraquI9S1sUr
gIg8OzeWCeZMxLdDMZFPsZ9H7UE4ax+UFy+L6eljw+La81VdgmU7SgjaQFOckRZoea2x+dChlJRj
3UYTRNv4snsSGdwlMQUnXKifVdoHCZXE8ZMeao+cm0aMWybQ2pUyO57NeW7/Z96Z0YSaMmkbLe3H
f/lqMTKY2W5d/smsebvVIFOAW27MuRGScjN/2jcExjawEkMXIRmm89MspznyHvCnFFBqcNhtrweE
tGeNchp+93jwFPzFWdiTpoQ3r04BqNKyjH1UOaSHfc7Tc/J13GgI98VvYRgOyeXtxnNVfnQ03VEQ
qFVG8wmBoUqUf7raJyqrrLToO3vFMZxNaN+klw7WA7R368BFpFyxfGYqfBys2+nem/mLLAvJv4dA
gJTDtkjDbdZ17RInZwXgt8Hbr5mWyuMfDhohWKbuhqixPq1XzkO1Mu3N6Xx59/XhZe7bhqWPMzPo
BZ59/Ft2E3SXpANyp1e5TtjigXDQhchgtPJZAUaMHimM7uT/FugUoSdXEA0lpaWoLY9pCOl+NgzL
p8Yexpl+RIisPFcJaz6hV1uEm2wocVcC9HwqvyiYh7PH/a8Lqqp7Oskewg/uR42hJP9nGuSrQK6A
xmAYGf/kosz5OUPWkhUuCpKc4zCE/1AH0HMUtUiCGBj8iWAj0nM6w0Sg3klPOPGZk7WE+LKw8ks3
ceVOtSaeZ0vRxOnWx1jNAnEdZcwbS0oyiDJm23aXEuDjpnhLdlvgc2hD4bOI0SNJv5cioyzpfuhk
HOIfOKqnSg+2CLmELVcXazN7zGoLLmWRK6e6b/i+V/ehAgAUInXKWHJM5YM6fvh+k66RArPrNDxT
ydcdsqf95rXQC56tIwT1YTp1iThFV7qHTOxIp7QIyupaCxwCzks69gDk8AifUYi4SFbs87ResCN8
dYQApknE3cK9thjNKpluA4B8KdIABnj1rLA82AnnejT3NkPdgostyIZkRcyP0kP27AanF93KaU9o
9IbqrD/N/f/2jq6fWyPKTB+xo6Q7LE4AJs3NnoQxsVgGBKvNdRso+R53tNH/7lsQIo/xRK886sKm
1RJBm/TgTCC97YKMKkRU2z5AXabvf8LAJrIOs7/xGyd8xY1WrIhr0/KrK/rgA2FHEy1RsiWVZmR6
m/I1dUrGkdMUJ2SJCTqFLx3KQBn5B7dqJbLKrIqw7hTpCrIAlamGGZ7eNhW2DI6I75K8ASKi3Eqi
KqsWm1YPalGi8ceKlbtcbaKZ0MpHZXbxuL6X/IDT8cxi/RQn/9Rtai1BN/FFG2wMQd25JogxDhSx
pKhtfmT8QPhfP8u393u4WJFVKiPnCOEy2szoNxbSQoEJJyU3aYIw0iEYSlIadb+/fNxrlJHJNrep
ncOgL17VcIRwTcKFrRjgPSQp5Z26WwDeIEJXoBc2WnErlFeAyLVqT94nrE4QzwyuuDysUbisakXS
oVea2T+3HZt8K7IVjG/93bfLyKcuNlejoju+foWLPXd7PQW4K4hb4cCUI3bxkKoMXlmVaqQPL6FG
nKWaqeVIGSi5rTSDlZCpiuUHCui0d90frjC9FVJFFe0MAkmQi02g2GSkSkn2QwLKYXnHboO6N2k6
e+1wBCtNf3UmsbXecdOy/Zj4+wM74wWp2rjV/b0/1MGWaRAkJ3ljbU/Sym6uw554A39CQiNcmaMC
rIN6Mlh+3Dt1wsdZy6nAFzR5pjtC57kp4g7LAnYjUlDPmrSQJHLIpw46IxoZdXHGIFUOwENJljpw
WiUxjLMSNcbszPvM4Bpg6TNPDEBIGsAKpBSXvZlSbm+1slVYzr5ctnWiWzEH1XEAxxBw+X9GZboe
MB1OVBYN7tIZUMbGwtWKDvTVULR648TbW8t/geL8JVkYN8/ULDwMD3iqLBylWxAnCCqdspYJUrl/
p+KTYJhbuiZcJK+5AHVhChSdr9OuyO8cEZ4THE9EC3jdcL7SBGou67U/MdCk5vmDHdUTiToH/OV8
TWjuaejpeP6ZNShI6P8cJYTzMXP+lpDviNY09Mh2RoheKfzVPED+PbpS85Mum+0/sp/shqOA9PNb
Lp1Q6usr6PT7Bg3p4wdXLPPF6Urs8TTIjpZ8rSrGLS8hRMZ874dHmFBA3BGERZoX2R0R7490/iOp
QDtEKcIUID3PGK/8jVQzbQFyTkZtGHgO1izXMy555NXS/GFxTZeSTGZ2nUg9ITkMOZmbDfannu1b
wQV1iO9TdKdbG5YEvboj/FMQGY8VT9lSQ48H65+FIznFfy5occ/KmJT521dx3ds3YC4hVRQnTWn3
CpybetUrtDuRGulPRUbCorHXYr6Peli+lWUjdoXjtkqvo9iHpIfUgTjGJ7SCjYIFrXLdzKkf0cB8
C79WDpXcozJ305rcXQufvKmWGBk+jj5ER6VfkSoMqlEGXQAc5rf7/x545Sr5pUW7JdbI/y/KPfl0
UXm4U6LiiL883e109Vp3ZyNGdVV0jLGuMDh755g0sO6KkAlJfNqRSSoBfjXuhnRYUhoTQhS89uj5
8qJuq/mo7Zs4EUF1cLPrHjWTwqjeDLfe0FsmEiw1W3xYIfnsEjzPwv1hFTHmjM9XKFvhqVBlAbFS
lMt/rmm0UN8nA/R+I7dZgPqFvGq9szguANgD3ebM1F/27jaOHuRATrMsmPvu3rDdW09lgXh71FY6
SH9/agCP8x/ZGfXVfD2tViWHstLXrY5/cfS3CS1vW0uEmsHFM5QrJwx4bDGNaJnursSMchq1GiMj
OrK7inHJ6ZhQ4a6w2e4DjQX7vlXgE0cavanvN6zI0ZHzD/3HudFqPwR4vZrLo2bFjMuZ0fwVwiQa
UkYebvFHpgOYJEpulFev7YdPy/VSb+phLXOljx8c5NN4Br9N7lxAVJf2op8Tc7NbRJbspJiPl3Z/
O39nqSvBcS/d/fNPOpoyZP3tdslWmijf+UqA98n5ScpXsM63qUZmcTMgrvv0FrBAvulqPhxbKIhL
9StxTfQAaxB2y7DG8jV35bVby2C3SPpeLL6rI8QeDLQpY+hLhDTcIVKA3ssyVdX8wIowocx5KB2M
DbjAsikZtDteOxnz+3Mg2mYOgwJ2CZ/Xifp3VOvJChjOIFSy5pM1QCxkUp9zXubQsCP5JmeMxCn3
mJdFxXyD6t3k5ADIIBRAhgLnC+SodSgTYmjoHlEMR6gH1R+LHiNWDEHR5bdnlfQE9qLJOOGV3Ggj
UFwMrwK4CFI2KcVt7uzUEZ/72o2e6L0fmYDSs+d07wo223iF2DNycNW9VL4wifHX37sG7o2LOdWR
CWW8XaZaQF7s6aEQ0m0A0FzHuebTBzzeR7z61h4/dWabqKXthjJr8/eczhYzzBWQyhDSlRNmvskd
j4RhvKISRcTt5Z4qG87/fqkrdVvSQyHHHgfGps+M3xDrpNukONJU5/KiNnsO8Nwc55Yj7m4RJWb6
SgtHNXRznVwQDecCIwv+C0Yd4qftLG8XZkMYkn31dwu2iwBo3iEDY7RK9fXRgRWkQIkS93+h4wNK
mHlkg+fMAnUgKjMVF+J5EqctfBQFZ6wHIYv2Zm4auQr6XAQiNizgi8yKVI3eyjA0DT6+/7OPvLOp
2fUvz+TwvPiYUq3LmPH+YByppmpINNtAxpLYrTcVbcIZkvWBdDC3C41yG4UKobJHoF/bGh2pjbZn
XFHKWzkUh9z9naSUjOwVt53nSln+EaP4mKUhTMDTiigZ+T8TeWdv5nBxLWdYt9LzTB0oEjEQwdl9
0Iw9uOJPj5wy2k4Z4CrWPKx2iG1kSe9hDT1Iij1mADb2CJiDa8Dti+DPxAo9hqBnVIlV/hHN6WAI
vH1HEBM8zaArHlt1pP8aNaHJpusowD1ba7tCxtHsyIYrEKmFor7hQMlZ7oLnM120tWTNJEZDdFsK
Ys7Spe5CQ/drPM+US7YVu9R+9PODBWh/CVDaLc9QumbWJ6WMVSZZXiFFf5mt5dY4AQ1sRERDLZ1U
pVi5OlgDb5BR3o6GCvrmwO9kUhnJ+0MdbZ+2x8BJra1LRl9U2ixpYCSqBhr7/9ybkdQFFsvhMhhd
JxnUbHOtBAg8NAZrFdh9Z1MPUPHzgw8dmKmuo5j2iLdRyImb+s45P9RG5cSq8dy1UyP1VQ3+4RxI
FmrfejHHYqO+H0kyBsRGH/nXCTaFCX9sTw5kI3hxpwayEPO89U/tExjp041aP7evMNLpCJIBrbPT
PMsMj803izylQPiRa00KYlKMof3zhaGlN4K7WkEkmqfJbahuiyv7s54LLH8gh1io7EZvWZLy9jV2
FFVYialV/9BfZ2iZQMxijNfP8LMD4EF09aVM9Cn1Poy147ssE7wgknlMZOkk8xcPFkp0oR1Op33u
Gt07TjAoKA4w6t+DpZbJMIfo/dSMYpWm978GbZXj7hWctqcrlpKbdyFPomZGnUE98hHsC0R7rW/5
6tFdVwGQ3RB5fbB4H/xP74VNVxrrkkx2zM66OUHj+sTsZdNGxj2SfrKGIPW1hea98faDFRaeT1Vs
Q2mzjgWZdM/M0GdPrfpG+tHTaOs7OeHnXMQ2lbJEXiqHSGRMQ2i5Xf5Zdr5ZsFoec19UoZahTHc0
9GKBnDXqPA+/SBPgIK307j0r3DsSBsgIGf4y/y+s9igJxAo9NVamQ+UfybRGsxCztj29PCx4nKBj
JRArWxJEkCStHGwZzeMD1d0VF1SzTGPPe+jBLY0WwM7zEXPhyErFNH4E9lq3wgujp/tqlcv9ufSO
UE6wrnkmhkFoGzkcTWzqskWippStVuakMxIXP6+f6ZOzec9r7uxWlKhQpca8PaaNCxEx5PV9wvoT
VwyrrlrCkbNMW5y49mXGINIvxYOAMERCdx6O48WM+BX9Xls/jqrNSzRXa2EtrrVy65f3HIvjVOh3
4Yud/Uc8ugMA0RD2NguImFL3lV7eKDcVWYxnwoBZ4pFrC1AKyaAi1uhGWA048dx7mOc36Dc+hfSs
lJwYBCZ/G/5M8/QMJKdhws/T6GpeEZ6QsOIRjH8R6ItFXQicUywYbyRHFejIFqBbmm09HMOtiXZX
RU3JMhZhW+/OKHYJ/MgHIPZNt0OB0+5NoufOOrOxZCrey4relgUD8c4rH4EZJOQgM1z1d5AtpKwC
OhTOpV5CUX6xywbp/C1qpamUVF29o1DJaT00KzgYK4h1KRTCbEtx/hPDN4FmW37ZkL3x243nE+Sm
YleZGMmHgBTBWw1SLiH5i3e7z7+fpWdYNRNjJ2r/OeAA1+YcgdTIyg07bDzZxtof+S26gT48BH8o
Li0c52jdTGolcICF8F6Ogi6zhrZYToDy881OOswWxoavQ67Fg+qk3zQpeDRt8PLQw5mK+HYaC+bO
PKPA3h2mElj5123p/117JiML6Oxd+rjIxNiYrOO3hQUTB/GDYtLVYdz4JZM3J1onWVPVvsEbHH8q
0HA5EbHHYhrhsKL8jmRip8XrxXJbCi8hm0dyHO6omBEGSikD+Yfm2+Lm/yZAXIJMhPelfrwIVIC8
4eHqaGL/TzS1f+lfPjM3IYefh6Eq6Aar0P2KzLFcnSY0nwoslMHNIGI6MNpG5pSA+6zJiurAs3Ke
Jfw5gxqCuVEoJSZD/7UmIpOujTlXRoYGMOA1r5DFUdAnJ7g30eWayPLxDMzXvCbu1oSrz+sY8OfY
sRDRIBxU8IUDqMDXTioijx/luqJUU+bR7gUQU+F+KPYaEQGRZFBthKsuw4R7fbsd1ffbt3NGPozH
3wHqYuQMGTEpmqDlgh301eBNdCydWtQIu/ZfMBKN10sy6woJv3REX97UiCrhlAGp+VCwDLHkxE7v
j0+NsLfmUZ1C5duHL23hhDrVWrPUaGwqd+j3aP5lToB2W0Fjv9r7hC7g8g/CFRzqKrkfrPwYtFmW
Rq9f/773bbEsXbFedtX/amkNhJe0HEjfzx9e4dQ90o59Otu1lN81DV2G7MT2veIddEVQYevV3XpA
iq6D+u0wM6Rkjt6dkyWI+NiKU20XX2KOAKgFvBQmxoeZWQgnoKvCbKhW77KRQaE1ZKe9QKd+GFPW
U/xsTnUZ9z76JANmswyp/Unt1QEnJVEWCzon44eS62+yif9NsQ9mZB+fTcBR1RSal5BgbircnTyL
9TN+vVsAXQOEnXOwLr7raPj2RpKYJ2JS6VuZQBzbQJEQEegFnI/nP9RDMIwkn8NQkVGly8iLCWGq
8t8sx/vI8VjCDMORLAo0SMCNrkVJxfSwNIBynozaT7Qwd8xVREn6fgF9sXkvCFFdqDGUdAdD/oXs
zDrNyPVppuvfCcWZsUxKtwDRL460GJ5IR004y+ocQXh+iceJm+vVlg4TDE7PrxR0iwI2Rec50lIk
XVJW9FLAbhWi+O3q5Go9u+Zk3zU3j2VXpUBCl8/ZQPMQ2jUXxfvmeNPsc68AXKsxL7xKr4P375r/
EMXkGT/NGZ9qxPg9wGWemvPIyVe8Dy50TxuptJ7i2IBOcBIcPCbCO9vWo2GK4ZsOQq7WfuBNI73z
X0AEhXGR8PFe8BPNn05ZnfLdVSxRT57DY62W4kYwugsQA6/hvQ3FaAijuCD0S5E5t5AyXXrnqakh
/HjOp7YOt8AKjHTD9HMm4SOK1KcusWcJDkgmhDw/7fsyn1V7ySXXhi2pBD5zgnZC0Db6gCz/zjgx
+lVmZiBHvZ59LVIcCdzZhAWV8V1hJvWcDgNp2ALxc3dQhbvdiAzhq/cDo9aaFa/7Bss9P8iDBfup
SbtE8pYr3UbKw5pblNDOgGiaJocVf/1MB1KQ8Ynp3X4dGN0/2o8HRrSSIbmmItxSlk/p+zVjsNbL
Tr8COXvYiSzXCsJaWReMQV0gDzhemqRVTUaN5aOeh7ft7PcFzYH6IJbxLeYsLT+S/doz40FTD1qc
XOrqP6hx3v9rL/ZFSZbT+YsULndTERVVvOb+cxXYqUoHHMHoWj6Yy6NJX71Qg7aEzR0kasT1aMhl
6n+F63JV5kj0SGNBMtHbH+XVSU3weLD60qvNXk7AC1ElUec61LtQ94beTqLdaSE0fmg34ol4lsvk
9xvpA/VLo291XhIQ5fG7LM2niksTIPYj7c3AejkS3QRCXjSi14vlUWhOBnLWvGpMpbM//WMGL//9
pQCZZnvQd8jfGfR0P409PyB/wto+OpCyAAYwcyu9GL+ZKRl4lk+nF9fNq40MnkX4x83Xdf0bS/1I
x9nlESgPsib0iv8zANlnqiOx+CaH+SAVCGy8l3u38ssl3nHZQ5MUCA/IdUCXNGBFlAaRBFAthQBF
37I0VrjskMYyAxgtONhkFqoa4ReSpd0j53Wpn1gB+REgSzYY+aiY9UVl3Ybs3niZFpU6T/Ix3YjH
VaGM/bki1Zs0Y6pq0xS2oxOKSVlOnRdO44gmZDVg7tR8LcLuG/cKt3t+5JyXdezMOI/0ixDnEaXv
NzZS7v8tm/De/GS6us2NwysHBD1iYPWlRTwm/4J2hJvvNAA43M2GqivMKempt1mOmaPqZ1u+y7TL
zbt48GAokADNqFkSqwq6JGOTL0gZE0OugVB2hycCHZWYH2KYk4ENGZYTv3TWW8BlXFlw4R/rvso8
hOEEUSkKd2yYrA0FORKW7OuLP3V6VJDZhy8ISAIRxSszWwABs0l/60iwVW6Erdw0MAKzAvS0G53/
xL53J9yM1fVzntXq5NX+jmOnYhxTzgkdL6OKkZf15397fNwNzjhKB44gAWBWUmZedzCkEbRG6zFr
c6KEi834pwDPlmbM+tgkuYKqTy7Lo5wkMntrl2te+NY0syMfGx1IsstBzI5DxcupC4dsnzN4Ja4y
WYJlzrRTwx4toB41Lq5IGyZYFe2qZWjLLetI4XvJ2UnkyqWcdyQfXBmxTrOA6ihKndBhh1L/12ez
5+I+5oO2x4iiaHdzZZJzMnA1h5IhSjxbcD/fh8JPYOAY5MVvbnNxkB5DZe7tnP3g9a8wnE570GJm
JnMBo2FeS+ywBWUGU8xd0LLbDzyWxJLeO5W4aGZr5X7AGnjUxjd8vqtXLrUDdkBEvfqnzNCFcZ+U
nqGW4VYfxN/SeqAJNgiXzvc/V9ceciSqYCDXUjvTPqJi1NeZ61wG/v2C2rZ8LUa+W/UBcXcCut+3
fo3jEGZf7V9WH/l2PbDOgt3FFGSvDbOBzmO1R1CKqPnEjniJ0DoByYoLnj4J51zHY+Ai6J7dZzzH
5JSsupkuk2i4SvCaJqlFq5foZY7hUIzkU4PlTDUBdtwrQSJZBHeNIjp1RQQs9Ma8ld4Oq7ftaSE6
ycuDY8CywYxc39hNvuHKeNmmP7mwgzbDAQpZhzs2xg8ndUH2LTvJYsq/mV6CRH2p1Y7NsC9RI2SG
nLRpDzg3a78Ugprg97WQxM5oHnBQFcDbILe3xWWADypUKD75LztAney+22XBNPUVhB+/3RRQz8/5
ykvndpKaEXre6DB23HbGmdHY/6x5QSyC0uCE8VTgAbDR7Mn+yFGm2fnX2LNGrLfOZKrY7Ueu9yX+
QLvIdJVq+ElgAGnfOTuH0daA5IljRfgM6Dh59p49tll19l4mqmngWoivhgxJoSCjJUBAo3fDqSI1
mPO8kdvd/G2GWF3OoRuz+jsdlf6zvgvAQ+C8y/TZBqatmbbZhvU+FoQlHbOiCIZ+OcgDpwJrwzC5
T2hEwMOtEUVquXyGtlOqkB+b/fo0Fsw6aMgpIZKaft9b3PHYBveUMNld0LaU7zuwaZu3vA8wd3v1
GmgURy4hUDFCpQfhy/HRNqEDrN9h7imvdY779GG9WBX9hegf+q8+MCTMxF1yw3bWCiSYeBPevHec
om4aJmT8wfmuq0S9YXfRqUj6UzkgLji4hbkWXIMfYDJSri5DWL85XlIXJOaNR1e4dknMgLADQFNH
fcYU+8OOUwtppU6becV8U9wnW/uqsU8DlebWygoyiFVrqqaSgjOhKPUAZcCpTpYZGw+3P+oht0Y6
pUjejLTYUrEBch3ukFyGxtX4v/Bl7mdC0gKLvOHj5CsINN7DhHf3ltf5Zy8CH1IZfllny/9q8/qf
cOCJDugDKB0KvuE4b5e1Y5lUc6WuizsNi6FGYOhC8awC3VQRPDp8Xr0KJE1vZXpjf1Euk7scbEAZ
gkAzp/tYHJLFe1namYLnq8VfQBUQktYtZdpCN8vI3JGx3EWMigX5tNxXepwqtn9nD5Y1SzgcgyUP
ooy4pv5uDUwn7Mb+swXiVxf64srJ66n6sVpUitTPiGFuuNEDSjt2iyUit3cc6UhJnb5JuQ+5w8Gc
7IEqpuEfw6YWNnclMb4sLFcNo1hXGkhGrlSlhiWa4kMPgXl8Xi31qyGQV7gJ1O/va5HGGJ9Mzgby
SP2JRXtrY1wTsUUjxj1AYVMjcb9PQu+VnOU9GCLV3LhVpSJvmwxpg1w5s8eEz+NwA7rKgq/kdros
gzyaUMr7LYqSJPqP+lJ3rYqAcMEmYtM0T7ehOlvy+LcjOOJ9cYAbVSIb1zNI4LrnJalGyEwO4IdQ
DQxvjMCaFi9yRhSV/82JHi9NMSAQHe5Lh4BoyUYfJ8EPZi34Bnim6dmbzdcADy5L+E1U6Fmuu2no
Zr4pWhd9CU3PouDbn3ojYZmwAwzYlJihKU2OuuN1r1xYEKAoG2kt88AxGhhuF+TjWMx2InWse8ka
I7V6cisnyS3iFAGlMFhrKgviVFBb6dL/l5cSvX11yVFJuHBnwG9an5zXe5L3M9j6a1nnXP40vKMN
jdoz3GpwwCdJT+2S8Foed3rLNncZ5JNbllWj0ophN3DKy20KjFCZEpikW7/IAEbqQhyub6YmJXUx
uSPUYA/mSBM+5E4vuJr5tPYqisk+KoznCuVhl+qRlDp+fJ6tTOjYtuDAZPM/+BR2BPygEbWJw3rB
5FqXMtn6IIRWyXYSKeNwJlzmF7MUN9oHRtuRzjI775kcET79+JX+x8/vF9kODJxRqSQXpqXvQJC3
p3SbPXigTzq20iBgltXm28lInil5c1XpXPK9fgV2wRyUsXh8g0DaXBiOA3M2oY5B9EVvXxiKbSgr
3x4XAi4BPK08Tz+4Y4kiV2n65lM41fxdWlv4gj8Z0K/hedr8LaSIUmNrmVpf2UYebkP5kvZusT6U
vdveB8kNIHMWfuoWp7fXHbTUFPpmZOvoJofUSOv57LwgcGMpnSqJehC0KA2tBGOPq4rn09YKPBZS
a9CYCyAa20tV/J9qEh6AJPG3LxsFq3AojQi07TXjH3t1AuWDMWXSfXKdSWsucZIUPIP3B6+g2iQi
hxC8G9YXsVmdJ6/JBPXyiRdxNtEfJ8GZK2jW5o0BB7Eda8ws0oQGPIGSe9StzkRpq579GyZYlwvs
reNPBS06B3kqUnM4NLfzMdbtk5+TFCCQhW5Hq9Lt46dusSpkck4+ODyd6ExKTEJnxSoJABcNLzqG
9o8cMPuh5n/ffjaXcCxRS+SzcsML88fFc3fuS9POxW3D3YTlZFL48450uhbGBWorUTDwwt7lhFYx
JB+XZ85UlATxTKG8J94IXDnYlGEaLddkvDX2mFtwZYDZQKDXlnY/eTWp/d2rbgBGPC8he4y0b9aJ
JlvEyy7/S0gCgrDGJDNORv6u0Wv14uNItKuJJ4MoBHMkCPMUj1DAbKY8S7hGqS/emD2O0duJfFN2
H3mL4434tYnPxLLXH91GFyZRJgnVHgBQFLFwyv8jYoEgmFGoARc2T4++6l7kYorfCpBO+CbQb1Uf
ifu1BCAsRcqcqtGZbyr9IOVjP+6lm5qAS7ddGHTHrsIsnXXEWMo+nfXIwtsur5CQeLCITSqX6aCn
a+eqw6afY06PpZ9fJdYZEANNcRN2bK/bAKH/aWTD2GyN/JELJx+IxqFbKlAu8cHwYZsZsRIk1Y12
qydIE8F/kM3RMC5YJf3rOjjn5ZSRC5qUrVgJBEqfZLAgV93Q2JO97+oOAxlYfKHQiEPfH8cXJ0Ay
xjpe/Och/KoJAPFcCz2BuFnl6WY1Q3HioAd7TxA1kTCa7WomRyZtVDUl+eY6bpTp/CmkPKq9Dwza
+MzK/6Uso6XC/AWaXKufVpDf9V3Dh6Xy6RzDYNFKS9u3a+FYcEc3TgNjJEhePpzjTGQhdETCdG8A
OW26VUqnHlbdkw830YAnicGlTicof6Tm4l6kUdtTifJHsp/ndoS6hP2cpLdhryYr/nrYF9jJMrZW
GF5yGoh3TjoFeZ1/qZBGJukTN8/Rzp126fsaAxQ58cMhf5m0qcWfeI20JY/Yyj4LJQk6WckAeCC4
TdyUXZiL9aS/Xq06RLaXIiRveEI8aTmDXclljOaieTsEkaEdtKrLHpBRw9hlryMii5UIgeEtJO9s
dLgQp+8bzhWbPBN+86rCe7fiKIl+Sw1tRjw8XIJv4HJCN9Va7q9ihwVxTjaujxzHjllDhNEiWMJE
GZcC9JL8P1NIq7CU4EJit00D5p1DTjQaLrupvgrXc/6wwDEMHM2D0ALW8TbhNVoI8VGBk3gtGaDf
pu7VmeWTxX9IwjYE6l1Dn5KidYgedaUTxgCq5bk6AianCMZG4SJXyK01R7fpwda9CA2bOd7ewku6
3WSZyqzcivY1CegBeuKZ+mH5ZDSkCzWQZ6iwIA3BoGHjnRI+1rsnwuWCjWKUWIrhvgfCgu8DgGD7
AqOFqZ95g42+scuQc/IXtP9uQx+wt1ir+vbz7GJeVKll49hSrb7qx7jLUCn7oKog0r4v+Kfagwjm
uOrjKbWgHEuiNXDiRdWdMkl0Mw14ReqO0KcCsMnbJRB4FBBnZPlPuKrWJAdVWrgoeQXmMdfHZEmR
SYBMDjEPSYvzSuUPqxlrab26YqptSnjDYiHX4+jCPbFdxbvvNw5KG6oebElda6qWbfm/is2O+bz/
hrbKVo5fF3AO6WtReuM0ogF0+SqyAbUwSFKQN/nxmMfAkrzX/yrj/Eeg1C2CXAWeOvPHMdWXS/Is
tjo7TfvyoYOr1lpyJ6bWeRRdvXsk9DpZZ1+Qd4z/opy5xZIK1etawPCmCgtCQHkh+kcuUKK+CQLa
2FvzGWHCTv6Qy7WOvfLkZKnwdTfoBSfQP16A0k1d3JrrPQSsSaD8DFWUT+jc0GGI7My1Iz4ycbed
b4boAyTC+NvkuDJdEZJFS3EDWuG9bH7FtMJQrctj+FAV1aepmTERAG3m5NgPmxDhskM+IvoABV1z
zUHwcTh7MziclB52zLdh5BRCXTdNSzXzevvL7ZdTj0xVMF/rScXTVQAYna3Js4r+9S0F5mJi1X8Q
5CSj7PnLTSc125XfQiPCc4lBfw/lW9fTNrBN3eg0ZYf92bm9/1ycXclYClPO6NkO32ndqKnlKIqK
JIFnZmdSrXFYAxqHB/xlUc6vvHNNyR51bYUOYOswVm1QD0tnFAtXiOk4VzYlTaVa5ppcQV7vf7TP
W0exc2iMRLC146XeSU0felNta9HiRLZ7fpVE6f15HdBHOXyUWa7WEa3bgVzmW/mr0mdzV+Lf8bvW
nc24Vvyy/zTT5Nvx+gNqQdStz8fsZHf5CWHfKWUeY0wy7LUCjZ3Y1M8m1Jo3s2tofp4ubMIMm2J1
nhJ4rF3AtX87CyScbodRpjTjnRVBpuEjeNmY28c90k7vEgQxw6UUeIOvI24ATxgR7LCLDg9SD/36
J4ZwH6/dYgg+OPynUg2SlUR2b0BHQcyJBkQbmpF11TkNoTsgX6uT50Vj5iwyHOLp92OuoyPTxfhA
zekE/xEUWjnNjJTzpo9yKTG0epRquuKaOGHNVQjwBHnj6sszPtABaibT1AS2hiCvHL/DtHGT6r0T
E16cXYRovrJwXfBE30cYf0XtcsoOrl3dXtr8N8V63JJYAB6oCj7AdLVxpeY9eBKbVZPhFH93Kzxo
iP5RqRwRfbLvMP67Xv3VthfQsIT+RAol4Q8m04PBRnIuYI2shbn+rXNdjLh4RhqfgFLo9Kj14cjh
FWGKnV3NzhnzcO1DyyBw0fLpD4tbfPFk/jjehlNr8ZDr+PwudHmq7FyRabyOO+l3XYj21YCQfAia
TsBDNEv4kFJYFYDog5dQ+eMhCfcPih4BPM6Tet4UX8MtVKwONodQ9UeJeZYDWeA0TkPKdppZ2SeK
yrs2IrAAfHja2wtz9Ff/AGzLdsun5iPVm4akBSEI/UW9AHRyy6JBgAaq/kq/eiAXs0FmGEm1idKE
+TT56Qazwi0Ubw0IqwxRlRdDaoUlc9NKcFNnDbvWarzsTs6JVo+ZAeQTEULJExdHhJaHM2n0XxSW
ckplCHtJjtGJZZjAR1FDegFZ4i3ChW+30Bt4dh7RS/VENm0gQQ3Ngs4+11Ph8YckeMufVsHb+7pH
A+LD8fE9A3p5CAyLeSDOjwvG1WSoByDvsjO/iA9tDRo92N0DOph7j1yfkRJTJo27sqwQ/BRuh5qp
aaFTXbwwDATJmyHdq+5VXIceNro7xE8MnMeksS3RGJJgjqPi9RXYHK6HTia+FC7DGKNXY+ySQyF5
eBRBs9nMqewVy8pbpXYxkDRs8ozNrYRgqZrNU+JEDRYbtQxeyLaWnNrgf3gB0Rkln7Ag3YrglIgj
3r1FVNnqARIVsxpOcXBonnYw+8+ujvcWrIvd0vt8pvfUFnuKxJpDviFN4Drw7vW7mKvgS7g9kQzy
j7tic91LOb5NJjtH5mjdWk+hYIrwxPTYSHNBNb3SbCkED+TUUXn11AHXDqU/68wZEE+aKkZoipj7
xo9xJkMmNKT6xWuBk2kwi1adc27WjP/l4oxLC8wg+kakTHARBIOFNvZu2r5QMOs5IiYsbyuvmg0y
VNahbBfMw1Z9RSa5Z6okZck5U+PH/p80tXVxOM7DRgkWOKQ26l8GUP+4HvnnlFTDf9Vaogo2ZnT0
IeqNhkvcuRFVWdgQPAEU/msx7yCdDhQqaFXnzPvKLw8kJBEqDRN1u1E7ewB3Ij45ygaUHn8vZBu1
hWKwjLLuDuWLCPIfgcKZt/jgZqE+NNl+CNyRpOvTfl1cvV+d73T8xr0Vrd9qFbqUOvqsyITxEfkO
Rgd+hu0iPxTwAzFJLrWigkRxVD9olIHrlOEvSFxGUExoy+0uWJtuhkjEX3GqMD3itCsszkBt+ZvG
9Nn8ZhYiX+mqFxCy7Gln0TfU/5Xakors4johTxmSPW3VSeT9O1Pp8O1lXPILFgFzPdtf6/4S1lKF
+30XPSg0Q5B3c9nFBBwEsNkF/ywnYzgtuP6IL04fT+zcUcQ2TgdLGdfj+q0jX1LRLzX/E9y+o/jO
uCfrQ7HH/56ehK0wMorVBd+bCAj6EVbN14V8cGcvhnv3AAIidugagBcu1bgLopmhgxLQ4Rt6sMTS
H1WD2vwVXaE2uT/voQQ4/xMuNLfTXvV7HUY6vP/4bG/Z4v16+iqHTLVrETuZDxQ9Jzjy2sFqjzt7
DyQsJeSE2kJO486a2UIdB/zvZpLuyZFkcUFw9Vw+jif9vZNMfw8W2wCT+zhZhOH7CearmhBL+xGT
smix5zcEQBSyOJY6xmyJ+bBTh0X63xxA6FeTyzQTCsHvNs4zzCk7Ymnci0M7Oj068FYzhdpEBm5x
vt0yLopalJZFIFEq4HkmIDpkvtFGZsWVSlgBo/mF2DuVFBCF5uQK1iYbP3Gj/6OevPVwqoph4XVH
l4WZDsSJLxvcKv0i075Q0M3jQisYjh8UJ6FVoVhpk406BY0Czz/hGpxTrNz5mD5/WojXdNy/46o/
DANHXDn120tkmvfuq+W5UOaOInVkMsD2M4Dr0fWTXbH0jhpPZwgZRqQQurx5kcJ9JOJDQj2OuTJu
h+d6DZMbm/7pn6Nzarh5ChzFdtOQbK90948IADYuYDFQIAsw+zi/MW2EsyrtN2gP/aInldKlRCMG
KbaSGfeZAiQLkwwA+9+fmax6YeeF/wLyaylri0jpSFbOXUtDzEb8LS7U3/KzkXCirh420h5By3sL
mCMKNZ9udW3GblUjHXgG/FPrcMketHbwSZW+pjfcww8K2QhMShSzjtfkGQB6sUkzxjiqMCwkwDLR
wqw5UVd1AiSl9CGxx/Hang6xUwhXVKZ6Hsf7NfvdFr2OCHd/bG3VzG5hq4bM9hddCvc5UDfleIku
IA8R1efnfjfFnabZB9QkR0mCnwibRcd938hHFtJWjNxN+NWMGtfLWFn0TUFFgXlGjx1nPi3Z8S/c
3jvTWYaBRJs1QCP18K83RO/2g/iVSBu43tDL6aiWfXYv504ZthVBkbnO1B2wqErtjayVF6Nvz2gY
xVNHIT/fgj9vCCYiWqxHZyev6JsL+20fmq0EtfZTgRovbVI/g48O8wvHUSyqB0v3UqN19D4Fu/ua
KK9l+n650xfKaJoSOdeXKatUv3R2fkEZNnkmTkmVFvQzPZVxCKBjOgYAhYWN32JLq46McmSTEfz6
4mne/sWEqZTH85DsK9JOyuyffFfhbS3QGKL3pLWQorKAFW0dF+bgOJpj6nsJdkLu6lM+1r9XCzIW
deYaa9WBvLvWtoK+MgXZFm3yGYs1R8f0VWOQhjgMQ+RlpZda/hbct415wNGawtf7e7Rk9cLaqo/I
Iju3DuK99Lpi/IcBupKNrPb8QiZnG4gk2lj6VxLW01xHN+aQsDqEOFTs/PwINoypgj5Fd3izdaNZ
9BzNzwe++eP0MfKW1TlhIwchZlcRaHHwgdM8sSOa3JYQ0B92zsDknIKbdFfpafTJhPpV/h4mBmjD
AWMK2zq3i9jc7mtfBSVGf51iPitsZpN/94HaXx904kTnnvXfEB2r3TUcryOTOGIkMQGmxmKuwjUC
Hmf3LwQfz2599eLGQYD1VWFj6/RzjQdpNs/6TcxHx9sd64ZQz3BcWcUXjautZOFNJyqItVBzS7g2
ZlsjJKl/dyesimD6nXfZWWw7xnbVbXsLJ3eS9laPMWu2ghkWrGUSTPFgduALhR3PJb9W8xOooHP1
6Ug4+Jsy3TsLSzwocDyeT+cPme7dDeMqGET+hXX+gx4VhOvy6GnJdhkzXJjOqbyxkUlvfqOWFdBJ
PiFeg2W4BWBWpwtPOZdQQKTRSa32xSZiumwNbFWGyR3bdXwmr5vqlkF8zyL9YVTo0ADCrNqeQBwq
w3Udd46l1eWi4/5ZmvtMdL2tJoQYSoxlak85ZOy4VedvYSWZiDpYZMU4Nbfc+GtnP0avqS+u7GCF
Ig9CSwBr55dajmIHp6VW1/1KJlq3W23bCQgf9lqyUIQ60tlXrPQhiZ5hYr6OZ0fOpSaCusxqTi7P
hEtjsI8CgwvyYtHm3AIvtV1yVw4Q27S2kUn6Im82P+NRASmi85ZEArBGGCNwgKuwktK9Z8UoQiWU
giKol9lJUJnLpimu0+iIKvZWiZXNa7g3XbyOQcio7Xe07rd/v7v5gRmJ70tOQwmh9iMR9y5Kab8m
cFrn5ZP7qz7CW9J6x1U7ivZHIb42nnrS50wFX8kBhTL/FqrMdw8Pjv4ge+GYwD8h9L1vhq/AnLx9
ikAq3AEgYSMgpoJ2QcR+pIA1kvlx5/pM887Cvsln5UNmpHui7OyMXPmzoKIV66D5WInDxFjgGGKU
1t1fX57vWXgk/5pKu0ER0AYqb77bUoTTBFYe7Rqv21XEy8uWC1wgK3YmKUW6ZAaMFV0Ygxae+kdD
H/yKw1sAiZEtTU1Bd2DQSNZhmVreAY7UOdo1FXRhPMYsIg9SoH8afS3zRC6EnfCPEvw3j+C9p3Xv
OzpwvQsbjYoPUv3FCWcQMx7nCzA/gEWpF/AiGBMoJLfHD3KAc7vUjd/tP76pn+qqcR7JqgAIk6+U
zbzIi3hSMy/e8dOMxXH9sNKUQjCtYMIONFwoH/Wf1lO2XAY/4UucRwd14SrNKgdGPWl1v+fabHDb
dcmeFIvYpIuAL5Uqbx5oBZfkhiyYQZrjNV/aJtzrKfTAFzeZe7gJgXAOn/qk4IYIl4NbbPjuib/h
kMuJrhDIWWfzaGotd1of+20cLAQWul34/LjEOmuspUDbEGFO2/OIruhAqFbLzn5xbXH3Lch5BnJl
Jfaqptr8vzjeRfZ6d9asFrGEK+DG+NfbLzs1gCIPCpfROYMZd2uBi8kOwGzaV41Z05+dQ2Xjn20S
3Nn2d0fBF/euNxIzsMEJ0s6J6iDt9DG9MAqEhvlUAPJAN60veJ+TvMyT2cYE9YYJkmsEtOXdK0e5
iMk9CmyplUc0kSDlbVaykPrTl9C7PqesKuJexe2moPFn1RLDqDomvLocuzqsHeuZnI2cyrju3MpA
BEvEt013vgP098d/P3G+6lzk7BLRvtHW/0hWsdHGzyQByG1TgHsOhcyIkrlsF53bZ4SWGmViAEgw
jQvu2jU2cZWGquIvxsXK3CvU+oXdWNOhBQJEQWGNbRHyKSRe2VfNLc2zv2l21wbl34jf5qjqA+Ma
DeNzOBFEwxbXmn8YvP+RTwR66OtSzWAskbp7xn4Bw8KQiNlI1RdMlV2bUUyVgxp9qE9RlGZK8uol
MSbaPJ+rrYvrpdxxPlb1XR8BIF1pePEtZTs/l4Oszk1FNgU+6cOB/XQ+epfGRo7up+ngU/00ymje
SoU9X5VJ78ZSz11avPEqIpZiRBv4H3b7OlBVXOehEBsJSDVp22ppaEC9kPS6oM3Lq4iSCmgrCCbx
/DNkJaZpUi1UTbjiInI1J9o9DfllqwSHQkT2kLEf3SLwy/CLJ60yhWGzadOixJAVfbsCVsgzz8Pt
mml7IONjvxN/eoBYVX0cjEnWZFyD/MsGMJMl3w4SH1fMbWImplcOWYvnV1+Vs4lJrpxZA0W5ASoR
2+tBU04O7kDuU5P3M+D+yoqLyQvq90ySnsdLEMrE4hmbx9bA9yf5TO7um1uRL7eJSP7QjOaHEXGG
3CSsuG/6jvk8fGZhGLZIUucMv3e7fRdbg3PrfeKy0TbE5WgpaKiB92+V6SJVyaq+IIBHsa3FRlWi
7ipw8uJPWzjLsCTlqTdOgqNDxhvEfxNpLT8aNz80iMNtT/o9fydMMwTTlyLEPHkxR5jH+Oymrgxx
s2vqpNAL2Y/DlbK7LPExCfFM1NDCNaBh4iSyuqP1hOUWb+AUC8tUlrIm5O4QXpBIA6WJCazItg5Y
+7Qxa2cvmPOXvUxzRG58RXPnPX3vM9/XQ1K67w0dC/ZhDvoCVgwjP/ioGmKb3J8AEdm4P6sDXXUI
8PHdhU5AUWeeBQmVErFvYoSMpqMVVDDbDjz0ZnfqDzogRvwdNackKfpx3W8vAYYs0Ew7wOwIFNzi
tS1eHm+QepHyCORMjdAXxNyI9PLdo2tobZJQSHh1ufr+76X78Dt2VaURQt/lntF1si9lbTCqD+sT
H010h4lJHYHIhoL7OoTYxxd4CpQ4PjD/NJHd35qkUOeu7+Jjg9P7InV5WglvChr4PDC8zepSowK5
+v4F9f7mxVxxCFl8Cm/EvCSy3ekiHmQRl6fhmFBKL9wOMMXXW453RfaW4S/Ml0dF6XDqTqI2U57C
AlKVn5yXWPkaSGtp6qJPxj72g3GY67Nlhnrd0yXu+e0dZXGXj8G6wG2TUKg/fKA6+MQyZZ1jzoxU
M1o/S//QCcyOgSef9Qbpr6M8OhW/RA+sO5xJM4Rmic3aKZq+XM1aNfFkTINz3j+lMsDL9qYyW6Lo
ZXiV8FALUHjwnYM2SP7quREwFgfYac6ohmv5z7LGxEN/WqkmCqJvi6pcaOC/viC8iatkviYeF/JP
VXm1xRaKQnO/xzLsDFs99iQ96+U5TGeBptTwFm7VcN1vmbdeB1HsoNogPeoqsY5ydl89zTnQL18e
+INcbSBGKcanAeS7fAVlgrztuJoCqwtJ3RDyqpH2C36zQS+WawrPIbuoQMW8tMd2eonmqtr0pgyP
lEi5kHaJwHCt/gz0OefI5RW5aDkER0Fw1EAVDTAWkT5xeNleglcrwDXgdd94lMTI4dhp/muQVYUG
K5H5eQbTnSfnHq+x6mC5nd0tJe/EvV2Vq8urUTOR73jyb7MnwZ8oVdZM+bFJluUR32ERhuLflZgR
YQjT9oLXY/QeSC70hBvx8NBuaqMUkLFEWlQ86nBkfiynWRI57iwkLALA/fktl3gmMBWYYTcp6YEf
fCxmzbFjLMbgjoKwrjiYjB+JVOWYW5YZVp+nx9SL2Fz8LabjixWIROYtZMhZ+AfVdqKTC9JIDKno
M5ikEcUrpDQTL6rBHbvvatfGbNYLDmLMrqYysIik52mDXRa234/9n127fLl8hKtI7I1Ako/W+v8G
3vqwTD2WKdX0RvUfPTCj0w1OIbNpCpZYUE2Ok8ehQrjqk5r59zn4vsV6ot+yrjzUfg1Wer6HzDS0
OHjz+2g75/K22TCnFBriNK0/y2+wWgqpZX+cWSux1nS1nbz9621AqHNwesCP3dj0oDSIq6D4wXM9
h3zm84BWbiXyim3zQl4riihP5Jw5IKabrFWpuu5ER13A93kSu0W/2WdATFtSWceeZInjeGnmg+OS
G30ISnQT+HsD13ZMFJq53KFiY1jFR0Do2CMWMx1msAFziM7BcsCOFYbRWSN6VWvWl/sdYsixtkns
MRE48kP8Xvw3AIDTH04GZs7SpyHqMJjAMXP1S6iYTVXrQio1dkBOn+KiyhvYJcyb0RjqSWKLk7Rm
ajWuR0Twry9OcOWUeN2/tA9vb+ZJyqkRj6Zu838tzI4UrnVtFHJ4E25OAJkfe8yYV55KiimWv9/h
FAcCKAZZn2Yew/ahH0QNbaiW/BCJD8htLpVKz5tvFEjjGtD6YZasDMAsB/DqvQrPoCmHJktIy7Ns
xF6a3OtZDYFypDME7LjeMS4cZrrV1cI2pp66jGrXEaM2N9jiw+nVZur2kcRyxWLmmAInj133G2Dl
zUACDPTitlHKqoz2Lja/7GvIVBSYSJEb3VsioR2ZKoabdzqD9UQQtFoosiVXPYXfUQsH4CN5b4mo
a33L39catyxIZm7C5pXEa3xVWnn0TxzE/POf2PylbNVO4Ve/W7YINY7+d1P/Fm4cjNW+cNsqv2XM
h6CKVJiGZKrBFZH4tTPYHOIs035kSeoHTcFoYKHr58kxP5PuwQr/BK/plcIUxxahnhzmDDC9WM5C
VrDouTHAX9z42KhpO2b+/pYTL8mwfqIibz4GcbHGJo0Inq7QpDi4ocrFEY7MIjLBq81pL1LUTl0I
At0inOgXXsPpTCae5Eqqq+OBgoYmzDkCIN6Iz2D/woH0DQjDqJaIPYG7SF0kwb4Szr8Kv1Aiwuyt
PLVXoQloOC0sO2yQglC6FlbZSrYECxBACmex/4+lLYBvrYdPXKdp/47wMCjj9Se96qaolP+MJ4ac
+Hgz+0W1/IrPIcKYbA+Flg8ZgO+wofkZwpOunQpaetZjuzXinqCmBk95W43Rjy+kBpxqGJKy6HhA
P8oItO0jxRj8cvMDycATJlAoB9PvnxwUOFGXPCTikPcbSpM+ncNN/B0TKf3zXak9c2cyqBWferaZ
Hybx9zCBGLy9FQaC4iXAEk9jFQ7HmoRezZlSRb8nbx5iFzZ83WjShr0yHZIJx+AIuSa6YWXXaUI3
XDq5eqld9B4TDJHpz7pJU27UP+ePgdBvid4s7qxAdYruutpe3uLQGz0QcM3M2jsEpQa3MlluUWeo
R1KeNQ/LhquSL3UqzgOjdA2ULNeQt7CAGhW/ZDleM5V1IRkX9NXLAD2ABYVS6Mg9O/krYepVnPxi
fIlSFNjLZor9D9VyLxu0lYIFBL4CQ0GiEFneB9segGM/e/0j49xMMkFtBbxctRJg0ThqXuObtgZX
f5h5IS6Mj05WewGAkffyldWeRZzaSeg1EM6SKeL3cMT5HOuBZza3uOQ4ThGFfE0VWt3zn14rx+3G
vxDOu16vrmoxd1chu8+9ch1EC7wSfwj+EE4f/MV+8Vq/Fj5P3HHxfb6adz3oopjZclKhob/yB9XK
cWpnC86u8XeJmJbfF4krYjyQ843dtPKdQl18x4Itmt/5N7xVqosnULKhUgZkhgwzsgng/olfWshR
7bdh5tGSzkElvMLY2kywm5pdNZi665pbPkBH3HJ3qvePYiv69yOHz0riIYVK9kBh0RlvK+yyCfsQ
gUiQZGkPq0FCsPNXwCxqw0MN/FtbTENuuHPnuXyLEpOdqHSAlyo5v+PUmBbpMbXVDnwZtvbJeTpV
N11UrdBD5G0+JUbtxuScNQS/NqI/8CoXvBNi0L1I8CCsZefEOa3nKc361l1UMu9pDI4s9WpILkwp
9e8AyLF93G1jTtgisaG9mjb3MnPLjD057TtjTmVoMEEFuvOUUSYW73WGibGWHLzwAnrX5Nw7N2HU
47GCj+Sctsqok1MT1sRo7b+ZIE0npr+q7A3AU3XEWbkt9WM0scufzq5lLKoJvJkqr6w01i7oaNcq
EpfoCqNGS1xY3A+o1cF1O3GVX5pw7TpxTHLVFbs0wwJCix+JADUpYGp9mMlrrHsSQOunD4vBIxSU
MUurtFMx1ouNo5NbRGeMp4qh/BwVhCOmvWcru4670dG3uJ7Hhbi9bPVNT9FwtFAtzvjM3tmxzn7/
HzqPibyx55Us5jgjYSF6QLB2IpKMFtfr8Rgmop1Zp9p1lTwDcGOmut17H7H4+78y++s7Odngb+4s
g9P22KYUuDQw1i9kCm2M5wVumQR0xJLrqQp/Gp+KIcSqWSnfrb2WxMulS85EfqkBRU+oJm546uNb
+yEZCOSegzlGAAFTBnkHJENwYoZgvdPDf3m4C54go/lFEg2lnfqA3Qt8w0jRTINyiqLwfEdIx8kE
9GP8BMvP/bLmsf87elVlSthDJZoNdsE1GSrqiamrIPhchpwmfkFFMpsclJUkdmWX0Nf4JTAFiKC4
6Nl62+Y7VH968/k84VrmIck91G0KqAyGKOnRXb87Fduz8X55YLp+ygv7yM+cW/GZDYVC7/iLmZjz
G4xfnTdebeld1FM9Gb+qcqK9GOqkmgEznW3eEzZzl26+/ahnwuw2fK8pM7ooWLdkMtBDdiujQn9s
YkFGfbMvZ5adu634ntmu6leYvzx72qLh0dxFXHLhMX7TKwQfua6i5V6Xqms1+sxG9VSvjB57+bse
1Wf3MyCp9CPsl5cOFpwE/6CySFNP5oDqMtb53rbKtRXNQbBulG00gKeqknouRb76fHgU3+xCULWo
EmWL44F0YJE5vcj/xGEPvSUW++NzQCdATARiMH8OR+iwgRoUPnpfcXjqjJvOXhL9RXT+XseUeIn9
3M2l2cTQ+kV7+4vSHmZ5lDDntqZ+m3lW472Qoj5yL17Elg7Ohj94x58+gXSjuNSsmjoypsVGxE1A
6dRGHgUMw5HZVs1TXF9G9U+FNhr8UWyGmdmXOrCbaTltnlaDn+DTotQigSl05iFKOW7hFr/b52Vf
DSYG8iDbix98FKPpyRO2jl6tqtihCYGXoRI3kLRAk2mJX8PI9XL5T0TreNqUNHWX024Qe7Xupo9y
e46y6JU5jnND+sKjN5sCSy26LYxSpNGq714bMJufqWCe1hCUf25WQKPc4ECwZ5M4CNBYjI3tugNu
4DxBZYhr+HXd83Lo1ZfhsyvvG/9RDAkhqTivL7No0tyBGdLv1TWDtzuOEerr6apjCI/B93ozJ9FV
mEMOinwBstbE9PryGJY+gMdUmg+q0UavjgJo3GasHGagfclhM1IDr+soXAj7BaGwk+9lN/F4j2YT
TS5gZCxhGUVw2r6Ghj4J9JEPFUbdHQf3r09wD/RPoG6GIpR2fgtHv8ZmWM4SGZp/ZvhHUesZJ6wI
F940OHaEOKcU6x4rCeHL+7brD303ntaGEdmUye6FSdGmi+rqMjX9wls1UTy5JOROxDbDLpmtf/vj
XuEM9dNSLoXJm9fKSJqJnu0DnG9ByaXi9Lqqhex5p+4pqInPVqVWy+87/CB7z9Nmdo95yWDgMbUt
QMBIb16u5v/MdE/qX+fZv5Hi7UbeQUVJqTs5DmJnmdMh4R98U3Hbq6CVvAIu+EXNtM7OK9f58a/C
KB0YqUaw2jRlsEk0aeik8o9hHjQpBGQ3Nl5K584OVkRl/MSPjVGBkTFCTxg379SBNSH7Y48Um7p6
ohqRB9ZGEfhkHa/nuuTfsCOrbmnzsnyy9DbSzGmx3bBhyCyECEGEe0bEKpTfTv9jFPh8RsOig9x1
DQogZTRs/em48Pyn23093+vcu8djBJakArrsku8VhrjTxQmBqfLfl7T0tulYBEx+1zSrQtoAfH83
uo+D6LVo45UjhwNT7FxFKT+Z0Rvlb10MYRLvnZbxWkaqLqlTFkkUGqEtKxHgVzIZiNdftASNVDPt
su9Y8CI4mCl7Sdt11aY4PY+FjrK8289iHn4IT7DWRICPoUhO8KUs5+plPoVXQ4A4/IwziWxMSQUG
GYdptP9B/8bSOjIyF9+TEbKCq4l7pBBbpD0nmnzohuj1DAcoKUtf1i3bMr0D1ivySpbkNk6vkcpG
hcCAm6WzCay+2qtLQEr9Jj88WRRmN1lu2LuR4Qjr8EEo+dcGvYb6VsGvlOruzPMtHsl0a1tx76+X
sUSlBEI5xX5eE7y7pI3N/FPXawQFp+HqB4e86aX/j3TkMKw9a1v3qSwQocH4dbClRbi+CG/2SMUO
zQEDe0j7A+UOLr66IrGlBPD8LFYz/t8/xuWF8WvbPTm1ICOTEvJxHU5maDqv8PztdHta5baANSbv
r7hdl0uCnU8dDdUIk10+phIsnlVJzSwtQ+vv3IgJtT85eay16Qe/wAmR+K7EvtNkjeHccwdx8DRW
60KdtWmc3eK38CTOHyHz4IsTv0wTwmrq8ew63wdLrw0Yey34/7xPb2+Hvi0BpFBVZl6IzxDf3o0U
iDVohUccTVy99SfkLrkEm7OyRYoOiqJDDz+1vvpJR5gIxBQzzpjN6mBLjWVVCFwrSJSbbr5aoGVf
zePx2LijJgB62FWGDJ5IzaQlDkcBrrn8v/Bbv/w17BEp9Cq6UWm1C9tSNGPr0t8I49pZYkmtu8n/
QDolMLletU6RxCvidbpIqBhbWhaP6bZJmWwkXvukZKWTCb5+fJCArxIaNWs1G/6nfdFktt7YwwMA
tJdy496GcBVd5D73AmOOyJCrPmXPI8xIe0hWhgVAO14SA9Ns47S4hFl1LsOIkOg81efaNNfWS+gA
qQKdg7WB8gIz8U5yBddtvT66j7bvirClTVnUelO1/qPHIMeCLi29A4jLrDg4Xhr4urVn1TtcDyXF
QL8Vx/OFTUKsln4VjovrG6KhtmHbkiyzHDu1rInU//911hLHST++RbMENnK+51xGLVpj2b/I5cYe
Srqpu3za1A75nQc9gIjEOadNhNocj0GzkMl+6D0IpRgPcQEAv9wp0ZCB/5dLOjIaeD2KIlKKzFiT
dn5ZQLVclAcu0/RWmKzl8iPi2ARdbWASQp6MfyYlPxs8Q1yO8Q9hyjRVzzh1wAL926i1e2w+8QiR
VvgOwvvNBT8d+VcJekuHN58lUK8Wn1uHN+ZtIa9BSNNmHlaRznLxuDl7AxguDQZXsBdV1zjvyFRb
i4+M3OZGp0QTY7b5OVhTk+kWkmwrTQhJEp2FUg1iMup9I8HQzGRhJR2SQbSKs/X36pE5vU6Jt2st
OmlA6N1m2EjSTxgVYL3PaIBlRcsTfzN80hoP6MuE6oNlqIkWFHc0XuYPwy8+g/wtVr/oyKtxsc9P
UATGGU4abX+3MIxyz79LIN39oDsSCx+z7fxqnD/0/vrN0cqTmxpLd1xIH170rgKaOP5SQS8UFtYr
uktjg8EeMTM2gU68TVbwL8O4I5lYaByBf7ZEFf73/lq837HEOhqPJ+XINgyXcr+ZqPnmMUdwm/aJ
gTPli9plcN193K47vIEpqUjQplj1GD8Yv+MyNic8bQVJcacPUjPsFNN7NMW2X5wJ68MjKvj1OSf7
imTfynRX1PDK5VCS+beO6r4/LrDqgs6QdsyBOdC2+io1G7YTvM2yKHdUseKK3wRwZSLJLXXVlwY1
R33T7fwZf3KVupX4rjQUIU0/VbvxS0gPK/jhS5mj9NOaC+n//KsfRz2gM5orMGLgQovYWjiEDFr4
D2GpnsRBZHrO8Mqdju7a7z+Fnuw6XQ8R/eoHDlSn+rZpoHHDRYR5/sV12imLkUj4twU5nyXFoNNA
hCU6zkl8jduHuWBjN5AsrNJD/h6W8J/M6O+jgWEoqGk/DPmb+SN5WYCoMFPNC2Set+BF2yIGNQOe
BAXEhLke/yaDGA/HSDbhp78VOOJnBNsFGPoMJSiVB4GsJ5Ahf+V058vK1ylZhxKo0IBrlz6nJ5va
UHNCb/uh28lP+eb9kKrT9c5Hlla9btyX8F67bcJ298SM+D8k3OyI/LsJoM8JynlxhkZr5h/gL8qa
pI/qaO8xorLP9HMjpMckDNUN7pq5Qv7f1uqS9MASwNsy2nkn8z2VodjwYcov4qin5kSuSTyBxjk/
g4uVdszmzyMmeE+Wv83C/xwIf29HlGHPKg8KTWvqfnJ9Am8kebaPwR89CezUsMvSy1Ho8QmCLu0m
kD1UTGz7jtN+MYYxAIzkbzg2o3h7iuuAPNVf6QgZ8t2mz6eOMm7PktRuvZuI4msiuL32Nqq8JOsJ
KvzD0H+6SbIol+Av7paJ2LaYV7s6qrxEhBvvq5KMRurVpQ+tl9cqSvAKVsHReB4Sk0pQ9Xs2U1+t
1iHQQdmA9LH7nCDxTlGe6wAJQK2ecOjTqiDWO/DUDgn6EVAG++WygXTOwLT2y8PPuSOcRsMZYang
WBA35xiODarqtNcqA95N/vuzDbZwUnC5Tebz2S2aEvJoiW/xeQ4cAUS31ISdkMQy9El4Hffwibsp
mrNL9sWk0rQQHaJD4nwjLLSVCLpQ07tlP9/QzGayq/TJZdHp4tYhp051Ak5IJPwdBRFwY3tr6xaL
ZHAjc5tKwPCusRgT2hALGXMsM333NE76f4pvMMMEfxTi07BMys3wPLHeGIyVYIOPq0PGniKK2mz4
XeyGYsFPgAwQP9dKn5a7cYJ+/3vgxlVP96AuZ9jjm7iHPTkKfoYSQqXmbhoz3W9WJoR6wToYL/ro
5fvkq+eZ4TmtpAHr3tFA6RZU5XAbziQMMK30GdIUSdz+jk6sjeGRlfrElD5lS75ps1shrveDvGjI
ssz6w4N4JxaOl7ISJoHTryUffEDehu7PHI2UXV4j52f61jJbczBFsIHG0DjEIjVAZlNFKu3J26IY
/bAqJ4Ar/LiIFrHeAx4pppPN3Q7hpF9SyGhwsM5qJ9d8Re5/v22TBMfNg0AkzyjC0K1DZAZqcrig
ugI6Jm/OlD3SRH3d18gePOoddoIjnqYuVMDozw3gsYKl8f++lR6lowY+VbiWzQZhMSiYebKqTgYc
8V3XmCcgcSPxrqtL8r0XiWsZrxDA1hY1n/50bg/Z+eRW4v4OA6QRMq0OaZFCJSILz3LcJWjU+W3C
Kifl5Z+gpSmWE5gQHxsVJuK0OzlegfopgHgU1pJaJ1UHlAQGW58DVVEeZIaFPyeTjMPAAQuqATUl
B15rhRU8Y5S1AWXZ7vTbx7d0dcjXMTKULbBkNLM7E0fLaWxphcRVFPtE9YZhdopPyhLcOhAZMLS0
3bBaSWcUAgksPYF4L0rECu0kyEG+UKamHETwbDO5MCMO+HZXcy4AeuIZ5X+mk8MYEyhsl7qIol/7
fJ7b7w5MCyNhCRSQSusaVkcRQHyBR0HyQjtK2wVnVd+DWVOf7WAaMGldglPfT/SrUcTFxRsDwQRw
J8UiqR4AwbfIHDfZUSpwCbGuSsFMgbGTiWWm7aPzNU1PBbm1ILqNB4dY4cnro5XztxrV37KW7HEu
uEMPP/9R2AGwnigclVoAvwrDbLEVNaJ/TSpZU6coOQKZMIkLtrUOr9MXNxY5vKvqKf72ZSLiS2sf
YWwq71OtxvyVUxa3CeYlDn3u8BpdhTyh561BGxaIsNkEPNLE0wUXzEYXdSOppl79Oa3i0O43WYzk
dVBhRUOqT5qJO6yWVKJvqpNtLX+75tcBf+75mq/pOmFtwGNxEF7QNpL5owDrqsKbtphP/GugO/tF
0saGvyB50916WgPyJovC6PPz6NUtQOXUJAfxlrDhFZnYnWwVRk0BQWcxHqGW3kEsk/Kzc54RhlY+
fNDSbdrgoyCjnrvYrhBtWGiRNW4PHdvdjEBrWPnZ2Iuxul3Z8NieffaNgI7FrYCv1Ub7XvjnXV8R
ok5hYwu/DcLV6lEEnmGwFqInXlYB0Vn7xpEBoRLSvVQgxcBCnnrojqkNmunwmWhawX8b84lmOGUV
kg9jjI/BC1TtwElQz8gSoSLiV7jppHpeuiBsT/JTR9nIhXelWJpz0ZbZBVJ40MnttXBfhCn9bn2E
elg4w7uVi9wE9ensmGMCL7/nSeMdfqiMHm9mTtxN/p8DukTN5PKxL0u+29GlkRI4sY4N9b1qcM8Z
5YwP+Pgy8rq/eOfjCKBFg7T2esLKuH8uN39VeRBJ0q+W10qkWpZjpE/fsnVmUuOCA6PKxqNVoM8V
Vjq9I6PoJXvpb6djR3/uNgAiTHuXsLggKfB3zCT+XAY1uTzmKtUY4pNRejHPmJ3jYgQpKnyQZ91P
xDROkzi7AiiDaTkzVc9D/Usr9peKXY5nbaal5iYCGZEJXr47S4WtOCOY+7MXFPd9WFtpHp0yRo1w
UvdaZIErCNVtSsoG0No5xpi1SMo1+VwxbWhP2ZtgYZpe0R3VbPUx7HEgMf13jEPOjxDQWywEGf7E
GKihKpPeJ9Uay3OnD+hstEPZOvUXNCKmgfc39tGc1ILiulGM7r/L3WaTFMM0yiJYeDh781dwMhEG
PfvRFw/V76+Ee2ThV/VVs7E5G+9ffzCls5Ea8CHFWm9ivegwNAtRK6h1PGj+rcoN1ZP1xZ4Q7QkJ
vtRTCL+qo2jh9JDEu/cBhmQ0Ejsxt5V2f+Gqnfl896E0h7pymdoixj0yM2Xe1fAxnNpJ/RB2S4Rq
JoNBEQ4/79PPk/v8jjHL5LUHDzvQCt5XPbApGMysPPQccb5stvkSeXEA0Dder5bCvdzmLjDqwc1u
JkIec3X/Iy8L6W9RMYucvuD6B7SxJim1XRGqG33k1wzJ3FcZpK6zOyddxbDWtSEOdyTUpAGFNEmA
mufQGHJ4s0ZOC46duWLFXiAJCowZzQHd+a9b5Yf4hfXei4SjMjYxhqVsxnxw89CCzH6Su3qvUkRz
kZ+qZngMwo6uZS6+QkZAKSvHeq5JfzlkyNChWdY3UltvuzBwIm2S+kLuzMu7LoDOfZf8J7AgVjmU
ZgHQG6xJEnql2Qx2a2UlIUF4FaC9WXrWFzL25XS4derln5acBJJEW4jtIIEe/gzpzSxaeputOIvC
xc1Pr5WO7D/uAU60feStPhjU6JLnQFXgbCMYfKXVw2yRhRXT4Kes2XHThio9t2ALCAnTJK13ZDqW
JLJm/xRe7urUdezeboBRnnNGBCOqmXwlCBklEfVtQHIkMoqCNP8s7Le/PJTFJHZkcX5JwAleBj9A
Bc8JLick0r68kRZYmVzHIR7mXUa0Mj/yqNly69/n8jUF9O9KlVUeK7llFioLpSda0fU6rJStjvqF
cVDEbnQ0pnhzFvC4S6R9JgR6CqAF/aJhTTKFtpzKlrERENhr9H6HswEujLasM9dcX0TGxcGWwnh9
PYN//Awh5LnkR6zqiVo+h0+rXrq3vIzd41AS5vEubz80MET8Yec2wZ294z0wlkzObuiC094XpeRD
nMWra7sjpsZCJHwLjPmeV7XUfNxdmfSRW+QLUHUkcTXEowHsDHsLLQHYJE3V8is84qcScE00H+SS
uVAg7dESOyuhfeWj3KR+j6H4Ngd/QpTTf0QykKqGUafs5U6yExn0zVq3DC+DlcwAVdrsLlcCdnnq
E+l4FifJwRQcu0YMOdU1IA24omyUOIkWus2+o6IdAJBL+7QMz7mu3JZqTjzAhSiy7HHH/3ut3q8F
4rVX8PorQXfy6tZgrbKivT7W8FcgNTWCEOMa5hDlu6Sv7PwwMEDOKmnrCMFVBNKRVuzRMkh1SQRi
mse4PtCOhwWXqLY/DxB18du8iOlfBVFRyZ1Rxio3pLcYdbUELr6hWKcgGU65k906Kbq0b+91QLrp
K9UO19O1buuutzaEgQ1hEIFz0+eN3ldpdiYKkcxOKNFWz6zh3ccYOW9iBjaPWj/F/3p96fZ47/25
BPw7VyOw+clskxT+zs+iSGC2r7iCIIfVOrTKPm21x3kdBIltrMaJ7C6iNQhcPiKadf1o6FO9dqWQ
O0Q38S8cgajKUDH411KKmdl31n6mF1Vo1ubKZwSwSKUgO0K/72Xz7Ln1LQ7Vvz6pM8pvNgMXK2Dz
JdtfgSoPz5GBuzWdSYYj5DATQWgI8K87efdMxiBlED4pkz+YMzHIwdZRudZO3V36Cr90LdZnkPNm
Gtafi4AS8Ur30rMjJg3L83Ni8oyDpHM6x02mBdaxjZdVLAV3L3plrvTOGyI38mJ7gWZSI0fFthNb
DuAX94M3KcnXQaFab+z/3oyEfe3/cLxbygnvEsLDUBubBADEiO1VsDrdgaT0t6+btJCOBaz0aG4/
BBFXZ6qLngefiNFmqX76hcvmBlXEtEXbK5gus3rNS4PYtqcw4bJmvj12iPX8Ah/JqIZnclSiFQmF
vAZF3idFHtqNHhESdYv5iZHRa5QJFWMQOMK1kFweXlbZMLLKbkrTAPm/aHnEMtdd3ZVgNWUrdEOL
yliwoekyzKK1aJaDATgwe55c2v5FG9ITDtbemSAHW68yWAvYh06RyZu/+hgBNBVzqXxYmF6b2fn1
foxx0Abnj3HnhWr2jUHXYMYQFChw5RRaOneMQbpP3F1TLUbbcUhC6vVRzj8vC9FkW4mu32WrQ57Y
qAIjiIBoOR6XhzR8WQ/jj3xl5BrppQ9nl93JAV0rK64pVjuRnTSsnFb2t2vdIQKaGKZ+iVb3id/b
9UE+MRWxWMOeDHhwr+o4v+f6z3r/i+hM+G7snmWMZXHFBRS5GN2oMFeKnc1Zb0jizaYI3MTclENT
uq2Zjq1Lsx0UgWiqX/ieITF014+7ZPet3HSvqqDjqIt4z+cNAlMGs2bFZ6vAwFAOik/ICmYErNnE
FXIITwsq2OagxGK3BYo8nNwkjFJjiXIEoji4Fa59uJsO0By9wdH5Tj+w+K0cJqEt+Lu6makVVTUr
1SmNThe0ZIs58rTAiS8SodKaYNJ/uC+v4YF0de3wKIHDDGjXIifWgI7aKrmEsFaqEcFeAlk17HHO
sPn3Gx5ytJ3X/NMILSP1ne0nqBO2miiCaliuHqjdTyzn8glYJ7T1jVFLKtuz9w7DYZwH4BYP+vl6
Fsz8/Uv/HKB1t2j7lDAD6zHHm+MlAxNkygaXqXqkhZEbA7TniseFs8AVVwWWVuZSX1PoueAnn+Bu
09fszzEzSjbBdwr8NJKxUVMG69sTqpHol2LOfz+Awz5XPkWAgIffoMfENxQl0ci58YOwMk0XxCvP
Pum7WBY8AGiljUO1V6WEZ21mM88LBL4wmzAYDmxyZUi9e3+VdG5DmsQFc6jFGhc1WXrSEtut4bTZ
B1xVtn6fe11GFI1Qj69F9SQAviVHRzzLoHI6+o0XQbSIm+M/a72V+1oQETWm0TJZBMUUYW9SdzRs
X6DL+HH7d6L75huM0FIwTOoDWKhSvU3n0mLaXbbUgwzV4vTjy2e9AWEAxle0QQic4mCd5CN8iz/X
EXFh0bW31Ebqs2W+B9WFKex3FmhjS3sB9J4fqEle6CoZ/OwOFvv2xiAkkawm3ZK+8nJnkW95smNE
fEyokUFbt9pMZCcvb2wmTl6OghaAwopSAsh3v6Zu0MegSf9NCu9jUPg+KpqOFKFOpB7aGHGIA4cy
84UM/DaBsNzUCgVkMxy7M/Y4OQslvY2JlwaGT7Af/OWToQ53TIz/IZbr8rYZGlW7ZdDBNGjWtY9J
tEgRp+zP0Jftp1ByxfTXRpqKeOF1t+wPceM60yMjOoYIY5tLrbjUbLlnp1QKuC0rCZhXISBT94zN
GY1n5oCJQ0P2g+kzv+924ochr5X+5mz6VqkgVWx03YJlJhXN9gaimSZYDDA6Gv5ql9SSQde+3vUC
HmiqLNman8r+FNRrXumM8vh/LbelGXm4kYx2DKUF4wU148YHpox7b3dqdEiOtOLWdHALTGYeUp9i
LaVuG+ZXSDrQw4BDA+gWq7uJhee9S3cTIMqFoFaPObmwvu5tdM97tFKZZqw+yvOtxrnrZEyf01tc
AaRiUDAZX6IGJMFEAgAkIpK9KmN1HVNfV0ciOMVQ8Fu8tqsoc82R77GlL4OxO/LnvEd4gjxOLGYD
LtYJVZXKYXYeuKwbfA2TTex7K+iVoha644M4nRcSO1uFSKSBZTMsQ/BsrmAYhs8FH+2+lESpj8ag
koOzDju/JC8+g3Wo6wcCbSZlwnVM6axXCeqkMqcc5xKLgoQiwZTK4THXLNomrvtvXPAV1GalIchb
Gid/9YyMFTZXC2nZj8D3C45oioU/o2sfreW9VmH2hW0ym8Ba/jUB/sXMHpdbAP9PJ1BdtBveM5rb
7pz57k1cr02NWN7nO+p0dZszS9ORowTnlI+JiNhss8YSBfFggyJsmZ8MRcK2yVytcl7FQ5pYyYbZ
EKK2pDPK+6z3Qat14a51V7Rrcm5PRDOZreZ02ZdsldHu7Z4BeXpM1xSoUR/RY+HfXe6dj+ZQNial
H5hJB+jPdD6OPjZxL5x73Wh6kCd6eeOXPOMzW7b3+YP80E8ZNmHNQaXW4fHvn4WNsaZ6yBPQ8uEZ
VhcAfFJBwO5udbp0x8dTYQbavtrkj8/aYnumw7AF/vCdkKND15sdeJF5vw7cnQolaFZ0YSOocm4y
Qcpdu3QWNl0NvJWUpkwTHuHJuNFMLAjmEUaPNH9OzLnXsNOw0kYCfkCviEhk+z94u/QXwsdj2ZUF
NyvKs6GSNIiyUNS5ko+Ut1au1Kk8BUGZehuM8M/dmwsSYrHF3myjTfgI0ck6WnqQP14H/tyjhByK
XilCu9jg+mPLfeXKz2Rsh2MPjmOvzQofGZDogfkzNMTufVmumLSPQmzTbWdhvexJY3RRE9xKf4TN
TYX1Ny3Uuiu5bdeu+Q4H9sHiGBEnMhKFy58lpA/GdnVtkiTuz1xvzmULAkIxuviJu4h5rUlMPn5D
PsnP5XSXqW1gBPwIGc3VsFYg5Ge58yI6S71Xc58Ibp6uu7toO1gYe8r5IKSEsaacBMJ/w8xo0CKZ
LFjzaSh9ZnkW7Ed0LbAfJVUyuif75l1SVSnhJqJDe7RlS/QVn6lsPvYrjwZZQFP53BYikNUh2tql
lOZqm5k4Hid2DJDsGSWc07IUt7A7cO3PUTZdB2b98yxDKX59U6AT5uVrIB0RkBSVxBYhc6dOgw7g
B3TEbpudUcF2FFhfL5NFva082DiwqOgjaKgH92kN3A7eeTzsiQ3y5vqFr9Z8Hq6nU5ab0GbaY2n5
8ld/NsQNx8+NDnsa49yBIJWN/ldNAp6kZv5fE1UefVg2cWi062mgA6pVJEtEldEKe0IRBWNEVZ7u
P4fABFOWlyuztIwnOYPf8Lbg9euQ9duxBFnHosU4oZalg305e0acdRlhsM5df/m+EoPCB95KMcIh
t/qDTMVTHsJAJKuyEpUTLS4Qdlj8PuBCRoJExIxa/35pcbRV/P53s180iyBo9aDrVsUYcITDbKpi
X0ABvCflKxb3OWolGAlIVOCWh6J2oUbtN2l5cXv0Bng3k9kJvljul5lYl6UQHMW4hO1tyW3y8jKA
FOndesUjA3R6eYUIqvaoR+pKhT8tQEuz1Cvctsi7a8FRUMDPceg225ybk2wpqiTcCwNLM2rR0FIN
sbIC2ImxufC6G3cTy0QHC7pmKrQkXALBGjkx54llIlCQMaT0VwzybsCr1Uhe+LxmVM+0SbEY70wA
p7f9PGAZ2awVQaQp0SV0CWOoyH272xRYJBTSxkERp435QbbVcjYWz8u1wUQHnKEja+zY/z4HFbXy
Y/AMn+FP9wCuSkDZDKtbkvHIJ0wJUWcIsCgV2tHPzm1NFAzrrMDauO7XZmx9Ss8qekzwTrg6JdGP
pQ3ZQNc90K1wfRHNoLDhU8O7fQuQF3Bpm82PtNGmkozfGv9lUgTud6UtKthHgjHHSofmbnSkhw0r
f6R+ccBxaD3rhwJ3st+T1vne94au+sl7iWWMFE9I3IqcgqFy8lZq9Fm1ETFxg6VZDjEwZPJWl+i3
EUmbnpdndvdW8pxX3EHslxjQN7mhlqmY20QRshzmlF8ylR3ytiOd2HafQDynyAgxe8Niqg80WwFe
Fh7lCAOeDybU98ghW8fmTpKQ5brs7MnFgGFxnPj/xGyrQUDpeeL5oxOZeb290UDMBIwoiq26Jk3K
5FK0CpAo+zKeidbXqQ6+ju2TpjdvdYUHjH2Zr0RVttRzdYRqAzqF1z3Yq9VH4SASvIa43867vOUX
UpOoun2CuZZH8o/Z4ZJaXrhH8cDMGjr1eyRPAlDS+tncAEqNrpefru3CGs5/2pmNqIuf7Dwff9dB
7/o0/Sd0DIPNwVc48kdeuZ00sphAKReQa2IOV6DbP6De/doV+NXXsMmFClcavT9exjCRu7DjEmTA
v+hE+YdAWvv+i6EAJ7+N9spL44sM5Lv9x8uI87BRO1BWVDG4diIJUH+0VUUFggVsZdDdiui16Zg5
+qT28iAtpkoCvI1Cp7HFKt/BT0MSHsiIMF+aiO7hnSrE4fRkbGCDZLMp5P+mhT57ScBtFR7o041I
b9jWfNN7Aj+Vq/RAurZd6FPEFDICO9R4VBYzm+TACCdRPKh5bWpbaTtwt0/Rn/ssK1ZF6liYMHr/
7OiSHpx+hma1VLmdZWsvDyCc0pzSBubfmqY+0YPwHx+y9HoQUDZH9n45sThLGufM57Sm6+Dnqf5Q
+RKPorcO/555kKjsRHIiALIt7Ba7B4gIbfmVFCcueLHn9B/WSgWLoUkkfivnExn8BQIbdEKEJV4Q
V+TCsUrpAHXddCUQCfyZ8ULmpS6rtaLMMuucS58psmJfNLdGC77562Si1YJ3B2088zx/cQ0Dgm7Z
pkuz/Aa3oXoph84jdCtvL9pSuQu0eiU9vvr3pS/l7oC+OZO2ohZ2yjBJn+6xnJkI89Z65r8YUTJO
xlP7CeOrzy4+2jS9TU9ic8dknpCHY1COapxjiYDKL0br44VBJwDE9PfIR71m79HICaoeKDdCAvXd
5ywADw+9iEOb5I+J9x+/AuCbVwWFjWv4hBg+4IuRQ4joW9D4CT0jkAipNw85euhbhlBAvR5ikag7
2AlWSkmO46opGhsqdfp7yJ1LU7Oe2mIAO3B+NC1QgG1evsf5UNOK4bpRWRS27TKCgV4rjiyYuqYr
5yS7Jz5fdsQUHj3+Gbt8+zaYNWKOK5bHSyPHF37HD+cLeen/kT1aQihkGH1Wk9Nf6+OEFvBpy3IK
iJFs6wjxTdGab1K1nSQTrvmoVNfhV79iR8DfS3QC2kWrJT5YFpIAQ9cYgAyascohOg0gkK/ahktQ
L8REPb6xjg0FO2coXURtp/yvMUzQwibDXVEy0gaHcReq2z4FJPoKYFsj0qC8lX6sgCTsezbApwBY
EK8rBXxDE0CaSkvr7vjkoZZaR8gSdcaC/frlL7rDVBhYgnMSySJD8h7enI0hDWj85eFWNlIEraiA
I/c7ZaU3G1xvVjX8MUoqL4vAggVEI0g0CWrlmPR9o+ibFFmAzeq+OiPUkEtaI7TsfaGfbXmvP7ip
1yLZf5DQWp3Urn578D89kgfNqS4i8/mkwY/Iq7UxwPBFBhz9JI4Uabvaqryx/SGucooJ4bqBqtqD
CZYgGM4R6u+K96Th1JVaP3JaomNxlRdLE1DHxgRnBabR3+/U8nPFJbUIm6TkmyniSlWNbyqg7bx3
P7CiZXXumMPdhJvbesEKze+Jl9Um2B4haV/sI9wgkGb9wEevW45HiUncVlUZ9CWmWUc5q7cYLCgC
IeBpk/jH2r6NRO3e2cY639F/Fm8XtJd8P3lpqvo/+jsoUbUlDAbD2oCBF9LDDQvaaqQkpoFVlO0H
HtYYI0SxA5zEI1B/wHjG6bBa3gHKPArYfOzOqNbMa3N02dihMASgBvuyvDZfbn1Uw2v19HXwtkZ/
DTicdkg1oY2ZNsqLsBy1NlBiB1hHfPqUUrYEbpW6rOHzDqZaI+kTWENY4uzijFWQmXOsbZIGg+E+
AJB0TRRbU4Tl+HMYXvyzxkPV3GRD+v445CHUaHdhWXpT/o5DszHDlWvGjRi865CQVWKZDkunjOM5
qSBi03EXY+exb+en1ztJ2gX5UWEShQDijfjbRddXHEMX2HAUUxnoncwIo5rKruxS2gnjkEr1J5AK
ysQB9nSLZ+UVRrQdJ9uBPdSAoOywMjNfrYQHkeCjMzT8XjlSBtqI67mCrFZdqM8HG8mn0n2cKl9i
OvY90CEEKSuWpRkB3eqjmpmlr/SUlaCA8EcdQdtjYkSuKZZ7nrEPR6FyRFB6MB3N8VFoaAZSpx8u
nbnKOPKzn+YhJ+9w6OzPGTYBlvPQQsas9GC9QAYbLLE74vOZlCNO1fckx8deF5t5YWKOsE+skTg5
mSfq/W99pFOMU+7xfg65X8XuAt7sKmRCnpNP2lMKfDH7+RLX4jNqX+jSwCQjFqUehWmR56C6Xyak
vPeMn+hXklg2KC6J5nlEI9vOmbeCU6buEjdw8LT1J9hfDwYA2beH8iJe+wThuNxUz+jCPZULYnYK
NUSCEUmfe7OZVJyEVWSAI/jRgzcKhFBx3tV9IGFV7c5liPKkSBdRPMDg3Wn7OXAZ70tzAp5bYa1f
3Dvm7X+pUABGxJmO4srLexVXi2LkLNb7hxEqItcJtSPgnbC/x8qUY83yohVjmFRNzyZvuvW55Gns
ITjbNOJMcbF62kl/dhADY2n/4GHuxDwNu6AS8AAZASpFlLF4lbgoqOL7N9w/8u5qpFWbGt6drYTG
TfkenBMthWAw6r8ynfFcqCuCd37HrUvEyo5W6JZ2Ke282KesOlHydawJD7SB4NLElY0orMVWSkiu
wqolXz749KfjQb6QdlKtFZFpmuEv75sap61NGgk9w961AzojcSxXrw7hN17jn8+xgLTR5qW/5+nM
4uMjVDBu+BJAK7TqjONAYQYeql87ThP7ak1Ty8z1mz6gThZnNYluDDdmhYyjQEv+mCctHdG2Wey2
VV3v1RiIuf9XleIie3xUfvhuPogYtd2eeqLWMUzDHMIMYEvFCF4hG+30dS7z2tu/YUKbAZG6UKAb
dWWuSLotJSChJtS4TQiTlehYRM4izN1bu5Ka+AGEGvrU+WtLmbSy2HiSQYdCW4Wn1m3gVnFE3V2Q
mGwhb3NIFIfIkFGCSbaUEyV5k8gLF2qzoGwZVVfYMG8f2qCk4QtUzNyh0OQrHoE+bShFcIEKrYHf
7V1qxoJVYaVyLXRCIooiV5e6Coglg665zUbTSv5Vvnd9oAi/8IhLcHjf9Dq6WB37T0YgQnnj8zlj
Vol7Eja7aaARTb6uzGQf9wVyKj+AoxfUvshEfTE4wh4STe1l6wy8clpzQMeqPADQldh3aiThvF0/
i1/x22eI+D6STCiRRQFLVZGIly0ItaPzTIMiOaXjn72AGOXB/KUF6YyAMBbn+6DEo4fvLtG0HLoE
F22uHllB5zZavv+dacSU9ZUfgK242bGbExKbjUOtYB0HCAsLfmoIlQ8fNBdS2hQsk8S0eM11hYxS
G8qIR9ueJFoL/GjYPFuH5y0nShW0QCD0dXlNctyeM0nK1SeFpvCG1DbZ5+tMzkf6ghlPcOmwuJE6
RGwIhEhWl0G3uNrXSZPOek+XGsR50LLqaQQd+arV6bAvIyCHqUYRLWmOHZeVQyf0I2ihvknH3n2E
dxT6ZZ7cwVGBs9Ewik640lthGzCOSo54kKnu+0Ri3BzKXoQ31gm+/wwwxoPK1jMmuRNvyhWmvaQ9
VmfGHXv7rjjCafiGotPStly8SXVISSuYVQW4ZCLg3N/uWLdzeyHSMxyckEe1KMzl0kAcijmhfS8f
Xd6Esss5SV+pyNTYLSuZruVkyMgyuW9pN9j4Y4emUBqi2nOW+btJhUhh+qCebQvLbM8DRCKWxg8Q
DkzAst/KhAQsRQkf0cjdeQNH8qmEKi6I/S4pB/xCnjYNpde2igBbtfCZcgdYL/8ZfDWEqLA1uUpf
gY/7SXt5un2AYq0D0jXyCVjVzJDOVKwDLZtPVJY9lKrmWCrX3wHRIGwB5QYBqLaRZWIpRmLPgcT+
fXsZ6mBIrrA7X3blAxKu/jQkAvelQj4X2X3K8yjP5dq9j1DzRszN6ytVUG9u8ZO6pHTyAGHANb/O
tVAtHUcR31RviFGv7Z3MCGt1YSXbY46dDxP3nJPyeM+/4nt6nXySgm4gBHGlDHSBWlmRjxR3L0yI
bGm9hnxUYappvF2WYWCpcvwvYrY/mLnCPQ3E9GaCsOK7p/54FHXnlg5U0tMgIWvMpq5gGWpAhjWQ
fseYRaFfZmtZt/3npA98wVkx+cr7XIeDFDorNNmxsK/Eg5LChfnKmFH40vpr5+wggQouxvVYzSN8
kWNnvWWkBBNt35InihAfWGvM2zX/XfT7neK0M1BmjxjCed99oohzz923upScVVniXjMcRGL5/+Gl
n2HAnKJB7f2KKZaDlBQLFtprCai8s73qm9yA8oVqvgXodJ80ykN3Qkzz4f0XBF3FBnTwVHCJedpv
VMwvxUNmoGfxqjDpExKv9uT94pWYN1C8wxh/RhWoa38YJSn3Su2OtkhMplIGiOTbX9Da4evx4s/X
o0R4XvigEYz28adQil1n3KiYKTD9mzOlZzRmRTJFUOO5vfDqJ9C7gilDxxH3lO85Fu09lx1KrmTO
LrKXdcYJCo9zlJVod5bbKCP/6d+5aGnr3olvqAldr+ywCehlxEbyHUTFLwf4sHAfIrB5xpHNCgRa
RWd5B7/ta53CWONriWtv5AXlPKWn2EdgSPutYycwVachJqNLuIigUy8acA/+2jVxnr35XZlzAuuP
Jac+IYhN66U9Wi+hV3h0xos34WwawG3Ni6etgFK+w9oaFB1HA9xI1iySydCGOHUgFfQq1l9lYjca
v45wg1b5CoqZ8eJ5muLGH+pMKQwa4zXq46bJj1OZ22Y/ryxStRbvo4shyR1FReOAyhGb//F60jCa
i3M33pfOLVq54t1w171qN+2wOgYKdbBhzUGWSP7bq8VxhYQkAXJsi/su3WbN3t1y/mqpzbS00ndY
cWNDaXmT8xw6eHkR/IvQeiE1N6eN2NNB30Cyo+0/5he4c2JEHc1IivpKMfQEapzje6eAkx6ymQ/4
clVjJ7hdAhgRG/R4FSMZPIUHoZluUCE+AOQPxCVLwyVzRqI75uiJrpc2QwVEFRqOjNwqUVyCnqLH
4updmea+ONAnOGpln9v844ADVgUN/CnLnhnXxvJkE1+zq1hP7ALPhf7lcDd0nxoabGEzu/k+1PrG
6gfouozxjqQmOryEAEpfkD+Ndes9tzrAq/zuKHqQSPPAGgQKRz5ddMBaTXQdLx2qhmdNTNw6hQfu
Jk+otApSnjOtVS6am5xDgLJE5Q4JmKVBrKSyDpCKlfaSHNcsyLzXp3QXu42+KV4IHWffey6lmlsh
8SjOFDXU1zmmRiP3FnK1vVIJ4ngytZ90EU3p+HI+7gbAban+pv4ES40FVGXuWAyN8G5akchHrk5A
KXAdvN0W+2epWfNSyI+ZRCcUI/HNBLcLfroOQFtpK6S/rmpLFFoS55fiL389NK63sCv0nQFhs7zX
ck5waXyUMCY9EW7yzOuzeE/SQpDtlb+OoltbOBzmTZEW6wdtDMp+OZfoSXm+BTwVPtrYTha4bOw4
kUif6tfTdDmdKPca8gm7OF4myCX7slPTbmRkgce44Daaphxg8g+CUyUKU5hFP1bzI2UpwWLBEAbn
oLR4BReIO4IzKYf9xTixh023N3kWL/pFI7ZLs1cgg9HCuTWLadfAU8UFW+Tj3MWlbyEy97BMttXW
Y/eBgbhKiVOMhkRkc6XgN670kshgqWVGumvUDqDkKaTDUOukIUvVk3PdFEAc9aGUfYpTEJ8WsGJi
aH62sQSEQkLKEXNeCoh/NIu5wZ0nKf1pwesSQjtsrmXWjOFh8uLYVGfs+MWza9sERzCV4pXbkSpi
iw2sgZJvgd10aJWxdP8vGFKaRtAfracFh0M/FiQvzfj5PUAK3hfTv43aVzpU0rpqKktyyQmvJLwQ
nmVT4d+cPrPLG6rB85tJGoAIiqe3uYSgiGfJFO5s9ua14HxYICDNDX2mvtGWr6KI0mnv4YDSdW2W
/Tt9howEwIkgW2C7RO9UAUhonbTcgDswgR8R3kM4UtwhiVO+tSZHKO/0F9t7VCS7JqZCY4N9UIxJ
kGETL0wcy8IJSOn3+Ktfm0uodF96tMVo/POM83BTVI3QbqEHgFFwKYJaNJibDWyAYKLl0LQL4gpS
I7uOG6eZDGiO6jjeHEMgTm82I4kqTkrF25GkbTIupdBWJt7e6Bu/QcgK4F7z5OGVqtaHSuS1qSf1
30mCyNNB49nqjsBV0Rkry/bR7HnpVD7TSZkjVow4mZpCoTQl9nhOUZ0Lmdzu78pNo5Al9ZX/llh6
iBMQsJ9+8fqTrr/JWVHvhdcsKNrx6P2X4gPOihKG7RAiyojLNPA5U6qFwfZorbYCb0S+6EyMFd+l
i0lsJ5Yr1YNTcsRpItGnsYMdXBB4qqHmkYrPVTX/UDwrepiwVZz8LNufarN2BSZ2IZxDQpNZcSKZ
hyspFEqAUzKBx1I0d2EA4Ebq17Rw32UuyYL510NAjMfhdrDnrkxXae2HGzCmQiBRcKpBn2ooQKeG
S5lq6xoZZjedyX/XMf1RvEQwarwz6lEpjcMHORlniWbF/gIgYbRfGRSnjZv7ULIUowLWhACayoEL
/lzxHxU5dGSb0agssT12RcaDO3ljvZFMT64mglhs/ZHy2q0P87Jv8u53rgBB3Ihr3Em6SJOAQTU4
6KP4yA8zgQGb/wBzIfVw203BTClap58ueadNFHKVH1O5L0nSUWkJJx0Im7e47Xo1OkkPeNGfHr0N
/7Lru9YrS/IFw0RDTZa0cNVzosO8K71gwFiBOQqBnMv7NX2eNSMWABrtqzIf0oM5QGV2OaPxnbt8
+/yZ/osPFSHnQKWry64TkdBvN5cn4eREISCO1yTwdN2P7SaZBA4MoCcf7DYHe1blgZzcSQYQuLc4
Pv3czpInSC3KUhNg5p54bHWAX5P8fX1Od4sRsdNtpxowE/Ed7GwAaNdDbSaD4ZgYkcKoQxHAHfFP
czLdcv6S0ffEmhS8V0eiOsBDk7Ho54HGVokCjDhFtBEVifMGTnwl9vfqXUaXeFx+Hp2XS5yBNMTp
EgFoqQFitqLMDAliJT6WiwkrRgwLEeJ3zSTiG7/qmvf3EgmphGtdnZee4M0R7bkg5EtGLKcUV/8k
mmz8I5fkwAtuChthbngeuZdQRA3HYAOkKr7zTGMsb65i+X3yEV/AaAEzqy9gFw/A5/CM97TZ6T2/
mKocHHiZkQTI3WSIje/9lBBTV+jl7mEawYWOETOKbPVLsaRP/E4gPcp8lmJuFtA6Urnkgscj40KK
YASscMmBy6fqvnnqTWeEOwunfegK8FqjNmWCP9yvV0zT+a+4sQeNZ0QGwqRwqK0YbK2VUktxg1tS
VUff1W1OIrHxH6IxrbpgjpZcInjwxLXmZujPhJ27xNCQvjjcRDzuogC6FBrY3bFELqVygzYg/yB4
aJI1SXHELuD/nX7qle6kYpwD5voqNwmeXX79Yr1Bv8Kfm3JQ5hPmUXMU5gQXgEswBI7TPzM51Ac3
SdPFEnxgAVBOsIHXhfrqxRSWtfxQvbF9XpX/+YzCDEHDgBaRddR8T7+2hhywhR8aeq+xSpZBCPqg
4xpKtBA4Ldc0TzJWzavLbKy9SPrIu6H2S8faPYpdm4+V1KpgjcaHS6YLIRqIbShpeRElZQNL5I5K
6/Ngk0p+EkW3Z6iikzsaxhfEwZ0G7J5JsaWaKYQszaXx8wUjnCimHMTQFUCWjv+z/BosEIMPT6Wg
z19ZMrxhSFInX/VjgnNIr9xRJ80NDeXQS6oGyukb5N0DhdL17eomEr3Wkmf0vsZKieN39yl37qKa
rmYLLdk0u7H6yaFGTnv94bZW/sUZ+o7xfKYpYhhaxRJFKN9qNL1KZVe46VFvRca07mhh1onEE8VG
E1xz9Jh5IyzuEB6B1hQdmGx78wyzTpurTyO5OY7OBSSVquiWBfjKWqqZnikFVF/kJh76T45c+Lwr
lY3hqSdeW42duKucLONnYX8KGFWpbgaK2icEk6PV4C3JOZBXjN++ZNw7P9ny67GpEhrRlyPa3oX0
4rL5kmC4o9b0FVKx7Rmpeq6vklIX0VwvqpRDnufVo6DiuT3R2K2/4Cdr35ljBnOLeiP7OBTDtZxT
k3j0/p3h42bBrdUgiEQj6jHAFY8CZ+XZ9Mn57B6+Qwo09/QSXYnF7FDsTKTYlO00LuWyFHxAb+vA
efx95l26DizlmPspJxTuIZsCnikt5N/hGQqfGAC6c3Z6WRNnTUsBqXEsz2IT0ZJEwKTIHJ2ZZQh6
uhuzgekiYIvS6GslYvBeajY5HWfinpmmsIYi9hh4dZw/U2aXXvFrcqb7tPGasgcBBhULzv/EefoS
yGosoEEsnGdfbStBiyOvi6EUuhhfRDvnlJUtdsO4XEaKZqLfARmWAG0jF67xp6raMYnE/A1XSMfD
WrSz6Orhi+q9MdRDByrH5tjl8EqE9HhkYDkgekGiKTj1vSOGivzMgBH2HSs0lnSQ9zhlCvPeJKPE
YI+ZzvFTjikP4PlKZhfxupBCqi/yug5MErK3wNL4Gklq+ZZYON3hDl20cbZ0i0G6qy6nQXwCG3Vy
SDlv/EmsteGwr5+teZAx3VjWFhIF+UXJnvD5XM+qNCQhVbp1StYadXcQJoMSV8vN+ftN+VBpJicI
unDbEt7VJlRps7ojw+a4EzUy6hkOPA8KWq61VvVMe81du3496mxLJPPH85INmD+qSX1JuQIS5t4y
D80Qy+IEDd4wurXT4CzFzsVOhH68PbxRmp6qA789H2eIg4fGOgHvm9shkRMNb1K06CS4SQbsBdI4
8kdytj3F3on6kBDJGQ16toBL2ZrsLmNqGYOCW/M83xZRbU7coO9ei4do7+s+AQJpVN6uL6RKv459
eJEWalwX9/6jxKq5O/jtk+t3NTptmbB4I+3BgqT4wVEp2nw74ICAfShr0KKuJgHSqyOvBxHnkGm5
oMOj+bbb1AcywHdn/xYI+w/LkGg7tAsV6saulN2jGGOc9JS1zxX699+atUjSMrSbEsSiIgXhC6Ub
MyaPorQ1RHxzbCjQl0TGE9I2g/j6HKO+Ymt2qGqxGtz1rxFlqO+ZStjSTDHRsLz0MU+JjWcHJ6sL
MsIUOt4yZGMg73RmqpV9p7frXLKlsMvzASGKOmSbObQ6mS8j3DxICpQ7CFP2bWNN+ozQ4pN467fA
13JDoJuENDvk2tBJ3T9G5M7TYoqp6eI9wzQVf5Zx9YxoVKRTuyZWvFsQIdmx/Io6xA0gSIcDf85h
2O99ZEqC2NZfxLJsltviJIGqExvkvIUrB07i/do1oi/XD7njiF15GjrA/NO6o5OWjX6LmSBF5oaA
E9ql+WRkNuK8TPW2DA59SlFNB4Qxj+7yZqo8yrErdrikX27QEavmBvMHXG/75WasufeMVBpEM5ZS
gr4qapXv3Ckcw7FXSZLJtbxvzR3rX3fn1tiRgJFOHz453aE5RZ0niLTbX0tWM7e0jp3G2w5dwlx4
3+ByusFJ/1wwLGEG83U1yRPaxn650grA2B3cGDV7c7Pw/Mn1VL8Bqju61en97bRb/Wi75Ugn68Xs
v0r34gxO/UpRCBLF6XyNZH3hZmv82B/JdXi+jSNQpApjeAsoIuMoA6KDpXdKtoRgftTkIdV5Ljcz
st8m6s0VCdrKUAg6RX9LkBAWFeizvAIpMz+1SC5bHxfYR2itUchB9ztZ9+zG9CX3Mh8vT2qgpOLP
+c5pxFbtMaNSmJoO5tFSVnKGG0FaF2rX5gBy65wmoNyhPxMqeRQ2w4dhLdErXhuld/rqshDxzVb4
waLmVf0JSN2FiSWLgh02bnpyrKFt55CTw9CifqtH7FjYOFFVb7BSfi7iN6TlitohJkzQMmItL1bj
8xAAFMaucBV5V0ZWTifpXDHDmWKfAOJIN2hj+f4o89Dxj4hSsr3Gj9gR2w6eyr/R28gOPzxi3wbh
fD/uRxJfbpNnBJyQqbOPlDS2teb2PSAGe3bFcq/o7mCoRT/mpGap1P9QZW5/pOR/kdDTeQtdGf+4
Tr8DqXIAhIvlfOMEvedu43K/g51wIi6KmCbiU5Q8spTARDwYdg8+hsUs8um7UaYhJFk211IXeJN1
touUvHCR2S3UTcfq5poWnAcFXrqVqPd4LYPtQC5TV48wKQS1M34a65PeWnXCN8wx+afU64B++Org
XYA2IR89NRgRYOO8clkzouPL72pjdSyKpZcJYd/MafvBhwY3CwLHeK4C2tHcFI+21tsr3AM0bxmQ
QtVH0oxFsL9xfwxZjl6ei74X/cpicGieRpQFx7qzG+cqdK59FNIbBIVlcTbgzjKRK7Vo3rlUxrLu
97CW7ZMX1KtM3vZNWT6CR7SatIioO2sCouoBnKoV42yhk5wt0oTNzHZm891SammhGq6qCZ5PKfS/
thdh1X6Z67fddQUH7kIKk5xCD7gpe/RzFdXieIfG19n7hw5FiV9DoTOX8Lv5/MsVHvfhMYDFK/sI
bw/lZ4bO0tgThmEmcd9/+dYU+oGoQp4xc81/BUZqsVORucw1SL3CteoUwyE5n9utQvDU5crqrYYu
TDrf9hgZ6rJUwPkteFTSlg3a5Kbf6Nc8Ok3JhyqIzZcXInQKYrHhoP/OKhc374MjyF/ajdCi+iNG
Rpr84o2E4OyVF71eQxL98EEFC4LJ1mir2HPjOWqASMyATRejPwaFwms9ZO4n2PMuyPYdbblAjcQt
29QE2VRw6H7pUQEh5oTNlrymFY5OVGArl8xY0SFKque6b6+cKsGVOdoPV6hwG2YEbYSqxUSoTx9T
WftBiKVvRVsYtDkpDUq20eEyduItWSt1FFgrTIYg8/6+cv0LEvnqGNpbeFdoMWxIuIVIxeckZYRw
Aj00eJvE5m2nEsikbIST0FeAkwTqV9b5wWJvZ7FJDRonOTDWXRREhr98SMTJFAoGm+avAQvtpxyp
3V3Xlc2loKIrb72bWB1/GjgaJEp4vYjPnypNo0bzYTMkEdgGher/w1+X5HPklpmJl/DJIgHLx+jD
MPS9nyd40Y2RUsXnnhVO5+ZtQmZlSpbGd7vcvq0MZGb0hLcZSZjfywcUp8tp0sCdSwO/j3wYF7w3
xYd7X6U85rVcPW3OzTM+dDM5MjF5kXU/KrNr8g/q0twLMWgvc1TMFBQCZSL7AvsP54zJpfuHIZ3N
//hnGYJWbqze3meHFIrdd3mwCUOMUIOKG1na7b5FYmlXwB8H/hm3L42/PJMZoKuSVKxaEDF8ocXI
JOJviT46TmjFReO9OkGpnmMzwjT5krKcDjm33z/trCjauX986sKZx3eu0fU0SrbqCNo6C7dKSyi2
rqYMU/55kvoe0+Qd23ezNoG43UOvoTEoBNWa/81BgaR0H6v4xS2RHy2g//U9YGIfADP8bblfKQO9
qglARnLF3h0luLTPUyx7BQWIUJIU/rUXAmMzR71JTz4KTYNK9+S8Upplse1jhXjzT7FDueqVSb2l
AzQtHxUCeDMW4QSvNtJXysJzyBMuEUuFXdzX4jmWBbjeXMyIvX4xC+3OdsglEs3ESRypYjEY2y+v
a5PwEEbUlI3cNIDMfpsfvVAMrjihrmORsGwAp4/J4aTido1IvLeQtzqTHHUbBiw3Ad3Bq/STaVm2
oENm5wAGqqEvucJHH6wt5M3ryS74zltx9z2smIUo7RwOo+zbnmcZE80blRguH8EQKFGIMLFO8usW
CmSrsPrvp+2hT1GNtpPN8ixfVgsEa4ZRbxv11RdBALcdf+VLQV6sRXfaXXlF9n5mRz6bKtBGDNx3
A2NeOZeH7hxscBgxgVCaqxq4YUuFB1HOT/3Td0c96san/tIYAJGBpcFNHJArnUUaJUbMMI3/10kr
2M8szM4R4lcV675BDq6qIpxYOPXBrZDSJLt/4W0zG4INFwSxgPLfVo63Ook8uKCfRQ/liULCPRJs
RwZ4Yj5Z2hJ6Vs0wKgumabyPUXEqjAj15AHjosT5QNFx8vPjXidmVTClGQuHl075m9uxFAQRU3fM
PWaatKjxMMOB4JgY8B3BCdPV4fDsNGbABcVL+GDX7jA5BYm72ZoCbL/BPGa56yF8b6wAwXNl6Goh
o5XUqC9C1O3Wr8da594kUCyO0y88dOXdBeJEPKhInWJS/gJrgUiuFlcc53tdCNM1hb2OGdavxRt3
c+YC3JBy+9F3A6nDYs11o2wCbspLUiyThgknRfxPhdwYumKWxICfZWhqwmNA0OKLzTtZXpEQxld0
hr5puBrg274PMdpoZPWXmS6msuiYhbvaxs8l8GJKhg6vqTQ1dPUYTQEax+dFHqL9dqAY/pUNRYfq
ziC9sm9aqn4dg6FC3NYA1tsvtBQoxnQ/+G6+k81FjtNnvBAeUk/HJZV6ejIyzzdz1+Tc3Ox3x6t9
ZTDjqczBhNqbGj51BJwpNTAuTjcb9uKI52kuCDXIxxvjTPTKp91BxBwj/HvcK5gWacOzR7Wc4xOD
8Rakf0z1UrlGYFMMFx+7yxSH6p4KId1B6octXC1xgKtzecyNs8VI22E4pfuWKNlQTnrI1AD4cX4o
tYPjfyKRcJZV6vWAegwRSlXW8PzUw+P4oVpIZchjGeQGOdHyKe1xNS+mzu20Ws5SwxhKIt/Y+ffV
Qqw5M0adMV93IdehCAiOkDNIq7iLw46FYVikDr4Hk9zRm2GZGWsUkNjwkAKvpOIittvjctp2Oz5G
JGb3lkcVaHqHB4Q8hVt2qp3G2zFlo4oLGCqdbdbUe6jXYs1WDuoppTVS1YeTzhmVeigIo974WzOy
ynqSWuAfQGp7hDBBh03DIFBCNZyqWsj5Ghgil+nmamR8HxqsiY7fLiffd/ERNaiAP2W8w6BbFaSv
zCWqS6EDT8pJftyJlScGBqvGd9e5IEYRF9lmNmg2m/i471Iqzmc1AD2H8Srq84lk9++sSlLfx/a8
fLg57yhGbDFsDaDtwFtxjxawrmkfrTITnktmQX8JgNdHxn2tQEpv+7eEFTww6B/lE5Qb3QSbEcLA
sIlSczyjT8F83nOGAawHBHfEAYPannFDYYctQ9Zr14bkcT6X/ILuqCfZjxmD4gmLTq/Q602H2Ruh
6eN/GQLqbnBWyoMSVagM42ccE1M5K+f5/mgEBAMiuT8DKgvDjuTO+T+z8xAxgqyelXhx7pXWsMBK
cl9iQFid9FffV7qBNxBW3e2OIYQsl1+xHQ13QnocMCV4THcClh0X3b/PPM+xw929WKriyuSzrUDX
PCSoQAY/jkQVz3Lf/RSYFV5Xd0umWxYjSWyfffipEJQ6nqty+/Vdl/Rcs3eGmspDliNt0owhKigs
uR4SzgXZCe0L3OT+fk8q3Rj0FxqIUYGqieqrOmrCyAVJ0/kKlD5jjVLkAg/phY3EhwJ9Vsgb71KH
mboR4KRE5ht0KaOsSANpFYeEbBXl0/7nks1US3Tynr3NMKQPNig6d4zBwyTTrLKFJN0tJX5jgWUx
qu3bKY2Zlzvq/0temHOpESWVWSa+LCNukIztlmCaoUAJTnXNgf0j8ehZPVn5FnMh/S3a956ezUkf
kPxa0n1A1+6xlfck4SkqE0zeXPHCc/vOcqsoQGHWaP9/D8vv/hwmaLtYaNENpLFBzt/9XAuYQRmL
HEeSVfzQGz0K5uxl4dyIOb4MtiwS3F0eWaQu2j4SuNd43a/DHw2rpt0DB1cgEST/QA+aprdL/Bd5
SpEz0cRSGD3vXha3v1nFTFSuKjKX+rEloBWjYf6mFFEdmak/otg1CknJ0ZYrbOdcDU6BxYWwClRt
RSCGzo5QSwhuXkUA/mbEMoEiYEZWQ8SjXcoy4fA7w/oCyzLM+sqyIOEB3dajcbysuTeE0R8jmOON
R7crDbjANLEA81fOEn/iLg1SkNNiHOa3iJZ0o6ryklyW5RsF4LIgts0p9gPaYdMrL00o3w/EdoNW
GdizFqexwN6fsNGTarp291s106oeRIvo0fKmSQpXSVYiQMJLnJ5sg9oaY2MKN/1fjkIrw8Tngz3B
9Mzy+tYU2HHxj8y3yxcdzChyuzT1f9C4RqB6b2yLF53T6cfk6ttyV3k7W0p9gCXH9AKI9hpgCLk5
FLzs6hJ7rffNzQCMJelKoCDH3xquo3yLXILnZ6EP/pUchAboGuiz0pz0bICOUy5bvsZSM2rNeLZ3
ufT7tVexMHuB8wAihbNL0l5JPFuIJogKDKSMfWCL8d6eI4DOyw9KX9+cNAVL3HXdKsQgyPwymZmo
RiQ86KTCqldVFjBW0W2IRiCNqt44m5Bcbg1UqhbNDKfeJdyJrDdNGP5+RAXhUTYq6X4rm1aINu5X
B6rcV7QzxOZTogwHFBO7od+COWFp60VddDvmIYU+l1U44lxmswmCKoey3akZMogG+SQkaxwyqLKj
eiU64+dHL9T1oCAgkVGy3ml9H8fkXtb4XR4z8KgxkhSFfJuZ16eA+ahUQgisHmNB2SVzbs2zYbK1
azyRjz8VmgllVbImGAqfw7eZSziFtjK3OO/qgWzuxIpk3rsFeVyEtV9IeB2WX4rkIMd/4iqA6BAi
5XwTJRNgEp3tsw55WvbAldQy1M6qSGHrIrJZSA+1adSCYzDNfnMN9n4n88++G3GThcNtQpUD9K8B
P0S2NVdodEpnNpWO6eKikTqlg3D4OUIY9DMZwWyFHAsjB9UwbW27f1eIVjukK4KBH9rDf2uV32XS
IlHRouRIKYnq4GBKKgv3qbYpYX8kYvfUQqKGj0ehhX11gJEYnXKkMOQ9U8Qwg5sjyWIwFac8JOjD
/Vv5uk5io+4/tojtAhQI5zi9DhJnq27Avgxwagf8mYRvJxk53+/OxB9oikTfF5mNqGgmfqInLGgZ
PR1xSUou/LMzFLuLvly2Uh5SLS0YXcSiv77h3BWR4k4peDttCn1OTvILAaNfkJ1mITka+jfl5Cqm
a2Pd7cZKsY5YTDl4XYzNl6XqTJAbLHYVgEI1L0k259ktZ8jGY1nyxPRgC55WLcO0y3yavPS8KHls
k6cFIlny4L1wO4vGSkZTtoNOO0Uyd0QYk/7JbGFl+QjHBMjmmRvdEh8m6T81jizOVdpuS/7MSDux
KulYkBTmcAIUruFa4RrAYYaIjMDSe8/psxtEWw7J+D9yQ2QcdXQXdGU30CTnYYgB4vblfOitOpoR
fmbJPIpWQLMT5/b2lP8ulEQeJNmd/Eq3H9BMFxIrRoERxCHzqQbkS97nCFHa6lf/GS4m9jk+F8/a
n5/TIaIUEhXeV/U+/HNUTM50eIvguU2rGtiimuLxBobPWULCZX+YGbmYbviv0RPqsPBGoHS0uoyu
sNk+/gLYlJTXKD0Gtt2X6/InIGDDiCzZMKysg8N8FZGb17PEo+1jLWVbQcXzx44LJrS0r7UM5SXP
7QG+uFXch84R8KSZBcefG+99zwWz7CS2Bdku/97B4geVKh/WWcZ/y2mF8ijcUcFW2iXzS/QaNXKo
zhXLwkQEupIpgkposwe0a7wZJgMKn4LMGra1Oup8fBCF3lRSrWOJ6LGRuaMwZxSWrKw1hIG1F2bR
ahWfVD8iU6DgbawaVTwaHT8bOoEDDiVI/AitpAn89DXH5Oyro/onC7rX0nhsSxbVLEXnj1HpgseL
aE8/UPySwunaYXvtZkJEFMT7OzyQnYAyO5AXUrM2iPc2GmAGFwNBwUHSCVJZlNgTaTbDZ9MnvZpd
zjBlE+aEHQ+hQfugdd8RvOl2uXeHWMIOA5nII/pnFRHUI0gpdpYEK6cD2IB9OXQf1nk4npHF1GDt
0ozPnahiMwOIQHW4vGp3VUomoF3nPxQxVroykUuBdrQPQDMnhHaImFVMX+12Nrah/34BLbMPwFu9
wDgfRwcRWnSHKvxf4MruuYkkKTlPMikzDqjcczYqWjcSaiRlHr6wQW0N4680buVLQfeADZzFbBXI
QuzoN+bTxuKXrEG7dRTfNImqBhCtOtWjTe1GL5ZC4+b3DGbV6BK7F3qPh2cUANOy1OBQxd6v4S2U
2SVjXCv6nWm5JDSnPLolAQgNzJxT6ZN10CK7CDkyFEyE1SKIYBOIo65JOas42Wh1RjNZ4eFx7hG/
Oeqsk8WJtZvoisYv6u0r38sTh6OZeQAhgolStPnGpBXyfJosU67tsSbYOBKlDO3qYN6Vw9r4tt7M
k71jResizib+bMUcaEh9Yv/jaIrjM1ZBYJvt+Px7G0bDBDFy4YuH9toYEeqJqaT/EPVDo+CLpSZ9
/wSZB+5vYKauiSAXXPHNPjs1ee5KiIzWLD9KPHNzVFVZB4OpPKRfslPpXr1xERAz3rxe6wDhsbtz
JUo9zVB32HZh/Tb4M3bIa6tfnmNUxIOV5n0guiP898C4Z91schuOxk/Tw80nmd2ZRjt03qDG9zKC
o/xOyseb5NpWb7vt5GCGGgHNPB+2nfY/6VepKTH+QKrnNgRLzApycW+mIaYo/y+W4E8BeS+ujv88
rFBjUUNFkyG/1mDwOLXeYGWMJr2d1h4awo2+WG8HcrCANWw6DEJKBwY4FY0REmexoCtLPdh3Pp0g
Jz073rEQ2jsVDJGAsAKgEC1d4ijkoftx6l3ngSw4J7wM5/HogV0YhPjmhzw20wjfY4ZdxxIjWO6w
46sTOiETkIGZmshPKk7rUEDhFvOxHotDkjliRCbnXN6+iGu4jbn3aj20EVrwQ/tnKk8xmbZz5qep
HpfQaVQ7ngG/1Ip5Pz/L3PI27pGKC126r/VOOqzaDupEITjgCTOhDN8LIeYcF5jvPoA7pxHPpPDv
YrlwkqDvEhlwStKNKa58XZSOSf/Id41TolEEXWImIk/6SHIgoRVHxiYv/YTln5wY2ewxFynIMgbB
hOw0ESZ3NIOAtEjU/9TrQPGcUtY4H6ecUhwClqR/yTQn4V1mnBXaB/IArEUvFItrkziOJq72QQ0K
DU5jWSXLHJs9sq8o8ZtC2AWtl6g2JD/8NLB2ij3DUZT98YybQa8yXIQ8VlQPJUhpnDh4bHEwtDx6
gAHQZaU9cJ6ftNmbvyouvHwpeao3tfW5GIZbxh9CZdq/cSZt7hsDokF5NL4XMxU/PjuchPNL4+Xo
fN16CZ9f1DhOHttmd+je6HB0XMmqri3q4BdeerkdQG8wCpgxkF9G115+kYros9Cwbw2zvLnouxe4
tflOOOvXbfpbyiffcfvQTtzb8wTsxkJcbTEnCinm+7J+CZecjMv1TdJKGVZcPjiXdTAfWqII60+e
nJEp+Vmz6KgfzaPf3+dJcD9tkOj4OmRFPWY3dt3pyKJQvHqnvUarW1sp7fOz1GHPiObZiHPtDokc
8aJVu7cagL//d+j1z6/Q3Z1YeObGlGnUoqT0HYzM/vXkwvFsognyfjjN8WrJoaeAhit3FYaOakj1
PviQL0JPKElGgpwDueAqK5AkHkgWZHdJ6ZMToTVlM8MtN7sJtOehhhzC4KcDr/A7k1Jcwk7sqd5+
GjxwMAx3+V3pca6YHKPrJzRdgDGlOQpx4AuQCOCIdlEUwhXVq86etiUvF94FvMCaiN9/OjhVkUsA
MR9wVyHfnmPSftP4wNOildhBBZYrm2EaZZFDfLiao8akyxbRxYOd4fDACWucam2rorjBEek2g2eH
yZGo5wPVLM8PPaT2XTC9X+V8Gz+1FZyBQhH5Eous1Pmv/0S3vPSSeJI9qHT0mB/jOA0ByYYO5RcP
cx9Cnd4dWjJ/Ui3UXt8klwKfmLlEmqVX8CmGBU5GB4wwbgsxwKCAUi94MS+YMGAO8Q8tc9WVjD83
QqF/Amqhve886A74CnXRipSqZYfe1NftcHANyN1M5ay1SLx/KTFuWY7y7z2N6wFUxE1AdWVFr92j
gRfEZqbh6G/vbeYVCtgmc53gLn7e9F2uSQCwr1Us4r5NB2YKvFL7/loVpZOikkWBI8dXwqOnM3jU
vwfmrdXgjDhHbtBUpOCYvyOFzhXlRF2rCKZtaTvOQHdPDt5ecFQSqXjaE/gM9VuXKqvZgxhQJIpi
AiRwwX59kqIx/E0NjiAzuzSE6u7BEnvsc3qy+UZmWpcNNPnch2r/PxDYEnJ0PEz/aLuktb5Z1RDM
UnuBifj8loHVFnuOyIfpf9NFDU8I2oVaL0UiuuDao2ReSe5lmQMWU7HHa7iq6cJGvL6pu5r7Xtca
ccjezS+tJo4Kd3OBXosMLQWRaXKjqnFn3T5zqGTK5c4G1463of9C/4l9yf7qbCPQPB973nEIEKp0
Et9tDN5E4Z8ObBJEJaFugMVusN4lbIywmg2PGOb2BjlZFQe/cTtj+kgjXOD1og0PZYK0spU4HwHU
yMZHe84Ph0r2LrAzGoSHQCxgj26KcfhYENjAVfRfHUs2N7oIBFbkF5hA5b4JgPwNpqwN1m9Gj+jj
VyZPxzDgxL9Csm2rP0PdAbsMGiFFNdnLpyAP+ReSSbY7Zge1gkGWRCcquxIGCk4LvS5bXNPhUAJk
OEDUsWF/cq31Hpl/M/KJs/aqTrAE7PUXYOTq2sliBRDH0XjAFuhtk2S72AVTS5RBtGFJ9bGvDsbu
KZI+65TqU+3MIb0mLsC9XTcEVWSI+YqR+A4fcmZtO3K4VAzHXuZvSKcs+NUYK+re/lOwPFXgbstk
5dXiBBnSkWgygbPeX66j7IBVWERu5GL1WHp8AvqXaOa09C1GisWWf2oNMF6K+i7teo4IXdvGlE5W
bSJ0B6Dn8pVn+qp0QgUXJrySwHEeX29Pg9q/+faK4Bv0yUIt+PBZjwrcrRc+yNI6kO+/p9vyjbrr
e3pQeAcpv4uW3GuyX0n+goWq1AL4xd8oxlDNjOkN35ZEJ5PbNDdO3cat6jv1fKOLbUkf0H7Tj1d3
fBhm4TPtb/a+PNLi48w+zSRAJ6i5LspsQo1o69wRVoejVLJWaoqWUxc2cY+KyyGqOevu/2RYoeRU
3gMh5BAiLSjaJr5EBZNtUZjALcGMyYpI/gQ+fHBeufW+uUK2gpQBi9CrQerID3vata+imrpnm8A9
hF47KDuIbatGRNYvari3Fj9KAtJj6yBb9HNEucH+ePoGMzr+N3D65PPiL81KhLt4WbGzMRVDPjyI
rG82pyqbzB4+vQmNYP5gAjgj8xhlyQWFGmAAPonHDh22nu9u5jJkutMp5HHk25tad0KWSQ9TpVbX
EpSG3O2iLlMpFHbnmUfzzOWqfKQfC1wUBd38gKU3zWtJ5RdmzVQAwgXFazb/0HIPXWl7jonHep62
CtfeAEiC+c37deCs1nskVSt8DwNAwztEomLVDr3Hh6n1YuRhW6rqkc8Avysbo5xayZUELeCmqNJz
0MFgsXxmYuk3KqlxM9v6qwZxQlhynQgHlkaavdFXJbtxgoXb1WtsAtDPyhbj5ehqXpvPjiQBcP9+
/yzxtDqbikwL1Ymr4vKQsD8IVtgG5/vgAvt3ZsoXI08cx54+ws/Zsugg9vG6g1E9355lyWwcLHh+
NWJd0jvbxZUpgcpwzDkDLPIr91aEQmXoiX79Qut26T7V3lnvaSGxQAGMD8zNZNeJ5pvHmEeMnIOY
mx0rCv2OnjuvyItKSg+QBIQjNqJiQzsgPRVvwcjibRbyxF5yGsBjXugHz/aLH1ZzaGGLa08yTHOA
0C9DEuoYt/wvTRv1Bi3kRceBENLvi9tHpHPiQWNGSdpG+X1nfGi6rB7wGLUd1He1JcVLcxww34Rv
aUHKUbvsu/YYgUoWS6HNvbFds46rFBVUq8nO+UAh7llJDQKvjVfvTBrUj0yxHP9CwRWy0ZKdOmTF
HsEYQ9iEJMhSjPH/V2/Am97w7VWix2sLRRZIUSbS88HayKePc5EJXEZYtB5O7r1P4D9Nbu5s17Sh
Zj+m1kuKwaNqDgDkX24fcQqleOyOph61688Yj+iEuJoMUkKT00rH/ZUPAHadmWQjNoMO4V9HfIyI
JNM9KQZYclgo0sfrvpu0WK1E9Biq3t6Hx7B96wQXeHi3DUtzYiiU4RmtwdOnx8PEjNcQK6JdWMdu
QDRq45pghOlDR5GBG526ZHksrcsKzkwyzkU8TpvXUFE4UGwMMnl+/0lup/ADyHt5nz5Ar0RHYPcw
NqFYkdisyr14AwQXIjRuM8tI+v4g03VY6d7svhrGV8dOdOyELyLE116sGeWWwXhrc3nGqrfGjDUf
yhrZgSkHyjgE5YNiNkUdriNkqDjW9su2Y3r7YwVYlx+g6pvif7VUo3P2BVnjNOGRjYZRXB4rRfNt
xG9XQSAvgB+c8hB3H0MXOSd2/2ryfJrjXwL/b28rPcM40ARih2rpky9JZ2lR3n8ySQYAAny/s9Az
xvfv+mgdAZcoqIsGSPipd7xw3Y7N5o+WHsKAkHXG1d0/zj99rGgxGzGlm6n8oBPFGQTVC0jHdCfp
KxrGhlwvcvs/hfzp5uTj2VDW2rV/Xu2uDJ51Yqt6uXAjw7Csg0ACa0jlV3JZ5QHa85yZiYoTewYO
761hESr9jDHF3BXzAnK/v4j+NFXV/2WL5kupcNRGTGl8lNlSBCZOQd83cjhvYynDpFc+Ktt62/yT
kJYy8psZMcrTdb70UP9on8LsKbWrGPVOH6aSocxHVE0T20yolAoRY4qpN3KHEapmzeTVb5NsplCz
31Dy+7q78alDi24Yb14f7nRMBu/ObGqe/S6D/fUZo2H5MgbNlxrsxo+kR+70XKWldYkVVlt5NQF3
Vdgr6k0iTCo2jGy6Dw0kgX1zytae/CDc5zS4JJe/QmPEK0MsN6nDmsPBDQxDLI0ks1HSNI/N3RvJ
HzP9GMZ5XBRbrmSQ/7TjLeYlZ3DXxAon1psu/i2djXjctwlW55lhZeQNUlKT16sfZWXxiVGzgfBn
8mmt24T11wHRyr/1NqeLN/qFiR4oSpoo95ApUvMcZJ+enYZ9vymtpbeQDYuqtchgkHqPivnxQdcV
4GSGk7gFSdRaUvSfYYLLAUFlSOr7bDHxxmBQ64nFYzifyU5YDuAx7okKlT+v5OyGT3IS7CmyEcIv
PKGqGWas/scJ6+QKl0aUfKcwXisK+MrFoEIr1ZMXS/EyWBO6Xpgwz+QhIvB8tqmDxfuJSzfL0QkY
r32d0d5P85nuqqfezgYL/au7JVpJAFJm632oHgkq0NKgdBgf2W6nDx9TNxMv/wOuOW2h4LwqXOxb
mawpSMwfjYW9X3F7ahB6r0bVoHZFJ1XFIibQR8RGCxyfLgva7kOhgPA/7YlKGD+LnsrRQ1fdn6Wu
SMMLLPHClEKwVsHfbSt5HW5YQbdHE4esrkPAHmn2sEWVjdGSt+NDpCp6Fbg7AgKe0iWHnHlPG0pw
KrVSSs43Z/JvmffEEDQ+zaBoz24PfuOR8Q/HEgepVCRvqfO0urg6oXeGWGza4i6DlUjks+Oo4uRv
647upnuFwP7Q4B+nC9Zf60l9Z2D9awYf0QJwqxFD7gHwZ9/71EmrQP7g/z3/9UEawnGFj9h1c94e
/TGVFfUjeWUVxWMvN8LHYFT8c5yjxtvX0J2joK1kS8P9vnQgqcc/0QE1O0s6vaGgpwQAdiSrml4r
pqv0pb/CsJkED84cTCk9Gm88MpndWCAEvcDtQ0Q3h7AP2CGxXGmGniQrfWB742Anx/7pn5u90Mdj
hd3F06Hs4fj9M6J9b6E30ITBnC31CgD1marqHKACWHtf8VHY37Jk2w8VKVMgnMKWOBPKz5yAPiwN
zaDN1f9OVM2M8xjkeNzaqgIQRPYP/f6oJG98aWzgcq2lASwiGncqW8jGsZO6+BHePM+OPCEFCriM
8YNKA+YWiZSlN/R5kWdvrjLlBWK55QMgwdvk1KEkYid8qBiVbcsZlmeupv84PL6XPI8r0W+J7HHV
Z6Z3zb7xxNvsaGWTa+m07wWQS4VORQ8uJj5s4qGuaAR1oAniM0jCpseuQUVio8nGfelNkU9xVrki
mqJSJ9LnGd2PLXfm2tUB4elRvwwKq4ZY5lYVEns+lfZc96Ih/JOEtwsZR6U+x6j3iCxOjkfxu96K
1UnPvx4EoLY5heyxIi83qsW7Omx6Awjm3ZLs3fSRhfYl5hpxXdyXoqz8MwlWdWZIRr3nOMNvE34P
3qtqH0S4jYOZ8QztRVQsRCyxn9v3nxm2HHYUTmp9cRFJVrMkpORiS4Fkhsw155eaIv0bXhvVkz2V
iOiRkO6WIA9JYcSp/UevcvTl14NaoFdww8lyXt+lWwRLKg8ai7rvWEeVye3YxZnRYD7bs2I3jSU1
u0zCSJBQUMMdUgpb04scOwKwFRDngf0pX6rOqsYNlW88rDTMm35EEmvTjxVtY5Ea0J3LII2c0NsB
TK53TcFie50JWI9iH0zvlljcesw1Fs3Auv+51xrM4lnXbihdPHE62poZPa7TUmhjkhs2BqymUXFN
+Fj4VbXdglgKbUelzH3Al485fxZ7PRRR3mkPo4t/4KGlolG7OsB+Ywt7B1INz3iGzuRfbYWmvC85
gwU0SjJ8piXvZpwAmOBvCCeJlvHZAlxKpuim0yf3SdfyryhEVkrbLLCBJtmOFv2x1A2mJdIq5gde
XYDDn1ZgCaKAotVJbiyAR06GtWjRtlLI0B/Szt90MNvXmjiO501xmqy8assQElLnZlTdBqZfuQHZ
Ivv7OblounD8tpKGcj977wZ25bBvrZYPySCP3tFAMOqfpt12U62rDOAawcFkqFtofI+a6veqMrKg
paOPjDVojnrTXnpBWpQa0rSXdbR7/0D6thbTrZ8joFd5ZyLGQxbE/J9v3AiLbNv1gl4Z4/lgjS2E
2t+h7fZupvg26b5flTaoV3Cyym4O6uKODTMiqNXIk1e8XeTOTOOKvFbNXtTf/p2K/3ipA+GVs6XH
11OuhKbLPjEawcah0kkc/InUnlw6T8/uPS29vzF2poCzJXFLwaMnNnfC/1ZgF4wLn+O3Ftp0GQ1N
apzATxaBxZOqxtAECF8Gwq+6V543OltyEPkxC9XyE/zWHAy5gVIncNqK4bRSGXcOO82Kw6HE5kie
F2ZebVp8pMZWea3G5g7R1EZvfp0fVIXRLxHhCVidHnV0/I71XJZNZ/9JAfYanBcZ/bmbNbx2WcTb
yPJbStXLl0t8bZ//xVy8dh8ykgd3HTa99fQz7aNi3QHx0YfM/pdCdrzzBAv35AEF/+nhlhMIahUO
9oB2H/LFj3nNxmGfTeA7/kf+9zRN9XgYGlf+FEqcLJjJ1aXAfkar1YxVD8/6Dr6CscWuZiaIB6wW
rcJyobcv9WpMltp5o3xQB2CSds2HP/PHoJu0CLD7eu3w9b1zOUIeS/n08tGxWVDMpvkz1UURemQj
t5VWPda/vh1SYwkeS7yqyKT+NDg2mqsl2Hl/svqeWaVjvYaU5g/i656VX9YFySXO5R6gXp2+QG53
mLG91JtKlH804q0LbxoJDzj/ennDBrbSGWLqh2HqsD4v0R0Bxhr359KoA9vEydolxh14MXxmIIRG
r5/UdV1k7PAQFyaQPsALxbJx0E0DlsLaI/eMDCjpJ1piQ6nSz+8+mDl36Trva1KLI47RepJxWz/G
bWfZyLMFvSvV7cERKjEqoR0MlgxpsBVPwX0ozhWkdhcjFP8cseUCDgJM0KTxFRedGdDX3CyYZBgm
ciupx/ir2Va1GDk29/wQCNSqTUehscmRB4wFBUc9EY1Td+WyiMRAe5/tuHyHJnYE23VAPpM9Jx6l
5J9vvM5q7la8JV6Wr3Fx6Q2ziqcXVQk6/rICoSjVNUWT71yDFeDs2cEFJ4JyeLeQbYXIlDqSj2WP
hzcf5IjjqiBmqE9Kw+k0ZyXNMkagNnKD4UNRh7qpHVDc1lVEbs79jevLH+PVTX1+Vb50RuLohFaN
C3iG+RMa6zkjKfiGraTkKdNylLFaT9709PdN3YoaHCKdVgJPq/GSUQujAbZWJcwRusadY/0I+law
O/qCm4ISUW39uf8blHqT5rR87opmT3QnstZFRkvZQVrTabe3rCs2oKPfKSVsMYY7S6WRsk9uSYCH
Cb6i42+qzIG4V3Zv2Q7CIEBE5EKAkG+V9jWbfmEzkhuCdT4gyJLps1VyL2UOxCLgCPCERy6M1DMn
SCh/2k0XyzgzclP47CET3Y4ZHF2ABswACiAdY6R6mYibP7SmskSpkym7sFureILZ1N9ALglmsX6I
/gvm1DiIROo8rhWc44+8TsTitR47kqKcW0QTQHkXY4xXFKIJ/ly/kRlT7lLRjXicQtXKsr1hcpF1
skxHmdhwF3KENqOkijCOEuRIu7G2/PLthN+2yYBmpARRvHAaVeAm0rcV1cYHGm4BDtpIgAWk0O9T
0Qae+9FQjVqtQel82G06W0O1vNXu8ZBhPUr2VMA9xXbqc9sOWbgDD0CCqr6jTodjqNhHhpfHDkAY
WlpiaKPXo35zIxqValE8g05aqJko8Y1a9NSB3PUaoe0Gfky7vhxodVgeFhDMI1nK3bYzk93fL3k1
1AW66rmhSFDOzb/BxJBGsQKLZb398JLFCzXy82+Fawkx9aC579gFwhaVxLY7SC5gxP2ZVBLVD+eK
6yf7RtEH8x7ZfYD5LZS7VOXOTHv2/C2pB9CG3hf3Pvdw10SWZqlOGlBNUcJOtbYfD5heeOfmKQ88
bHpU4EARWfbqIypV3XJuyeEMBnYU1ndJfvMFegBLb8Hql6akd2g/Jn7SYTYm4tU2b14OlROKlLwW
uvMwXIW4NyYg++uFgAfVUe17yQqWb5LK/YZMb/eMeRk8hzRNSn7Uma+Qybru1gkID62/SAPkl5Q5
UVID/4NjCTUxRvePk4tnH686UI6qmuskAo8bXGS0FxpK3icQIlE/fTwMYN2qPl4l34G8nq6tQQF8
/DHiTp0PeF34pHUgfSX+z25deDfKFl8zcALmwPUS02+Lys7YQMykVpqvDsoeVbcRfpoiAJQZJY/F
HQE8K/7IUEez/6EMleIPREuhy4LpTfOG6KucXG75oFE5Lain3gXLXpZ0UpqWocwM17lgY8uBvvHC
6z5omtKBVo706WrDV66SVx9HGzZhOc66oiamdlbsqUZcASxuRP6ncD24R0tIlb2fZt7Plz+yRe5U
Nn9/gIrUUzsEE8xm2178yOaXA6K70PU52NULe3FusaSQ1ABX3IM4uTujF1wykQUjfAd6F7KiIEfL
xFMVrP9m0d3h0JCmehHB7cu0PrITpm/tLWQ1JPaK5diMfMizBdXlO9/QfUVZpo26HeXlog1dO4gn
YZTT681R0OrV/9MJDk7/3OCinV3agjG8h78lamPtrlm6ZqkpUpdNgoiiSfUsogu7lxVo9+7xSgje
gx1wpeC9YGWaZY4CM6iMxmJcZHc79EjTj8PGRFIst1R0BbmbViOFYaYRpJJJjwPB5QQCSN58v8Lw
FEkT7g19+JBj/f6lSF6W0DJnAY2/FknJVIQwJpFRsCM58exJmOOk8qn5D6AEGxGerdOdzF8yVb1i
CKpI4GJaz6ag0PIS1HOKMtGC+9FjKYae/vQo0qJCDUSwbHEmaVdR7BOCw32qKfPgj8uqkI8fiP5W
qMKvQRp4oMTkEeQaqKLsdWFZ6yVgBrmACzGKPJoljZt9zx8mGnvy9v7K8OeVfjFvaFn1ddgHRep7
tFiVH9IdCSAd7WVH6rf9nQYbwveKsr5GA7nDM1MUYOOGPjOfrrhaR0VH6fn6cLBS8PeXhw1H9/rP
wnkZJ9QU+hEEHnYX7nMUseIDxsuE9K5c+oXKxFLW5OVgRngbaxs1lheHu6TkkX7hu1kDBlZgclxY
PDeTIkbQUqj0u5cfTwDXQYM0s4fjxgFpuK+HKyNAnlHPcj3VVierFqtx6C0V+uURNdi5+/DPYD9k
+BB45nPIXtghWMo0rqiSvJttFQVzA/nLvs7J+3x+SamSD2xvxYPx/XneBa1vtcboFRCb1tcK3Qv7
lB7NycSrx8gmdjg4qW6eTanM4kw+4gvSlt3xVG52A3abarzddGvQVTt9y++vwwVUq1aIlUg7o6rW
0ZMlYzj52aUvh8/TuKq5LZtwH8jP47Y32PvUC00UiqbzPr7ABG5IX9BRnnjN+7rqUtD81JJqdlHx
2eigsf4Pbsqqm2kPV4gt46fwNogYp/y+iOV4o5ZaxGPFZ1lzL+EUexecAZsoPTBIZZkCtYhDgFzs
OklpYxmFwXjZLd2iJcAcTqsPP4XeAFax2RH2OWzPTPyBsNN6PpEqA+dIX2yIC/sZ5tyt4lmfghz4
IqYcbDOIG369fFhu6fZgLn8D6EOSWzOTgrsyVEDIV0LVE8sqah+kPQxVhvexNlOdqx6AAQMyghiM
LZyTYCn0lg6L0bXGMjGyYfwz2PN/WeXd+hgb32x5DMLSwzanWRbaHFGImf9YQ+VpxYx/x9u4Zy5l
c2IuarwSBr3Tt3jCpFnBcYg9iUPZtRKtoDB++WQ+ntW+CxiWvx1f65S7BXFABd14iBxp4fIqoteX
dDmY7mjCRmSB3MIy+ECLGMa69w3n77SxZYV6x7LG18EoLw3sQyVmukbVDkb+8y+BB7iWF6Zwe3vU
KeGuf++QyATYdY8U33VWQqDHh1QCMOHWs3/YtlEsU3gEN6lIMgiqjajhxVyuPnHSPFGZ9hkTHGFy
/CH73DHL3NqONPuVNEiYGl2GDshBgRBJ/S1YfhyBvHY846NAMvQyLzFOwzBFXJySmcVGiRUakRcz
2hl522DN3CgxPJHgU3gIFIdnj5A9W5cq0pznb4yHhRB2owKLp42ZAAONyHiOv0sbAJm/zQs/5DiY
noDJIUTNbzWvspjje6rFU0ynGEYwrQckFo4sjRT5RiOIJE9TYJiNYQqVaqX3WIS5FPP6JXLNxnMI
9VnJtBflNTCyLrYperFjl5HCXnA1skwhXWYc6YF7gILd6w33g3qj/u+Gyl2Tqo6AUcxYKLkUOPC6
rLaaZoAPctGYODwVmxBghWdD3eFpZpWA9024+KwKUFKCTuMiXQTpBAENvZdYkyXKBzeL/XDQXfrt
U5sr7F1epLGPRRK/jJIhLlrBMRn22ScnT6io7iJXLWmwgClLBVU456JhmWPxhkfvDJJbxWhl7vms
pJqgqVkpF7kcXkXpd8EtFKSD9qevmneIo9+pcWSBlOk2wmQbdtF19hgE7sQ1J3FWDPbdSUYtjuMH
ac21SN/nI/2oC2hNBdtaYLanPhoXCqO8r5cx8jQ+wZ1fa0zdiTMwLv7s9ozRI/pW06jO4zTui8eB
/oXGvoM0foCwWLy3xZlV0jEVmoh4/8b+Awlv87lwBs4MibGfimTZSpYPmx8L9rZA4xRUUytgE3m7
ru+7ROFYj5WJiAHfM51XkfA6uR/+9tWaV32XZsuz7SiDUId8Jh/wB+FGjBgIJBuFDvRRGWf1+aQb
0fbx21A3SjWS8U86tkHgRkg1Fl8tSpLEuYJdKMVE64NEQZyaoGHFKslSZzUq7uFWUA1xIWWDqy2p
9c1LEO9ppjNzLLnhz+ltlaJLYW6hXIn3ZRYKIS7m4I5kmEExL3PDaU9jY9o10/RSvu8xFdeMmWLI
CkCoRRiqLfPmuAFFjbT3IjYdzqQDf7WlSofjZ99jTyZJFqSA3BqX4kKtrl3h5h6dCOxCLjGV8lpR
0uayRupPgsLwwQ6Rw2JqaPdF/ECScSZYqwEYZm4/znGGtAubspkIrEaf+hLCYIyqXfmKirmIs9v7
Zi7h+NNMMSkZ3+AvnLchjNO5iT12LdYu2dWTmUW/jf9pqFSAsdxPrmk8mPcb3t72yO5h43ndzEkA
92KNZINEIqlyRUoZZalFew1rhWwlWLbXzbFgEpptHASXZTerVVjDabdyxnKeVYcFQHDyHKEKBpVH
JONJWCEHc/nWxUzcE7ubnMWzzUMmJlF/S17VjH6Cvd9EKpYqqL4gPGuJECiqD/tRkxTI4EpQSVKR
5zMSp4jPU2+K2gy0CgztHSk3ol4IMeHlNJxFDdFLT/9dY/Omas0Pdv372fTRfQvZlsORAkmWcS0w
rFhtnirzsEu23xUguLnvlpfpktrjnMcJthyiR7yDryxxDvETNs29AKDQQTcc5SPPvLNoCDa2i/73
fKHGm3sp/5tLpnW4xMti52YE+3aoDaG9hBo4z87BvhwoUoDd4NzDk9z/z0u/82iktMWhoT8wnHhR
I4DkdYBUgH3yADDw9j7YORfCvm8wkwoISzReL/AqMwz/urUw7AgHuJ3yv5jaxA1hq2ljtx4UW75o
IgZWV312oEehHmOUZIc/UKCUZKGitxTQjXcQvOseJ3/BGP37j1Nonur9l148cVh4twDd5TmGmscW
Oy4/+pVKYkTNIEuHSzQOwHPArZA+T6mhuoilS/XuIX1Y0AoH60Ou5gKFqRg4jp+JW1UcVoO90HU4
w40AkB/vMtRM9bx36AsMd7rVm1Wg5CpO+samybSuKhJ1ZREYiFFdoQhkCrU69ND0gKsUbehbUIm2
hxevnUsZKsyH1oriutvDg+1SmjTS38JQb3w/USsgsGt2SBYcGEuKMm0ETWleoMcUq40ffIX0kV5J
ySBVZLeiLi1gyTFM/0e3gWMNCn6+uOBcxX/VFaxZPfRiqTHCQrLAs8ufSPJqwc2aXzznH446Atst
X54TmJeyJKLbChMg9Wl6AABoHgSXtd94oxcehIjgqJOG6furRf0pxWHODgnJkD89ou6VfEBloaUF
F0ZjCKvzt0Mvl1cAyJOKpTzbAhlRjWzCMyhCY9V8J9EE4NPAFvSy0yoU7JAv2kKXtiLRJM18717d
UslikKlKTb0mMCm9A6G0TYCqE7IZ+92rPqO+tVCGXa78J0IQYpB47EPMvGa5V5MWswlNguy+xLxF
IwP1zWhwTyioT/QRc4tX4wMS1xdO/Icdm2HEePSbA6faPMjffBIDZkHaHQcnbngw6qjtNqyg6Nv6
NSgNHjFiqxmKUEhlhex+Y8xF6rX41qXk3rGItTVjQGjmqZd4qYyJurgjkuyj6v//SrZlBgYjEFvw
woX9MkP0VbgFB3TJUvHoEQKY4z0fOLcz+WIsWnylLY0YtAy0wxRpWYEv+CuBZu3/hYaTW3saXNih
W1OaIqXh22MQX0C06X1k0S/K8gjtfaBpFJ8lYgDAyw9fYeVNk0NOup+MbZhmYkqNplU896zd8ND7
c3zMOqZGvdYVokerDaN4JSh+0t8vrbv5R3wWFL0lDWPvzjz5XRqnxuvRr0vGjaM1rHFO64776+iz
6qYw1qkxdrWx3/GtYjvdgaWX24kcrX/qN6LhPvGgAU0Cn5NCxC1QyKBf0x8K0BMly50c/tTeHBNb
fy28zHFMfwO3AGJI4OOI0WqmQhmNJMXvZ9Gs6KODFCOOZ8P+zK70/VM9eDSOyO7VjOYYR0zCAnV2
/tnoZz+zrcomfo2DOwpOJ6/xnmGzWxREREjTxKtIQgHsbaj4o7N+HC/TTKAQFYOfUawFthh65ITc
7pNuVsjgG4JSQABEwSd97Zz4fok0ckD5paAGxQ12VnL4nwkyVxv6kPQJd97OidbL68oTgREbi+DN
75gMFZX/G1uIcN4x1+lbbr3roubFBlB8h+/5FPidmfzzTIairMKYpacc1R9CkMgro4djCABAyv91
SU7QJII8yefdsGkSsUPq2AAD0fAH/amwwb+/xlPb6E7wXVTgdkiwZ/ynMVqyVFtW2qert3taen5k
0Rad5i9mOnX2mLQKF0vtCgTrSs3UMCpjFmq2GRR1cae6PYx87DQGy+ETJOM6ANHoN60B+63SxayR
iq1CNvxEDYlR+m8J0eBegXgXetBQVjqfEgtZP1RmdEL9PHDlBy66NtIl5Z0wZyMt36EnjXpqYLNX
aTwMKaB8rQD++tPXjX86chuJ/ES4umClR1lvOBzDiEnDW7S43+IlvmXzzxhrZiQFTahZlJaTdCRy
N0p+h+GPKnXA2YZShfNbK7l1j0m2ZB4OeQ+O2IhgKVuB+EqQr9KsQ38mCiE2/ahTscLvi3UC0Xw4
kAxzfzzscIQw92O+5CwQuV2+wFmUATO4gE3xhDH/nIDqSr2RjhfeiuXb+jp5lhwldyc5h3GQIhJI
6XNCYwc9PyIiTicKMdDRcjzo9mdDDfMcWAxW/q6+xqE0jzx7KrIwmg0GNRPP1TiuQvVKkoDp1Vlf
IHwGU0cVdNuoE0djra0pOWjuCXEX0hyM7Q2Do7AnPc1QclweRD0HKfgUOUFSSFJpBBrhOI0edEBy
07UK9Nz+coTYfhw/LLqgV0euPxz4JJv6yVU1cIP/Jgod39wdIhum/rlsgoUs0uyz+ir2GBBZDq3z
ky+dF0p6Qqf8EMOrob6kRK+p87iyaB0WcX1egF3n4UFHUsd0pAqVM7tibquC4BBY/bJM1GDngW3B
0D94tjSoRoD29yDYWNJzmpar5vK1fx/3cnJMSH9ys7gxqbqxSL7wtXX5pH1Jg7jK5Ar8fmcUv1lv
EQ40LWlISLUVhlAI1NWC6d5HmRl8OxSQhL47M6Ca4UHw+o90N+xDuAKzlH65ok6FWKc/9miKrag1
iWupxAXPve6eJAcZX8M+xK6ollVcvL/pZQO3YkL2dBuuokdoF8i9FbiQ5rjVujaVwS0J44f8AAHk
SIaxu6BdC1Ndt/A7sBodGR0cQ3YNSSHMeNfrINpJWhCZNl7kOprFnAzYtGNtWLjw8s9X38A+hO1M
0NdKGIGr8w3OR6+HS2rW0D04+X0osfz9/pZqAKCwazh2uzkKFai31zGhEW9C5fmDdLoAC+KVQn2X
bHekXZPg1+boFwNBGasqUUPIZ757hWBaanhM2lkT11JD/Y7OQExAsOeoXA6owv9Ud2CXcM2OxdAV
9m6qRgmbzqCAVQccbfVNhenaN0JVFFY9chLxJiMCAje85hICiDpga17F07Lb7yWTwyPr9Prmf+cS
KkdLIikgOKb6CMTn78DW0QGOxkdeh7JGqoMUDxqVbeQPRMtMvEz7CBB08hOr4SiIzgyxSPAa2wCQ
n3epA1DTNrbpLmkPACA8kxmQVdk9vBrKz3DAHKr0Dz7QmRzeEhHGG3niWMBF/eF/T7DLIZQlhQ5E
JcTEH+3aI+gwoncJVxvgAejXZFLpdhHnZatQGsim6ugXNwxHZyeP8RKfA6dmpI6ZbwXqv/OAq4Nt
it0hka3GlS6hBOODzywqsajPsWNjYpJOyd96FmvDV0K9pyKqjpXEIinjrLGNG/25Kgrw0l9Z6hiv
6B1GA80gkTMPV2giR9py6AhK0G4V7P54Cw6V1OmlaXdQytw9hL/R+F8RjfTnVq0Yw0k//cJx6sis
T3I60Y2QgXsANz/pUFdR1gjlEoh19jRqcRQEj4KUsvBlAkoEiKTmGnQhQ/TPqDMce2LzqA7tJThk
v9vJiL31AJLHrYL+SD2fcWGwXSHHt6jl4sUdh9gWki4tLCkBzG/ffkIrZbarlFTb8xeHoeh7uOeF
NuAOS0T7m+5P3MOVATY6UCxRzlbI/Z/39fri6/l9fs2aOAgNGv69g6u7h6ZfmgFt0ryTPSf4yyu4
25//68vTHbCjUqMDdLyAEVzLZyjs3DyDN0k5YQCftyqvOEpyLpLD8E7y93aE9veGw258qOSvP2z+
UqavFlI0FPa63QLBf+WyLOoaSFBw93ZIyiWmZTGEfrvsLgFrAtXL8okjXrA99hHoUQ1Zj8IPaola
sdUD0AkyPuSMCBqK4DvAEgwHjLVZAUJ6fMNKzkupqvRtAIpTMN9S6i16SgQQ7tYr14ctSzZJDCPf
31Tcfyc2ck1hlZOCDj9ShANP3ROFEzJY3sGd2HqG4RqmH2e7mIoV6a9hekKPGoTFPfbtPJrr0gEy
4SrYnuc5Klc3R9Ex3W6VorGdZgupFfgHJMYE3Mpk24FKsK4fMIV+JIsgbs8D2Wcdamjq52RsONIO
jgDBZ2ga6Yf3gWyHCmJs5piMWznwfBG4WA6wDjtpASX+qD3DSKhCwEbe5bi+lB4yGWlAjFxu/bS4
G9CgW8gZZaxr7hkMJNm2vz5XooxT8UAquDh8+OL8zpaG+j+/IdVu4i+ikycSwRm5aYmZw7hYxQM5
TwRtG35wLfaHoVCFpNIbYWbc1g4wq5BiNv1WdqkVmTFAwyWMXo1bqiSy93zBaBQEjKV3bwv18XOF
cxkxy3ojiaftkBZuh+8eZIWKnqXu7Qouc6Caces0/hKR55QpGG+cPfk6QX6LSDLPvnZY0tfy6RfG
Iu+J+/xmvdyfbWjRUBSspyzmOX7eHtTq8zghdbYcP+GuFKZtIkqxsgc3oTgJX943k7A+eJWQf0QT
hHgryqwK9GAlfbG0UZLcwGYwP7fnLA/2BjsSXqLgKNpUi/uAE2Hls7fhsbDHoq9WzZ+fVOeMhOux
q/Z637DV8ySzHy8m+9mfjdw67Nm+PHp4TMCoEqJa91qgC7WOIPTQOeL6pPbpHP8apOPR+haAEL+D
EuIcwfKxUd9gYGs0WLeMuuHktNd1qB316iP0UOjGtEbzFfn446cIgUTZbD+OInlxGqaFq6q1UZ9w
irWPniSLL7mj6bxlYyK7fvlOBhKlujF+6CPij4Wc+yoxhGhOxlISxFt3Y2SLsCsPEt/MqgrmywR6
N5vktgU4RKynvOxXa45WRpw40dElcrgcMdewsoo3cMv+aGN15TymLyHiyj6cb/kw/VeN21dIdIFL
tChY+b4lE4F4K4HjBYlGdN6MU7gq2DXdv35UQSd4Zit8AHcGL/aoOqCeGwQ1YKeRbswsD3Ezquti
IPLs+AJSEqIhWCLU54la0JLaxw1jdO7HhAV2H3/M/ycoobPU38Lc4FDXsNEgDCTjgWP4+szH0WUY
h8iKPNS0Rx84PuvgSEXd+bb/KMZQ6K6KoeH7VCy+cBjXMLK64kBAsgWjDtszvBz5ydLqYJ+2XUv2
/F/ibrNHAPr4Uc6sM9MYJwmL6pe6UlfOBmFV6wD3HxsHiqlSjOoFJPdQe9wO/pvjzXmb8uHdKkeS
fOAlUGbqw0h8wdAdjwnXrbKoSG4oi/Hgxm22lB1sM+LBI9s0Qp1S5wS0/Y69UI4zTSPHtLCFzCRl
LfUceuS7F7f7sUNohGuQgeDjT8V1hCSXol9OzetX4Mm4d7m/CtjZRDFVCTvcsoKBTGvIqlhA35DK
bTohe3vJuOaKX4//nM+aUDZmmeILFvadxld8oUpWHnlNvDNXH/MuwZZtZ96y8s9uC7qok0WRDfDo
06CptZllaIlcvENeGmMuuq3yQA55fT+I65eMOt4vQ5FBoentB+7pJzZqkEuBPr3YK+k4NQmnvXiO
zFKelJW15X3EOxpKrioBDogiE+kSHRq5jv4AwGwpO6WTvZ1q/+PJx9C8nSmA7OSexiuAILzq7O0G
olGPHVHH6bQ2z7rT0EteEH7v/ZOB2uZBli7obg+qCItbwsjkiZk7KkabLD0X8oAYByErCwrJgKKA
91Bk3ykiUqUhouW06kQhs8pEigrab5J7G5Muo7eVdxak6xAGNoaazd6Ar7I3+459YSf1J2rDrVd0
f014Dnsd/Rm5cl22rMKLPG4nubjZhJYAxjS7XaEWOpGsnJyAklEq/+yfbjDBirRfvuN1+HnmNP8l
Ve1O+PIpN3uik5p40FYbqhaEuWFmpqOecX7moDtj6ba1kLnQiSfRrU6wPFaIq3rM0N80VuZlHMBO
bGmHvMx8St0Xaez8TTI4AenkcJUEfCLEyfFBgQvcwcDq6Edlg0RErVfU7vp6N8mt+Bt7JOQzgxEW
BjtqkAde2WH1ZupGgP5zgTggzWf0t3NADtHpw4PvhGfnELK0Le9BXaJZm1iXi3bjsZEOzXuS1IYJ
GfsNFebpKCRsqrH1Cd2sG7illHfJNrUPMxVhFDs4yuCHCnxiAHdYJgEknJ6SxtDzeb7913O2/G5H
qLbll1Mkm/HlaCK5/ybsIxvI5sEeEMiGpS2uNYmdN6bIBzoJT1KvVF8NL9onsTApPq/feaqjHlYl
AiDIw2UXTOWkOD33LdGreK6XmgU2j6TD09V9WTXX6LaTxTblxtaM0qWXrRmIwUMe7qxF0B68wF+5
Vro5+4BIbtfRZd98oZT57a+4/SEHkuITbs9TqRwr1e+t+GxnZz3c9Fb7Feg+yGQenJR6YaX91b19
QGCuBhoSwBpphbF7s/7aJiYG5YUSkeHwpfEzfybEROPJuKiaKmpgp9223W3ZXQaglMw5u+040OI5
GQ+Z7BT6VEePs3iwA4wA941PzbvY3I9hM4kFXBRuobcT1chvjuWRtyvJEFPENZFUGv4pb3YWdDXR
/dUd/hbOIfzPBLDVEfUzHFeb17IriRcTlWG35GBvwzx07CmfzyLDrzhtajPV23f1CIhpcvgWBo2G
dzScWF7VNNL5WXhbbuRdR5VKES340yFc0YT3KaJ0ednlIcP1ocsnqAWUQrK5ibMDqTlqkTP2Eqem
m1mucy9oyWc4HfPErILJLWXr9vvFpsBYLiIfSSVOynjChVHJIpBnBep0v14fOm8Qyb/wWhDF0Hyy
62/1fZ447Q+7HHttaXiEtuVqLQhRsB5bNe7zbOT1JdxxwCnh4XVICM96NinUpUlE/4fjDsOF5PS2
d0WVWseOJsgYh2J37VRklTkrkfOXUYAUlX1KEqNvC6rPveADrpubCuksvEVpQTztZTNYBbHhygth
i/l8kzqcjREY97K86eD82NK0Ti7VX8fv0VO29Fi0LCgn/1nCiw2Es5A2hsVn4DSfbNHqksFMHhMr
XAFTpWd3J/3MBv1tkXgAVemEosqHBdcWNALcs1NvEyLldFtcyfVB+JBywfwufiQXDayEEw/jzs9X
cT7rUK7BcskgYdAS30SuYocUWcYv7m9AlE4E+ONtHscTJzl2ll1rwj79zmyPMRue3xPohfug06Gc
X4Hji5+5j0hMH2JD4djh/0KbW/ZpvmiB0tZKQrDihNqjsTUQs8WPmaIwYvszAv58rJ+emA7O0QSY
Epd5yxVUyCGfjcsajw6oeU1oaKP6uqeQvWrfIhb8zYXeUZadJ3p6Ug0R4AQ0ZM6uwLgerA8rP/q4
P3Ti7dUbgCO7c/fQZONqMWNjljfPRL26tznJ6lGSHsb2QLzGvuxxwD0IrFXX/dTYgMJ/u2jy8atL
lOwgC6X4bWEXQLZqhZSBn/ZgX16tbFCeUCqhPgSrWDBPm59g3DmUkkAppxb0T16h/J5490qIiyu9
/+xCARQiXESbv2zd77DYIjpcvdIdEqCPy+ySbFrCw28neODW0Nhz2qkqSIyUlj0dQeJs9IYMIti5
He+cAwafbyW1cIele/Lbo/MqchqzPc0L0hqmhLaoGjiqq/UGFXAl3i/QmZNQOVr1I0/Q1e+z7Y1L
2ajS09Lr4Jw4GJlUnVRahNkQuxyMYT24dzXY0hFU+12KVcVfMyE4u3BsBCVJN3t2ni9UTHRlvRpW
PMPaWNq4x2Y7ifmYxE3f40bmkE/hNjvbduE5ZjPEYTmIVHXKM1OUXvbs+aRQr6uIOrCvT8kzGXsI
Vu3ZQQ7Huba8KeM3uWSRUbAoUaIDsjaYLJPV7TGKhpXPKO3GuOPz7O42AFCyCe2GQoVAzfFtpgXW
xGyPWlUkG+obCgDATZWly30NKVV4QFKKm1vhWVE6WLzG2oE+3W0dZcV+RpyGR9xB9tS4tWYS4/Ae
XGKxR4ULz97uFcKrpmydrsoje6tp+/EYEV9cRWjHEpJsr+D+r547R69FrLDxsvCI3CGaWyTTbfB4
rFouwYDEgIeMor8QqxkFlMCAAZZotKjZSXhYEgACnlopt+9TfoyIV4ozaarRrK2B0AL4G+0Q+f30
+hf//QOkO8M83DJV08EcJSfeOFDDhd9FQzC4pTI4IJmoVgfetzuOuCcK2OOwtUqZLG6wNVzoihMs
kd6cb5IhJ+whRbTaV50qkYzhN8Mwb8Y5accTgBFWny51PWmmB5rVf3yGTK01LFNa0bwB6wGu6wfv
zgOAEMT8fwK2PT9V4BfSNLzmg3V73JoNLj79lltE4POb8tO/qdBERWitJ9Fvb0CtOXghz7/hqCv8
1lKhGkuvu1NZdRuZ751kgS37yEjt216K7jKtbGgU5P+LIrOwheS34Xhe2A0bkn5v/LYthgUtSiIp
cmO02rHlB0WCwICG4gmy/2g5kE/r716l5lYSj37Zf7mYtHZE5CmZkmPndiggFRuBjTz5TI8bigMC
+tWz6TgoLRFpp4jEOne6H7bsSQ1/3z4NJ90IpLAlEmRH9CDgIhpIaVnOgH4R24iJFt6bP+q2yZvN
SxYZZr3WWoDPemCy8IJzE8e6sVa9iMLu+cLsmZ/POS6Cf0P6pwxmi1+3IQthDcoZlcr0VjMOE5jH
T44Dsol4sCKNP9RurhBAHdUD5W3jN/9NKjxypcZgnBs5CrA5V27fMKDX0KIm/2CRn8jY031qcqgZ
DLnMnlR9hdvdl8UhPRgosMntsoF3XwmiZ6G49nr96kf6jMWEipPV3pUr/TKVIE+fSffnekO2M3sE
oMRzrZXGMZd07Gd0sAggRf7o7xcfsjtAuos9wHJLhGknaY45tXsF0fq44+HE4vV6ZtDW3PIRZ/KX
t+7pL5UH8dkTBw3BpqU8H1gtG3DBtfZqTvrJJCxlAUaPJJDNiwS4btGkT2crgiIoGM4wEgRoN+d6
1rA9dEU0gencxlYktKhM/Jzxml5LI19ATYryU4KHH1gU4qJDpAhobfcWS+p1jVYDzOUGWufO9x74
eeUaZBPC0qhexzo8RmC93rzjPuwTXrOF7RBXaeK5VxKDdgyBPtD4pw2Gyx8Or44mux/VJX0/uerq
zAn+iMc3/wgCLAjYWnbFKVb/ZgKknI5hoyGaQsCylIRtcD8jCCuM+fCaNX7FaFJdkq1lqz/suafA
cvnHUMRtO2WrasTxbDyxae/0SNqrAPUv5lUCqmxjk24isBUJPu3rr6xpdRNdgf6TDNxBljDtXuoa
/Peg2h6qVCE6lUxuLNUWKpyw4S63uDF4F2IqE1v8s2FTlozUczvYkBb+6kAMebNZF1XrjugSt7Se
TMA/3hpatAH0jrh3RwGfPTv4IKUXEqFDol5QWOElRX6KC+WGtGCWa4Yq+W28f8i4yYLTEjtoqlUg
fZ0wY6v6FKWpkOEs1KQRutfbEE3FmbdpMtgPz7y6sTifrkvHZAZxvUxcvLbXmNKWWv3z1I2RxS3y
UMGt13F811twR8c/stdYbiJJ3Ulk9lYrclGgsdUm6KSE7tBLLqS6dr6TXkOpRAqIYgaVznHM2/4K
DCGoNiLq2aVTS0TKhEiElzANaLqIWQa4GzkIQ95cb16C6BZLiw0pzFvKz+05BQfOfe5zaShJ/Yy0
EtwMbA3vV73xLyRacj3O7vHuzCA5MwN0cwozJszqKYhVeQp31rJ7UdUN/fDObsIJmnFBNvRCYMln
uMSw50jZ7A2MfMgOu5x4sv37DR+E0Fi9W0IY0azMMZJZrJkPq6FRTEeDKYX9atp1D5heVfjIFzt5
WuvoYOPLImLiodyxFxH3MOcDxlgSxTClnII20qhtQv2AvNBF89+Xi2U+Ydy61OThWfcoz/LN2Z7M
yZ7pfkQVBmb4e+r89wsHLO5STnIUFjNPif9BMkofIM1IL4mwmcd0pECbnmfIBjA+4hRsKfaHqrnT
DNTq0z0zhctB/uoND8EX3dULgTuUpDo29292MisHOUL7dsyW1ZY2x9WtUk9NAk63s1C5MsCcqqsD
u3ZBvI0r6qPKFFkPGL3STBcrcpb9K0ltrYfk4pIfn60A1UF30xyNDuUUnrMNsMQOvabx8T9k37zX
oTQz7RYvQymYS4A6AkyYCK6lT5g80t/yiU+jCXxgywM1HRViEDhvVtNYbUKLNO7PTazBSKwFL61n
xFHoaWkiBqsztV9JRRGeqy/GWokuZFYEBHz8wcyjGUGAMVH0k7H3dsxjqEiho9SoOoBkwrUrx+Dl
mI1uDQGM3iigk8Rsmw82qntpyGMe4NZf02Ah+aSD3+73vhZ+T9LZqDMVhfNJ/NG/H9618F9eZ/66
dzBM4hxrAQSZd+uSWipOEevRZaC0EwA9hWgpaMtOhhC5japTq/ilMB1QB0bI69UCL5ZRvdhMQ7XZ
JtWPqlovub2MADru/aDhS9trupZT/ZPdpw/fv0URiM/lxedrenXPCd5aaVYWxwNkt5Vc4BuHThrx
DH4yP89Vn8fnoIPa/fxLu6JQarcHGFDBjiNMlpD4B23KfoUFRRgbiM8SkjGHtaDRAwdnsvMO4lWI
bETcIZ1y2WmGmjAxoRkITFC/HNgD+OYUKD3dfOJGHK50bydvv/k+cWBRNzinvfwpSRzziLhz3c/P
89DwfD0EvnJHRuyf1chz1Wx7Tce463SZ/B6QXvzz1Bi/krcRf4xFbV58KMnhVEAbkh4RE2bQIGJX
o/A+uGZA0vMZWbcwpYWwxcswYtgFSIYZNOW/+afxISMjRyEa5gq5laq/UWiNx2dZx+D4eRNhvH9K
waM4k+Ge0wYZ8jyTbzKU1QpMcdL325Xi2OGlfnZ6c0Iv3SdJgbYluk6eiq5gHipxDP8zrGW4JDoW
WMdUwsAk6zHvBd7AKURADJ/fg11mguu9BJdZpsJsJql1FUB9m/eCJIFLrBCSiEZLNWf1/JyrWa3u
lpWa1ledEAuOMGvnwMCadU4342ziHcesv6Z3qhKbnfVAnhK0LW428C9bwj+ywBLaJSR8nFKU/IHs
q4rTolFMKLs8J69zMJYsAk7MEZYZ9lEhvj432w+lSlcoZrNsjzk0RsvglQx1ITbEENHb4ZuXz9z3
ReR5lprhjPqVpfu09TuB3L0SMSNVjn23iTxw7Htwfl4TQzukHYtXhcvvAS8MiibII7TsP9+IjSQg
5k4iQgQBfAYiul5YI5eIgdJDY1k/Rvg4PMc4JmtqjsLIWlFxrwZkxKAfVH6u4FbkfsnNYnO+bzTX
Wli42bY8AQ9QcWW8UeyJ+ps9FFim1+s6/UIqjVPAexvW5z3wLrAzjhY2rwhQtTQyedJ9iZVzWf+v
XBWgOWBJhyc20btNbta+3UKvyM7e0KwIe5dR7aPk801mAXOuLKdSrD+sQ36aAffES6YzXerDpTaQ
9atgVgC5uJy9on8JGiKC7xYBAauBIKTk+J9Z3VE9QoK0kO/0CP+BZ4d0HqmSKLwVAcQG8OBed3Qx
x5MnRNCQtkmF467eogFOj3PYqWtCFQqj+ut9TkeaTGoDHFN/VnQGi/bz+FM6Uy8dBjTcAe9ryt1l
ZVAH1OmLBJ2+qefrEIEGIu3Z/JTXcPBex2MEjJ1gb9sw+4/bRQ4NZZ5X/zetFa9OS/+6M37srdbK
cE1B1XAKXgeLA60ijI4zRn1Zo/kClt4vhb4BhYpF8zycyjdJCkMDn1Z7FyWS23rgaz18U8QYLpL9
UTEnW270zod0F7hWNLk/d2iuQOPH6uf6s9LCmFiIitbPWbWJ8h04ti6PnbJxt8cpJMPHCEm6wreG
jKgFBjVwc11Wo2py51BDZMhD7vVhbJFA3TOLm9b1RPklsxrrauWOhWhDurFR/cxQ8LhHwtqrzGSV
y2xBPLly9uBPwXXvZKTdCtV9jAfEXEF6Ao6UJ0tudfjEFMpW4v1XIOtgTWIEOjqCHy1ffY0VJy7B
rNbxRpSelTe4PeRA63+oBIfvj4phsRvXWfRviw2RFggFn8z9Mmimkv/pSIwPs5lCTiuJxfb1udki
eAC7/hR2C3BWYQHTut9BA2H/pzCU7qHYgRp3mWzqZAd1N1ekwtUgBArUvQ2J5vwFFcVwm2KRN4e9
tTwRiZ4Kw0hbv6XL/c/UF5x5U5+lSbb9HqkXpGPrpStLEuk8NIvn+xeJvplC636omdK6DNqeY37I
rSLt7tIB8MlqCblYowh7dkSwkJy8wkSgHPJSDyYIG0YzWawNvHa8QtywigKMHETs3I90kjuhkutI
YkX39L1cXrru3u/DtMdYPTmgi5VPfio5X8joX8qSbTFzpkkw4Kz1gB1AYGlm06m8AdE9Wj4kooma
9eNiwXZNPJZQsbEQ4uLpJS+chwrcVkWIW9Kjs34rLwz0Tw7zGV0qiyduFFIx9mcRvxF6Dx0WfkvB
jvglrDPs9fCPPFl023qVTjk+odUOYhb1lr1WI/1xZN8Df+bwVLMMu+IwDi0GY97mwDLOzf1i8hDk
7V861TY2cjs2s1x1UrsbeP9S8XJqPyjPf/dTy4meYZEWcQzUUFNHhgzhvtxB9H0o/jmar3/wpVLJ
czXP8DbLG26Ohxh7dDZqOFW8nmHzHrWClWAW9pKFKahYeRPOLu7N2Ob9cod7T/YYaytzT5x6QzwQ
8Qfv1eeSehzmPMhEDF7KHvFtqjpkWgf7vP2OemyPqmk8D7NgGL13VIAselwjJi3Jm8qYke2B58/7
bUsPPAcHuNcVfFO5ZlON6EqaeCBfhUZFi9fE1+fMeHoYbeDpadhCZKi2NxMGwDc3XkSEVOlekAqN
lx1rEv7pCt4FGyYNylgvNs3W9EtpTnmaPcsXGwb8t45A2Z1a+AAXIPgwohaXLQr3VCffTTMfA4E9
b5DfwiEom2NuohThQCa2/RVmgqu9ONHL3fo+8BOmtic/zg0NCKIL4NE4I5W0vAwIYEhDdMPqIABO
MEepWEjnabb0OARx7W3d18epChzzWTq4zLcbTtr1VsXR1I3JyKz73Ow4dbL/CU5mdyCW5fx5U1FL
LX6Zy1zx3jPVanDZozt1IBuiecGbWGZjynK57m415nFgq71wp7idJLkwOT/XFw5xlDPgwk868myI
LQ908m5gDaIqIgFd1tqGpoxgQWZQ6fhOnZflURjh1vqc3QW2eGavzrVVPWb+uObfIivkiAIEhftL
024xzih9GmOyBk6lqG5avxt2vCYgsxwVvJ2mYTYWXg7O4Xiws8jcfyMCCtFTcMMsUeOe2nBwwsB2
ZKekg2JQLa3GxX0OHUVN6RxCUvYjOhuv65yYZ0faVhx6441fckeoiKJIQNpf1eRWBMuGGy33pPtF
nEfrosLW7LLdOmhxMQV1esfIqUmK6df9TsEzyqxqqEIyG/YL7NszXRV25KEN5l7m2cqf1nROmTAt
IIFGJPhQqfrWTCRJJQLOlNSzyEeMvqNeEZCq1O1BRi10Dh917Oey1AH6z6NxFviENSoaxLbbsf+q
KCLzSihdhcW4CIfATK5s+y18+hF1zmwwc2lLOhRvtvJWws1F+o74h6IVVGV8aRwn/kUEhtDdyz3h
F8aksoQX/tzcfsa6Ietzh/REV725xqCihcLk6bFiYgGcuAG9pRbmapbr6i1gCJUtSPoq+VTwF42N
zukzQQTYiLUamrxgwkGH8oI7iz+QV0fhEcRQ9oi0xdcrXENdYdV75cmp1roz0VT2UIj7IojkwxvT
tBRfxBTkAg/bbIX0U2Ez3s0eLftQtdlCjcwwVUHAt+HSt0ty8jKfxuJ3vHmLR1ZiG2Gy7U77klT9
2pnalm7eBGOKAa1Jm7YOFwRGne2cTk7XR4NswpzMVw9TbE4jAMfoXoC3yjKCoS7gIK9lMOhMH/kr
P8BxeKGFKGd03cPa1RWeZGRCStvN7F4QB2ZqBwSBbJ/PDZ6paGMG9WAzw7BAqYM0JeL9QnhzZI+l
ZqPzBrZyQDQbHzdrT0E9IgQXVK1R49MlqJ8v4zqPHWghr7oUpPTvrV87eo+d36PXtiNnWdkPq9w+
jQ/xtRa2UAx67Y6GMPDEKi7nyElHl2ZjR7kfq8mCF53NGiQVwkmGftZf7co8A2onEPGsuOCuFXqv
uLs0/EihNZaGR+PCH3ZMBO3UIgURuImuIcZbzV99xasaTi888Z1YDV2Wl9MB3lII6Tmrq+dxMbdQ
YvolAAA1MGBLaShFayGU5pUQ6SoHc7tKuhkS6ECYzgdXUkMCOGL3QeaXxTMQ2Y61+mGRJ+cB72C6
YZEcgLH1Ab1ayWm3Ghw7yXWMej/MJIA/iLNYmR7m3CtGd8hw4QqFIN4uXRyHelqSQZ571ThzUCOD
sdr8khz2YkzsvI9BbQz4/2cUeRnGo3Zp3YuhWiwqsZ9eW2hh1PVx4ZztW2I9j9LKC9MKwwhkxwuE
9R0tc8smVgxZvmRus2sbF68NvOfS4IGd8AM/Nwul2rGaInwFcRXxk3jgm29fFEZAr1909wtHMd72
d8p7NDkSZhyV0GZXIpnTN3reuzNyYfjAvV/cCpg74SysjQwcpTb8+1ze5USGvpIeAlSs87yrKYsc
ayNtdRyrMihLXRGdBfLBVnwpKe7D3dqXnpbzpGaus1CDVxh4VK34LL+lBwFf288MeSsRCXJ7j56h
qpAqjil1vz2xwndkxIcdUGKESGiiQhZc3q7cM+5N0Y6YrNhW6nv4O4Z0pMmGC+FfV9ekLVQVcKyA
G3umJVWcVzmm/kCLmAebImaOMZnyDAXlPtqbmXADofqoWVc7Njsmpe4kDi0TyGKkyRBX28OMAO8m
b4qv5tc5ckhYBM43Vt1WztmbNXAR+MvdRd00r5zd5IReQ4k65IGPgq014bh+tEcCvtjgcbOW8Td+
H0FaZMNxDSt10InGcuyeOC2HscxX0LTE0EwP6NUR5SShwRgu8vfkTHIF+qt9BDuBNxBsZR87/9S3
NrWbqfol/qAVvt0j1PAmX5NqWNDIPsFExEcMTUeM85NrU+J6VJaEz931cawT3e8aAqc1oLSFq8Wv
+0rcGVnOSWfGDQl1KU4m0YOumz2b5GYdedKnxQ0PRAjpipLHzTWgJemO0e0WBw/YboI4lo1k7Qa4
9Lwf6nTiKwOr00i5du/x63IzNWEYaXaGezu2AJ4tuWMnfp1D6Sdc9gMrnBsFzxyLt3mM3woeGYkn
sgBjr/PG5HFHQ0IxFK77HA9TfT0BYacY1JkoiqCEJB5qtqfPwI8NvN+o1bAE8mKZbHP7kcz7HSaY
NJMRO58FZe/IFybTj3eKsr3MhnsdwYHX0GHAuzwNqG38oA52R4pCKa3RHZfN3PIDMpVaXgXfdGcp
HnAfWRQ/CF2vOdTxnLMKuO0MY4fdqx7mo1LiYm4o50/8mM4n93uTrQyKi30VsyG6ctErTO+VPlBK
haHiZsh1PKyILLKwmluvbm7Sm3jdG/aXXJxBUd3ncIWU4KScPd6k8w+/8N1lScJ78GaFCpdpOxd/
Dc1LUwwxGCclN6EayC+kethbOF5bYNj2jJRDvnqW8sARLrZQAhOn6ej2M1WCcDthgum8HV6qEzMJ
Ev/DKbVnYZnRrTx1HMYmxTWIzUfics5Ma5+5Qyw3Od6C/AghVWzpChuG+kxkyclsycHYBNqjUPme
mHokAXmdYOSEvR4me7IqpCx1r+jpwaAIJVk+bI/M6Y0XJzcSChTwD1/R5zusi+vca7Pa1hcl0Upm
TKQMcs25CIgmr5OndXGbZ0OLtDWSUJy2fJPp1VxGBBXoo2dwTUNbgc2kNt+tkQ/u8x6MSQhE4uap
SmnMVbqPtXKQ0xCs1gW7a/wx2eTh9tp2cE1IL0r8bqhnBLyJzkTs5VWpQr4hk9HoVtQa9jXWBxSS
xzeFXl4hRVdzM0fr//S7wlZUTKLD5XNHgOCGlh1VyZELSpfh7GjDoqUCNwl757Nbbp/os2k97NGt
KIw12smCMuIi6fFGqJ/KJM/UFdaoShAyHj3Ra9TkbhSxgL9e/7w+SdhDQRavbQ+rPJ40tK3T1tZ5
iopCxSKDmRCKwJAQt890yLNPiyKf48kI983Mgkd/ppsiERWnamASD7YnH3phzWSRBmm08elFhE35
F7MJWBVjOWopjR2uunnWILigFe+F1G3N/KRmSFRxrPZBQARIqlzazFa4JaNnbMCLjiyBTvctSmfH
lBbWD0PBHkH3acipcZwpxee8gYSFptY8p1APK9MJNo4eMIuSd4J5btxRetTdrb5M3velrtyUzH9Y
CJ6w7CQPcZO8xC3wAo48Sjx3y1oQC3EkwzigeHecepGVRSQMUebY9de/MezBozYfpBUEkUTWBwAx
2QOUDVfECUy58ZLfnLwJ8YIdfkcnEoivu08iGtnkXHk0NVTW2PpQ3cNLYp2QI85T6Z9vI4MAA6ae
2Bj9EMCw3GccuneOjV1LJj83MyAFBi45cqCzvnG0VrOt0lugyclPxZ715nEISjaJoPHjfi3m5Fl0
nyZ8u/PTHvy8XWuaK6y+LEyq6B5HNwKV1y2gIDyCwds0YpQdQEL8bzoRsAaPPs+y43vJU1J4rU3q
QRhDgQPLcyy7f8uIFkCHS2n9M5BEkThOpHyusrY1yDHfjAE92S2P5knSgucwvX8LNFds2lgnucwW
a/YNHBWfwLEbJRgr7e1/wRoIjqHKgtEJ5K8Icjuy5Gs2wl5itEV048Q+qaW3Ma9jWa5XbU2M8A5U
6+lYcnhjNbun211OPLiKOMB3oPyofLtV/YaDLuyGK6a4bxhHcCcjWifw3M1v/ee4IynJ0L2LYr1r
xyYCtHwrAwiDmn4L5qZjXl2SNcMVn6d4+tX9v48yPX1+k56hdfArKt4FnstKvcnzy858dVezW9JC
Ut+e0VTrK9p8id4fXOSzkak2hqW1m+rJDKhk5dzsN4diu9xyXIhrH2jRxfMc901C2BFWPL5Zjv2H
nTiACRWH6eUCZMiQtsSsI3xuJtSUtqIFSr+QaiVP/yAEx3VpL7WLPMwaSClpxeJA2ea1bwy3m0CT
EKDx6ffppSyWbO09YqoNQ6bsHXcu2czoUJ47WlxN7OREUJzyhmadZTt+T3SgfiaKgWDnIalDscR/
Y6RE/PipmvK8RJEQLp02Blzf8PXRLYqT8ELMqzH47Dm6Sh5DRB4vOnlGIsxNLTIC1tfgt8uNMqQC
L9Mv3LpI+U/6/yuuR0Ev75V0BXDoX/lEMJrzIl5xcyQo1iBBGS+ha+8x/w1Kwp2ta2BErKonGOV+
9kxCcSeq6O+IdZVU700PyJ1PkinwQUmwws/naz8xl7di5xM7aa2xZCdFJKCkDvWy5AWDNwMv7FrW
PBW7ALM4Pd2ua73EYRr0qQIxtjI0EEsMhLeWnWjlDfNlw1izsfB7iCoIgcHyKbuNGJhEHnHkKUtR
sAHb5+YzMOM9PRKOQ24c6X+i9J51XbMEZGxHA+rqGdsIUbOEAvLaKAvvFtCBanGoz1W1CICiQEkC
O19HA09ibLwtQB/6EXCbvDfQW8w5XzdyCpiQkM3/FiMKMiQK1V3EWWu0L5P1MdBzFCJAH15R/isa
NGR+KOuzIL56cIncbbsMEzzHWAhYr3UyuIqhfBi9VeCJ7kPvaGY94kTVEvTQKBTR/AMoxpqxa8OD
41yH6KzYxKaqswhLABPhm7pxLk9rlfxVKIO2OsuakVdvBVP1vkCgv0gsHuEYUiwmCHu4H+HLO9P3
lrazaOi5t9D5DpFG3ZlRiYMxxb49EEq/hwhyEdjl2pa0Gpd7e0aTwcEOcsaN//IJK8ek5YgsZ1S7
dCM4XQ84IYa3VJtUX+7d4vRwkl5BNhi5GG16lkDpHIf9lfwDnXubAxez/m5St7ulSSBQzTRz9NJ8
ELp0XKlWUvmYb0Ody+m8Taoubl4fQeDffO/jNkdA6YIW6LQCOFu3IYL/9EqouuJUJXFv7xn0x959
GIrNcZiGtvNXQzWbTFw1JIN2KxrxfU0qQ0wt8S5gMfWB3Yq2u+vxxPmCrlg6dxdmK6QdKN6hEhde
rvPaQa0apWFXebkIzxcFo8yp+uP+iqUq4aKIzh4jfqmSgrVsOCxOWZz74oSLAJT4GwllgPxuqBke
N0uFNM0/Mjy3fLxFk6vEMa9rN6E3+5e/FeTwtfts89ngaocw2UNzK8NLrldeifl3WwlljG/S+bJw
2d7+/pahMcMsojWJujzyWWjohfLJWDYMZIU+geeiEdtVa0HcKI4t0PJPnAI999EmLJHkR6lGhaBv
ISzsrM7p/S8bYsModxq4m1u5XzMXQSnEhg5aKKXAZhec+kNeLWRuHlNR9pLw3mM3pAuQnaX4WAC1
BHaJfs5j6LCVpz/U0rqlayzLl3vH8xj+MuzwqHqxyIStScuA7usiL7ZYARA0an3CvZnTMigTqrCK
gjOHDeuSfpfvPghYE9IdvAQEuqhyO3hDWtHFSB0TFeFC+kUra0KmGIZQ+DFuM6G/+vFLyfLJGZj5
6LcWUCmvXqIlU9WZcQ4aA/pIMQ+jqxEzZPMSIMb+tW3pvgkBaIkPq2tAtaB2Q5llzNmdgOKZOw6E
VQZxr1ohOpZ1U75NW8RV9tWQjr7TOECCx3sQYU6Xs9UhVaNDwl8JDE7rEVTiVVzw3BTGYOj/UbOB
gOALy93gsdvCE8+f025t8qoUwkYXpTFb6ApiidHbf24nLmarCkcD5MrwYlhTjzU3kprwhC3lbi6M
Fw26X9adEQLmrdG68ZmiQQHvfjoojMgwn8151mwYZnYTjtRbjnpWjYPuti3swPuAEs+81ABSBq1G
zamtR4ATQQirSKbSnLS0jXyJu2HoCdTcRSpIQbIL/d5ynGvczaKQCkEULo6E0qwEG1jLnMxrlBDX
X0pc3QB0uy2F5iqgFErhg/BccuvX8Sv9NzulmvWP1zr0lPv1HUmtzoboEhBoLHzWqD95zNizGgRC
Ornb3FGyZnJyFASPoWlkrA0zfZF6ie+y7sQ+R4xvpTmyhuU+jt50eNCzqaa0BAVvFv6XNQcpCBBr
nQk2qdFxRe0lpHf2MBf2QQO9XuuNcCGART5UjESFu0YdvD2poqkooP5r5aDjXIafeCVg5xnnjqLy
BZCbVU3H+VnmZWvGOAYVM8dRzZ3IXzN+ONmLEVC8Y3CBPbQ5iQgJLACXLiz4N+ZJXL3ZMsV7PObP
aQp8tsqxVWkWp9vOxpiGtNQT3QbBmRoj1qf4uXT5EuYoimgQhExoRirs9WxqaG4d3AZPMYA71Zkt
9kVF5wCgs55x405fcbC3a4qnOJMQjuCBHDN4uuBHjW2b0kXcYH9qKU32Kb3tRuUWoEiNBV7vC1Eh
Zf8ByHb79DmNiygGkpHCfvq7H/nQJtgynM5XLFvNSJ2IH5v//TxIpMw2090l/z2148MTWuEBpURR
77wOY/u7hKAJ0uJ38TCqwy7f8auau12UyeL0p7PJGItwbRUw68PR3KWbx8B2RKLc5YUcildTUZa8
BHdH8VpDPN4H7zXEslRPsZyQsnI5tmAiCco+SIqtz8cUswPRbULCVUE9BzvezHc+eLatvj4M2TnG
nkJUWappfMCQURaWc+coRN2OuIzw2VKWASYW4AJNyO9z5zo7YwE0DPjJsSYO9Z0XZHf276M8BMpH
jd4Yvj3/kYbszGDfa/HV0aGwlPxcsJ4v4gE/esHsjruk3iMEYLdZrF8fLN1xzyh0qNjdACbbHdQ2
YB8QCY+OH3e/yPnaua/Wl+TDmMSNvPvdbkn2wcLZKXlASF8Rmr+SKrWGmrfBAiFQVcqxVp7ops9l
rbnGUAf/U7n8p4nhFaNz9T8Wb0P/Ljy+84PAlfxYvd07Hs9zvu2m/s01Z4kH+JEz8/8b4SDhuSJ1
k2eKhB7M5oa1eD89JInTZUiEw7tLj9v/WOPMTy7qq8/LKUk+WqGFb0S7Gy9h4owAz09yoxCLbun+
2ML6j2jTamGAEojY0+BaWrbKILyxKLSA4iV3K/yK1sG1MAdEOWc9YU/1i7i76VWovuVjzAyGMKx2
YZs/mQ2lvyeKvgTG2nvLuB6Eb9GSjymJk90EYCjo9HDa/Mq9lpC2cKeH1DMHO53Aw9uPlkSQNJTo
zAeP5afzmNsvFF9AVuyzs93xP4nIiGx+eO2HY4B87eQcki6+WccyU4tWS4kIo722503isKUPHbtp
RXiJL15jZJ0NQ8nqcH+OyzvXfaRY2CHCXbaDQjoWukuolfEvgfwAViOBGg6V0/ucpubJyGVJzmuG
YMQrEyKiaWRTwAJL6wjtIFCbVmUnaGhXZfFzLngtv2GE19mI263VrBUp8QgxmGLgBjwnDahSwlNM
tiGjJK8k1kl3A2BiNc9WL06NjSV6b3t0/YaBJlN+nhmRcg9p+/tnZZoK2E+oVIQs2Qh15SrNk5Km
h/0yTd/jr7Q87IJRk06uzU0/NPWDOK2ew00Bavz7h3jK61UA2xhXuH4p0GVBFzAT6G8OIK3NGEku
y5SAfTU51g38uXC2qVK+2qmfggQnyxbnPECuZ9bgSz3GKpN14/K5X5sFKdx49n7rdNEodfH8MfdC
UAw7DGtWprB7lDZmPcjfV9b0LA5SEsAkewLkZEOlv4FwbPcQNLld/7Mp50mL3Txc9d8hwIH2B6FF
HY/xsn6m4c/gY2g/OYZV6uiFXuOCkEqYNX+qItmsoasSzzMnRrlQb2L5mi3ZrnRU+mKSxhQ4sWGB
c/mAxfFh5HSauHAIG/wxd+kPfA+O/UWmR3pAJUmhRlXy3trtxrabUk5L02s3Qc1TqhNWDULFDaCS
ePnoHmTolLae7gD1hs1ouAJ/yl0msngDnUF9ogTzgjZg8VJaE9oFRivRBmVilxRIZHjk3Z/iorAl
FLlZ+yUHMgy5a2Z1DUBAf+9BsZtdqsctaOXR3Kab1pb0s1zCUIwE1lboPERU8JSasoTvqyPLI53t
u6Nk4pEV0DMGKVdc60p7SbneaF3QoahrjCZh4xlY0ofZzQTC8AcSu0K6Yhlkf72NuweFJqlmP4kr
LTxnkkz6ZDxJibsurEYy9KiuUsDHaFH5wbmf+SJTCHdc1XaTqe+aQ24snxX5bSmH4XjDML37Pxj8
dsnwvWi+J3NQ5n9nWK/goSulOtXqtSQlQgG1xPuixPKLToTWhpnGzdmRN/aKEuj1BoWar4lYgda3
1mAeg0AP1r/RIXgWNf/fa81LBQeD010877Az2OSwsPLRO7sg02Fa0djWU7EHvupRtXGCccA/vsnR
ox5v+Zmn3YYFwVWDySWpBajXgmbzX4zBJwmsuILRRmpZPhUMLsfEtvnjdAIgOAgwot0lwQMoqQuY
9gIncyBnjUPkqWfTyGje3dpXb65VCq8lP0L9RsePSmN0CwfYwzgK4ydEmJeuvJFDDarS4o6Hgqzr
OUs5APcxD5sedaXUFnS8Zsq44ZDkru/nSAPSGFQw/fIey/kWGavtCFQ2YI1Tf+L40mBgPujilizW
41iQ12wOYRjFwS+/T3C/YPjuuhmOh2/4iilU0VGRZZsxvmtjdOHVKxnmJkNOMov1A8Rj+ZYJ6kQH
gYVCBEGuH4znjhSvn7xIGWQO45wROLrXiIYWpFfecwa2vGo5mqPb5iztya4R7IUVikO7KWzto5JO
/oLGEOOX+MrGvN2qk6UWps2T7JETo5tNJX8fSE3RU9jQydtHgOPFPEYVhtkzHcQzIdvnKJ+a1hg9
BUTpslYL8peAyFjqZepFVH6S9IKONepI+oqEydqa3HP29oFpH0rZpYcMgglr5UD09d+9QLRhM4si
3rlkDUlhhBEqyCWHLlZIAXrKtGpXkR+ai0Kp+++FE0yCHmb2fx4Xq/mWM+y2rtKSeRHvLYIOMc0k
uPY7A2sxqke6y+5OmPoaXDLGGN9eiG/7+WJUYue7CExk+zkK9MkFjDxEUYFVk0EWcyFMJr+LXNtn
uWxtk8lcjuFLO0IkSMoWNHUG5Edj/DOPvsQMQdYCSFQHBonFSrEuPShi6/ZM6J5CuQKXmFUWeNBl
4z+HAlep53H5HidE3Zk8RnrNz1mCF8htSl/ckgNA8O7Ui73EEQQNHaU7ZMSkVV8YHSxcN1j9XqTD
XW8jP79AlVahHw6hmlTKRKG+X+/S2fn54gBid1lg4BrrnR8FeghRrcKGlCDRI6igKHRcD7GF3PlJ
yDNzAj3m4KxYvOQb4nbueoJFMddbB/Y4AMDAhlB6bUo3juWUgOhfE5MMH7fLdbIjLx6A6ZvYYRiC
+v2QY7BeVteZ7oW/qFQd0Mnu033YPO1ueFCJSh/qSFLwwxUKy1ne39LTjParZmzR7dae+zInvGHP
IDe5LAjGJEFOv7B7WnP40lcZgl9TRezqkjo/EJePWmQ2SsgG3Kq1v6hwGng1/WfHZ6VwRzR6HdH2
JeAFGCpcw+/045q6IUZXQLOb44JMRXwhE7Q+wYMk5Sq1wZR72a1aLE1+3ymOcYthUwjyUIyR/z22
oWjIBLha0kAhdUOWT067zQR67+eXOg8Xhdgyh5/s0sOSjrcEsKq1N4ykaT/CYgGM2apZ2kcpobQi
7kSdDZd/QTXSVRTjXiEG7rCaOX15qfS13D9MAZbwi+lKmouKkoMBGu6HNqmlv8ICVJ8k51aKugCi
bE5vO2VVo8KUacHuptneCBs5DeFmxTbDDc005z26MFdsXD7an1LomRpyURF8Tqj640d7cOtWYP6u
pcBBz3jBWw+BN/GKKxYOo7lw0CpEpiIXogix82sb8Tq/04I1JJYNoEpurJb48e3fSDK+V7LWhUMI
TmhAjAX8CFWRHgkMeuLPRXfSsKUEy2GdZsiLJsD/01xTfP8ajECGV32oMUNiTvYVMHmRBYUNhC/B
tJ79enCWrzzwp49WCAujNz5bXCZ/Sb3C9DTBdM5sShYf+VBJsn0hhXqaa45sV4LxZc/r3ymojrOj
eFOe3IKgZklHsr/qfPz3JZ1oEjOkuyDZrsD2EdqS3vOXQAqgXZ4Sw08mg2owfeBSvjM7uNIBFaz5
VyMLIXhwAwF1b+a4hHzATx9Ia3Zu900wHFwBKuWVIDah/fg92pkjtM+yF3HCxolkvkgf023bvfMC
u1ZOkzL7HtR50aeeAf25iSUkg/rkfwpR5AItK/S3iPwaSJ6afC8O03JKusnI9RyruK3BOV2037fm
oUHoQ2K/UuPBKKPh46a00Qtu8Nfq0o157YMo29iEn0x+PempH/qbBAjKoNuEvm/sOSQrppPij+aE
cBP5/DatUJhjt5L41w+bBrsDKcgis0rZaqbX8eiIYbeyMb7Npjedy/HpiYNyhYzicpdWK7pgJF9w
fpX2lCJ7UgomLM6k1EGzSqZaqW3Th0Vmt35gsMKv54OvcN7pUrn29HkE1fqG0FclmxwtruTPgb7B
ywdCJi1iAneLx2JXgwww3WCSTGOCfsSgMwAwNZizwQu9RKl3oIcxDaOHYqeZxApJTtq9aBwgUUAB
0egCOWACjtQWc5L0uq+ZGrlnPatXcrUkH5c3kr2mZU+poWkLLPyBsBwsAQcGxTPV+nXq4uDIhYn2
ob73CXSNJfl/FfmM5s6hAEZuSCR+umrY1hV9tNttM4VT/FMkHE7LWaFGuRB9JluJ7jXGyJsjFjHX
wrz7Ii0/H1qtAnTveieRXNkE9QWA9XzFpDCCdtyZ3hgPr0sxt9L1UgoLRK9UKn6+E3M9AERQwAk1
2cfNZielV5DrJbFhr6QNAofGt7jcgsxdp7MOv9LBoE6FlTueM7M+coyInjBQgXrc+29Xl+SR6swe
8sIrdqXbfKBSbv/YK2IzvPXE7QsewLsu6y18qCGZtjzYXGCDz7SV4e41PlkXB1hS1mLGvJrfKe/K
qkLY8y81IjqdvPs9erCpS8FU1Yd6JVPz443Rz0f/xtdTN4eTD8/XZkkPOJ+FgFj4D4yjKyM62cUA
JbbB0ZkXeaD8rp9qlDIc15i83XA6C27PY15XnvGhdjQJ64KOhWgTId3M6OST9dFOyL6wxCJBjQJg
rjGAFCFL352p6pvM4H6NxKJEY3K/bVuf8VsOjqD+dDl7tLw8xPmSqX7Agj6cRtR8Fr/XXvOXehlL
C4KqjZ5wmKuUTk8C7HiwBCWsuvWRI+o6S3+3VHTHsVyn5K31yAF80NS0Ipqf5aWD3xTXrf3wNDFl
iC1mdMPAI9ego2ie6ez2Ne568RLtybM3tIQAZkJQ61980LnEpWji9fW/Zm4MQafVDreR9Dzx2Kuy
l6pPAGmS/i+bI8pbF+PUWKIsc71xo37tWdTpSe8dz+FhtG0/S+PWn42EfpkocbBkQbIci5Vg3592
AAvpkVlVdr+AVBa/pBbArxT4X2X4moO3kUrFLrCcZkz3AIAEYNwNNitsdPSlgiPSRGKMdXxO6Gkx
iRVjUlAESKwNI/6lVJ5pvn/dGJRW55B16M8sPOXVF/jak37Pe4MzUZ5kcwrcfn3Ay8aZmTgxdNAx
7b377f31/tzlxfecEUt7tBhcoOiLzsOkXWN43YO2tgkWfa7U45IBykB9qSWJWKM3QJwttgFVPNNr
qxNIcnsM8whfOe3WhZw0Z3c5WAwPg6q0k5WobQ6fiVjxwabyXkkNmsI5/2TLLrr2HY5l5/qKLIH2
H6OzqNm5jO/C2RgnmIZI1Mi+KYpcJQldVLkX/HXDb19+5Iupi+qJCeGyj72Q+k/qIYVH87DpJL7D
SsTcjJXZ3AHo+6+LmnvkTe3tMDbgorIXnBCwWbpl9G2+5F4r2Bdr73zocfF1+uiXguXMxn9yAJFI
jdvXHlVJraF7wGUvm0wwOXy46NmWpL1O7FiC8+wYmN74V733nBqwLHTUzkMBmcozjNS/mQyMAqAG
N9krtQrOfqXto8YogiZxrItlV6r0Qqx2tH7Um8+Q7LVTAO70oCYvgFCPNzHK1OuC5YdYNLsLOSDA
JXKFl1SA+ysz0SZ1rzVyetmEfqy38Eke4vXmU3wuYKyI3TkW7WMW5b3wmPF85QZ3085f6IdLUuoL
Ycbd9KiJSB54PGKRgJj4WwevsPiUofjH4fLCTdKHefwXpKMMHjNMssJqXcJRkZdsuCvIjJG53JFc
CYVIdPscdZ8QblUvHdx36lg7CJK87sq4aZw0aEsHOmSNsI3kzxJpsqGcGEgRF6CEpasgOm0eavFZ
/3DBQlNsIXVgTsdsNWAWyaqUf3i30pfZHwB38tvOCT7n9jRXN1naizmwR5HbXdzA4f1b8Q9JWbk7
6CwFjg35FTeJmaDz5ec6/0iRcVWJBH11y7FNsXdlni21yV640/mpVsI02hoEx2ROTtjrZsMopjZ+
H4BZEzwIkValtNpxi6bzrW+mUxUWClsM6hsMTMy/e2pDeMGnEdNIrR9FA0NaBBi9MWF3WtTBqa69
ikPGKjulrR+Xr0MbAjN6mlb7ovH/MoUUShBzryYhJdcrXtWRcTZkDJjvlECpngOiGA08yyiOH6FV
EqJm20LzQxVZA47ldPK2/F97SGpxvgecQBTvqionPADbJrmVCkrVkudXxFiZQLezmnMPcsbw+HYJ
ac0dZctnBEncp1qQG0uyMAP4d7HjdZT0syCwPMJlKMtHobPUFJ7tBmeO72azL6WBht2WCFgak+fk
bZrrO1q94gEncdNo7URDL3b24usy2FGFlpVO4Xyg2oTVlpsZ3NOC7xSIYrezfs9K6Y8GqyN22lOA
tTBqswVbXITqd3hpBHwikGBIRT3+23/AunuOVYP0pQyV4bmNhWS72yna2eI9SnNba4LUHmJGEo7U
5LxD4Tll3BvFnN0sYx8nNqT7YtAKOTLfBJ+0P+/1DC9laeHO6KgTU3K9byVkVEbTnVGyViod5gAR
Wsiv7LFUu7eJTjXF86qTFo/RI4g2xlw93I93NGo8O6b39jv+KTPLOPozrYtYglC7oKYSup5cCyCz
gKnn67AxOoGuEomn3GXBjAOxzslRokVA7nTlUFF/RpGJv7I3zEUIx3mUBmcQhi7tJbhAwiLhp1Os
xqt+t9VtILUhqspH/GgOFMqrPdFQKBknUGZQTxpRLkznrnTkNb5GE30KGnAj59Zls2EQk66eWQZf
LeKaH+u1i+kfg0tW9z1FQG04A7pnCZMSaNjsOAACmZQ01voEtlw5AhYq4scuZ6AzN7YVSHbOG3Su
efhfXm8piZCZHS9p0FZGYf3U6anfH5ZGqlMRKzJPs2CixqPLOEfq7Z3mHPr7w62DrvEkZUdSk/bJ
mhNiurqlycLpPWbZxp2CQDzFP8pXKeZJD/AfCQ3V6rx0648pp0N4Rrxd40o2qSNqTKPYUFcBT39d
ERECBXjJKdj8rPRAMX93yJSSLUk2vPOlPG2wdZ0Yx2QX/T4A77CwHVf05PjFgS+VnvXreCrrOa5d
YaROgQfzLoH3G4JGEqlSxdgupUtZDRhD8fBZRpdJlarKgIvuG3KkxuxgWRJ+nQW+4GuINRP71yVN
eKFfYYZtgEsCSyqap4mvl7cyPPndQz+sGHh2uuLL/ekIZX5J7/E974KX89ZKNVhQybvhJDW7npsf
vM3SX9Qw9PW0B3/+5hyLhXve8FrKO/2nAahQ1yTPoPea7qSjcU/aM8rX0yn7uCOQnnAWDFLXwl21
z+CozB5AAddGQIHashiwuMS1mnuNRWrOzC6RE2OUbmQc3cxx7PYuv+ui8M/MfdgOEPVrLaMgbpJ8
XoNugaC4IJ6bfOZWYdJ8kpyVbtzhD549ICLrKc8Ursy2fEX5p67+4pA64uijSbE4ZqZ24d6mugWH
r3W63pqoi8wSz6GLcK+xzT7QLSnka4k+lleWhLirmdSZcynM+dFFUrnjtNjYT81BcemPX7LXWH5e
YK1bsZRkjn7OwZhvJE8X6bzttHdRgUiLaHr0ICwLxUiLksvNnTARhik5d4CSRA4HJwEEwcM94rQj
hm11XblAo7TVcBbyYiQc3QCMoNi4VIZWywxQOyu/KWXnMMdSLCNSWTG+a1q2pTT5cGANFVZ2d2UA
iQuW8d7YQTWDn6+7AZ8XUI0la3cRXrgwxgsc2Y1lQo1qhod/nP00xNAp1aaA1T5h9t5XhSR8uSEU
N+ielvRaoNnwo6/3250KcklZIeurG/0nODiS+M0+NGIWVEfzQH8G1Pm8YE/XPmPO+LZbxIGhDayf
DFkG24lJK++yNLlFP2yUymEFMG1QZhhs/1YHFN3kG6u5Q7W0vhmcvlNtKysI+uMAbXyAxIMMi5r9
81tEfMcxEkso43IG20ZrnvnQUzdK9TJZ0BfoDOt1G6N5qHKLzp01aKWGJbaZRq3hUmsc6337gHQp
zYPiVvKB4mj6D8Qhw9rqaZPGo3PM5pAV3MDFKlOzwyOUBWxbLqBjxOlfT6H2172SKSoUfk8NX0RL
9Q23L5XR6ENS2XnIS1Mf5+Znal2s6BvcNVEtYwtpEYmee4Cl7waWF15gUENgONVd7zxS4fuc1MSC
/Svuvo5pI+2gowWRNvnjI+J9E81qmcwjRMtc79qhTB4uZQVvhMXFIda3pFqkc9Al/PMzwxlkZkyo
Rpi1I4+lrbI5GRqVeClf696VF59ro60WVNjzqFSvJOX623UpUBwojJa+YcaWq0XEo6IE6AtAgfhF
dMKL9o5PUjEEMKzXYeZqTuVrg5Wn6dC/FsuHPU6vbIxkAb+SUpGjwfRBM61mCrEjFom5EXVXwmFh
QlC0zBu7bvwgD05CJwrW1QnnUHoPqYHKXDeGg/SZ3+D092Xr2wHBBL0w4Y2GHq9EhvYJToM/zhFm
st2y/qRDw5MvVsSEHT/nUTEQCKZRFxHHaAgbKR640tPJZGwOxi3fI+/kODlIsmfXSHPxyKiSWRuQ
mO1Folaaf3kXq2lv/yot4HW84OsaEAY6V2xf2cDJrsEuFmnsMCygQ1qhlEg7jc6peSDRNOoOX8Fi
TuTlKjKtw9NUOdqd5XNplQ7SikWWnc3DwDQd3w14V6n4ADdtDCCUmdM2+HHVUbabeJy03zHOake6
1hFjXVdccWs3NDRca8qVSZE1D7N7JoTwUUxYwM3A4JlSHxHe44362EjMzXh2XEjUY7gApDNYaxMY
neZa8CIXjNlt8C3OB8QXUlS8/10xH48o1/FpHfwBRwZURL5+NegWKXRtLQyxj2TYtIVTFOsYlNV8
9FJyuPpfF+49H21QCbyCv8mgc/H7z5iw/9Pjm6wwe4Lkemf9H5Pj2TXmebQ6uf9t8RgsPL71Xva6
fbiKpTeLMypgQhtvEeZmUFPTegeAOl5OIS72gMf925jWd0Ofaq761QyWZtR828gpTaOyxbYpMpoD
kwBOAkacs3ccmQqNRr4zxyOe7xOPulM0ekt5MGpnx3HYpilUBTNZOfx2fvRkG0Mm2crjBYi9yT6o
b/Gwtuv3by0WsTAm1MZNxMdeqm9aByCXbp8CSTX1BJl/E/n7bkBPeREdF0UuaXayf6TXKG1cci+q
YQSNFOwosnd4N2kAcr3/nuzbqYuWEcgJcBldXYI3xXoU/eo4JRmdBH26MxiTFNCowb8fb8suN/Wj
e/B13p2MlMF1V7nqbwqYgJ3feZDSDnsC72fvsbm88htnKTKE64B5JmafGmoiPtVwxEFZpYDLaD4d
acBgLpSjCLGkl6eJrH8tW37lNtCBDZaEcpWPFBJKCjOWO5AXvLt5cTcE7RVtqnF3aKKUS/uNCH9M
coL74sh4pzUe/1p/jyME+XEtFOCKAdKhxj3A+N6neEsMOwvdq+qjweUnArCqdfhOPZrSALnJauVl
vyEz9Eeuxd/gRVA1+VJPCAPj5F8DKY1PttGpZehYdazB/0ElLYum3S8VqRojt4t+nuVDe84OuOpi
CFerKXFejxpdzTkOgGVVYiOH9mgpDGoLfgZFh2lpcWoyIuG450X3dXeeMmBekZ34anRijAmYNnRY
4+Ng+eRv7IZNs5SMgW2IiTPii/NG04qUrr9d27gkz1UFx+ax5myeDpOENZcsfLjlkLEiWMmVu1Rl
ZXqJaA/97zrdfVNlywVGxShbtRghvd3LISPn9IdOekZdjKi2rEAbbG0bKNoQpArXGqIUc24dNQbI
P5cqKslFsm1Hf/dtACW18buN+kEPc52ZpMxCWq/tqxwe1BG/9cJRYrob3qu/WVRCkPNhfAAGF3C0
ck4xaZVes8CJT+orhKZBWDnr4vxSDnZ8NzJVtWH5m30W9JWTENJLQ+/QCai8T8APQcmmIB+RcAt+
jyO3NEz8il/+w+A5LxQw4jeoB2NI+jIeJAjwR8llcELECDUSqTEUpouba6kQ0dmyeBrlQhYt+vO3
nTVnvxtf1S2gpVIpRYTQ91E0yK13atgEXyI6MCBO+M5F3FVirZ4sMVVVplBBauj/8HmQe4HfH8ah
u/cJKoct3+q3hPavkM0V5p/ZMwqAYGoLI71p1xVefRNybeTH8/Oal/Z6Pu8H0KnUzpbuo4FZLH/l
qaB4lUZw09EomnoovXCNMPyleSGC3eOQ+oEFKwmQkfrk9baWk31GFV8R1sVyvhU6HBEiRhKTfpUe
evQIJpviNcagtsJw1uSiFkkwVUaCSwBS7LUJxMtigwHrbf1sEBoYm3a4ss0sFfYlH9Q1kqq5ZjHA
mUon53THsT9dB5N2esSAQtOMD65IvxHXA4Ppqf2tDRVLlZgSIVI8lLh8/sGc/sWnYtIMxydfE/2S
WLMp8Eq36OIv2Q9P0ds3OEFI5slUT5KKaK5aWyJkNUn7dLJCY0juHiRE0Gwiv1cklD/dRRb7W2we
sCc0+ur1ykwAQHGN19JclJiZdBcSW0ECcNLnQyG96mNB2DXdtI6RuZBYbL5dhURETrA62DU7BVgY
wMfqO9V0sVMXArciqT3un0x5qiMQaNZgFvHqESsnSUnqjuX17hn7kofk7bmLurJIA7MddRYgugjD
BDOFJ7Ei5hkD2z2E+O2vV3Hl7bjT2FsrjEcAjLbZw2gpJXVvw1O9NKw9DJYGykqNMWiiNAfKTaXv
OCPt158DO7yW9GxG12IAKEogmquLa1+hDkDrFi3O9VwoCV4KY7s9UEECdX4FYpP6rUR05WfnruW7
xxIrFxT3NSO9nmnRnKQq4r1OlW9vTOnRGPctFvtTnHfUjFEesBEeZ6XapwQoelpneZFYPpMcs6+a
jnaE4RblFY6K5Uk4cYOE+327cREOLynqipNW5GDsEeUkvQWjrGYjJyjdVyc8p2+ksYRjc2LT/7cc
oLojlR63mwyyCWYk4kW1KcjeOYKbEYLDOOgrsQ0em4uukRcY2XDdOyu4lUPSgOLno0jhszaGJJ1D
KXYULgdxuICD71sQkb2nmzobhvIU6q3bxJ4/Nm4DVIuFgLU3mOYzZ+EYcf7GiRTAIQodMd7v4J9U
k6fKp6XU46DorFfgKWSd+HPDx2tAS6frdx4LJdFa1wn86jmHZedTpYFaX0W+jYaFtYDAcWCOk2MQ
ht+e4xMe4F6XaRMiVD6RtmHZ8wZ5tAkbTr8jpGjc6TlYcxmNtYDVVsgRhvSNtm+A4WI8ax4gAebw
gGJkRvz4zTtH3uWA07ujs4bKS0oUt9bH/6MUvba4jkfvzur7zRClTXcMoaJ0zlVw5vTLHUkV1bO1
Q3/6AjULBn3YzYkq34/M1Gax+BVnofdP5+yltf3HPfi3QnMIxRa1ZtD27oofpl7uyxEUFD0BuurR
WKVeLaaWB4PUgeGvNivxXJ3ofKFUp+0ufQmdMsObd7yQufSdvco2w+MHKy2Bp0qLCbs9Q2flv+Bw
OgI+eHmUGt2hiLuVB9rBEDF+TJjhxD2oKs3OtFeXVzYtXgCsljd8zAavJqWPa1W2RhypsNTJ69bR
ahY48Cz9nN03zxxK+UerEQDRbOU2xTkdAGs8YB9wvDCqqD9eDOe2bJM/35EmFI7716jY7saftOaf
IUuXwM2O6iqKKKfGFUzWg62h1fQG3g0s6jiuqGMSQiMXGxm1UogaC8d8rX1KmDfNqYiDzNXuawqT
V+1AJei17myJ9BcdtQYdTi4c0dxRMHVtMYEPWFh9X/it9DRorobcjYxx/Bwgh2N32RSaavJ58nro
lhoNLHadcBf/PMkaECjvzaU+oPbw3yDcS52QK2vCZ+5Nwab5Uf36Xm4BBiDhkGPQlSmKYiVBY9HK
AE6zrTLDHnLbf5sBfhGiu03bhf1SJESMZOgWjy8e8+q0GrCcFjZJqxqfE9AMBQzx53uRizmY/z+I
mG9sq1Bdnt7owG7umFHH+9Umue/kc6YaIyZ79h+8t72ngCqK/cQqydBpRbyQ4yL5R5H1bkuyRdyK
UC6NwsMTTP4WIo/6hY8GYaA6geFfDHsqZbjqqyN75tOhAxlYeW4Ac1b6c3YUcfKX4aglKJH912PK
nhus2OjIs/Vr4FU+RUUesiQarA7xR/A195D1uVEZO9/GIyo6ym1j7FTybAp+/DxuqT/rdX9q+O/b
CvtT3l/3tnAkT0DtGziT5tHCZan7rlgC1XYTckaYPu2DuF/nc0OQzFn83kykjO6FYD1HzuenAu52
SIytPjs7zwRRdA8hn3C/AZubVy5Y+Lu6WWSZWXEAX9fwEivV+gP9RjHG0/gYH7X8835WwFziV4uv
6gATJxFif0ccpwiv8DxcDtP8W3ye13cuovZT6e2yjaN1HI2EBFk8aDUhA/izZ94J4/JRXiXxR/6/
hjwpXIzxF4s5giVpq0F3/XMk37EksMaojn5TnRCvk7hMZl6+26f8OwhHhnwrmjHixMlPgTjiRrXr
O8OreezkeaDP3qAMqKPWadmK84p1TPQTG6S67OxscYm+VBpdx/WAA5xPReqSBLT5AJAFlQf2mqJN
DU5bhcICb7VTNdTWe8pUaS3eYim+u8cAAAEDjqJh55eA0+xfF9mdiKEwPkkS7ptTxba27S9FUEXd
I1qBL2CVHkdrAkpjAhSzjRd44410hQMdmvF7YRpTsTh112daxd4i+wkGegaVMJYqguWEOgcd1FwD
UEKQtzU+AxV0onRmrkikOEFhVpf0j6nfsQksC0CWBd0Jw4hqSuJqxP/pG7XUDz0oVoKXLtbc0+Gw
/RSqxZfdaw674O+pkjNAwLF7MWl22R4t4TyiiEa6R0HWbgcxwM0bbFc/uY/Yo4mX6iR6wj5yV3kX
FzxIbrbnWax2UZj4oD4jjRRAzqkFyjwp/zXsl+6gpTPMFF+HjrzBg8VNu/CcZWyX/QolcJewPo8j
/p+TLN7zKFTskMXDOTMQabrk70NQ9XJJn6si5tKA974FFUFfnXxCPy02LAE5IvIoY0qlNS9li5qY
a6ExXQqfWxCfvaILNsDW8Ta8qo1Qq8k++R6aUL1GQnkPe/jTrCeDSLV/cskm5N1oZ/fuR7oqNdxP
w93Vjta3hG3Wf0QGPdiALQXnNjFvtUpJED7KKCmQl0tdd/cXSNjwVntJ+XBxOPKy9LeaF307fMD5
n8uL17NyepSkCP6E6ra2l3SmS0DaASiyl0IPcbKHYATNyJPcx2ns170jcxi76hC6B4nWjOApNr85
IBMG9+ssJoVgM6mdDxK/gtwWi8v05gTyGtaVwx9pX+ghkKstS/IAMeRnmWxPHYgLO9NosOKPayda
P0VcS3tOdAc43ZYuY7PxlKYoaZtuHWOs4G84VhR/Uf4syQ22y5Mgdo87kQlLMug6PQa0VffDqcgy
CRKaz23wAnWfjaYEwZRvy86v688sbwQi8xWeg5GgxH9Eh7K5TEMTKX1FQkAq2+ctl+Lg8M56YVoI
7Ns6iJQ4B/8/kw2JhCSQDOc2uF9bcMV9Y4Craa45iEoLn3cAecXRjqmYSgeKAL+SIJ028wbC+j78
a/C4KrDtHXHIbGc8jl/6A+iaJVGdqQ8KWnNkzi7xqECoAgPmsQuqdLwMkYtZD/uffKxMN7YlCcoI
lXQN4LboOBHCTTsw1HVuPPWv/6r+9W7V+9J3wXzhrgb/c63R7dNGnnW06BQ2tp1npbEHG525s0Et
vyWXGTqslEqSpue+9WK3hRvJns15r3papUtR6kqKeEkMLdlJlkxVybafOKD9Zna1l309HqGxQvK5
Ml+gXLdeZWqzOH9FBEUAPBvvBaY2Gh9ZoVODgmR1VdD9qL7/kaSvvzIwMn4UZWHIKTWPXXeW9+oY
S9uwUjbBS3kl9tDRMk+4EcfQ3C6YYIa6c1xbeJOmJFWAvlRdPzOkwtIo4vOPDmwO2YLFrM7n4PR6
oJPAZ3FJ+ETtFtQQz21DiBCdcH6t99Jv0ViWN/s7tGkiotwDtMOos68j0xy/YGF+HTqIvxR+KVGP
+eL7IYjGEEXpFDDuYUKmELphfV5nomOGzt5s8dA5qafCmcGHpKHA3keEq1SmXOrHsVAq/6gg38Uf
/Etxrfsq7+2vwOWKR05oXovXRZ3GbcXediP+o+cWsdq4DvF2F0SJIrG+vNyh5COHxV0kQGoFXJXs
480gyVq3H4aOYZooqZ8T5O5nyZnNzXHPzxs/0FLv8q1Sl/ua7oAVLFAv8pI/lTmwpEcOTP2SyB3z
bTCzIXFH2uCiwLbFnYxQR7Bo6waXWjfRscxYa/uT/59yzTfp+4UDSIOhxrj9cJBegXEKTWA8Z+oQ
RBqL31HIQ1ClnGuktRegrs4VxLKjbIbmCVR5PwYzECpOAXJWybmwCsoB4Xpr5O9tzViyj3guONcr
YMc/VhWjTlRO+PD8IKppEGjALPNJUeUCovrmW1WLWH0i2/3u6Ce4tdPMC3344z0L0TDLakwLkym5
2QO8rwoyk/xXlbOk0/X5yUoAwuG+SoUE+NJHxQKQ+bcZwYQwDq8VOc01p7theB7YwrHGrgOcgIzf
/jMADPxfACE4UB84hC89BvFKNfKO7LC6JfztJwJpJzdKUBhxlc4k3BL/LMIGo42UqLb4XjttSYuT
7vQutL7MvfCwu87wf81pbACujV06K9SVl5zrhON2oHlfmMrZX9/Y/oDbfclbmXX34pcLLpij90MB
H6+p2Tt0tHwgxM05xtBEzVkCGLuBa7Sw0SfpKmSqMCcZ06d5AXzcEE9XmS4D9eUxyZohEpZ8pZzT
F/shn0F/iYvxBt41z3S6h+ENcgpaaYKmH7LMsRWXV5hmLruBVW7ZNkeVtk//grE1AYoYLyc+wNFs
pS5QD8ieLSEjfdi8n2mdiZffYbAmSEX7FJd0MvLaONMlC/a4/Bsd45G2lEKe7Pw+BbCNFh+rYM0x
1ZAqxprwdSiY748YuK5TmU54MUzCpoN/opEBKzmfNGplWGY03e4KF0aV+zXVV9YX6/38kW+dWbd7
2QLt3oWNco92L65BJmA4SYAv2X4/UdRsR5axs1YQBmKC7rfP7JlBT1zMzhoXpvJ8Lq8/ge5zLGrQ
tL/JZpm81iiY55/D4H6Et1NRXyQcY4JR6UipmqB27rUcnk7U6ggX+ExU2hN0OBULsBizPgv3WyC0
0yiAAo4NhEEKsYwK2mou8xUW55mCUKia7twIchYY7z+wLW9GU2vQV+yxjbozbYTxLHO5/1x+noKS
zqsGpnhVyvqxTj5yNVFX3hSvAXosS2Ayf4MhKZnAb2qD+9wi4IH93cApFet4XUNC9Ivyo6+krQUQ
YU+0NFGMUP22IxROC/UqPvs4k85ZxGzwx3owdWuw0z6z7bzmm+rjD0VEISZDcz2jbtCgq8jt5QmF
DjrjXaD5u4baPXPmxCfKYBYv1Z/pvUozgRME93S89Lv4qMIQXTkuUz/vSqbkT1im2Zz3B6yaRmxO
hpGZqaE7xy77hQ9m3UkuKin0yShTDsj7tSvxT+uyj6eFCs5QU2dur+78YWFGZYL9NfUJ8U4hyOto
D5ny90jVdYaUtceKVM0H0r6FDzbuhbodq/DfdUixM7EtAlB2F8FpJILowmLHywRm4QydIhalBndJ
NorWgUQsd7DbBxnYfJXrcCUywkpTCLBWIUGgxsSPtPIqpf7IXiOB+kl8izSBhPT/shs4kn3Zdgyl
BtjS7AEfY2kzygJuIwf9qZpK8QjJkNlOjtDWbtQHzfMGb+fMYEIksCSGcCfGPp3fmy8OAzSa2Pv9
F3Qj/KJJOBW2ADHvkf9kcxeAxnCcMTvQSdT//QHUWSokGjyyFMd5b169f6iY3B08YezgS1GTX11Y
ldi0jygshyh6gb6otFu3lK7oCEIB7lsxU/iYMh0sZeAMWRdWx0SmMpkprjDy4N6MeAW0Va2fZzg6
hEYvJFk26TEpcWFRQM7Y/RwTRUkveo9lS/teW11RMcK+Jzu3jX2U1KpUfjFhQbzNnFzqOXvws68r
2PFJIuOR/slVfhmL3ZQaqscv8WCMGEnvLvK5cdmMud/pg3VjhOPpl4YhPCSa3NIvnpcJs6kEGMsV
+8pX1k5oQ3dgLkq1yJfshtsxlTKOpwRSP1TlLL3eaLbtIf3mel144N1ubjR/cLHG8VR4LnvnuNym
s4mopDMACRiNcG7I4JfjZ5LwxjoJpubDIfCStW7pMNJcS2eGZdrhTC0fvcvdbSnZCQuNZ0pkXPqm
SJl5QIYRidpvWqFyULXMOaIGKgHFvGfI9uPNEtcVuOpMlojnu37v/6arxvPMrJQAf576VlC2LJ/F
pW3qiueemOvqXXplZ2zCuuu+C0aivex4+YxkBTYw7ok9VGp1ylSMXz4mhHl8DnPvP3Mu3ZOxkN3m
nNSyTsQ704LLRzZK752IoKaQSzONPwvVovlDHbt8lAXC43/rAD+tIsJa0DdBlEXjrgEx/BluTvDC
p85R88dt+x4lriv8bHKcRj8s95L2NZJrniCaqGQumFBf/nyPn+6kwIo3CoN96saId1lLvLhtJwcU
1fxhWhwr4tbpHViliKsaLZyIvYwbUekpAinDaNmjc12BHG1WxBqi0vPWaRvXJc0nNXtmkhXouaH1
ik8P324F3u5lAIGjuPnt8ypk4zGIiHBFDbI+O9IROqWO0Spj1ZGsGkGA5GkOkNcN4+PnnR1J2oMj
29b+e8Pla89xnCnJx18cNmklI8tFesLf7d7wVp5/oPJKlzF/ZE2fELuOnwdWXw1VsDN9jZyWK9A6
NXIqUdZJ3lDxozLmPLJtSPnQmSFw4J8hV4pgvA+ItM2s43VB/hOME0TrwwSSRwg0mmkYM4APEb0v
6V263WJ5f03Pu90VJM1QyVU6hIvOLfxScIymwscb7q5tTPmFlDRZuRn3MW7g6N6y4NRdRshJJuu6
3+BfdQ8Gicv7DvuLBNuBwPOr6LK7Nzd+UrAjZniVjhoKHbeAcYfQ9XzklK/6hB8rzIKV2qcDAQ3m
xQ9XFjHremjgdTZyYv2ho/xj7BPsVGcxhKiUPfctNl+BuGh71YhOatt8ZryRBVAJXVTiZ1fxMZSe
Q8t7yDQN52BXvi0QEIOOCPoFW1TGKKL3hLtWgSzpAVUKfFL2uvRsXQwzq3A6cJ6pf6DwqGmfPfh5
fioLhwl+HNxnsQWTByDZ2ow6K1PCik6gOeLkJ8jwOAsWj5Rtfs7Qw5FjHLgILmgc3OXRvxZ+2ji7
MotN0TygMXK7+gSj18VH36AXH+qjtm4b/aKZZgUT+qwwE5evV36tIuN/fBe1JFZh6pNG66TfvNKG
3LAV5fx2OjrWzvHmNL3UiUsn+IY6ZTgXkj+2xUoZBJj49uHYGYDdVL8+bf7pyQ8zbFelxMFCTEQs
WLSLc+O+5Imyr+jXX6vps4CD6D3V3hx/mDL07TRFOp5a4cIpGe4M4cPvMylLNDGgddIPyz5wB3uM
TR1V6ik5MPgUYToNmG5GtDdnNBARARDYXsrm/oPs3Ov3hVynZDIKwIiFDlnY3LHDl6biYdbUNHb2
7Zlv9Vfzb5pS7/MlYAmm8UtdRvXeJzCekiDvudBeebXPRGfBqhtFnHyHRC+WEYzOnn8VLTHPciHe
sb681tIYWocRe8JwNxh98PKadB0Rw4CvV+yoL7gKmCAmbOV8k/rjaibzAJLOlx6pLZTFNg4jv4xf
FquXuv10GkMETO879HjvqqcsZOAombtWQ0GVR0QeGoEZnAJnuF1jz23Cv369I5OdR5LRCW2olBMF
G16YWqMGUPjm0j4EHW+22xO8Gp+dm0/2/zRf0QrglN9Alb7HRs9Nayzq4tZ7jFTT5IkTUV4Gtp6g
XacbGeaf9bSstRf0MbqSWwC/5oaMyIpit0E07V97G08PohvcKVBL23Wb82CRvo+wQ6BA/0JZQoeG
99H06PZIA//t5HG1Bt8qUps69bsRAngFEDNQK4ASCV3F7832KKhcn0htJ8NQigtf9vWof38emqSC
2qcLrvql7ENY9Rigm+kJ/J3JBG9hOhtUdZ3aOuePom7gdB0jrJvU9dMemZtno8oJ5cpmX4NlLoCx
U9nL698yd1BPsHpKxrJx1WlR30GvfwAJ+XVGkKp9v3LsHFGeD1zCr5HGWKXBx8bziETS0qRkbZiG
0Sjt/ITERSANYUxvv2icsay8hHh8Sb3jHspo6HGCNSdQTK0M9+lnQZJAOlj9NMvE/MtwKf6Yzxdy
XmCUx0Pd1MaViL+auLvb75hjqR07MLG5Gqvi+/PqiKDHVpVMjIlXJNM/w+VuWcdnxBiTgNFV9acr
d0JeDX9Og+mwofUs1M3YtciTpJsUxOcQarKIPi5wCjO9Y8OBSBe+Tg+R9VyCYbBUfvpvrCs/yUoM
LTuTaqBLbHrpJY5uNRTgtQasTixob/1oOC7czikTX2Jt5MMjDzNL+fMnuTMHGFFLcke0rH7MVzDr
NPZuJAi944O0F75ARxNwnsShpm1HXFlgY9Fx1c1jFQDtFTvS1UKXgCGkpni2+r6rG65CbvwfHT1r
foQneiRS6L8jihfJtDMqJyXvZqoIufgxk5+dmGj8/vV81/IoMqMvwVG1V/Q+4dSKdpenaDJwI9tH
9mUmepkwkuPtnLpjCT3SIVIjxuW5X0xaKN51m5vlWPupJe/04vdlsG0WB8W+R0dvjxklARp7Uvdp
hb62VSpxZK4NSTZxQ5+nzmi29AabAQ467gxW7Qj3mWGIcL7wQEFBO3uxX99FjvFaTx1loYXZ3Fv5
9Bnt423WgT3BIHQ3VV+PxLpQ6c768F6zb643rI0Pd8pkqXvES+8rKNPPs5q+kp6orQ2XLcteA6Bc
PlvPAWUVG3FAmVSthjmYiGJrQ5ARLsTs3BnAuI8bC7gEnqHJvw35QDmBC+XesQIq+/5vPOqU3/cX
ptCTj3m+oxX+Q+7EVcQNbLgzJeK3mT8kQB0uRo8ciN1FSZRaG6vsk+7ICMuhlsDmOkD9RPwckMyX
yZV9ROF6uNwLVS9VaBe+p4n8ZKBIwPiQvzqje6qqcET8Aln/HdzS/A6BYCCtnqDbL5QDAN9Es+LA
tcam3ibtaFJ8qzlYecAOaJurfD6O57hMgDchvPrfPbrGPMXO6RAMDVuj73EUrBpno+I8fXzsXBoM
9RyzZAVQ6QQNMgu8mmORenz6V2b99brG6xo+yTlgHFAxyllPyV2YF3ZY4/0rBz0Gg2h3NBW8Ii/4
scIX2S1BIccytumqolAaibAP8W6HFJKJjWYdsgTjLfRVELl5C/1z8jB8IxH3e6DVRy2SP+Kn3XAL
id50wSEkX+X7fAWk9rormuprg9ecta0dvRPmwfqmsCJeU0LB95oD4SLtaiW0wS7U+Cn9N0Ha0BaQ
g2q3dxSaBXmNoJCLJ0kbJWY7wOsQaG8koK9d8tGILww8HC3Cfszmv4Y/JlQWGPqJB4Vprobhepuk
9gAnBY+JlVZw5INXE0v1oU1luwX5e3rvZ6hLkZRfXurSQDMi8ySdm6VXMFitccaAYOuhqTestKkt
/18ig9qcfjIFU7stU8WVfqHipG/rIsVzaf1N93NDWOjzAntGScq8SPfbraQTwTnxaSLl13xiV1Dz
tQFQJ/yHHDNO+qB//sb7/7HHLfAWdeMMTcT1nEm9MmaU4z3WX7ZaAqWjNgPjnS7uziavQnlqPOr2
aaE9EvRN4GsCZjK47uSyQfdlOrYkOB6mDMSB0EynFOQ6t5HVUZVCK10jFzYyUt+llpIHQIQJKZPC
csr+0aMpQH5O/T7ddGUOCeFliiD/ZkAZB/SqkB84GHi9odj7VXnEQDndDmh6qdq4rfDqU/Vob49g
llE/PFmuCNGt61K31P7kK6JN0mtBUoXflD25EPCcsmYCSaDJqTPcmP0gnhDxlx9lmgJXI2o4D/Bb
b7+V0Fdyjj2Gv+7/k1JaN1hTBCgnMibhzer85iirSBNipSbbwKTLhmVlEt+cUYMe8wiCQY8XtyTX
QysxNDBTbntHeTnGO0RSwG96vAigmYqZ/UOGUyt/b7AJfHzjAkbCYrFqxfTD03wuBm+j6Dst3O7H
xaBcQdoGbFCkLYK1IbQfVOnR3LGkVnNTZzCEB42Z4NibxslXzJ4IWYzhcQI/OxLvMXoEEBz2ZPAx
eLv12S5Qq+gyPxiwRbAPjAtvd/JLwxxOen21g/wznzt5Aa8xQqxz1NavK9dW7Ze6UIHfV3fnvkbU
p/VBLrb6PPZojYGoRfWC4bYrKaPR2xUsosIBtbzyRJ0952owG20SX7ZwnZuR8Wmfc89dhjyWuZ9Q
0Li6BVoYVLY0UQ5Waxe5/DjMWqjwcjMFAEnpIrslOf2kQGe2rIzElsHNwMh5sDgTSXIhJr+nQV75
lpoX44pnoNriRzmVejkXw71lS5WxC/ryJJ//2vqEVezfGcEtbzmuDUip+rlWlkmTdNGfGcT0Q5vN
GFU6zalH2ha/scSA03fcfi17vwIPlnvdVSy44R2yZL9AaUjL+gMGDPzNH3gX//h1FUql0gB5dNhb
6tgWi2iYV85eOFYzx87Owe4Wb55ZqZ0UhGLMicF1cPBwj9QwwADrBhXYCm7zsyVn4NYRkmMA7kak
kNLm1Cqx9paTSeOOvCsVc2O1FTK2kQzjEpP8+e9R9ESj6+bIDaVCF8dEy1fc5rImxnNuQhy7SZAO
dfYoMHKtMYeo3ny5O+A0Dj+19WC2CCMz/Cdd+nOWT6/oshutWmjPcDPyHP6958OOiwXRtkeNxKva
udrOcTnarzPFX8lc/l0gqezOD7Z0zlzZMPRXGYN7CeYvIB4H8n9hbf4guCf4MNypg6kSIbR7WzFr
u3cdUNe8Nm+BA6TC6A0MFOYt5+69hx0mJ5LjTvwj1zq1V27+8wfo4TY1GE6d41iGhFa6khNFBPTr
1bXRXlBUX9FSA+18Aa5HnVUWWDMaIMOV7kGqtL/5pjy52BSU9uAhbGuzwU4UL0fA3o3UTKX3lZtD
9b5IdchGMbFtNE3Fs2WV4zx0e1MOQ/jAFZYJvB5n4l82XAo6JFH19A9Exwv+/lqFIktl6wRxbL53
HKGK3yG2d3YIR4HZuN+iL/g0L9ZzIF80K/8zpyYudB3aT1VbPL7vmeBET+Abk4URQ/pgF1Ys2OhB
KnK01x1i3EHEqfpWmXudHv9xTq96KCEL8ZJWXQqr4QkIv/ex4qlhZZ6CBzhOiE/Hc73QbQE05kqq
pU6ao3TJ/K4JPjRseI8M8HKd5WTNqbJlZaO8shQMkOGMVaNneQ1y32jUpn/1UxZs9ha7GdEdSyXO
RvI75VqeYATYkgdLXjuFecRNRGeTZK6Q/y77h95SDwQMbbs7lOkcJ1VZLuDPXmXCJC7ZbdQurF8P
bmGqsncTf0Vaw6J9QmQUdzpclKRbnvqeriYs18miEfp95ZKhxDp81gVTGQ8NSCby09iTb1A5tNu+
eK2X50bsF4hiRTIeNQpOQc2fbc29xXgdoWQ7Z9QZDMOpakZ9m4iTAIjo3VhiAwJoIQ/4fOAYxDRH
yOcNhGIiNVB66+zob6goaKi0Lr+gAT4SqsNfIrmRO4tY/4fO6BUEJlvJrlQFkUo0AqDhhif9MEPg
FBeiCw+6yl4J7ztnsfzjsE4OS+kE0aJkqmGszjgEyMrW01OG4hxS5XCXXsvDGU4jtiBfHYj2Wdm8
nUgdR2tdBMA1uQQnr8HM+Vvmv1vjpijBlQS3kKDWi7Vo1xjNy04bA5RiEKmSoRvi00e4Q3BuBJdf
E+LoZcfPtIzhIvgc6zSV1ea+e7tINeUvvUHKrvSJSFH/Sa6+yYw68h/6QNa2dIRgp+FleTCK8nVB
270yHzoO80t/wp1xshnpVfTdjloRPPakZ0X4yCmiRuANOu3IIKo9P2N5Nq9FHLuWyTBCk7kkHYFb
d579slNWIghsMgyYBJNpz2/oOa+U1p8lj1SK2VVkCRnnXTRLd8uCC5ErYb63iHUl0Crreym5f5pu
iOv8KsoNbBzXivmQdn87KaTCFJdX5N46ufuyGB9UMYVg+zEtibydyaEv8EGwta1NbscMfpZOp2+K
n5fFTfdwUozyT1ZCwNPzy20W6J5GwddABESeCvRbcBha2gIUTL7D8JmjZMuJ7Yc5w7VMW7HP7kb0
hAWiqPfSS5+aeG9XSXtM5t/admSBMxJgwEVdX9bemGGcQ7whN0Zrfg0z9RWkD2Lc+0NodUn8x2fB
nFUQeNryLvwrw0hkCL3N4W/dtaejwnd/zrkTCRFo2NjzOLKoViULHBebZ1++o9ZxXYb2UFCjRqqN
6HOpKDV3rZN643gN20OKc0Aaug9Iu5C/oBFnYZuEd62Cx+g4BBnRs9wFPTct40BUIP2vLGKdExbM
kV2RDsUGUQUOS1LhEHBP2AAL2iOKiKM0M/dr2jV212/JuSO1O9mOiwiNmLVGkHQGPYOJeBXGGjXd
SmqFznKzwRWlUDyMVHUnJ43vV8ERFH6VQsb89oG9dJg20WNySR3IPN0/Yacwz2HPG9HqRIgjmoCH
LHqt8ixpZqS9g+akUuwTjLq7KyNWUFNkjF6VUUCaowYwXc5iC0SA/N8rxvZD95ihr4HCz1Q0p7Y3
QFb8ImZJtU2Y+f/hnK3LCqT5iEsD/mFJ2dldHJtp4CUdb9KZYHaMJ3xdJx4DIAy9RRu9NgVWwNsj
G04bmYM3dCAV8CzhHJpFx5OhBscQ2xo6dKiZxE80jA+5F1zdnOW2Xtu4kVnBHWBkA2ueifdew+Zh
t4uJou7kAP/dhJPL623XAZlS6UzC1ItlKE9B7XNe3wocw9iFCI0W/byxtQsCLWcbO4qYq5/5m1E1
tsiwTFsg6wsuK2pbksSEWnbP0Bx69uVXdYi8t2dExQomsuMRfzymQuB79ykzUOOTJwsigSDzLEoO
JPOBNDb5qa4RTho/Ef3ZZmYSK97cZ/gjkYdd+SlaLUxGlsmObW9MfDn4NFuigUIxncf1eQxjP7BM
e4pXRAYz6Fxl22mUQeZs2wRaPMwSTOCXYQWupaYFKZSjnO/CmmhC4UclWXdfbHmjP6OZ7t+kmvNl
4VDo0jTkteVybDT3vNfzhmRtavAaoSDAusTovprAdAqNd38QW1p+FHuWkZoCTidXUxvxwz+meC7J
hGlM8bjK1uuc4Zoupb14H675xcwB42+r0kNGZvNn1FHvHaTr0IYS5ZtDuOBHplPj0vqNxZgdaI7x
1CWP/X7BuLKC8LDW8NsYXobyLtSH4+RbT/Q9JexVDbY9J2Ehhb9YiOXrhS07FD01XwtJPOWAsDpz
D/jaNjdaPCewpQL7SgXG1cpGfdZP7QOutD10EkrbqC4IZ+z0I3Fkjqwtv7P7WWLyX/OX8pYW1CQt
qbe8X0ZLANfhEyqRGwvzA0ByhrzD6XUlNM8x4EKoO/XhiFc4GJ93rNCYOI1jzAomYOK92akr/5pm
g5Gz8JPUg31ZzG8mvfNp/s0pcMcSqugCEcyvIyTFsWs5YUKv3KXfqWcheIYiT/tFJ6eBwf0m8g6y
1g3RZrY1BQMZU6ogr+Nah7QGhzqx0c7fQR/aeKO0hc4IDd9/32ABRj86+EKquVibMI8MNgrqX9kZ
WCzAeLUTi3HSvO+NrLE8YmbPW7rtdOUaZKRdJcCcjr5vNAEKY0tv8GNgJiGfC+DnJepfwyl6SMml
GGjwW6/D5hQo2B0sSekhtAoeFjRjUf+dFSQolNENQPvoOPIWF4/HE6rcs8C9uxsV2uK9a9A6BMKe
QTChWKpOSfgGcaa1pCZqXCK3gS88LR4YUPg5C6n7ORNz7hLcemwNlqSkvjGk3mfVbmCexlAITJvV
6xxXOFfQdwS4jLovs4gM1pu5TIVQUaN0aXv3ixeOn/R2hgXlBPjjfh81c5dPbE28Kt4B8A0me4QP
vJe4etdMNdgJhjPZrXIXzW4ZKVLwXZPTStddwEBpyy2KNaSpo3REv8OUglxbDEJe2otOjhCVDOcL
YNNAxoCpLi1o/aAMX4vTmmjt3ahnjRYVS63HGoG+ChFD6b6y/bkk6q8ajQEtwDTU4zIly8pdYsFt
cm2mbErSaecjdz0oaxDuNBHeAyxt6jcuoqFrwo4+/Yu9+fVPhK+jqlpPfWiuPgbtuTect3RV6RhF
6PljMLjtsTrnjdPxfj9D+3wu4XhPp3yDeToP82rJ4L6NGmj03hKgOIkAG2yEF6fh/BgWpxkGcrqY
+7FSr96PEllhjaNBy3/lyejJK6KEP0x4FmAATglKocRPGsC3XDCWrVcwsnrBE7HoK3WtAtcq697r
D575lj7l9/mOJ43z4J0UU+ULAVRrJJWJONlGsUebdIajm0eQey7G3tnI5dlej2gwtTcN9F7ZyrrK
2AzHLPA2ygetSt53zwEkbQnL8EnuISzImAQWEeWY799zMy+aZoAdGz8yJ9WBWWLrCrdyDAQMaGKp
hfkvipAOqgBJIlYtyOTdmQW8zTDrVTQXk9rPUSGS4/9LO7pwSel+MajENFG56TYkbVVaNHzIibgI
W7uEd9BNdLMZUkdaswe3tDdqEi67re/xLukUEAEak3ueEbE1h/fLnXrRkuMAUn9aqM4zC3yUyp8c
WYU2bUZDhIegquUegTyxRlOvRY9FH6qaYv1pzp/KLu2rGoKUUTqIEw/KAvG7yyddpr48NoUmKwvp
TWNDi/AthLgOko4iOt412+nM1NprOq1oQ4BOKvzf3MKW1hMH1vXlPrTvggfYeALpIBF6xyYWjuT5
8JPdJaJQb4zxClovXTF5w77FE0Pj6+bdW+FUxSICTeolwcuG8uFqCV6KjRJMopbgQMR1vhJc0A4+
1Cum2uHnz99DCzgKld5Kie2NUlKv3cdK/d9no/9ry4BQ1FLJTokXgMImc+0ZK9DQspgYZvxyTZAN
X4AnHF3t/ww+w7Qwm+5uDeLTn8LWfcrBGe1HcSM/7fSS1Xd52RmlhnLq+JzCWT6RW77Y6JgXfraP
KrxB54tLJ2/xbrWkSa4An7jUh9VxlB8eechyo5jqpdp+HXTH40A4Y7R0xPZo9vptDIxxjPOwRgaw
HEoJj3oNq0yBnyGuM7dVGQbRu5GJSPPoSuVQCxmCdHRsO/JqWNjAB379JCaRSc36QK1sJjg2f14k
yyrXTTAXut/BOLT2mPr+WVZrGtcouWG9lw0tW1DNeqgoIiEQIEVTNbGpRva8npRjy5HJ4kAFM2my
9kjkUKvwrlnfJzZiZTNjxgN+RDyX1goLLUJnuxha2HATzy1HdC3l/uusd0ziSpJFCQFAAUFbmUjY
kuvF9Yr00zX2pr00pbdXaF+KIMKdgAol3hvdSXhOzqQ7vAvisuXWgOTfzwH8nsYrcIsMDZ66t34q
0Ir8zpNL5EPErrGvbjzrKCTig7VI2SevoOKBHONyfn6JTzKvXHFC5nmbHgcf+AO1PyrdJmpUbG6t
7j7MGYrOMSusVkjStJ/pJ7cBlxZ6o1hjgIvCk8JQYUF55PH+lrh1YozpQ6YhqjhX/10LjuucF5An
5KeWUXA05Cv8MTxjsJd2ChNJL+rlDeY2jBpaySBuioeOblKiFds+rB6/bGyO2vyscX/mfJ+HOxi9
qSpmYCNLSNR5RKh/hjEUmw8F+3VS8s1B5DCI5MuIaHxWxd09XTEeeYN+xo/nT2ETBhZM/wHO44hD
oLu9ybxlIC4UCd37Kb65Ut2p/cRRx8ld2eu1Nbo6uQBSjPP5ODOAfADG3fC103AimIv16M6PDz3d
51mkHrEj0PQrhAMLfSAwBfhXkJ5whB//aRqn9BxQtTbfUz/U2OL+B8GA770HjjkeTVM+eOazK9Az
NisdQeeJdXx+ZpkRlraJn23AXI29s6g3BOvPm43FVcIz+C2LXpftr0GXcSKNAu0UinHNncjR8CCX
mjVkjufnH+r+uW4cB/bN7VX/xLfYFSqY21256fV69G5+YdzKBGsykzBiOSbSQG0U9T1mBmEwzhMR
rdzj/WI/GtMBktjhLD7iGlW/9IKBUYX0MJ7crf953bP8IghtAMQO1xBEpCpLk5+pqiX1PQidMQ+I
54VTByFVdIYq0fjuVNqdGcRJVUtsxBY/LebIv20lZ01MM40waJBs4KpjJXHSqDVT7M+luNVyZjfj
DVYYtDc1IYoSgMILazq0EGTkuJPMCo3oeGctUxM7FcQqJ7c6+XCYsBWIIbuNoIQd+nPCMnu9/4vO
DasH2XjXX6ygk3lUpXlB8nieof3K7qxGDV+SYlYBQvayTegQl32m2G/C/B2T+BtxIdgp0Zk6T/Ri
MaoSpwxpdZC3gdFhKpZTFlzqWKUbWVeHCXwANsHOGyWn3+D2N0wi9mfHX0Nzuh82FHsiDO12qsUI
6KSTT5RLc4uXddXwaVLS50cAMMn/VDTiA8kha2QSacyrIfcKjpeAu2YaY/oX+G59aahXU9XnfGur
5M9JgjKXdNhtRs6BqJblPOZCMJaDF359bblgxRTMCRIjxbFQYtydBx7NjDKsFwMG/4gO879kToim
tTmwdVKb5vpkH2UUVoGonyBWnRw7y/Nj3VLpIyCWaZRwGKyunAgi1/eayePwrlqrvSFrbxglMsUR
T8hIFFcjrfrVNWcQ3K2X/7kb4GZMyljgqEeKZoIgUFTzZvC0Ycu7g7PK6IsxHfjeyIKaaQ8N/RjM
qo06rr2aDUO+6IqhsNNLfQP41yldzUNzUXgJLVJEzYuKNmTrG8ztUxEFDf54E3k6M+M82lJtB/sj
xapDESF+h+llMOWZd8Xx/mJRNQU8TDIpVy4lITwI8XhfsDrwowGMBOOaDsA+WlbM9YNTjKObpLte
yrqpRHbF5TCDBKCdn2wfDHJ/TZMMwi8G3D+EJCThUuAfeeAAPrgJPIX/uSth5G9vVN840YKnPPZk
ckTn58Cwzd14+hBOTYAedrEQVQvdWu/bdEbpPdbXJNiSeLoCWpmU+ZfxqOaUJxbxU1eGv4fMk2AP
yS5T80lFQepr+rtIw5DHxriz0ElVDfVflTFbymHa9H3KEpsE+CAHDmAtViXhSU9WNRDv7AeslrMX
mrxOq25m9V+QGfmPRxwuxJ6A3Rt3lC/aovMMsobL8AFVkv6VY1Eb9E4lxCyCQZg/Dl7qQDUd5m0S
pyHz1Fx2WVkgnSKibojss+ZA/OGYsDSkhT1f02O/yM9u8m3uHxGQH4eWfEWNEHZhHkwVugIvahlV
RI+Nbk/YWUNLHqusRKlrFH6mpXMWhBui1RMal9loFRQwcSIAcqBnGIf34HxM1KQDaLB0SQiA+jx5
ndHwMj33y6Me491GyjvgxvcNqT97NF98ygETDbCKDDjmvm0DSv0872GaYOaX5f2JygvVeHuq216c
+ShuUa/3oULHMj+COzMs8VuuUQk29U5BTEs/w7Vnf03A4LbTj6KC/TTUQ2Nsd8pud4V4DA6VAJEa
VJYtp1mI4kN1UGpKemChobIT1ujwat/QEbVwUty9M5WWoPitKg1JYozVN3YPrmjyHVxWy7bcrEdk
EQt/Q104UcL8DFIbO5GsFJpmbtBUgWtVgHQMHNRuH7aMeimsxTko8U+skrpU3PEkNpIef/SYVeTn
bJXWSCtovjFR8Y48bAf2ITIDHCqT4XCgXUU0UUZcZbjqeOXIP2o5ACyTsqDZh1iezFBrhaXRF+6x
1X2VBrCBp8TA/pQoDoj8O0k7bCnWyC2UjkVjBJBvlW6/a6AK0kLg3JJL6t/d3fu+A8SHaYu2YVgF
Rcbd4m1KSWCS+fPF/B9298vD1SPM9bZrfjOu2OT3HbNsiRzfLCLDqOBhM9g6DbbDHjfDVlNSLuK1
j9Ek5pzLRgYsBjRnlg+JfxCl3LhZrLerdsqltSlVqpV2+vxFHQrAvMOKdGhv34YIl8yPwAhkILko
HaEctTia21WNpWvSdcF92bzpPXyn0yhK72ZAyuzfkaXzuvLPbvtzK9JW08BSYm18Pv7w/8mY01kk
c0KdU1pWayR1oeFcoQv65cbrF0FRa3DBeFn3Efp7Z2Y+fpxqW4AmTyELMuqefxPSydSdl3U4wN7y
55Q7qQdNWQ4vI05/qK2Uathqrj8PHTV/bMxrgO8p0p7K31EVUR0+eQH7YSPl8h9148IWHFwtAt5o
3t/aHP6WN7k9RTszUhZQvjqJWRfzxu7bRXjbB7dG62NjH2f+uO75KA/Ssx3pyrgToTXkXSdjwBwm
hiwKup5tsI3w/tf0l2a8kvHao0sA3NDRIrTxSE2pbYH65X3GjLwy1PIK++b5doybuOAJQwkn2/NP
f+GunKEgffguanUDzyBgj3Lh89A62VuIoZl+nmGdPiE/LcSpfJy99FK1kZnDiDSRZM2ICyblouiv
XruaiTeWIOVduGtJNAzAjyZ8boSf3jFhBWfDohrpOkwGrR15a/K/mpf0dpVGl+E2MoMMrq4pk/IY
DzEWM2S9+2Q8cHCg3VS2bfxEV4OCZTOLJI/mjidf3+cRnL0pAHufWsPMWA/ex/i7+kDLzGgS77HU
tf1rLmMpswS2hT+E9OPiL4OpxfEUdhCFAnf6AfEJvz3Sdua+bso9iIB+HjQBXMIfFB7CDEi2cpdy
0b4uYJVmanNBJNJht4onvyIFRNOQeqzbtYJtBNGaq4/+DptkhUZuVtN4AU5jMHV45XY2H4TRcunl
14ga2XwcGRTJznQk0JIGssv0JylDiHTwg/xqB0a3xZlEJlbjc5ZMmQ4AGQiaolWr7hGXgpLFebpZ
GxcQcwhxjEPscRtvc95sx4Bw6S3f0asEf6TpSptlP8s4/iMLBWy59VLgQ2whuiyV7oVGbA/NKxaJ
jtoCLIeeVMASqdmtg7PxjA+xCnidLaUY3wjkost/TR7lyl+psyAAzepIZiQXs0QSnL8WTwmi3/Ob
ZyVWbIzOvRi4zeMMgewjjFTTXY+jVV40zOiJeH3csKLKCWqWJXZDmxIAKn/yQ0HDLMzTqk35ZYgg
jWJj+VDRhITs79+milK3xOXJsGcjlpagnpxCVskYBBOkZYgeuSGI8Sx79nHXgsaOddqSpgLRYkKF
I28CJRdSd8uD4BXvjl58in6IWF4Mg2ojiYz/f5vJT7dj8/a3hqJo/jzsT9xd6xo0fYOstztD6Llm
2nq0qe/xkVGOsfgJzTykJ7f4Ri7jFbSNe7F/RsXR6YwEawK1Dg9kJ5YBxp0Mj1X4U81hoHxsPDwP
DMp3YxL+sWlQ2SBdrBMR50VYyYDvlj22P5X7nqQGNAXFIjsMhAvB5w6CVWvhS7ZOsIl6YH/qC/TS
EWlwJkq9tafY2PyrPPIByZApAJKFq2rTDd5Btgx4DQB+6iAbaG4QiNuIB67QUE+Bs2ajJx6Y4vVS
eS2tyw/t99Hcb1rFKGU2ZqryKt5AIwiVZ92Es7C818XHcc1N26fsrmFFo4YfgDKUtnc07dacz7uz
qKoigh64sDxGRQShfpKgAjkuAFXwjxXjp1HiAID1Brbe0bSLLgCKRcgeTwOdTw5I+gsjWUw8TQwv
mmqGoPVCm1LM9tgvlvs+qH/MkGwLTnCoZ5W2mSnIDRCEQuhXL9ElWN/azE1NejiLJFBgG3ZaWpVc
Kh/hjCfFT6Z7E45y8heLsxrJdEowdslzp6/FY6R+09fTLHlBS39/PfLLhwQELsBX/44yN1sy0uh9
hxNXWsJq7wR24q5DcavS4uNTV41DpLFelBexePv3uwzhSAjSRJNVSHvvPbOAAPCGQzNdnuMPxWtE
oRtzjFI6WhC6ksW9N7TVdZfC2pbxtuLSgdGAkUTf5MzCCa9/tPJiFPL0k9v4zkypxF1VEDNrcHl2
mwAyPAOn6DYbqcyh7FUJBzGTzkGtmIjIAaacV45chi4nl7fZKYNovtuytymyxs/RFuzOJGTDCbqb
a9kqTmEByNr/Q28L4yJE2tzD4pyUB4yrRHy5sPre/W8GWn1ZgksKwOFikvWY9nb4LUoteo2I9h1N
ywmEoxXsG0DzN2OLM7oHBP4QFSWrXxBoJ+cgEM6xLlKA06Ai49l3Hmx55dv4B1xeO63DE5EP74fU
qnTgYwLCoqTFi9rhw6NpESALkYczdVs63TS72GbhtEiIPqj9TnRKAn5rgbDQZghB6dpCPnFVuQsr
Rhslfi8ZAWxSW+FxfS+AUnD2hpcdjjgQ+Wv7BNjy6WBp7W4IMDeJUyWZh7R/dwzoMZkISoVfOPxY
1wkKXVSJ8h4BmNtLUvY5+wfCTMi6vsEN5VOEpw0r5oCpv9kpbdyYmsfSmL7Skh5fuYtx78aWtwFV
v40WRE/lkhEo7GS4FxEH02ePE18/QfZn2CThTXd0TpNOQtFDXoFzNVzb5QRPZzjL5ryu97p1cat6
WhRsM1/UNgcjZV8aVjbIt5uFVecydK/tut2xvp1zV3nNEBy9Dvq2WUyRlHDV5uRmPSk5PpmtEtQC
Ki32ykwK9ry+ROQ6iTNU8Pbb4HeJrmJBNJedj++AUHHTlQEUWxUZ4RGhr4EjbrhbuKgPkpOvmkQ4
Hd78SKEA9FSqfTXmqCK/DnrSWn1YUc+kLXxhTQED5fKlcwPpJt1J9zlrwjK18oMckrYe/2qlhS0N
J6KCJGpiPANbgEvbOxH7QBYrfP6CxjS8iLp054IeN8kUHA3vrBAjZMYHVR/cIZjQEtRP/qUK6p+l
wpwA1C6lUpTf8/pnCcP/eEF0E3EHfkBFYW9Q/YnPR9uvN0h/xX7An0CdBUNEMQa0AUrE0fJEQ/yV
hloYDuK65Dp8nE6KHpl6+Ut6sgUs9vbohXp3fhKDX8c9HEW/CCqBDMrug3Cy+NPnnEjY03Kks6v0
QbBpMZIMYJaeccoHFEPwe7GXFigFNLa8xPUnoemiwpPzhwFAaTFEDHzAwYYkslj5fyY3eP19jTSF
WObMvkM4upyh6nOsHkjABVRq7IIPFRwOeIDwa/Bi0WITwkw6PhgDM70ICjSKU2G+6I8eHK147kK/
tj8+vwj68ltupK59KLwsHz6pnChKKw//Nc89Z7QgdlB/3up5i0d7A++aunEZQIiEDL6g/7IV28OB
DvcBu3vwx8Ccs3wjw30olu7pKdMdE2rTzIu7Qs6nptC0vlXfKIxNtZQnSCBslawsYnj9IWGUhT4y
AhYnmNkztqaEv59+GWOekD0hLIcGwCwWYDf2F5OuSTSvnTj/xspAPjJXgnobGAVk3a193KIgbpEe
LQuUOmw+utLNjh43l7gBsCDVngPYcnLYPeRt6NmhwXG6RlS0kH8z5XFsMUugpjjzMOWfOWtllNA5
0l26J3B2wqDUwoFTGvN2+4KDswBs6zQixbax7cNEnnrlpwF5pVEG5AMPr0qzXscWhkihOkknJ7Ni
tVmrx03cXw51HFue0K5NNy2tmgNotWiPHsFFdIQ8xtQNXHePd65hNckTcvy+kFtlnKKgqZsD3ak5
PuW8/RqG5nQlvuQ6JVfAmSFH9a95rM0FlShyhKNHZTFbXKJjgG1Do0gr6wijgFeiol6CEPeAEOon
/cDaiKX8fKltn9iIf17T6YV+HmBkL0ULnfb56kptn1BpCQN8b49MPh0s5kiqWTclVW+VfNYmlTe4
0SLpdYrlrFfuYTKiXDA027BMn+n//EE8oW3GtEfe44eiWtxpOcm+aOBgUESEM4Fxo332F1g9b8wZ
4J6TuELQBpuTyBSTT8APREIMCTz0n+no7Zl7RJSA7gq0aIAbJ9cRYcMUgQIlUbSjSnVgHNCdu6D5
VnBeDqum82RetrBUihr7oKDyNpWXRYP7YLEzkQSoaPlX7umNC4eRktMVNqcZWqSj1Cxleo1tSV0e
2wg5ZGpwFGoz0S8Rm+F4nFFJOlSosAmXBFuIDuzjbX/W5bD9GAuWBAFwcOlZjRF32OjTxQOGJkZg
9w1IzQ2E3XzTQ6bfF+fqmTAyFb1S+vvP6ftIbPDSdbwtM16mClAX6D0uNsiFh4VtQXoVse3rUfNM
0St+uS/tHFi/3K5xSbBGIIYEEyoe6waMUdTfObxafX83BxLO4DZayDjJ/L52B9pNr2G3r4s+K6AA
B4CYcDoalgU3AyS6W21Zs4tiKW8QKf3IW6NXoXoRAtJKOHrZeK25HdSo31rcaAYDRmgcXLF0K/YM
Hrut9fTfZqN0VR9ySgA8CBvxRJrnoqOgHMuJSFaSwwSQf4/E9CVNdRqmNCG5/V4z8shIQFVCN0DM
ETQQu419FtWfFwy6rZM2L5oHTYa3RkbIy/hynwoXF3Tdt09bY/zuNSmapfqWUuGCq9i1xoeuntU1
8R0bd8ottfUIrItdlj8hJmMDsmi1SRrngueQ/dQmyDlSwHcMUq/Ph4dI+cys8byCSrj9F2QUZNyr
OlrzY6vE6lmOWh/SXisto8rAnQNjNOJdW7c5+c+EIV+s0P+QNRvXJEuUxWwcp0iwftu8Hu1hW1D0
axiZpfhVFDbs5nOXeqj4dJUBvNdosu+V1EqkVY81/HSlCdZ0NhjKRm1KirDW/hf7m6RFhus4FkX+
D7z6cmG8CatSP2tJwPPmkdHZW3K9tK+VRCzj8EsBhc1KP8kkNI4HM5Kr5EWZObjaMn5obVFoWcGo
eqOWbWUAEUJ0/YAgZmKywoolHv+tSr+rgj+uN4vSVcOIz9pHWQePh7gONqyNpwslXdoRmspBISpN
BIcyie+yg7m0fcOWAUyhhw2xNix70bCFYfpX0JM7KSjkEwY4TH/uYb8ZDUCwqAF/8g85z4Fm2l1C
p0ouK1AS0oI7XWUzjZe/hoa52YTS7MNHGWuz6WZ7BkHPmSC+m7qyw/4fjbRpZPUeQro8dB1jTKDw
uAxjM24NG/tSSkWz7ho/Kf2yntQtGDIKqE9awHpEqISOmdAkadFvoSRF/KC5vOwq/kYC+qSrmNda
vWJ8spPl8vJCNHrvPHnCdeJFr5EjYXVg3BCf4wdmS9ZmVDDlnfsmAX8uLQWQ4Je3Z1L8KxgbDwKr
GaU8Ty7XkMmY1zuk/uvPQ0WwR2mrFGrKExzR0aZhK4xdvYP/VCEeeKju1I/QoEypt0ofyo1u7qvn
yKo5/JOGVese2sMBHzuQPmyi56DABIBmjflvrzdwQYa6vSlQf2wz5FQNTF3hQ4UWInkcN5Xt9jdA
JGduDnxgn7qFIwd8Rm5M/WM/NZr1bidGRQHHIWLqfGraHIAtnYnKkNlWMfEQsfEu38jy3Opdz1Pq
ZYANuLwt3cxNb82sX9vVXVR6sMWqO1RXJJk5hOnP8vPFEnxpi1fdfSXduksLtwBihlOkFqRjy0YB
3HCW0lAxd2zdGjda92X4TEPFr8qq7y5JF80m5GepdsMmJt/5CGWNltNrP7OUAAOxCENMAS3fkCFJ
rAyse+2Sdt+zW7IqjK10fbrFPOtcA983pOVIi/+9PzBXyWrDJI8qJ/fqjmAmdak8+zznH9j6joRC
egRW86gFal/wy/XTiuNLFFYp2bvV7+bHzFf7UnMV4uYGWjqNy8dJxtVreqhPoRmhrBqMIYYqUomw
F7ArTcq16OQ3a6wTiYZoF1KJZjTlpx5vkbQmtczS3J+F2ycREtzTtKByBi0FdlUcdiJaSz4MMjMR
6HNRIM57vCYDTc/hrUgu1Hub3oOrsG6oSqFXZ7t9ZRbf8TlnkkiUoU0hpQdQYITOc0IwQsFHs9Xg
Y42zyVD/jS8FyFgJDTC8wdpSCZace40mAzpaeaMIvdbO3ikCWNUUH9e1tXHYdBckWSY4oOqwq2dW
y46BApZ+ZxybnsVDtLlWX+CL6GIAgCpVUM2aBm3tj7/dXqkmzRWnuSojDnEw2bjNFGI8pYyRMNXT
SBjgp/l69xOeLpt8Jlpw5hoU/0RK0K8A98dcJY8omV8gyNeSDm2HRXCyaSi9PUyiYOX0pBAZ4vow
hpLzff+kDv3/6KE4FOG+wYkAhenqTbGbaOTQbovtRqN4myiOpl5XAZ6ImLqMxDj4+X8b4nC/QBDu
3uSbGdUQ8UDW1loc2QSdapGragPFe8ZGIJTzll2VHkyqSVonDVmhAVHB7Fc3aAV2FKtwhiQocbxz
5EYwsmVoLFEHXW0Gz5YhrFoiwJ6AN+lBphDplL+yDpvzl3TgiMHxq1lp2tAyo/MWEnSI6erTzPIn
VYhcMcfNfPR/0+CYWn1BiP/AZxpHhkAFWN1jMdspTm5POSH7wnlNeHzf1N63P4ZxuUu6O6NLwWX3
adiC15nE0bbulZ95xQDSn1gnYVr0kvNIbMBk54RYbNFpIU4kU+TWAwUWy4Y317BVmD3YZ24ds1Rx
ShLblnEVO7yv+zGMcyAVSVsyu65Dz71e+oWRtCJUl062oxE0rw6CPpqc0baao1m0iBvBVXxS5uIV
yXkg48jyphwwzqOkUSinrMrbNI8h5q1qPdwK1w9rJ+M+ZScfmN72NHpsUQqR2O4cx3/61YL7ZIr0
lt+XDsQNwkRMeD/1LHeaYHmkUlvjAnP4bn070CZu8o63nLavPT76I2i3+/htpl16PgJdDeIXKWAi
363/3auIj5orZtMc7e8isam1n1JkzRsQyDZoSfN2BSOTl5rFKs/LpGUin/8ldg+/2uIJFLniaPdf
RJfUl9Yv+RDIvDi00xJ193yM7nZYpXfWFjlxnYRVUawlGAh9adRRkiwEE1IwEqpr5p8TElJKia/J
tazRuJysFPG0x9Gn9vSp78IG4U+faHP5OgLbImCQQgoTRAy8+CTUuvDYY5QoV5sesAbXsUjzV7UK
xgx2O/GIHpI23LKOwtiVxPybrdcf4bhFAsOHzjLxglGkke7vEeawxKPj3bfeJPZ9873B9jZq7Onk
2KQtIixvxoBDY5AAfxtNmwer4INLdXqifF8c6BsziWAo0CgqE8GgAKaC5fSk+ho/A/llOqH3UgP4
ZrdX1Twoeiv7qFCJA3Zs0hmT5HTY4dU3rDCGypuuwsH+olt+E6FjrwUKbbgkzo8KiUyEnSmilAeu
8bSCxJrQUyFIMRcZa4xnWXgNK9iCa7q/zz80vRwXMPPjjvpfq7LbY/K0YcZXcpXeYvaICZYWWHEs
9fF8jH+Zgt/Ao52d021he8o5rp3Zj+J4BH5k5PgIttfxBcQr9uFx4Qjy9Gf+YnXvV2ik223zroaC
EOyhdRs9NI1dIvYIhn/fp2X64K0ldCkkH/Q+WD+kCRG/KN3Yi9tVZdYe7UfnHPOAsssDP+IVzMQR
aAH3HjGoaQSdJCjwutVvwXfJplhNjNcIHB8yia8KTWOx1ZXzzXtJvZ2fkTAmJ7+NhbU0PGrG5JWf
woHEhxsc40h9kU+f9JzK6Z192sfrKMRStmDiywCPxRhpD8KoPYYwGe2ydwAnlXu8W8/XAScYOSok
hmV5EdVXKG9iMdfyzqpbkSMGgi6Nm/rBtpdQLcj8OT+Q785mjo/nh5mXWU4gSTfnGUMv2Reh7kWK
SylhvPV7i71UV8ahJuG9j2jxGf1v1rrOpZc2CRpGFx9nxqoH6YXs8Nj2wVo/fXI+RjuzzyYqAcNs
+MgVnZlxNsBlJ2IC8rn0uNXgNW9GZQBX8NKPR9thXgLjXbYbxuoQfyilcByyU0gdNVAAmz2J+XJ7
dV/sdb2q0idLcXd8dR5p6b/nYlwfOAEa5D5mvIZQm6dTpp8zsCydh4AVhQ6gWHobw0N0Rie9RIKs
yxuT+E+ZwTo7KFyEBE6WqLxr07W9FfgXEqX0k3nv9ltbag5iY3+kxy+c/DdcIRUVrNshZBZflYxa
LlCXh6AbjiSfkz0EriDoEbgpG5soqY+SlfkmQUlQXLziNWk3Yr77XGj2zHv0mvWrr4sLeh3r9c87
I0NnG8WH1szVhJxpUBJKbcod/6jAe58hdLTs7ql20g/0PDagebUBue+VVmAb9+V9S7nQP7OGM/3T
/iK2bfplEZ0RKHJeDiTg3xcBxaXkAZcS9qMhGhbx0ViK12o9TRuMK9wFBnQPUVyQ0qfk1BMFxp/e
gGZxjZFgZrcmDsHtUzk+nQBpLJN+qKrGvVC4p5anBOOthXJKYqDIiI/Fx4MMBfqy+9MTcgz+UMyW
S8+wrZ4VwRceWOVwHqDGzO2JrrbQS2xdEeh4dMf+zNMc8Q6VIin1DwzemFlJvRlamoDKJGe6raE6
qk7aqJKLZG2GrLk7/euNsjKeKoCVHfm2qnIk/4du8V6OOr1+F37ho9dzS7z2VYFaPCJAylXb4v/X
KgUAZUkLqFU1c4K0BUuNBFKwi5ZNJ0NB97hh442QeNstCegPTfJztFnKDvoVrhomrD5VA0NVnoHk
5Tu1NbPlbwPPH15aWRjC2HB1tRrfu7B4TnUk7Rt4HpLOgFfEsYnvAHnNxlct7RZlqZlCD85imWMp
oAdW6IaSs5B20quA1H1c2up1XBhIkwqtka+PwXde8YkFb6DwhuEEqAceJ5rWANTFi4a928yCRnuq
9TI6WEYBCVlLwtFtNs7LwEJrtl6Zk8BUUGzFdIpSLXXMPkx5t50p/d6hVZ3iJb5c3P8stVnpWiDU
EWiQIqkGQHZBrrVW3emMxjR3V00LsCOObKvg/V6lsecEvpF8jk2UKqF8hMc9g/GloS1riM0QHGJ5
eYxqAX2dRGrMW6lRNaounWCEKhi5sKecdiIckOcB+8jue6MsJAVSnuJsEmQYcpOMCYEEJfP9evKP
w3OQ35Gs11sTEGQfZ3JndFZBq6wzwB3HkMo97sz3wA1bNiB6UmI3A76ZIwZftsTm8I01/w9MsCob
5qnBU7G4syBjY3u2S7kgS2kXR8R6d3nnlgwaAM7/HyaajloxKtm+aRcCwIksu10qLfD7DseQziJu
s8EVk+kowgzut8X+t6nwZOd4Z5HSGV7Avc6ERkrjw6P9bBDXkhd6RS1nXEsofPnhlLWkdXQgy+nx
Lgqg1KT94tWeHBxhLcWz8g7GFUDQUBOBk8ThxHcDzL0MHF9f+uvn4FDXHw1rHJTmG7ICQYsiyqqn
doxsZ+PZ6MR+78sINIcRhGSup8shl0x4YEvsVG9CteMhiGPEb1jVfbvy8OOB9Yc6Q5reZqpoORmn
u4lBBjANnMdESKRjo76jyJeZ+A9Ec9657i4JtsItb+/ouc7eXQZuNRTz+o7oG8Dcq8e8OxnYDPpY
eVlT5eM0510n0BW5IADQBc6YLtUGV5nP7PwFN3xs5M1YTtYRmQ8XcaN71K5m0z/9ifeRCZ5yUKPm
CL2UNzJt/hLsp+UGoCxG3skt80xfPB0pAxB/7otJxzZImcOiV5KVMnpwsziaSWQsSQwHgqw6TsvC
rb/gBxnxMvYqcl+jbeMWY6pJ4SnrPsZAjTUWbCltWz4URTL7jZGQ5fZxRtAR53Vpe+4HI+Zfvedu
5fVS7ieijkDYKLBf/Mw//2FP6oR7NPg6swVHN+784UAZFSWAQZJnQ4Q21yMjAMP7LEsJNcaTxlll
Dr31O7OxY8ud3NzDi5sHI7z5139Jhp1MGAsmNiT9MsMkLIECC/1yYA1+4JhGPfbkDhUTCz3bu7kI
nkLSQTAFURrFin9TBio7lAKsrNCSkKznka+wPoPeTCW+Ma07LMZkx/AgsgHa0UWx086zDTKqLPKO
znF7MkSi2ADjT2+0+dy3CRr/YVqliG/ZouO7H5St1kUU7NL4795u2uFfO4pJTXzPKS7XzYmKD1bR
obJIaPfdwx/dAxjtG0WoyfY1oJhuLMdeL693IS42Y8dAd8Y5tkPmHIPezNFNjuc/l9iCWoa6cYX4
H8Fah/qtqW5TuS4WAnkKiLRvb1kcFYM355iWbjQp/GrWXbG4CCxPvnPMTKssnelYRTX2XpTa7F4/
RGiyMT6VQVb6QkH+lnOdife6iYCI9clbINOyi1EiqiPGnbulXCIpHvOlrkOFTXOplHTeSLFYtsgL
tJnwTWkeesUcfmzEI7C4JNWuhHurQYGQZpioxj9KN/sCijagKdcGUvcfFcEYWYZDbUJI9Q9zPOYs
w4TwlSmBDAGYZQkKPOAQvWHWZf88bQNorcEWbhkNu06OhtAA+Vy+5ip6ft+5WCKJTIQjFHenUKc0
z5jBwnOoipTD4TcIYTmDjTNuB8QBJB0VXvjM8YSL1F9i4q6bX6bjajmPEedqUTighL0sK7rUPOYc
29A89un9XCptLGxRfSE4ql7XFOJ2akiPZEsq8OkMOczw7dJziFVbN58F03nTV+/qnWST5kQ+ZMtl
vMl0GRK586PpDpoO8thV2YL5drfr4FGPEwlalvrkujOj3U49I2pxszxmoq9QS1avY6KVx59lKIPs
0TVacJAOzg9i5yq+VjAoc9/EINXUm3APEWiSvKei42657R5K6BOXEPzHXN/Ot4rw+pa9FzR9c0Qh
2xYdbDcfN64iRTRbdmk6yhL6sIzlhzCjvdgU3noHByzARHRz8M48damUmaN0bqc5Y64kJ0OrbAuT
jOf80Pk4fZEDOVmNuLIohds4sEW5VzusBvXyVOFerYdEESWvwQrfUFOdRj9pe7Qo/kyLiCWiOKpW
b2zr9+Qw3gmVpEHt7BxBTF4FwCMXuIFjzEd9AraJ3u0JVsyglfQHziI+N3Oco3i0RkUsOk/R9o13
G1J9VjodR+xQG70NZY5MFY/MUKLfzEa98UNf3djvB/xZQexorBmvrb85X9KjpijOEXMPx0Uv6lDG
zURiwizIE4p4+Phc6cWcWnT9eCuXYxQ5HZNBNy4Fl6e5QNFd0ND9OXX+cI1M09cFeqzwunop6syJ
y76LHAkVC7HNQrVHMxN3/RINAS21fzrKvaFcFTXGUFaDnWKWMsAD112kEaerDEgZkrpXHLmbmS8L
7SDbK3PZRDvLWee2x7R11s3haFrZKKfbIIgTmjsBLC6gcMj1mSFt0sLMwnWziadWXPtTbCbiAa5D
WURAW4y4UAitLcCG2k35ztWyZRuTN5posMTsGcHajZvpzS4WF3O5120COtrm6HRuyBmTguogqd9i
czH2HVARJDElVycmnppLDbxzKvI81Zbdvpp6VGBKgVHHkoFpdzHWCsgahUs3yzErAVVVx40EM4xC
vuOl4kOYTV+gkb6h4+PgyyCDepJkVu5Fp3k3zPdm7iMYyUOErLAFQZwnmQfeRvWpq0qoXLPe3jCv
escRGJDo/C8lPjyWA6Ptm8n05EXFg7Fc95yT2av1RdFjaHlL6P+6v8SxuM5qD/gGcBpsKb4Uk6dr
Yg+YmGn/6QZjXZsTZqWnrPb0qbIMLMb3gdVFONPgu4ZncKK/fQmNKFVOoI7PHTTV2UBI1peENK6a
0o/GP5KDVYrJnzEvBkrp0Wc4i6o958PY7vQLue9zsLWnldLrgjJn9e+2cb0+TBpHWd0kBRVFIBtc
2uJLzE2hX8GRAUUtJr6erlMto2QWGPUNwCXsBKcAkQ5LmxZd9ya+PaJcWEBNrUNjW6+Ik5oondRg
3eYQ8AJX/JHZ5IttkUpOH1A9nRNVF8QITybOQGoOR5b+WDD3qVT4FmKjpDuFySHiyaAI2rGuzgbz
0mSLT73VmxdsQ/h9HgWHvmpkbru56VuBlTEK+yVDo1cHlH1/sSXf94jbtwVRekWCi+cvUTb5LjOU
hVb7i9OhqtPmXj2oVeFIaPptXk4ou5ncFIkiLIR6KJm5glYTfQrge9o9RQ1bkdvt52IU75KoUZB5
TGsFsDRdUFB45plCud6N6e2YJEG4RnVeGQmZIlZIgOzCzwizh+9YZ3V9iwhVDjsl9ukcwtiok3We
SxA8RegTSPMzAYfs0iEPfPhhZxRcgE6u/Bqz+SxnK4XZvdTxOLUrBEXgBXKLMrcdUHb343/5pQav
1WZvVzUkFBWmy7KdzNPkEhCeKm34NQdXWYMausJqivY5uK0glYmapoZVtozLKM88F7RquHOReLYc
DWaLDtMe6i+MU9B9sAd5OJfV0w2whNffp5QyvXihHkgDiMAOgiafeNbvp/bKY7rAV2uzEVyVaFfE
Zbtls38vXmNfdZoocfeXV3n9t+1odG9ZbAmVLRwduvxTsb/PsEsJG617JAaEnpsJXK7mzAfmuAOW
RK5WWZnGm0olBjMSFfibuwr2QCdaH3foaj7x66rdHjMSEd12YXAhFQ8K0yccyos4/5KlSkHWYqey
HPADaNUAx5XePm5Wjt4+w+HhN/6YdWVtoEHq/tbj0HiPqG80KmtrXwXiRf65AIxBkybieYPVKwe5
N25HR8NA3cVJ0RYz89Se4xd/k+0TpUY2alKiitnC8iWQQ7hUGEOp+4h5Lllo3eqhXupiZJODp1AZ
vLflpTmrhO6NaQwifAhWFP23V0vlVhgvrGPiTg9tUuglXHEbflhivHT6RqoyXZDCwGAwNMuYbkWk
pEOTlYdL2yjTjuf3Sj2uURDAoB4TXBK81H+7gekNrMRXfaz8O0LPZlKn+pLGCbpeEpvE2I+m0gMX
jW+DThxBpND+8mSWGxuDpH51/nxnSwA0KEHqSuNO08gBwb1bQ+NeBAhQukwzGsAYAV6uB3RW8Njf
hSF6R5KHjCtzJX1qsrHZz6uYhNAmHr+dqdM8ugfGQz1kq6R3qhOYMcwc6ivwbAYApE4SqlZrvIoW
bVZA5h+cHqBybiJO+Mnw8btq/093cR+nxeVyPCBnkLMqAxe3QQKOxceZMnFEVHnWZkTRcebwU/7L
pTsbaLLc2XFHePHsqrg/ZMb00IZYKo7A3m6ZOp9xXq7AMwjY/OgiCWzzvceobHb9jUckFosRRyiu
vMXenjybULF/NLvnVonTsS0LA7EpXJ8JE1myXBhqmK3/cqvycs5SRY73AJOukCeZcuW97XWnYjYp
taHwAT2ETQAioh9ePap/KI/LUwx8UUW2ptX9ZpJFcDdzRtRfsY3Af6kUjcR+C0WL4Nm0/CU/u6vh
MPVqkp22zXMOI4bwDHXSZT3S7IXpvmukpulaHKGkUzkB6DK/mp27yra9D4dWYa3WmYq49N7EkBs9
tekKDiNVbeOLGGGrqtaL3Q/ohGDhfZTcXuFvIf8juhXx+nmPo0KpATRd//diSVK7V2JyI09Jjy6z
SwbBfyFMT0LGISjvoAY8FwkNOp7aP1+BUcPFDjDQVKPH5pfTdQnx4ueJC/9IF2hGiP/xKAju/QtF
j/EdG5Tpt7j6WPqufyzfgyaeo1Oo2Nt4mTNpTK7uo9KDzemZyjPeavWowFhUq2sLLvZzc5rAwPAn
hx9RQuXuuv/yMSuVFxKlikQ66dWBCEsHpysLmzY0E9Mqve2ocEHDR8SlleGxMApG0xYRafDSS/jw
vDUGSTDOEvzoDGRGdQlGq+RuFSP7Bc5Z8CEFsHbsd0tPxldXWryhvTz0NI0H2M/KzatBJ9Ai0onm
v9PHmNgsl9MdltvhYy4SZL87rwjwaSUtcQBcFSaykORyI2wyV+pCjGK/p/5rPHODudnr0oqieUAZ
X2mTKZgpAh5mkj+Imk+HYcHG36YBv5dS/RIDkkdgAmZOv0N+fVcB3Z5px9YDTEeHA86SJGGsbuqH
prB/LM7w6Ue0C/9n1D+zvyb3JamtMOScqQNS5l4tpGnbF5K1RB8J9Yd3s+U61a7qyxNfsV8u18Kv
b11JXiy/BRknRwqKmEt2ueaEgJzcXnIPKxMWKrYMxpZfznBRDopAshSaa/7DDS2koODpt9IystNL
HTBB09VxeBq5Zf52LxI9nxwpj4R3EVXwgYOHzO0X5KIjUeEH/1Rh9uxJRPSyxofotcwXDAUvtA7K
R0LHTWLiHubqZRU55oGLkwsEL9H1pN7ck+6bEbJg9J4POEQCemmzwD0z/+sUaQ0iVoqgmmq1J7vt
S0TxeOibeZNaQjyskuO612WJ8x98ZVHlwdfmJ22hh/bS3WHgPm1envk1GqGWk1XoMWlle8RP46J+
E9GeS3jyv3z0z9qHyUgr7o99AobrE5BzzNcVt6m+Kvn9Dds0VAj6OBXrpi0GGfKIh0W8VdRyt9sm
U67pPIxu/nhqItRc793P/YdY1viD/P2wbEvbQGMQtJuf3jk/ZT3Y7oIaQcg6NKbUp2YEJEmzW6Sp
+gNoGUz3dmnARGxyihFMMAef0cBKN1c2nC+sAFzjg9G0sqy35DHRvG+N+f8bu+0MCRORNAy9GaZ+
iDldMuZQZlOG/3VY9e0fakd0nIYdsRVD5u90AM93aD5fZDIULRWo7mmgcvMqsH0QcwLTs9jvBBLR
jRYmWaLGp5v17mhvnn4Xafu8bYW4oJ9XQzg1PRTexUaTX4RVyLllzEG4LSpPKUHWbK/U5p5Hyy1H
SdfMVGKPXuXex+VXPn14t3n9y2l2HMY9P+SAYAhYNczYfsVXHlKOI5bZZXU5BSxzFalPFJweWV2M
kQ7lSsJ+1mF6fZ3Fk/Ll6gM8FqFZOQnO86esSpuAipiqf8Dcyf6/VtMwoLL+gWbMREOpuWEcIcs3
adkE5fK3nrQpWJG0eF0KmZG3zwfF3DApPdlcimxFyWbwznsuPmFjTS4T1yJUlnGGIhEzvscxNTSx
l+58d6mietu7g1Uwaw3UpHAuNIE0W/UYBg+2BjkI+MGAs6ERagiHW8vuvuu1NELLcNayck07f/QK
1xIBb8bfhY7kWX1dh5D63mI1jqnJSnGKJ2npP/7JN1zsvZxINetu0HbUYg7Vq3JfsP4DGcLCbwCW
9Gt2SLFyq5Us8WA/qb/IFOobuwAy8dorKOWC+vkCCHzSeXuT1jIA9pk6sF3G9CuDtJXye0mKlMk/
893reLyT2DCrWT4KC0UkCXjXkEsZKwhm0Qbu1QXAWFGyH15dd49gRwLOdRVEoLGqOM72Edaf6qji
ivrZNbKhOlFNSbjJ4WEx4AiyiKbw0Cu38BDMvoBRp2+96d40F4NfjYOiTqqDNRtCcozbWnIoZlcc
SfBZXnFMJ9V08g1yS+rneDTbz3Qwb16VC5235WHFlR+veqbQr9fwwSZ75JbOY/vhWhUtmU2PyMgm
aXbb1vYG7VU28HtmprwEU9kow/ftGmt6AAHL47zAoAcpctPDSJlIxIRzf5lIWe3CXTvKMYvUjqRe
I48q29wM8sMOOmrFT7qHjTcEr25E1KoUjSYU8U7JVutGM1MGA1kDhzvbS3dA3/+kr1NzYethltDj
DKQ7u8MmLm1iQbKpz1oHQfWfT339zQokr4c50BBH17TPscGE2GUoSFKyYV98brGJ20fbATMwY3aL
arQNE243AYslLELnRSWl37qfR1ftUHTwWTHN7OBO4NIcA2nqjOHTE8aHUQVrtT0ntwTwmL0e+exM
btZTTlvfyDurFRwT+P0+6w8LRE3pLbSdaSXrDS6unJl+oqVklSqS16lW6ihGUoA2VvY+kRfl6Mc8
KhCwvYutAJngtssjdHnlP8tZ7Hbsr5CxpJXD+FjYSqKocs0WaxkZMXexmHuaaIlnez/qjsras4PL
p0SaAeujzjR3cDilWb6K0MSNsbhIY/UTQ9qZF3fLr5CY92nHix/GS4IYZUHKh10kZemYj2PPvzZ2
mV4WFk1ifptiQPdPWhJoRWaf7ryUsQsokkWkDcrjjX7ceX7Qxli3I7FaxTvAL1HNzNbBprxiT482
2nvleAn488Qg+eHaFSUUMzQJQ3yG01EZAK4qZpssp+lkoKK/1wbFHHWtyFm016bXxs0ghhX49p2I
QdfWZyrw9JHTatnhHlmhGU5S+qgMxHPNvP6Gd7Ov/+bDkUhP+ZDL6dwJycgFYrDQOkWO7RVQeC9v
SKwFiXax0u+0dhC7yw1sTzQ00MCSkDJoQaOMYJuHBlX+B7CQXXn9ngir4CCSBQCrDIdRAZIAwmAv
itmiS8PKtnMpsCv0vMPDPXdZXvTC+zoS5b7rn0u2nRemeytYG3xvQJzTl8g2kVYTSlHtNGnCAZzY
ggHmg+mbPzH6Lh7j7V8RFXcCWA3Z9kwkI0J96nms/lxN7YSm7OoaK1W5iw/Z4SIjSs7dA55Wfjay
Bt5xJXnYm4vD+7jx1B9W188W1hUzOEIsp1+hq4Rd1PMDsiiEJkcFOGEisQSGu0l7jiHYKo2XgemV
HuvXtjlbt+BicTt51+M2OuVTu9F9i5G9nxHsDrZdOSg9mgSY09bwx0SyGOCEyQS3J9fv4YAyj2Yg
I9KqG1/i4j/2dGe5t4mHOgfhcAmnULGRH8OwwC968FRPRHUFCOfDodnjfgwrw7qG6Opb3Mqi4vjn
gNapOOiAnbwP67Zy6gQCdmqCqMWK9u1BlVcqelmxvpakYecuWmFZDoXdiZ41mriOrPnWbJAfQazD
Khp+hfoxh8pIZz+QEjcmRnPzjbW1BI7R5XYnXJn+Tus5L0JaHMJ7E6Dbg4NBrOCtSNRJ1HAADVod
piZHwT2DLrF3lTo6cUfvr7SNCiEjqJ9Bp1DjUnq8G97nQoaFuGKUuygpFZ5qf/vqW9pT1Bf6BpF0
fIBCEfocO2YCrf6Nb6ZKFuGBpXj00088ayUYuh/kk9TDHQQBYwm9dqi1ikbGqzwRHSNIVMwojkPD
xpEWigZooQj7Hzic0V6FZGxCraoyzDP3kHjXFVIzNCajgeVgVLYWkA1gcoFJ9l/o5NDMOKA+3gqw
RZNKFD7kRGgy9MjlvnGvjvJ6gTgU+Fj5zCweRKlnfm8ebRL9tbSOPUuQSfdd5tl6ph88E6fG9dVY
XIz9o8DrYIPW/3kroWAQY9KHOOy2FZTtx/VhnbgqpAGYGlgbWZZkJ3WUSwdaoQdkWOOh4Qlbargj
1BDzpZbq5mRfWJ39x3AyYAbByOp6c70/CqiyPV5OeNU9L17LkQFZ7I7me7SP6UOegICGRWZ9z6hs
WOJGx+xU64OfMhO+uOW6CB6fwxnT9V38/gPnj8VodO9qfHcWuRNVJ4yywFRDeVHASgGedViDhTDs
pRc/UAJdu+sa0qCXGlx0pYO6Ov644fFmMQVdobvC9PGeAr1BCOVWmbYYzWD49+oU+7AX7ndDdsAj
j0jckwnL0VujxPXWjpp0AAVqnHhTEJHPpviIdsfJcDiCAxc2rV7fvSqEeto7xBV0CqSPV6euAsAD
/L3dlMKLUy2YmV0eqPrSGLzUhE0mnE9a1GxbEv1PTwG5rjoXzixzGhOs7c6iEiy+osoibCd8ruTL
xu+uiQEan/odvvHdXTTl5b4tfIyjoJ9fnL1itfx1VKw+Ou4wch9s7N2M69+AdDrDsksT2z647QsQ
2HE4FTWX9yHD+vfKyTjWx7oV2VY4vUoO5QScSzUs27qHSA8X6K056yzAVMlDRqZtxeOswgSZwXHs
Y988pJp7BBYe7U3udnNXJcJGJKbDbsDcjGo/FuD7QdoANDxZlChQDLKwLTYOqXuhYSEjyZEvsXbo
7xn+8gp5+3pyl6WBSiiDkzbPsRapu/VqIvdhXhDCk0bjEECSZuvVYYOr8vBbabh115jBqPikm1rf
LpvlZ9/qQmBvOTLTP+LtvjbI+frRf5B30QRfrmTNVHl//3rwGDFpWR4+BZkIS8adLCVjXxpGkEc6
BzXwKDm0/xxcbpV/vEZWhgGzExlFgbHzKM3DloM7Wg8pSclGKM1EDeZK9CzpIdIpAWrt0is0ajSZ
XnCbN21jWCngEOyqoE/PLn7M7Gwrpq0Vtr/8pbLpa8RPmlTal32hh667eb7tI79g0/xT6fHQjnyO
v/IgPPfbGnmGtQxso2JhPt23uieggLDp/5UTji3UxfJfb/UdL2MtBm1vNwrlQun7pQuOnhfqy09x
9TqHRsV6koD8ajRUOmZmrdWYXZkMKGfdQ9IDRLu2hpab4m0nln4WaH7Y/EyfmCL7PeG24tQRxYHr
Z2hcUYpa6VOYvtoDPUqet+c88cV8gqR5XyITYfaRSJz7lPjpV3qemPb/tcrkS+H+kJDj8Her7xj7
OOghRKvSnSfNkLAyQwWHHjLHNpLsSGsOdXBRaTYOxtsSuy/2UO50XSqjNHYHxOmwaCspFoAnWFBj
VYLZtxyQJsgd8zm5pbA5qqpxz9PySSkIL5aa06XoOf4yLFNdhoyNMSJY7fZQQA9aO/AuYR31gNqg
AsXJiXAQEMbohV/WqGiLuuXHfOeXKNFrwuzIQPr50jtEZ2opL9sKikUQkoPOmmXv8B23AY0xEZ6V
9nPFdmeU1qv7D05zwTRmE8BvBfAD6UH9PW3z9cSyP3P6aWoUEciF0AjHApxw5Njqz1PXbLcR82qV
866oTuUt/6d+T/0k+aVIzOzcl7xfg7HfsMp78TCoYIISxKhMaEWFh/WPz8A6iPNMR6RBMrv1mxyH
nFNusf+BtmXqD7Y21VOocPYI3cywOOi7OpCWslq2hXMwNoH4Z7J0rr2cqV7edRzF4nrvGCXeCSLS
UfaYmIrsJhzMJLu4DeFrd1BOIZTkxNbB/UFj0UwgCIZmgX9vhBBf9hJ6+DPRXDucRgvIenm6oAkY
7ET3o4p3am99gdj8X7CKUvV5X4vTO7fag9zJj86LboEqnfM6SZjX040YZ9AR4/ormg3Rg/DYOAYU
ZSPibzvCAUxcGEAuenTAkz0SDVJnOKEkAtxrojOmuBd344qJBUciQN4GCgSpYeAJVOdurj/B7DGo
J8tRz0r/8QME/+ntQnv0T8VjA5mTlS0fIR+ZHSjS5Z78K1tTOw2CCDgrLTNya9XWfD+MNfV1Fv0S
VCG2KKHQs5IEVHTQyL1+OGOPqNQOqZAlhj/I+gt4Hnmtu7DazASKm2ukuhuQqEe39MqpuZLEHdEC
7JSf/bAEjf5TGyIjjjeWxedCzSuKaiXe1+xtO01MVZekfchjcj53qYImwzZRtFH0Jnf2XkvpHWWd
Eq/E4RXqHkVx0vG9OqaX9IttDochU4ZCOZd9BHVvD7Hi52KdBxPWU3R2vA0wSkcvHQap0V4x9qsE
K7YcnoKNHyhgNCiKP5Dt8bjel7ijLFtsgbCLJfVkZTcuG983MmtiQ0OKEVpCiZTknb7FOoIxY+BH
T21XRymwabNKjsxKEHcqmP+QSN1TyPzvHdtLXHD7eweb6iOjkMTouqYGmgb8QoOqHbXfrQ9oJiCD
YtbDVwUVFx9nUyuLLyJQpnf/BISNPE6hBvvVrtIwRWG2QD35pt5wxQCiIcy11mNa5FZF62r55KIq
9+wmpgD5vWmiKemVf4rNI3JB95mbvc961V0021gY9ltXqp/ujzavCY5P1gj7mKfKMde9CQ5q0sqS
tL5ks++IawpLerZsX9k4QSgqC6wjvl6GpNqM/fgK75DlKa3LreA1rPTXWZpR8CkqZwbEcudg6k+l
/FpfYWl5Sz29BDLtpIw4i76uVQmmXPPrKhOV3RuaLrvBoUIUamfH/afR/0nOak6vyTv+xg/QZO7l
sQelcmi384C00WVFszeve59ctpYRJVa1QWq9vvxIbexjER6+MwQNShNzy0Gh2RbYmvlB7NxRhGHD
n8qHaiQwXPSIgdLcmD+xbroHS+VKe1A22NcIEWzRrQT4QWdyPUOFlUgYbUgvyiwouHgajAJsXxcc
Ju8eBl3FjURXfwrmUuojNT56/5GXz9dGLBLM99gz33Ls5Hzu/xLZbnda3+GlernCO6hiWpYlecYn
iI+K2mIpWHNQP7Fy0BUNWhrjX3MfQyjw7wNkUESIjrszFinXjQsuAX7h9UYHm0O3e+pXuifVmgKp
qU45rUEBuec68PxCCNNpBy8MnNdcsytUCBF0piLZK65D2Epfa4CL3WJx7hK6bdc6J8APK+Y1qcZb
vcTkvoDQyI5bQTy/rQqoxZbr2R78RaolAvO7XHBfzQnNTQ9daPCsNUbnra6STfb8CVfqZrEFKKmP
1zOyf7n4AI9uzUa+HUiUeYpQ5s8tVuRJLSwulnl8RniAFc1auzd6g2hevqIQ2/LW3J27T9MA2/vn
+zQXMxojpdRS1wy31rB9z2SjQVNvm3gmXLcl/pTzCU6CR42S1lbETNNy0m+q/PSbp0Z+YOXkoWlY
0DJpI1JKWqFCt0fBj8PfOgvnjiQe38FOVPbro5acJ2tRwDBchTxM4r+6xNVbOgpprhTMN6JjI/yZ
lTEp8kB9X9q+kadfWUsRhFGq67+UaWR/txe+uZGx+++BuGQuRHO+5j1ECSJkjEY/ynfBeR7drf7w
+JOyZOyAk8KANrwZNynmljQFD/VNqRJ3y+dxJ0ZZH142poHftLHlzhS65cv4H8aDs1t4PQqoTwmJ
7Bbyu0mIWCC3yScBVyjvv6lpKQ56HvNfxIqNdm7YZk85OUrVn8ZCA9mRnCiFcue1sXl/AYHiyQmu
rwTDSt9LecN3oj9YhNVj7BtMKe+Zlk7VSkW6/wPjPqGbinQTKL5/cJQYp1mI4OO/TlGXQxft08iv
KQcJPby+iY9oMPSHqyKBiWc5Sy/mAt+ejI0mu/Xz0Nr/kO+DdtY31sqOT2vVlpSpeZcV0j5UU3Yq
QipgH+Wt8xbNCBsj0PK5HcGHo1Ym6a020UuRya6GSSIdkDjHmw9XIC1SvoUIdEvqi9LP6HOMZM97
sk4CwxzPbxNRcGA6DMRiArYSHmXBnkKsJVqciUqkqQoEf554nRnESZGSbkbeARPrOE2Nmy4qVhQk
d2jPZib4lvL7YafUrVo+VZNS3PYXZeBt1lu4qzzrZQ3sTlnQlZuP/3cYCAshh0U37obA0L+jLuPb
a+8Fx82KVnyQl7IbxqesA9iBje0EYWvEgQdsrre69dT7k+elJpofivIbUbmeY8NJMMj57BcISaIY
tSf9Dm+hxheNH1ZSNbxaImnfCct5spUzWnboidze7KbFAEnkK/shzSux1QsyXUyJIUXCHTq9H9s9
/8+aHbWgXS3GvNKZo+lwFwIet0FMYpDS2RkkEbYR1F7YskllB+fXkNFACQI8egDzcR1IsL9f47WC
2ROmdhsjGXPy2VJh/jQvYZm6/3UIGYQXJrxUbJeo3HDBY1oRcvK3i1HFVnGGSds/Y/QBgkeL1Qme
PuA2jfLHoG+hTSwS85AiCO8h4fp5SXSjzGNNNBfcJPCQQIj7kYOxgLpQt7MTEcfCwnRRtQWyWvLj
w0O8uoUNZO3/jC6LcSl8K2D2LxPsl0O+1fsGkfdU0uW9s0IIunj6KbW7VnyGHZl/pNoVPCFPYCb5
FayzKuuXgOau1ji0Nq2Kn1F6lw1BmZLZBJ4zlHIZlHGZtlBkAtP3AUWVwL/Z6d4Q/8EswQBV0+NK
0IDSf40lG7PZOq1reITULQOwbtTy01WLqNszaZY/KvNvskN6ub6+XmrLoLuwWLfe8CWS53loIZrp
CUDzAfmXkOZspyVR2vzmbI31lo921jLYUUycfelsMM9BhllFBAMOtUdMmZrBScIisoimjgohC+Q+
p+mqI/3y76hSSfTpwHrNNLbTtq3nvqu4BuedhIkNmhpUX4pNRhq0qkf0GDW10fkWCCebI87iWsBA
olbodnU4D9fdci926nD/oBw2vnl6N8mUezM+ulOPCmsnP4pLkBMWU1TEWX3YL950iEJBIQ9OFxPR
SLGnXje6zLONveviFdmVmY1MYb1oMjkcqR4JHVJ3LtAz3OkQ3j+AcIa1TTCu0uL06JYHrlswkmTi
x3PsfrOpNmsfI6P8oEjOKurIFugv5bAr+EV/n1s3kQZC0HIIpvX/EQVSxXzTfsnNTsTzeiT+MBlU
sQqwdEHbUZH9tR/2HR/XeP54Dwqzd6aQ3ef1Fsv2oD1gQyy5YKPFEfEjN4OYXzZYafFya+GYqpTB
n9A1t3kVMuaukdiyA1hotB6fqiGt/OLX4FpKTu3ThiISeKSX/TaIicNu4oARBUB5DXAGGQVlN9k4
uvEfrdyTq/zlz86WRZxtNWTuKH8mGLGW+M3JQotfHH9E6gVKVXqNBeZNwYbxoGO2OiiL7DeYxSX6
P4wkcYMFNrz0XVwgZU0tG/FIERoHXa6qWvbcT+7JZJRfm9gKnrAq09/I3NDeasju0gJUyxP92oz6
lAoe0eO18nDXcrHDglZ1CcqJn+hFL7G8/0g8nGqhbJONPR8VkjmJrKQTBnUfq13CyNOrlFLh87hd
6mZ7o4qCjA11v8LncXjQ/QiYJV0hzNecoE0gDGO917fn613iaXIh8+MtDlAvKRW4KTKokwUy9eOa
8JaoMKyNbWxlKcnC9+nGeKgSkppnQmy97ulqLGLYWb8Zmhq+AYjbMKkfedmt7WWaY+vJFPcuEGnR
4UVW88e+9L5N5U3i5RaUKRBQ2jnxlAtz009kVMpK4wDxncq7Tm3RJWkwV2I40TAgttJ3OJOxMgGc
h80GTpY+uFTmx7v6O+9YxnW/MikhrIbLphMywhabzgvO8xLyrLNJGDQmCwkRn6Msbp97QIL+uUfy
fhMbU3/Ja6Ao5kLPdo8cNYTrPiiQ9hosBgTS7JqyTx5peV00WO92UP4gmomz+JKhSeFnrTcMXSVg
WrW1GFnMvcsthmLAx70kKo/Zrd87gHWX+WkN/JKCCUPpNpK7IQRgebP70DrxgFF5XqI0pwkFDIFF
or86p6crEppieF2FmGicla6Aym40nhXB8ZaAuUH+tnMWPgmYGxQd256wzsF0xF3DxeWGBqM16IJu
3Um3koX4ORyykGWTOW93iLE9jdyL0xpN4DG77ZLROMvfl6VD2iv/OIYICFcKLZmg1qUXmdx3bnmY
FY3xbn2Jq1DDmsmi+0vHvzxsG4S+RQ8wj+G+7HHpb/DES4PAPo4or2Jm0Q/eIN1EyD0RGCIPcLP1
8rQYyMQ4U/CGoxoie3J+j5AohpG4qdyAoProY7m0weafMLyLgEgyla5tCBE8Cuq1CcvP1K4TbruA
b3qxkxHw1LC6P83bgZ37F0gRaqSSijE9TMJ4A/Mjfq188LxTJS+ruOsPxgBopk8Itm8bXNZcQcuv
3ngRZ8Cr4XjCOU1eaMazjVqd0KqSFAT8fTqKlvkQfq6P1eCbnTW8fpcxN2KtrX7JcihpfyQX5r6z
WgxCYg+ouxBu88DsHXjFVkUjyCA9d5rOKXF2wW+xFQAvrgPlw0n74/xEG/58hsOSoQSvL6Vj4njE
JMeo5jc5SdOfI1xJmqNMYBugN9rIE6d5q3Nnj5M8tRiIsl1v5pAv3oBig/bhOpEP6Czf4TYEFAM0
D6rVV3YUNeYjpud1/YqjQR2Ar/Xy4/DKnhDY3/Bn27/9xKUYii9yBhKCPlwdvCQuaXViUybfpt93
T1Utc8mkuNgokj4VpHJe1NbfczwIkwQ4Tca889d0uB3kGg8HpJ6AKEqKpy+/VrvCVTyhl+RRJd3n
f9zUSqwpqH++9B2tYj1TODGGzypWzo+dZ/Rp8fuNzQr/8p8qKx9J4Yhrur1NZmj1gmDrVC54/Fg+
RbihQ0fEozgyMLd5dcHxWBR9ky8fhKEjfkOjXMIodwDyxEXiRkSUtxo6vbSov1m7TuDhcqZK60QP
oowiOR+zdhJHUEFdNZ9OUflGpu4zRacIUuHAWmwUFxeYEea4793o0yNdIDU7c92ru7f6Sqzjnn2j
mwz4dv5jTb7D3qBxGQEs0G8zx1QdOQpMYUWmtDR/LmI/qNLs+OSLglYRdg1HNSUzkJ731OwaGK6r
j3fHSHHftjN4VzwBd97bdgI2+SnNh+o0aUxtURrHuD9Clv4y+NyZot0TcA+Uc+xkL2j2d6L+tILO
F0/H1leOGGOqkbeaADCyfc9fv7Z+qhc7vIpDE9ugDLiz58bDaVaLR+ZpF/E9/w/d1/XK5Us27TXZ
mjqTqia03MF0W4gvV0d1Dl1ruKE8IARDCB4K+nXXj2cTEzZmGKMN4MVxWbJpMnp7zYlepAc5/rqp
ftZH71fdGJnTP7kS2kMoZ8wjDNh6aIn3ZtBmJGFTjS6wPT1OHXFNwjGEV5E62Jm8GwsLo/dbDQZy
Sd4jqRTfoegUi+DtdwmIuH++PBKMWZGpzNy8VsEu7oZDL3DRcCaSTyfHKaoiTzADYJgaFPDHmq1e
iv1h3Pb/PYkZtn8hZkd6nIx63pfmVLUJpWuOJpUpT/7WRq6L6NyPMwSvKPOMSxXHU1FrR2+/Auh2
FS7mmGzAeqe0zdOCKMTNV1MWBoOqopGpQwru85EE9P0Tg8CoTNBFNdlwtOxF6LNXkyHw+bQw6yYp
EZ4HQB64y82f8CnqO1MWziLClSFac14p9qHRZ/rZkRMavhA98/9DUmzvDiOM12w7alXpewN3vlhP
3MIByEE2m0pk431j35iuyKBN2DdskSboZR7XjXr4XMFcXaaR2svM6QQSB7hYDEE4S9tomkuZwlhx
3NYTyxibuOFOV08EwDDGU0iPYVNir2KQuQjK79oW4Qv31b3G21aAypXj56srQln1hLMWJpE3fyoB
CR+9f4rMabJso3kienkip5UrKjDgPCocdI3B43nVQ0uC1G73ZO4LGqY1FssLl8Nks6d85E/H2B2l
BEU+a0s2V3rqH9SKFxchYlq1yY4QTXOWivi0ne+4/V0T13IB5L13S9DbbuoCpQoFSJztPjunC8YN
wI8Rd9isUcffrI2mZSFKj+Ry/pFWN/U1atfUdYIFE/jlFZIaO+HXaqaGlAB3IT3hGo5vTCNTwd9k
BbGy2dA6qV/Mx2fv2AHo3wuCJJlGHLTv36uBpKiW7OQnIjuSsX+vQ7wKK73ix9wvqcQt7Temvv0m
EbAs14Oy7Tk82GVnowSFF1pX43jsr3x5fBq97kknfhV0+KVk5A+NQvK4pnVs9usQYJz0kLFMiRa9
Nu9pocOQcOejabEutopF5i2el0JdN8LB3epkhaK3Z3kQVbcxnXdwShBrqA+x/PPxvvBCEorleKvb
HNcdSLNbd8Wk9u9GT4K06BXCNbiLY/t6diEevytU9a2FkKXkF+ieAIbb6TT/wwZCOh/hMV6hG6PT
M/3jOhOJqT6kiJxLMig4b08RSOHLn/d/NmR+1jlMIcQ7P3Upon9YrEEsmoqiGWBbvJEXE+qY+H+i
NXtudQQarZ3IgWvZxY49cj0YU4zR0wJ3svWlWwnHHuDZsUPfdj6Cn6+VJzvIeT4MW1ax8Kco6jSm
weYV8xzrkGHUhtdjy1bUlQbtHdiccDXzUwixlketxkUp9AGmJrKBu1xvpkHUbNDwEQLcE8qfCO78
VKPsSPDstK26NeAgyYqNKfeUXiquTMWWvvexs5zA6C7fupQ0wD88PEo0NX6SSFYdQirTO2CasXDQ
TreyhYyLQc9sTrIqTqY+y5d5Tz0A3Pl4xNNNbDLyXGxUJrKgUlgXWMUifl+6Bw1x8HLKAN2asIvh
CiWs3bPo1n8ZYoVpYIcmSKlDtfiX4nYXqNv6g23x1t/LSNM8HQkTXraX+70YrT+WyreYQ3cUhl5b
MqMkEjp0CklaA2uhuIpyXIiLE3CtgwNGaMbUjvoinhGwkNkEvobXf4ckyoWis8muoZ6OjHwJcgxm
22qRP3SlSlt9cI6f8XRG2V2CIqpbRdSvWoLSEHbK9LiCK9MfDvHKT4EQQBb7r1OEUiOJS7B0iNf3
NKsdz8j4C2hRlUVZWNHwPt2APLxP2iiJFSd6ksqSLzRuh2VWZCBJZEvjA+PecTGIpMD8VjL2u8F2
/aLrH0TvdxG+S71BySAvX0bst54eBTRL+tOIVYAIXgZRA6ajnGdZRfWYzPDLt9GTX/i3rjOvdunF
cqqMjYhAQNp1WCObZlMrAWz0YIYzLl4IJ6apDuWh3HNM6CMypJ/nWaSwC+VnNpt+9ljanDNnQuk3
WiVQ/Zje3x6HUtgy1p3HvLX28YdnXYlU+Hy6sme95O+WQPDFgYsEcXvekhT6hiKCtSntg21v3Qa8
Y8cSn2zV26bVP4iTkF+CsDqY7UcgMPV/47o4V18r4Cojq7e8H0jssTMVNh6UCFQqcCfVhuc3AKDT
tEemXRs9qgJef4HQhizVPaPxJLR568EDuuBd+nVohBShl3IDXdK4cNxDmqrMH6ksrXShqaHYCWBr
uU8Tk7owafae8txuQqduVuKb2dI0D19RFf3jbALlsmrxWthcfTl9YhnyExkQD0pQxwCKP6zejIfx
6UzcQrPbIkTEzHG1BGYAlmZUbc+nn76W1kYGXUyEoMgDIdZF+gAGitqa9GaRxaHgoyWlbkzzm4Mc
nmS3lyG1Ig+ZGNCj6+gukWzFMftLfovi20XYsAyFLQsQz5lGeumkjUKAvWPw3l1RNQxEuc2vWRr5
dKmUI0r2ASKnPLkf8bnjadSxmN3yst8KTLgbhZLGjLUg0+pODqb0x7d8rblJHAkuztd7uugayTh/
defv+okwejKANbZ+wAy7NZMm4zuu3UGvFBpEpEpTe4ZCR04ls2R4bc8/qq2JXT6egjHr627Kv2wo
ZMTcbSj310LLD2Hya0Ga7pbH+ehp/vTQIvZmr5lG37PGTqM4q/jIHUkCCq+NX+ub8n5cugyVZQEK
5CaPeVf3zKScHcrZuwjQ8X1pFyFavszaesnvcMHYARcU/D7ZAOu3l0+QGSSe/A7irW/aG8IoydCZ
2wv8gHUK4efxGOEwSn/zwpVm3nhW99aCSbFeUQKm/MY2Tr+pZEu19QaYCdI+30HI/YsrDtm5t2T9
bTaSWKr4qaKfsn/82Lbw2DwEKZcw4G4EBjtud1uxEa0RzCNwXXNLFbiuUGJkoBgFd7u9J187eish
v5vwOpHZSjqD1HkFRkUa9kSyUD5T8+7zEUROrB41R+2dAev2W9TxvDkxOo24YvqffTiGchGQC/an
Vg5AWtLFkZpnvWbSXRKhgFkmC/untOwIkLjYySzNvmhDSPkrj9qk0xB/Fh6UsWKyj1Tg8SrZo7J9
4238m2oQd2wKLDb+X6K4iLQRIbJnLCouzCcmUmy/1mW2KhiyAHZO/wrxWH23w4GYU8SFVHYNgOH4
LZoTFqBjs2vq0iV1Oj3WsceSVHjl3rOTLD4j2lirQxmgAn7NmTqSn2+NSEFssVL1uDhTXLe/WK3t
+qhlVPKmmN+sYS7HgY4flOSbRmS8AswcMWfZAJoiZWh8dCMaJ8FqShEOXrYA6YZX8iPcmIeDCYH8
mSlY1dBBAXhh8S8ZUoZ2Xc8eFiSYjfFt20bPJ5p3Cotf4yTWXr0fRWNTUsbWlt9yxBD/LHKjb8Ql
zHgrdTpE1hgPh5QZ+riJF9r0azfn5Ex/5LSTXCbBCLU133IoJGvFtH4X9BbSg6+2/RcT2KuFwrKZ
d52DO4A4e3PhCc0EtMvr09fUjYtM9BNwUO20pCIy5yVtoMeHkk3y5uA6LmPkRqhT0DR7C8LtWiiB
lZzvL+JMKU5Fhy4Th9Wf4ELX6FV2mOljYHpYV8L2oz9Tbo3aC0ibVwT5SfhTPJhraKVu2IquQ23z
nlaWrBlu9dqo806qEWD5afG5yg24FOS5tmCcAW4z1UdxYiHCnNjmzcSf4wxiLBsVsKoBR5sbD2nE
1ZXpaviaVaPxZGf/4VWHzDZ1EDgrU+RmFn8yVvqQc0Gjubq+F7Ejb3eHfXwynUpZPCzJTCvxTaXM
7aPSSYS5258z/qFzNdn6UBhccMuZBx7orXBzLi+67fWw3P5D1X9tE7totfLHmHpFnYouQxKkZOYn
Iq4Y8VmpnPJZTGtfI6KXao+4Ao8QERT5r5OHt8KPmWXtb/rp1TtOlZEQmxFajzlpSvFo4rqaB46e
zL2zxjkaF9AJmMEtu8rKxB5288tCJSHVOP1ZOxeW0NPJOFw8HmJ9HKY/N3UNbRl1ZeWCV+LVQinH
N57hLLSPGp9LctCeWJ736lBZGMLYmr/YtKJPMwfFKVN6Lc2Vi4uzE8T5I82IlhsXOs3DveYQqOW8
Wk3tQgChjpt6eU4uDhFFxxtoefe3KHsRK9pdTopjEP/kVhpDCgdKlaiiBID0a3SaXBf+63AFkvlx
E3h7xrcGEk5AMr2FJiafrcisWVAfCTB2Tji+t0sGIo/tLSsY6pR3SNE5MF6NJlQhJRTjo6NDFXkx
eDt9SVR6ERp4r3OkPpK4LFBYSaP/bUdk47VQwyhNANJFdXVTUMPJG6i2GLFdsiDibhZQMuxhKO7P
lJoE8qWqff4VIKgLwsoax10D+k9T8GOupaLzKAwLLCsM/1Xj/UyuOVCz/AbulaokCIp4mRr9V173
VYpblhcYsCd92HMh6WP5aWJ/jbpbmcDUn47p3c2J10kwcFF/eQM3PJwNjNl2XTSB/TvmE5BwYc/5
O+p9xElQlIkgBTXBYKXGc0UYGkFNtrKERj4FdicSe1DMC8/Kptab74k+xA6BfOE0FQXoSqkb0E+x
HA2O6G969mkTXMVSM+KMYzuUhWQLdzQ6o2jd3wTsjo5+xh+YeEaTLZ0+MRnhn9EpvilpOmEWJeKh
6et5Py/7vnHs5ZW9R45nfTfMiHWoTRn1kJkYxoh2Le6SRaYHrCxPEiBry14nmTubyVAK8fwEy3jM
Ni7HyOoK7D4FjE+1qvzbeOZu0M+pojvBIzXquVbvqZBlm+hl+X2aUOjzqcJKy1rI0YZiir+XZ0B9
55V6YSo0JzDNUDLQsgCW+auqluGq80AWEHNnIObScH8ZUa8PvG30S6dkN0mnf4Vra+Qouc/TOPUi
8EBjwUkcpxpTiOcHm6jcQLQqG5xQz+YIWAp/G4l+RNgMnyuDkyFgaUolbL0QR+6fg+03qk4+2atA
8XMM/ZNpYlCrL0QU7gWdLjWWinZTLAYUEF7/xnazHCEQT28S1x6/7FSYW90Jo9OQLotkVoaavtym
ETswJ5cOvFQvs44dtzPLJoNm/ar984jcTDDIti/9ys23GtucDQuFMOjarjWP1Bs8agHW9w7Rn3rj
wY5ZD8rWaggtf/FK1ODwM3ssMx9AWSt8juN/DdySe2wUzzGNWece4+zj59tvw1z8ClgxMTwcLkGd
vHTpDqPMjNoXJd6X6EfFeo+yIfJraVvvEplvWyaq25m+q+cgwtwGuacfOw1dJ9tH8AFRP3RkNFZC
WpG8vEsUU8FDFsFJTaQVrZMzLuhq1PikzgOkMJJGyzvdXWB7D6aR9ezSRHmbNDBMWCC89jWpDXVr
P6eiMI4t29wMCwHUW9T1fOt6/DCmbr6FwZBVUSpitJljhxFSGU2xYm/dmz2G9CaAaRJuuUeutoiw
phYhC9ZKsY+pJ9zJHvbiDmoDtO7XiFpJkTfA/nkktQBz2W6GInm1oYbnKSk29OLNCaMZ6ILr63EN
DeRZdr+aBRbpCfUk2H9RlKto4TLxMjbd+kUVTh9gbrGD9Yr7AVHtLWheNyzPwN00jWFRIrw8XTiT
dP0JF1dobkh6V3ioVe+Tcdd4dDHzambiR7vvoxItHtdOf62UwZFlCq136iMswJtFXGRiJTBnn4UP
aJWnLM4Zoz4IwsqHoUB1A9vzpAZiwm+r5IvgJRIBKQJTGMArSHHIgeyClikxOBcLDK27+6NLwb4x
9j7DsyR4c/cLgHt5fe/+x/s01IoBFm+jaoSALNc/pCgTj9JSVYJu8pLYzxOfxxPXtda8gxbca8Dk
8nQK28y25LgucrN3fodYM8SnaJ6sSFEXQlXrmVB43btNHN3VZUrM9xBpcA7Se7bMOaVgVHQKWALu
Uom8ee1g82uXVoppMTCHiha6pOFzIXFOo8N0vestl1zU1hfcIcJcM6YB1+RYN7Lh8mfZi0INnpH5
a7TwPHX2ev70S2n4cbSxksfkvpz3xJBs+xGez6md1OAW4FWGPgnUqWXEG+GRCNjapP8X9tPDJxSI
HUqJnBA8D242Ugk5lEHdQ4o6ZoUfgul/vQ/Ik+IKCrb9C7WA6mypNTbaFtNBsN3DnmZwWLuMuqWG
kcmW5gfr4njDilTx03j69KxswZOmy4NBbSEbAESLgLbuARudyWcmmbKrf8YEqjIp/bIVGr8lEX/R
FQRnIt87Efh69O1uw9ypUckSxO4xpyYhAD8x29G8Hb/ekrTdS+UL+0Tk8BwFd5/O/TSVlU7wMdWX
XmD/hPv5ZWJR9Jnz8wcdF7MCwvfOPWFmj4wgYE8/g6Ewe8O0ESuayh2OrstDCZ2aauY0Vf8z0SyK
lQHTkrKMPzytA8yCbpnG6eLkR3maK8ZaguP7JzknNnMWmMh852xFxlSvZvQ0W3oVEwadi/tOdQSQ
xTqmD0racd70X89qmsTx8JXM6HMN0QrVTIPH23oZNm5qi8r4ipZGCXVQl0fMAWATGQaRfDXtN0sb
3c3N6+L29KVu+wkUK/9bHC6iV1aDrNJQEt8cbr7eJdDo7V0WGgxN9kKjRF7KTWQAjf4URo9iH5iN
aP2ak79RyWvxiDcfdacU59NOUVh5diOkyG4HJ/MQ/ZXhFr/TVFa/aPKdLaPPzyM3ZYqGgEQUgxcu
x2DEd1d2ujL0NWt8WLELjhUCjFCIKD4f+00rdSpVcZLKJ0vnozM9VVKjPevhCZ2n0HU+095sZQyf
ZIFWUooLdiXHuUUsrBg1AfFAGfX+YX4XEr+yxz7n0ZR/wd4dKQ27LdslGovCVoAdSh84rhwY3XkM
02wmIspaFCFeGljoIZZhbbZMCuetyjV6YrtoKIXvZUmEiSL1QEph6LppNL1f+FYW+pJ+qzE2P09b
sbaIZNxCL+O3Mtch0OHcAzn5vYuy9USA7Z1ielW2DpBbWw+p9PprdB7NID36vNBwuGH2U6rrzZtv
FDMLA723bKoXMSeXpGTqgDZQ9clibwdR9NaCsHzEJoa86kHY6LWpyiLOk1llBu0n/gk+FZK4eHea
LZXWI4vMT/33Pyc2DD107c7Kflse2OEh+8wfhYF+UIDIWtbpMQtlgsqOiXpIALU87hs99Rc8YCoD
otOR8YFE4f+0ayB0MjFyXQ9mshtSpUP9uceiEiC1zYVRrjk0G+JlJqVfhhkneg+0uBN4gV/PLUKV
TjFvd9WT2ffqfhgVjdQhb9H02bY+ySgkykbgCi4yU7mZfSUSmUQ08xo7gnQ0TO/37FGC4AdN+P8x
Hky8fQippTw5J3JDHMw4UfS2ApEMOIdJV21IItbj/DtIu9hKHE/eRCL9JVog94N74ubDScgZ67SH
7O5RPATdq79I1bHfiy4V/b9EOz79Zaanto7sPyUDy5nZrNP6e/wfIwuYXF8c4PyrPsqVpwM9dbmb
gCDhz2m+zLwGEubo3lERLsfvjfoz/WBEHz/cUPi/1GTt6KxdCi4YzF1yTfDz4cOjnBR75IAsUWLH
G6IhG1E7QiayawwmeWYDkSfycxj62kaTOzR3veVGe80GukfTrJet/+M7QnBG7M+Dth1YE14uTDwd
4X65IEWqLxP/8eV0XFZ3Ukzwx/RYRXTXARxciH4RgnMIcXUuCnB/XttaQsypfhwEsyzsRrHuKA5q
IRsesRIZwp7aVvp5EUHhsPRl8DwpA4sE0yAnDcdUigVZgjXqKChv/aCH7b0EFvj1uWiCoVs88QXV
xGXZZQimluKCmAa3Z56tHIrJgz9QoiuA3N0X87Xyzrt9nJ5IML8OqXzM3Msk0jSDxRT6PyP3VRXY
L36HHDKJG8YBQiUvx8+Xi196lBzi1NMhSTibEpEHJ6AfC+sIBMVL9iZs5dqG69pnBmg/MOBPfGHn
6Lvy87WmPG28XW8s1t8M38Y7e40awVzAAJvLAzXmHuBTryfWjYdlAfHab4evACfxiGYuipxEFke6
iph0P4Px2eSs7HOGw8KjWE/qP3qx+pl5bvCszRFDddVjxzN8BO+58UK7tyGM0t1H71vBjW/13q9J
1oWj5ivVBlU05fnhLGGJfO62M1/2+XDq2MqBBYjSOXTLAIA5tBZ+ZuEWzdZ0EwbZNqyFhvFnOGAj
dLslXRX6f/WRV4lyfuZAhv4vps88WNDeC8QNKosLquhnC8pAKuuHjKFK+RIHYrL44egaxthsusrj
e4Gi6hq4tsWjqOmhhnt22O/mcFFZyWywocvjP7JbRjuaPQA+76WBGELMLiO7/n+GuxPRym+QRefd
OivyDDWpzS4kI8LK5e/V3HPQVGRL/VGFDDlXM1fQQFx87oAX8F7mptm5zXkKWmBg4xTjQ90cswMl
W2Bs734eKASmGpkWCzUVpTW84ohSLoSo9Q4aoaMqyKxnOUcqfp+GZKeH98Z5d86LXlshUSZkpJLz
YeXNik4dfSQeFVluK6ON5/vhdjLtGrLHFHvpyuXy52cWP5Hud6pufk9azWe+ItrDjbUWFQn7gn2T
E0PgQ2Zf53sNJDhlJ9f9MLwaRJrHM+UGUo/dfrXndpFKYuhKMGvHWLUMAJYXiIHI/802GN/zYBmC
ArvbcuyH1GZ9+LqKAHoRowyVRWNvrLiNsvge7hWgIL8oEEU3kCzPXiTr1Ut1sfVP+5j1o19YZpy/
FDGucbeFhk1dT7rMAea3gzUaZ2rG4/ZmxxEkg4jhQBgFTjSYFz03gCX9oDYuOMXDfMfeNpsbNu0y
5iaGHfE8HKvS8OtMBWKscduz+enHP/PHld9EdOyp/rAQdV1bRcw2DwBwFiD+O7dIaMfBFHZOr6Am
3bq2w1hAdhW2E5tmsWkNXKDibZXcGwy30otfj8NowYUgxningQS5qsLFS5LuIuR/YrlWqBhXmz+s
KLhUVW5WOcCeatURhxl/Rb8dlAiCSCAGoJyjGuli0KUdWqgkX/okMXp/xNpFInEf7S+4q12HfFEH
KhK0dzbg8zE6jgy4i88M87C7DlIKy89tUIf4Pa8xZ12krf9sSMaRimR0dAnVVCW8hvpJ077x+PRw
WLLPJxIPVDUoomg7dlUD8uq9Bgfp3LMvN1xnZ1JsjWfhqk7aAO51FaOZwi4rudbsXIS94wDWjzFw
Af5PsMN1I57QfzkqPwiGYymtmTP6ex7nXvvS9OtfXMVusq5XoaTJlTsFzH9cSZKegEz/3CJLInMZ
rWeIgOIwDnWPwDO02nWl3NfofnJndbJVPrIZHrkyWakCJPrPmuuSe4pGQOd9hqWA4/m1GukEjQWp
17vVpDpgOsHdVLzHrfShZY8QmmHxg2+CAfqvazHUEKmX23S4ZNGWd7+wYMbm8gO/9gWLJFeSERN8
zoSaF9mQz1EGKdGZocG2WQblycItmk04BJgFDvaLNqygFxI4x+5DygG4hYcMSJld7BOvbURUzQk1
OnkEt2RHY6C5s4MIqGq5kgTgZwEDSufMOd3qcPOKVVSUCg2fGOmatezLPVNajOXhf1bAndTq1211
yJR8DulTryI8z8RvD1rBdquGeED/KBNBw1VROshIIX996DXFw+7nTCmE/ZZ7k4g6w8VyXWDUO5ov
PXauUr0zpl+MZWaWkmmaHd9Ku138r0Oq9KYGQLZ5vwVB2/6AIZIQ/370l5r/ftz+aL+hiFM/TM0c
AWfPlNtbYa/P3YOcdClOv94gVEHwLGNsLVL1ndERByjgoI+YUYzv9ttsJuCWovZOT1CIVgCadgcW
yAzt7MsWJUQcsskAYh6VX3O/3C5az7dXvqSSJ6e0g+v5FbFYyEInZKxYM4HFZP10L166JNI7/7oz
KuG3SWCenTv2MzF8pv/ZMGNL/mRIzePGETHZprBXuSiE/LelvDzbHDOZhG2lPrRtkyCgzL1lOa4p
CofbmOnLHBi1zMXi7xg8zgbAoKtFShJdFEYIpj4uXghIYq9Qx09DlgAJVByfbCUFXSNV4sG6yaqk
ZZGalO85oTTs0eG2WQSU78d3za45JsQyth9omFcXpNas0JDrnCb4RDpS79urVZnnQJTWQtPT3jj3
393t2VbqjyTIyfAcadj1VvlQlTR83jLltrZ4KS0anhK1WsQIQ6foRe0t5PzRNdSAEkcfyWDcBx6D
fnnK54u7/OmNirlgC0rwxM63NI/QXSrl12g42rcAsz/vhdct9ykYFaMF//Iu37rVZahLBjmxIYTL
mVb6RhWkWcwztOiW0gYbdUEuJ1jE/v/ia20P2wztxuX3SYzsetrumB6+lBrSiRWacysoN1yv1nMK
RCWl0oIpX19OZ6chR9OZk19vDPhPnnwbBIyEZMj3xcbgoJ7h3tqOXahHZGOy/xx8DkJRjTb/tge7
S5gc5LFYNK3SXtYtO7aZL0S3+DjbVPPjU+REJcajR2y1aYHE26REatdVbcEjpdCeZnfOEq1LbhUo
6CK4Uoo5H3C1MvktqdvN5mVT3YYts3Q5Waqq9AlW8eGfzJ/zKXkU59OJS1BbPsLqZOfFY6WBEhkW
byO5N5eNyJFle+tGfKcGEdNqxDe8H8fMIEiOdybeEnYWuslJEvzmuGMrnWXzxCGy4YsJElUivXb+
VUEN17KvI8o/0tUKPWqdwmRxPV7GmkhglGv1wdgfy7VzkA/dJhXh/tIdVtTwQ9W7+pBJLXOGnGpC
pf3QqAZ0jJJGIiLem5PQIRoSwaNn0gX2/V5e69ueCTtMb4hu6//JCrI7nSniIUCF4ncuE0StAexn
hIQDH5wTsZo58uoCxSsGRj9Ibk0Vtfp1fCoRtQW5haLMP8dRC/PxCoiGX4o0119ijimnyeavETjr
9n0zhl3GZBsS3BNoGg2uVIHLbuyfLoaxmcogy66LrdFYemXGsMauI+dvz+HlJAUmxLmWpFDjkthz
FxnooB4ju/jhou2mBor0TDLH3n8f8jj5qjMkK/g4PpEjCGcDC8Hx9QT1rcm4q0d5pEp6vS0GZFIr
uQtuPVLogf7+jsqMObAQvx06tt6wPDWU67rjCpCO/O3L5tQaVrAcqGDzZpFpqFnwe8QCVklR9Ev4
D7aAIwwjffySOXPHqJBZ3aA0xX13YlVdJjnocdFPurx7QZ8fi76PIN3aMateC6yhIvIZpPlWDR83
ksS77FV1/z+zhcjZNMZu9qjRQay4UhT1XHl0g3K/IgchY9x8GNcn0wlF0gW4gaK5tfNH45SpdFPc
RKbcXhAy7rtYj8ALZPCgu1FT70yl/o5zr2+ta17F8+1bhLg2+hjKW8oko+KzX2Jv7SUKG8wBMcKt
vgPa3FygldLCODPvzObqOHJEnDUcKM1VHp7TW13Le3iJKYf2ZUhcRxTr1cH69nIpoKXxMqkgJrvi
DQG8Pr2Zar2MOrgzmXfybXOXp3/XFTW8+frmv+WfprQdbllcQUx3Xm0WE0eUEXT8HG8Nba8G44u2
AnAT2tA3JVtVKMP/JjF3wfvngroWMbaBQ0ANUuKSLJYDFQuLhDXa5CISWKUhHEWf/ziSbQLyo7jj
5rgtu9RBqMYbGISXPUOmHF8/dClu9QYxD3S0tPLa3JR48kijnL6xFYWtITl2S6QYyvJxzOhAtBLN
BKq32fTsdTgEQME2Vu1Ecb3AhY/taeDVGZgJ5EVdHkuw4sDZGNzqThiBfmCEYSb8pGpC5SBe4ykq
7RLAGaXyLEf7dRsp1VZShXzuNx2whGcPlLLfPZz2LGPWdLjfZARsTfrcSWzzwfWqdgAL7zRf2mBf
MHLDFZ1ju7yLxFtMSOuH4Re0ivdqbxOSgAmOYSgvCb+me3dhSbMvozsargrUwFAI/tiasCPtsttR
b2a5ItgNuC5pUFfvIL+w9cYMZQnNK1TgQU0VohJMnHfPDYkBiaZIwXCoIdm1truFXF35fXTwCesx
kJEZlKK7n7uP2ZdnqQBQTOt4eRWjwzyzHAnRlJqRQNHPf1hhYj+ILpa2vl4S83qgbA/mq52IS5uT
xCuHKG0AxY7u8rlVfYPXe/jRUJQIKUp7PNvE4kIGwmQj82RJ5YbcTCVfcVo0k4yU0gqPnBDVvnLt
yEOJeG1WXaGvtHA6ys1ZJbBLHWoWuxAMZocpYXyG8EJpmqnZXEfyW0ChwmfWiEW7e5HOwq2pW7lB
4QqVbpagNykXIjj3ou2bF4cMPbMCtZlixrvg/07uWVkcekq+t//8EiqAEblPpRW7Wf43ucVuBGzN
vNY78MSwBeBEjPzSd5gS+9twtqe5tJ4OzwjgtVxBVucHPY3+QuUA7BTgJCa0vIpZKRi756yK9Ofc
Q5JFRclhLDAPZjKxMsVSEfZksc1EIvezTtT8yfmUc6uUU3KAd9Q1eoHhwPYJDVxJ0vvshUfxr9+d
1pbFD9uLH2FDKdYbqMhVkYmU9QsxdLRN9J+vuvTm8TwDh/mxqi4fZ7pYTVmjUAXC7qpWeuTnKy1C
kZ419QTFaCqSV5CSxNGksrxCqKo6F1zOKtPr8UQpm/fcgXIg0O6pisJhaJZ9mT+x52VDqGrZhyCF
Fr4oSY6HyyfG/aRrIzmNvBT2Qrq1kb9V+Oiha+L59eAUyzj8MaHaFUNs6yO3WCEFHQGaqWJ8/wpK
FX7S9f8JX+S8M3MIHcV6fdgTrgKbodfEoHs4PdZU9XzB9U74Nuxw5C9H/eFXYsOoSw2e1tiuwzvp
jpMoeEngFaq+ASy84mdPUzZJEi3ToYiBR8fgrzSUempoboabFbo/QnVGwS7YLgEtrg2PvABmBlpk
Yg2IhTG8GB7CiSiIRiuRa/1tKcXKliZXH7yr4qHWX1/RtkGLqOzK5sXMb2HFNUlmnNsRDf//YEI0
BDcVffqQPxPGkNHW4KEk5E8Bygo3N4lxXTGN1Q2VEzO4A+b2mP6mrfFrMaLFDmTFHG6tZm/nX+wA
UM3fSE84se4XoZSQ46/ijfFpxmuUBnB5/tLwbr6qX7Z4yZszoHFF4yvaA111jm7pNAJQBg71HT9b
NQwyos3xH84dXgPeESLzCJcqmco9t9TYN0Y1k/G/OKsi8dMwir1PysKqEwsyXTaPmynvlyoQet32
KAV4oPcOyu48RQft+Pd2UMsCOFsn+b+dQsT7JElDqi7DDBA0ek7OHhyFnNi7rbA23ufYUXGSUZm1
5A7yasMd5ZPwfJlBvAxwtwj478pC6BOkLHFJembftrPAOFTo0NdtVoDydjmVfJUdYnDDxCZPD8AX
P8c/p+8iZrx9oH4es7f0s1NtA9/eSWdcZuPVbA6hP6eotA+wno8YQx6H6MR4KW+ZUr01TWXVg4iL
ELFCr/8zMV2KwhFW754mfmlkwjjNNeIJ58ZcvEzfAvc5Lr7Oncgm0pmC4u/YkL17J+tKBo5Fn2yb
maKeMEtgCUQZzqoLesG/Cg7xR4Hv1vV/Pcpbuk8euCnUQ1kOpSt5Lr7FknTNGiLdYy/ZrXgCLfZe
OeChOBAkauvlJo3MFqMXKgeuV5aANq4O6SFoWsnfTI0QUU08NTcqx+ER10L4L6a76a9NrR+icdSw
7isGnoZKSgF6yc3jKD5G8uuGrpz5dgnvX9mB3jMa0xIKXymoY6HKKHvTBkll8ee0Ia5PApUcBOzu
eGz329066iP7TuNHU8TDWWbwa+xjxk3vj6PzGy0vNbWVJo7FeQcyECIFv7Q7iEGEFVw6g4G1nhjw
yG6z5U5x5zeRB0xSnK3+RbYiw7u6vijRrIQMjpQ39gHqJMviyAVVSgQ59pLT3zcwWiNpaDGh8GBK
RLlrsMWboVKNQuf6gzRcmamuKkCyTzT8o0GKzVfxW8sb2w5r2z1V70rwDaef/denoGx0O/PemXJO
aPp0xnCIPCuTAgPXXFfSkq5e93wlsFla3xGgGjqMBlKIqBMM1Clafod4sCaapMSNvBLvZb8am8R8
/6rxrrMJJFU66+whomh3O2/4UT5I/W7iYu7lyIQvSC5UUWNkkQppg7wPliR9rv8eNVuJAylgHJZv
F3IajC0v2MCmfwQi8csF14hvCpUXTsHqft/XdqzQaKb4crqhhf1nJmiZhr/mfGu2P8M+Th4MsrIL
kC1mD654TywmaresPubdf/U9jPDUAaIU5kB5nVtDM5b70EPKUCzfGtb7prXX38m0SUvXfmIpPZEe
F4dwnUUIjy02t/o1wgUdCMfC91Q4tQl4X1md1bIlsLmJrmVtKYIxyHW8DTDx3umVT0SneDpSDhiL
eDZV999ObPNhuW4p1seEeQaox7ujnd+P24iiAwm434kPMjTyGdzXiSQjOeG7De4+2iMtXswzbE5j
Ix+JnwIbWbC+94Q7qiJ4tM5YDkOJc7Astkzkkz9szcmPe1xAzdh5nuqqQy+swtoETi8visAVAb6f
qoegUjkBpYVoyL45il4QCTcrvXAa+4/Ocf0w3wz3zz3BJ8GGwL5Y4TAynpy3pUIEvo6S11G8pwUz
7Tz/J6upaiL29iAMtsf/66alLmhnkwlimLiYfPwimNNrKjmhhcrETs9D8EQdG4wwezyKVOXVxvTz
tqtgFvBUGoGAUo4CLf48xjdc150sG8tqlo3Zam8uo0L5XGMT5jeuD9K+F2DNpKL2yUsZnzfwzhkI
2jTVhYMyRMgpj8duC50hjBZRs/w/9OsR/ByHWQNAN9DiD5bym5Zlw91aMq55NW60HvGpvpLxYQjI
cDquxu3OmHrtSuVFQS9uVsjy4tkL0r9asFa8YxDpzmdlcL06igQB8CWA+hfrVIxv3EBnnkvr4Ibt
aei4eQxjPntlLxAlLKQxmi05QiMkNDhbODO71q+DhkQl5dIGFGDIhsaXAfFRs/rksSlP3jcwUusO
Vc1ge6KhVXcjGAK0aLmHTIMLSZwhr3WNW9SQBi+KY9EmJq6MPInNw+7pUxvPOhg5Zh8t8fB62WH0
RgAG8lWUOkoBqZBHdeUxT7zs4/9SqVRZHbE5wTb09ou+Iti1v3N/Kmk3RjsYMToLs5DaVlYLMpkY
Yylly7H6cYktT35Q6IDfVyuqKvBxiffZwqya1HaciNTBrFr5qC8DI0P4WBeqoCZXSEr8IlrMDBe/
Nrl5JhfD8qGFvbQv2YOeiUQxl2zpCV3+BtmYDv0GVRkeMdyamE1gqbou5x1YyGJMIA+1JPAv/99V
4G36z13pKBUJvMU7Z+Mdbi4vpFbxYcjWsIVEu6y3u5Pt/Ig58mJiJtI9WMq7axRW2X2cOtWTP+90
Z/XokoDFOlCta5HbqE2wsqaRhOb5r36hUYLdFUz2K2T+Rfjrizi0/l6SXQmv6aVWhhf5GFK4foMy
AOqgL6umvTpJrBZ2G3cubkTHRTa+WMbtwiDctdzuz7DVrF1EKDSXqhW25Szm+lS4D1UMl1ZdHyCX
iDvtLu4iLZokriu/wFLKIWemWKVxjHLtLvtE2v8+hJf+p8a0PTT5thFOYvRy1n5Pzt68zd1Ko9ZR
GACmI59i2HBQXY8vqbrH5SMWSQhYwelX9uPICVOwm9ziL6seeHWEwazYQAD2MP/Uk8PgE03gYvv4
l0k9X6D+xjkBUZVHpZxHI/JAegTP1xG9cOXEYyXAV6cGTLAf+4k5RiSeGikMQN86x/yxHcu+QjDQ
PHCHpiY/EEd1AGExA0xOmtO/mrEfPvbf1DsMLLcwI567NznQq5NK2qX23ZTbtdXEjBmF+Ucw9IYH
nglpTHMCVoz9y/KXNf650zPlgP3MVrmmahW2EIDMmvpE/daj1WL/VeWkNQ24vopCWXpBJD57qo1w
54CvCMQ+4l9/t4mUZ75BBfk3ub2huZFDJHT8PtGJrsG0kFxbNBURmsgdG1zBptMU3vv3xHE7vkMx
Nos0GYzH1xhxkJBcvRa7NA8hWYZAZ4BQw2NYqRQDgL7WcV+xk+W85ZuBw0KBfneq31xjI6EWiLcw
7sC75esyTdr8EMEI1L2T/i9DPcUjCPPRVPoWWcSpSF8eHDr6ppsx+2ghikzrYEQeZgcYztERnNYM
YZUHE3mPPMmeEEsWubBJW92A/1PUVQG0Xfh7pdn5S5eKt4mIRki4HmD55VLQ1AWu4Sqfkudb+QvZ
gblIk7V8X8XAjohTm1WOm+o7CiyGkrWEuoN85fPA4gZNonFFo/Eew3ZJw15yP2PHYxfQ8IcEZwwD
NhFNoCKDbGxCFKFXYpf86yp5qFnz5SKbNltktAzanzK5Qwg01MoYSmgPqQOJfzhrQWJMq5RwuM4s
bYCRiv9vAcWCwm5lJjMOlblvldWTlHs2eeoBurPRROld/s4+l1AC7UrvpwKTBzDnB5he92P/YnzG
ICiECZYqmGUXZvDyw2tfVCYc/Oi4qRpY5r+Qg8JFo9oMnnX1hMB3jU+bTcQhRd+zXq1bfxlaXKQV
iP2m8aUDhtNGCi08Oj9F/KRirJ1lbd2sji2pXxF0snf6FvHqGc4UvqxcUW3frW07rUnQQaOCST0/
FcmSCGjzVM9bXjsZJoAi9aNIGFV4WMtZel0mWzc3NcY2SqR43RRYXEw9DSwOdTs5DcsZc9AUizj1
dXKKFLD61rQng7ZsIRkmY2oqKDV1cYqfLk/sZCzLprA0WqTKf7+VoMLYT2fnskfKjlmLcZEYF8Np
8flM4CRSZO76gi7iDP2LklQPKc4MESSHBmlYcFXz5S6VkQ+qmRq4jCRCZS01ukptv1oxiUq5s1FA
9Yxz1msWdhelZ4siVW23mA4cw14Wua2rt30tO7xZmzcosj/UHXHqxuScHSme252bcXq4UN4C/bEu
N0Qqx6Rl1drieh20Jm76qp8hfwqwS81I17Z07JoROKOdsQfEXiQL/IRDVvK7SQuAcuA7v0e87jfc
nhukjkIj9dZaAUseF3PCOtPK77Ul1YXojYZPo79HbFW37IsEmDxLk8/nL4Iz5/QQN8W4c19fFrK6
K4kXXD2yzRyUaM5DLOg5U93s5/BBBLBwNl8smeKBITHxcbXK7soN0mwzyWmv7b6ZJ0ICX9+4lXeJ
jpNkDig53oQvhNpkvikoHo/NVtcQjoJCFK1pQW1sRBoinrSF/9KUoXQ7z/AfgL/dGYVe95Zr5T2w
rWxZfDihckG31ssgKFmriS8+ahDdZQyxe3ZTuQP/TAgPrXgk15gsIQGZUrjVdTmcytUwqerwvXw2
swuQAukXTMizf2Lr0G7CRs8V7jmsroHTnJOlX2SHMgNcbn9/Xow1CesxR3FJWbdgpyQEwWRnorE+
5hQzFvobU/f7nxDVIwWWXtLm6kawRGOr/FNl/jGRYaDIraGRtG8kmXI9kyHI1KnTIVgXQrJUqA47
BpQDzQgyie0Nza+33jXDQL1MKrqOXEGBmIi/+juZhxvXuVFWWnGQRSBcd3VlfeSfgvGh41NWfsLm
Q0ExcvRRnbSknd7ujJYtoQNPFHcGC3/wjnzEM4FHAe5z0mIFgLZjQSB8CV+Slt5m442CRDiYZ7Mk
dzCU+HdUz9FackeZswLTe8KvGEkvcauamWr4t+rN+8OPbJDtnLfcEVPPWQVeTQToqu11NowPkXqy
4CaauXx//iYhEv5JRLFyYGFSJanZXlXqN8w46Y/No8VOmMugkAE8VTHDkCo4yfFhx0a9NX4qwpjh
TaYFi0Uz8uPoN5BoaNFZCExG2e5XifEdUVKa1g7xi1epqISa3OE0XBNs+O/ckysytHIjD0MHu+Se
3NhxrZtTaJFYkv1j5sQqBhgrCOfyAlGfgiPoN3b2gXhEuWM1EnDMPrcxIPdFnO6T50R52WLfvh4D
hTc8Yuk5QQNk32/jik+3tLGudgWs8CuiRGvcMNCJpoSOvKRnfDVtDOtLrcfugjU9WJ4Cwrr0ExKF
RIfy4oQSoxj/yPsAFO4sBraPwLvaCtOECMmnGsdpG1sRBv0/91dc6jgrhhh2Pw+Ib0WnrMG4SEDN
mPhy4GkhMZx4uDlMvoP8olmXy6RfxPh787oADn3s7ww5xHfTuZ2CE5ogpzgf2DeA646oO1kxYfae
UdHQYezR+bnS0OXHOSr54YXUxY8LSf747RbPFb3m0U9C4YMHBKDq2Jsw5XbSihvytaLY+LZcciSK
HzuX1hjCtcsDWoT2i3sg5lViSorgcjr41xcWLw9tC99CH0UzRJ4Hr+Ne4FBGYJ7an0HmNZcmq6jD
NLx7vUPXXBAu03U1CDbYqYhy1rHv31F8K8sApd4wEzCwm0UjmDEK+ygakfIEFkysFZqj3/Dxc+ka
1vDHCEazvG5lhutqfCt0K70+5PSo0Lb8n/kqkz+qMQO2Lt+tBbn10sxhoY6QiYavLrISHHnYURgd
rbKcJiXeUd38YzuvIgGwYzTGaXWC1lmbssHO6UdyQ8aS8kbXq3NlPUB7VKlXnZUmVc1QEm98YrYc
9vUqYqld1r3aY2NPrJk9enFUxBhoR0tcnjznCI0JaQisttqfG1NgEI6PMlBlUWgsECxErHflaTAm
FpJbUdsfW7lCQTOJ6gc+c5qdPZbp1XBH7kECSRHf3BxcEa2xW8r5jot0T1s+0zCGUKyg0uOjDQ2q
7sInM380i6sgcInpMPzMioGlzZZxbmE1C2NXpfURe3tl7N5MRzbLNF3cOZQ7qljEnluSl2tGrrqL
Xd6HSjUUAy/mYZIyBnvg3vwidE/LmGb6W4RxdaL6TI/NrAFjJLcIy5yfaE+bKRB0Dlp/44uGgtZb
oH75LRujIoJa5YDQo/jEBf9CGHz8hqw58urE3oN6XavisY/zKQXr+RHihsYtZrlHhnhG7v1KL0bB
UvZW3/EqDrn1NStZuX7D7xuhhin4L9Th/Ez1rXzEStUJwfzLdE/uTIUmmyogOjMQV3VqACm4Z8VZ
SVMf3nEZvkyTvRgiZWcQhKUocVWFI8neTsNpEZNXMqlt4A1D1seqi3SydMLXo82AHQ7Hs9yhMZGF
8FYFziDv0eomnmA19NHzqSBZZCO5yXOQH5VAi4QT7iorLxcV8LmGTxo8zX1+4rtOw0W0AowS9QJZ
jvuXoSmTiSlmKh6KfJPRSGWEkWXWM29GTgSq1byLvYJe3C2ZrNzno2FTw9N5xkrGu69wZPRUH+Cv
nrYW6bFcTbxqkRhVoT6QWINR+HY4nD37lyVQhkJRlIAHFS+hcyFMaq0VclNW5LrenkfschNOhv5H
vrUXBjmhPPH4G+6w0gYKexGb6ArbXPXJc9TAVffgWmb072rdqqJCnDrVORwJ5710YIHJp10ZJ7S6
8B5WeE/wwsUWWke54zlDd/cu9LSeFeO2tvdpy+ykiaZmdt5LafVc97UeAFTHTpfIH2myJglkaM2+
Ikdh9NZnI7o+XffTr8iS0/ffLCRcRFiVzV//Hv1gfwR2blyDt/0CEtzu2umc6gy/Wb31TyXeqNfw
dDjdsbS50DplLIUVoKHNEGTyZuWofxGtt4tuZNyAJ3B2avgwG25JuTlFu7KILXZ433r7EqwOzZ97
U1GC/rEJ+smE4wWxOI78x7AtA7oTbkbndk7zJRPHHYsd3FEfHZcVJt3ffTkBXDF+blRpwRMA5AjR
f8Kf6xqrOrhUXWbSTX8q6U389Gbc8jH6JR5NAjn/NdV3bCZ5FOliNXmhUcCa6cItBwPvWQuRZVdZ
iTEnPvbtdgDY7EodO/SgiSDVOAnR66DQS5pqkABGH9mXUPpXeWeDcoukQSFjy+Ncdbcvct8XeHda
C7fTWdhSzlsrAW4gZ6inoeeRn0bixPnMu9P9Ku/HOO0gRyZxcuxQ9lRUi725zVvVrQOLPUmpbo3d
JfvLFC07KlSJxJeFTTkJMbexk5uFO1zSun7UJIWXCvCFebCLNdWbngUs+Z7N4jWG9upR60zXOAcs
DmYrXdIMFU34FubJAIQS3ctEuSmekWyiupAl8tRikV1Zxcz0sZXhsIsyYcV3RU/84SngqMUTAfUy
Dhu7OLaGmAPuQKGQsZyTQsw2y9pr1WcNIRktZs9H4sUipNfAFB3Sxqg9/H1bfOKofKcRoudFPg1H
etLTNVNR6m5guIoFDYQViOY2oN5Pm/2WM3MUXoz3pxPktOKMPR1/2wBz7fbdSiCxw56X7dYpzUd5
9YJMpeQInSwpCxDvpRr4le3LVPWu7OnQytdiU1bnV0rVSA1q8FweEurg1QOZxgm26OBVk7KZrY4g
pTYet1Oxdf33VgkBl1aH9JLE3MM08GZTFg0/SefOuckoqJFBk934EqRrgyZu2hB2O47EFUuX93lF
4UuMT/nSGPLNiLmc/PTpgPqZ+J6s5CyMbTwV8TcQ3IHv8HNmKHLM5QqcVwvsgf5H6BPsjdJXhfmn
aaxr3Rvnks+JWa/CCvji/iB3AW3d1T1NVg6K1mszXtxhefOpwA57iPPsSKz8uUSik6207Xhi8Eq+
BW0t9xBh+Pk9+pRyH8vAfNl0BIjxEnMEG+v6Du3pdGUb4gdhfWmBncbPID/5oXKacEXi/hehMA+W
b8BYDY0yJRWEnsFkPFkj3/vqqAzYEjGIx6bjtUmDPcdbxskZS+ap55CznXLg6oAgaoG/x6kb+6Xd
OYs4dUtT0m3mtOdYKx5glJ2s9ygOaOBH3iauJbUGwM4zLZNI8yQuQTrfPyus1wtkyJwOc7uLrTXL
9gvMosEdMocqUH0FNMESc/V1jjSPXqT1w0aZ/P2yFjWuRfs9ZVCCqLRKk1FyotWiKX/UDpEZaLQ5
pgmpmF89xhIyZnLlcYOKHiitVB3GzkYliK9r3Pv8AwcnWDXInv9ffE7JhxOqFpGuVVTcFd/KkGL3
iZ7eEANhsvMJWRu/I3EPH4BW4Ym5wgzLZC8vknsEwUjzHDKGn9VFahjbgDwBoD14rO3CUlJx1Bv3
KjctKnsX86FXDj2NteBZTKWS8GOQWCPdHrwAgaSoKFRwlUzgwId1M8O3BVzIdwoud9T+1yyH7A6z
QP0DwmoBO8mL1xYyJMaHwcH4EJW+eiHDCnNvVyB4/Qd3MKqWVSSW5cG5LY9Ay1x2phLhxL9/eO0A
ji3rjY708NaYDeu/TBFL0CXWPiag6wYFXeOlb7riBkyVbI3+hWmyZCPPXm2qJKRVpG4WMc6vPU9q
WLz5bl+W0y9N2Rp1zm2Zn2GC/J7OMxa+T1EZcHwqc7LcRFcXyfyj67KBcydrPzuvsl8soS8gGiTd
OI6LBnUPMSUpZXclmugR6S95fsVc1ugwxLU/NHtFWNt/BbXkSEkZKC7JVFOydG/HNUgkz9LAApZe
xUT+QMH2fMwHRDOQkELml8b6gA2MM6qKt/y2GOSpxcIguhYyWUxG+oah2CkSew2wEPTrGUfsvFGU
/CHwugtIhHX9J/RP6Ej+2sZTEW4kYPx8+N5FPIsGWGJkejgXxQWXFyntdrzZ1KQ8KgCQmVjR0cPR
brs0lJjQGOJsmQX+Zj+vJhEEDYQlbZOzZCjMhHgk14ByoaSnDAdxvsIgKGCX6VwjYbEuYJyoVLLs
tqKCCK8/HG0ZuLAg33skoYQpU1mlHphbPhZ1409Krnp8kgNqvkbmpBnPSUZIpALXYGNPl/3YhwFB
LjRJWQA6TUOENBiKG1t6JoItj/vJ21W4JwCrl0vL/+9h5H4zyozeY0lBpDI9iBT97xCtINQHfnRq
xlDcvA172m25IatSI35srIWGN2UsCrQceEWVbCoyjSCBA1vpfkO+eGx5z2jOqk1q72h0ITb1YvEU
2MwFlyC9AGswZuCXJEUei9BwBDnvqeD09uOuv2CSuyZ1pHayyGHsZS83MBiR0bj6V21qKaomRoZI
/BOZ4tnuNRGiXAgYusnhodX5dzcyhQpG3Khxo3jzO8rIWYDV/EzR0NY++j/7uM32Ao+hax0l3xbS
O8EgoWcg6ql5JBCtnYjpvMpTLaVEBtvgarbQSWunj3jF1Qx2/M9p0cH82opIjJya4NJaEXZP7bCU
qqKhqNofKQ42I9MPay4is/bGbEfoyW/MTwFCj8SNboU1rXD7LHVLr/27JB+98I3G8bJXNHaByeX/
QeTs/ZoU/j26ee2Y7SbsiVQhU7x+hRA4hIDSRQX1sitkKGwJBTuVE2ilf0RDClbwhQ1WjCPSdu57
z8NVuj/I29DRM///39WmWpOab7FZhN97wRcZ0xo2TpBxbgcvij5j+pCroyz0yv+kw8ZgK3EzxGtC
HSjTD5Tt3Y5mGWXZaTShwv917Nr0aTSO3lxAp4CpqOu4Gpa/0TlIkF5jGYwJcz8pe0JKQczXdTPq
5XRl5SJXe1uw3GIn5wc4xepvAfoH3fI78i6DyDqQsIolX2D5ZUtntpBqU2I2YJma6cPBAZ5jyvFp
o2J8vmaZz6xdke14oi1M8cvMyWfAOlf6NewGqZMR/sFmX5uWyQ4H20n0SmsUm83xCQrV97V+heDm
PX1KyFpKLmo/P+P/cWQECD5B+XU9uXBQanzA5Ox1HoZZ+9lCJHQvFQqv/wvtP+bMehWo0B58NOTq
vCw3pxnJZst3ZPab2nbUHsGcSUJyr0OmnW46CqT1z1pCw3JGeahSvlwbqF2vt1ZuC2godIOo7pdI
LhmF2PVZ1zbvCYxUiHoBOwXZM1TiMtCbSgWrB4jsflCdQvMiFEeoRVDLxl45l8sbFvQ5JIPUlDfc
A5SSA1UjEDlVyeLu12ZSp/05socOrZvOjt1YneTPleW0X0+Hbb3y0gV5JcFFiec45oX+B9ves7SB
WJ5f4Q/dqgBfkb6YIq8OAWyCsAQnQB/0trrJCTs2Ian8bZR90rvrtB9XvNjr9c+yJw0Q2j4dtS4s
KKpQ9mj1mgyFX8a69Lf+mrFdK2E37Z/16bQSiBGXsRpF3FUjyAn35wT+XdO1tLfRfUv+M/+i9FwN
eB+iusqVHNXP/pWcEvnScb1Y682E8EHSsh3tAHvJ2wjHcE5pkHfj6Sd6fQ9MHDBbROy7TFlscc2a
C68mVcmbog5cpuWMuSX4e6ey7aHEGH8O6C8JClftx1QxWJfi0/4qjwKRgymkCKd2W0RlPLalOgj9
M7UYUEFA16SjkOsu2QuSktrZKUfqRs3brPDBGp6kWuTHnrXrh5Gf0zMLjqC2PJPTc3iJweI4fBXy
LRtEOsj9mr0ZwD6tSqQM4VNuCROJH1BkUemk6dPNTBlL5k2ktOUi97K/My2rwWPUOUQ9thN2JeDe
bsMFJ78lbq7CxAhoWFZp4xli8JPNyttP+QHLdj5SKJmJrdcQm0NdTr2Kej1Yo1lgkw7Rc5zhBYad
PPRHqgUUkShlLhiop2dXg0eFrQ0xGew9pZO6eDRG+Q8PZmlLrOr6XkGfwlZaLG0a128rHy1b/VX+
VQ9wsmoB1ZH8zcu1FLfvgt5FVU4aMbWd8LKeZ/tLLAM5qxseMNSgqdLqm5avdsA6yrZf/Ex4LlSs
YkWkIqjiqbcAwYuOcZw+4fmd/Rl6d7MH87Eyo6h3+TjNkad65DrehqR5bMElEMy2r/qHTAn6DQWM
rVb7YhiPGVfu/hgIJ1pFjKpCbOxaOkw8yddvJANzr+TAk1sApW3uJfI1orgehp+PGGOafz01b2d5
/bD0LAqNnFMl2iN9TeNo/aaR3XF+xaMcwfCFFVU4lMFEQNZTmdFw5FGNSo5NTLatp0wmh607Flzt
Nto791rTam6oeOAv/q+dKdsFoSrLD7IaxTwgSFRQJP4xq8oqgMjg80giHHhB1SM/lp4ye/aG+1cs
XnfNuUMKdeFIyIC33p/rm22OrGiVNipUZBzsTfKhc5ZMKIIKx1j53UxQVgmwRBFoJdzD3siBymPu
mwK8Pk87xwL3jrd5+GToql5Eie24TGbx4JmH+vdsNUZcZzpNnf6sTdTBFbgTdQMb62GezOKhzlva
EvE77MrgRa287+xjGpB4UNYUgaQQ3Feb3R6dT5Sd+7LNzeJ6j6dWysUyklWaQ2ZfgM8R6mgitOY5
VnELP55PpkBB1k7J16aOcxmq6teBPTTge13gbfmvLEyFDdbmegLJKZ7KRFLDWFm68LTZjVXh3D7d
ehGi2/g/HM0WrXln3VCE0mC6WAdd6rSdbWh21p6sum103aQJNqH0gz+Be8J27uDyDQHZqam3ygEU
aMlHv40vLCz7KF7jJ6wTeCw5+/z0Y//6Y+6p+G4gxBfwnq3UiWriFvKOB9C11IK+TejqHNm68Zga
cCCcuMuhjSuwa0stnczW3LD1aIDXtXsKgid9N6gEZOXMJKv2MbG5TiyOyZ1ezJlJzlphsvecruzg
z2C5+ymKHJLlZ7gkFknLobr0UUy9QRW+DAinxeVDYwh4WFeGlyuuJXF9VZ/elxq0r230xI5M42e2
odNe1uC732hTLryNNDGYsVm7oQCjWxCM1F+zH6gNqaLByXxJm9/Y3X/e+yNd7Ix0nuz5a02Q9/VZ
8UvWbe1AGrmbEI4S00dbUqjKhB21/fRuc4RgHT8MAAJGv/24BFv7dlL4JZ31d+SHDLI1Yg2tlas5
dx6Eu49ASCx9nTqo3eqrQLTvtrgatl98WrEU6wCMjVMMRGqJranjqvvkrM4u1wKAreY1Gg6o0I4N
80nX+viFQcdyqBJaQLFG4dgGbXDFbO2z+UlJd6avTFD2yae5U098i9jCMJrvCuWhf7wYXwAoHzb8
heiJJaodGJwnoo2zGUxxOWUMwxMVzNGRw0OqdsO0GjnL+axG8ai/SyLutKYulW9/Ap2HaVWdcX/I
grya2miBTr4F2cK5IAVQgYLXH8np4JC2T3WWMagYk270tehZeNw4O5rKNMolmfzaAM/PR0SrloCP
0hcHBos2lw+1fA1Hbz92BCAwH3soyWio7wVc7yWpbuHMJ4w6mqokTYh1r5N0GKRmMrbHTDS0H4IG
sKonttruhR8Q2/VF+9R7neFT5udGYy+AMd+c8FlwHQkA7XxWUPl/6BqZ1wxNSlsqOL1GxPumixGm
DtGS+8o2h9S21HKVToh5oghG2ZkoI6/PYyavFavtVhToJh19H3TrlKkHHohpHGk2OmPCiUm1XWnB
uQanhcfEgm/nBVB9p+5YREq9tKaC27DyPXqBzXIKwiN914OQqH78vHuf0uQqAJ0HmAlt5Zx1BuCq
0Uhfn25kE3j8UxNgF77YmEL3rc8oXOCcjgpW/K22wcIOM+ej0Ltf9Im6l0PWooCAO3PoMqxPaZo+
RNkWIgXT6kUGt5z5S++Kk4gOxAY1hrdvHUVRP/iEE/yMoH8JNau3NLRWU1yunYHHrahWT0A/OL6j
XyyFn1ZWobwWaqMwHG3BJpyCaOPxlNmZvjidEozXh9r+Q3mi49lIrOVIAsmjcXr5gbwB3a2NQAIo
c0ScHHzbU23HKRxBWNQT/ORV1RnJmmOq60gDU1jPp5OrHmbZOLc5LGNs5yHHE+5ul8pAkPhRDEOe
i8IIt/f4ApJWzmfmuFvYMxkAMN0QS4qI85Il4mVwjQGQ4MmOzQZ0sl/rTvyhbiTWNO0ori+Kkp3i
ryrW0DgoXItHWFozie7Y1PsTZEaBpFRy7mVhy5fLKotzm/LbmR9Me1kn/wC3+DEkTvZd6908NnnA
boNWV52Q3isXIgqLACT39bpeMRPAOhnCJipZb39e4NNstJqoX5AsMFDAhM02iWALB6YYFxzgnYUO
yMqbTOU4W6QfLYCQU5YOrO6PPqvNl4PupmfNuaDHDGwO03xvlEzKYCbIUF5wglM3Q2ADOJ/mukbP
XuNSQaKNQm5URDEf6+efRGqKOd51ctY4vX8pRHPPWOGd9xcENd4W10kSfLoDsdIvo4z77fUR4+tC
vyDLzoOwgCAlDtMlXB5mMxa9/MWAowfg/oT5pfWhFnaJ5uGJJT0E3ydkOREl3PyC4MNXAaYnkydd
4hAjl0uHSTsMNe/SRO2P6NZfZGVky0fWn1uyvY8/FUeFQNEx9zWYk3DhoQ+Lb7OD5Pxr9e31l0pf
bQelIxJjXrnf5pmVPySfC4iDwm5tqT96j4fX3hPrT6uKj/QY3HyeqXYH8905WPvQ+8EgFhZrfnrf
1LGQSvIwY2NpyyQyDvsPU0f5Jv5u/XjxrebzvujjCtNRPrD7EJVu0aOvD57vw4ncZWe0I1ftknXK
9V9NGYBQuwXaMb2WTWzfExop9O3kshhHjpKHMx9pMYd4GxXKcz0y+KtEJSuNe318H5nAMLpjl9zK
kWKRYPIRTMhY2ukrUMx4SUJEXzrC8Tp9lpVKz1UjvMj2x6f+MO1T0PkOTxMoqc0x8+D+l2ztheBN
M4uSIw2tL1qn5Wfe/leTDiVVmv7kdLUPfEXi+zsSMY+rSIeCXZj/8V7tjQpovs+hyhMA9pjRLCQL
tpSlLdtIMhq9I84jMD+lFbla2hSw6BoGp02N+NhNffspwN5tieCSWNPUL6+GA/u3gPAOBnqsqh1X
5xF3VY/MFdeZ6aFbHiD0jJ1atG3tHz/G+khkI7oa0Wje38TQnipVmihCyosLfMbUlirLBzp99r4D
dWOKNzDNzT6SrBOIJl6Absp6mJ2SMvB5TDAxWNmrYiWQsUCgAnSmy9qYBV+MVgUPFOhN0+yT26Q+
ofboTI10ygqvU+u9VqjJVp7/NVmUXdbHLcNBuMYHtOl0DC9KUJx/FpYr480R4B3pzzWdb0BIaz27
JC8lZjGhCBWgWqYWLUmHfSMQWREBSNUaM7WPjBzbgZboJb8/zFrXT0WJLHjAEo9KjWsoOV5R738f
2mq25n4aaYxlg1AYpJVNV6/g9ls6SgtZ/LOQsxJjnXcqhnPVABSHjyCP/FcPCDiLe/e7saMZz32G
yRIdv9KW1MvX5rUH/M60DzV/50+E5QzgB4kpP2gkebtwUbwu9s8CYmMmQKr6Hne5S8uT7U1fXRm6
qnmUAMOqFl138d483N+w6ZbxKFWYHGFnAKgvXC3g70Eh+Bd6CpAob+ZJEtnnutnv25+7qKLlKpxq
RK+xTHOhLxrIeLERfvsdo4a1EYz38HB25DmeuDu5++9TQ3HfNe8LmQSvV6uiD29WUhP0G56L4j3m
/XJmRqpxeE2kDfsMvOCFKfNq9gmtLuQwUUcROGNU5kbPVhiKyOWlIoQYPOofcsCCT4wxqm1VzNbc
k5cv5gzmOUCH6wNZS/gICbY1KeG50pP3jeEHC3QmuA+InJtW6JaBzyILHTx8NwKdqNZ+TumDE3Ea
+3f0xuAs6bJO7pVsl/gGFTCG6j7V8uXU89w7A+K0AhLcuWSXT1dn5l+N3ijEkaQJI2c1aMF8Cvcc
95sg6W9wvmuAION2wU6xBbLL1h9a4vlOUgB4odyh5FWHkILM9zUm9asPcFVjt4Un46DwOoOo+Kr2
PWVYKrUg5TWsCEwQHDwlXL+NINBMAlIcT678zFiKejqQSneXLEUW/BsbEHaNlPVozIuiESGV55lQ
r+MIfNmou5na87cgXLAc6qdFQi0b3P1vGG4ERjUWYoCWmhRHM3EVhloDZeCOuwXxci0ecI2Pp5DI
hxO2bw2POG0ES5E/SIJBAJHpnnuIIDa4Qt3MMrGUXUnqTB1b1I+9RZkxkyqGdMLBRHs0sqpwGSyP
EGctaOhqd1ieqKrOJUyLTo3LjLpZDD39HOrsVGhrAm1acIV1qYgOqqv5UaWl4H9y3qd0b7m37hXV
55i9s9CkOJS9+cA0zPJaSDHT3CcOS613d8e5pRj0U6dOillJdDAq8X+c8Co+Oob/qzqCnTrgQ19a
U3eUrd8Vlch9Y0ASbKM31y2eMfxAYpcg3TpMijiUmcivaHb40I+raXKuI/eRvabN2yNxEY9BI03k
OBR1JlLRifrZ8WVOMCeFUM3Y0xtK3l4ncuzmlzMT6OVLynW2ixk+wBCzDUC9pVwkGmc+DkO1UqGJ
dKBCePMPAX75iYsOd6+bH48gMaFbNqUHf2cFLFxvztN1B86RAwdrhAmrrVAXIa9rg+rtEguPdJfZ
VSzwveKDtdZziUp4wmCx4lUsNQ95LQTD1vgzqvK9DxW9bxQ4Bi6pgKFiPTaFQoIRdji7uyOfx3Jd
zXUp9dYTHE8trEmwkSkNG10Mo6/tyUQg36bDI+FePj8J98eRyX+OGie2mG6eyZ3HBtEtRRtGEjV5
XVJBbP1WiATw6K9lIjLkBSqk4q1JLPYciX6x/I37nhCvJVy6qn4nvsx15H7JlE64fB1ithCjFfrt
0GVCieVpekqyQE5GfVFz7QWqrvIufTDg5u4rIeJhymAWyTvNhO5MIwARGCOnFUSpEyUEAtAsuL+c
WV5O+Wfpqq+Pf/ioMJktpDTjOj6sSP816fDZVCukAB0maeMe2PYx/UkbWJYVjBLVpPw82KGus4xP
0iHL9kcn8kw4F0EVyF1/QXeX03FTB47dHRw8qjcpwRvlKXQV9ID3Twh+qV6/Fs1oMxpq/kViI5Q3
qisYgOgfqrsFboeY9i9Ra+8f4GSyF3HMX471lEi8m6xfi8+kWTz2RGDP/5F65PpYVnUR8H+OODjM
W1Vv0UbMfD0xFBIpmbfigydNEke4niKD1Yr3OU7QrGbz0zhGePOMliySy9NMM7OWeqT6bCfF09tv
ftzYQZY8R8hbqcCqW1E/rPaIm3g8ZK+4oVB1z7r7YxGicda90oSvbXsOP4wTpYgSXbsg5ivD37wZ
1pivRNx7ET55lXO+4KmIX2aiu+bDdSXWpocQ43KRSkB9TNXfTFxB+EezVLhJmIezMNyKzZPoaCYx
4p6YZhvf1Pob34q6QHQG2GFxQlRG6OfkD+q0b2ZQh7fmEhMqFrWxTfcGLrVdFEfBWU0wv17TTglY
rFzn3IzlbwebEOApjnDhyp+leHaqwhMKBOlafG/vnGZyOg6kSxs4fUu4B7VXsyZHBYzUHsDWorqq
wnpnCagwhFvpQOnfBxgR2arQyk4eqzEN9R9HgwLRjPMe/ho2DhbC1dXOuWOJSHjCyWiLqwi8576U
gfbFetf3/M9Me1IJKqEwI7nKXg9iR8Dm5iEMtLITI8J8YU+TXdI0+SYi30LVm+77LVxccbneOPKw
fvnCwvGufufBQGpi7/6mPnHjcnckjyDVpP5mOWGALRFtFeyknagHcfLuVl3lhOy42efng/TD74UK
dzYi/UIwVwCr7AUnvIPcQaIbRjxB8yi3ROGbRkePXjvENEEoqPM469njBtYB7h1Zi1A5GZlurZxB
IGUJoXm7aI+S+cGd9oAm54wWSenEUez46JMJ2Q24uBJkH12L2f2fvfzrlJq3LAkA5PBMjcEgF5EI
APksQvlc8jh3cH5KtzGaOKyJkToKno8eKiFKbLLAdB9qKzSpX5qDOCPKVeO1qW7ZF8b6+O9fI1XM
8QbByW+2Vc+J3ZCiJAoDVmH5d/5QtuldC25oStKTNC9i06ak2NrwmA0WrgUhrZsaHS6PbH/5L4BJ
FC2n2ACw9yY6IONyq6NwI7Cm6Z5WI15DbLa3NTACDogmKI2BlSvh8ClTsHIOEXjG291RpNo1I70S
gvMWL2+FnGfrWhPEa8INuFWUB+pceSJL4ZAfrwb0E1XWaZxDNYUctEDOQ1Nk+4nsw8yMRQCqAlsA
iDdqvUY29xIkLVT9DCxrIQnNpXpIanVH+3MZHDxCUuDVxhbDKM0T7wXyTmgY6vowhFzb65TuVkck
/Etzr99WMIj9UEBP//B/ve/R976Je3srEJZnX5bWPWbkFsdn568VIDrIal+augGg5alLW1TLL1aX
zaMuwzA90SU5SVN9vZxWBTBSI5vk9ZA8ZMPjFJLFrmBDaHY6kP4Bew7liaaGhFNYaEGj0tKmUvwO
z8MSJG+Jswa9KjuRKVOVfa8VzmxWrKWyHpCmPrkHxoHrSNvJ+/R5KFrMKd+ZnGVjp3x9VKo6m0mg
+PgHOTkdedDdbvvPhFQE7Z6eJ0BdOlArWu8DPM3QRTT0Ul3KZBBqxpfsFqH+AnWBM6aGeAsYXsKw
C+R4v5JF++qecy/bJQNa+uEMLfRIKWy/S1n5kzAf2fY3hwsPSzTiZk2bnziJCFRsYlLeOKeJND0U
sB9Z9hsk5zSZ1SLPyV7pxOVtGUrfD4SIgLhmT7CyQ407etavFoSFPtupdf6yCfAtHjbd353LJe4Q
+7TzeLRzlUunE7jc2O4s2l8cIurNaMo3jkj0qpRy37QfQYxMLIOaDmKbcAmSrmrBEwiqmKs3GqGg
WDnrDvBcLcMXuLMt9BhgjaEMoOPzy/ssCNKxtIX/ByFJLTDuOPAREvvlRlHHzka3Ksy4KnAngnwF
64i25x9qxdLW50LpNRSP7oh3yEyW1lvg452tJ6ZkrKGGe5g+QKx2HPdXG7Krjt+N78LpHJsbf2KV
Ycz06wnfHmZTBu1P92V9O79I4qFG/5EbWGQfyOmgXgMTZrRaSetlVdvAJD+Me5pIMGMbTNmIKcuG
6AgsrogEWEUkP54yJZV/t6ro6UPqcFXBI1p16NKfufd+U/ZZUj5iPt/z3CY7GRz6/RBZTLrL0jln
H99lbDFNC9auVT/+kkoSaylC5plSsHy6zDcmrbRG0OQ1PL37SUy4H4UoDuCrgkXOCZfUJEOL9EuR
2WIfVclHpEsA1PnBOXCvqaTFU9+G8RrEmdZajiyT3dsQRBUzHGJ+J2TX6YyRUxXpQ2XOoWyEeN5r
Bk/5iLz33CBW5+4UlXa18Y2INC7Y6vDt2R3+JuB7myEsO/cs1r8jJo/F/rdO5ghJQGFIz00caV5l
8Rn/sde5g0kAXGcKToAWUMyX8fcKz+5cHdIMBuYVMVMCg8832tQL9P1ovIKdYjRni3qDSoQlEppR
XKEva/IBaqXxiFRlU4ZyHoYDxqAsyjV8+wJc9n2nRHyoLFLZgn2PqNWqCy+o60oGdi0XZmES75bK
fTVtl649U5AwfQvYIEaGXPhvSjvWVGMCpHu1432agtsaF2BndUzEixPEZRkIVqdYzObLM4lWz/1Y
GYaFdH3XboWHRBoMspSaNeQbkSiDRYBl0u7dOpn+Yu6tW7y14XsynIoJ1ellDKSac2dGUPqmSepg
Px5F9jEC8wtMUrJu8h6+qgoCISZKtL8n14poIyBiYmCvfnt0/vIdYzz+VqiZUXYBCf2cHdiywodZ
4MzRT6ZWoGziCIUJ2CuR15qgRSXwa6ZfS72lZ0KT+EiVrVtShSv2O8w99CZhLzjLH3NOFBtIDgxU
p046Qnzoub9D4HHbTVkLkZnFWnjrXjkVxrz7cwTEcTmmMhm6wHlGvkingZ8pFYFVn+LA9dFtN2Cu
Bjaz26j3K9f5u4AVcOcq+WmozXa0lKevi9eZsEn2UoU+NirW59ZBgPVcCbZy7BZbr+/h8bOPRdNd
dcBS1hXFqtLbe9oXOT1CXCXm8o5WJwHwUGQHKw9CE6DlKI9EfLOXQB/E5uVQUxkP0ydC0Jmf2+vc
Q//30wM+o15cKgdDfqIn7ryaGwIEZLvIo7UjyPJ4jImXPi2P90jBr5kYElkjhMxnpwYinnzcQDV3
k55JwKL8H3npJ+D6Q23qV9BjkbyYWTEOhjNk0KPB+/nSVaD9PhPTqtK7aGYAEZ1ynn9nLZ4zW7t4
hTmybBCUrkg14Tni0b/QzjFxZmoJzWuZRANi1wmTizozTxhSXNbCpL4aYelE8S230anebBJfiZRs
/T8bZU8Qsg9OGSzs0of4OahfQ+xMeM5/S9avnyjDVgI/1r8sBDOh2g2HBRQ5qVuROosSq306gan3
CzffJTZ1Z6woMNy7UwKfHWjWz5gN4ZZAkyIfm1CVHpxzANXoXQXsaDXnWl++yKndpcVu+imAVL1k
717v1JFs+8LBfw9yDj6RoqM/LDtvPP9kEhswIthvjwcS/v7PbUwQPPYSyTLvgnqjWMJ/4YxgrrqZ
wCo3R6Cizdc8vgu/YuChZHkhXqCDufwjsN+SVk/XY419gB7yN70fbAFHdvmtmg/oEIn4THNyMjPY
09cthluyFtJNEfWDZicv5lNXD6U1onwZ3a0x0rs1m9Kfr2ltGBdBz4wwAO4Z0Tp8JKNIFDQX8Urj
Mb8zCRoCMz8YdRWMkEkc8/EB3Uu91me+0016SUoOSoq5vZ2KB8wuW3VW63YoeUY2qZlZT7MOikUX
cbDtqmvcpmM5tII0l37Xf9WfPHpTGD6qysJcN2YTik/uM3ZVIdeD8APRHJ3TfLykNbl+7aDPLuTp
tzY13gQBmyssGp8eN4FrmlDzHB3QYkQAWTxPyKOKVTGuAXkLJTU4QH+VLgOXqUzdmTE15FSz/RmB
1IKG2yAlE1LgNARkCn16pHredcuKl12kPPbBKm2HnjrlS7bErvYwkbLviXSrZYcM0CsqYM9BDWPc
3N1zYgTQjdKKSM7sTp2yynmeKvTG0pBc65PkDCP3ipqhRoz5VI4rvXQTLkMBYUTEGXNEsC9Q5B4T
SDjCda6BjHy+w19MufWtdDTBzUNhm2VabgXbJwe0zYJD9hXKrKm0RsPQDCBdBQHmNi9rlQr6HtG7
jmYKOTG5AZrl/gVz2sM8KcyAaYINnyhlWPV21ewvAxQvQrZKPxOhcid5B2dt2w5HY1H4OTFmwDiP
gNskJ+wcyttSQOfj60qYGnGrhFPPyY1aqZqhXJBlKvZ0F21Nn9E69K01+79Q7ywdka6ixzClNjaK
Z/H+b1hgd52q+zyrQEYlrR5hEiOpz6olC2J8aTTI0rm1XNmvaEwp0XEOymOPEUOg32Cv1fr8072K
n2NgAuZ7/WGtgG7kx6MBim5+Bz9EjpD4KWSNaScIlOkz4E/iwAE6UvBuzFubkAbdIu6LM504wRoA
E+75oRJOU20Zympkw/LQo7igBatLbJQFvTSGybSN5egieUtg/wBwpp4acvITPhP10pkGvRPYMsau
/coRrgPYBFW0PeVbRIJ7zapOaEwQi5VP/UchHUboItUSDRpSXeBxXHcDMwWZFhBh4d51MjJuvRtw
oWN1KF0J8HRvaR7yLvXvi5RTpQfdiaZBe+wXozJgUMp5Q424JjqfRHrYip77g4gLK59YhpyW7TMa
1hPRbp9deIB4pas2jg2v/3IrkbCBnJ+a8bIIpjM2aGKW9jt8MiJnYMmixSfXr1Kpmoa85PAw2tcK
QTxhqRGRXH4YAzjBZiG6IBmY4gdJdQAsUg6icsDJJaobQkhxI6hrpgVcx81lR0++5aBkC9qSxKmA
6/K1JUXgO71qNSJ9IooNIlP74tFGKtL5EEaoaR6IOimiBXCeDzb+mt/AbEq4tc57VlJlRGVT5SRm
wa+7relUymDO+CrWzb0FT3eeCizmze3n4LKJXdtEjj2hi+OHgz2BWtDtxCy9j0O2CWGImdRqY4Th
HXQAiswqVr4TVpI8LwSUvTGhkGeVfFEeH1SuDoNIX5b6RdTxmaVRjSwb/1isrT7c824dnOOzWkMG
Ox5FrmEPWulARG1x+S2lhWhWECN2IHsis5qNRfWoI3kjIv/rGLrVSOHtCNG405Y1hvT1hsujG1DL
Ce8N4YAEAI/Y4hzj1H0HYboBwfHlVcVlVp0qOX7ciJMkWvpf5htAPZWl7gDT+2UukBh52jWJwZLS
SWcT403hLsVQCxHzLzh8BYSeOTFZoPEhx162HCNQnalQ+O1Srbj4MVowsSVKsSsRV4xNTTxdXh5y
rSn7b5PpcVm1g49zJznWwAEIJqykWdBzNXR76cg5D97IASUzzSmnP6TXxAlQUO4ByK9vF8LBXsRB
9TIPus0uR19kfEMQNF0G93BA5osvlihqf6+Yln7eyAemKgEH79U3JR93rRvAte98diy3FnxQBnF7
oe3/p7DhubKNGE1f6SGPpEVRSvXIRqzCDaE2xhADtgTZpnZCujfeYy0cWIw72fmJOSjx6UWhqdH4
QBpCrZ7aKz1AQDSO1ZBEgofjyROPDjuOLaF5kKam3Yl2ClSsLpAEaiO0liwEhiqUaDiwaNeJ74zp
yAowNGS+wBBzqsQSTZAgvWcdIVDREQRPSMmPIbghmRGNFX+ld81lHDYmM54wrkrJg2RymsCV+xZ7
hKmTLKKVovffNC3Bo5oKtyt3wreIraD9Y7PFwu/d2Dg4S9OJFupQl8Tb3RQaBwWROJTM3Ou2CUNF
AfMbW3uJZXiAnYvHYjNalyl/MiTpEVQ3zT4EFKTPAD0SyPdXxzgN13TXxcz63XYtp9AHLkk7vwa2
jTK3WphvnKbV5wETjvFSCTuRJn5kjcpTeB7WmKd1MZgQ5kBiAfCn9OP6ZmRRlRKdaY7syJ20lUQc
AZKkPpvT0IszrD+72YQ0ONUftBY0R6yhMDKqdOW/95D89iY5eQZDspwUpNnvqj2xR4ru+fNLKxAv
G+C26wCu49baVHV6apk2SQJ9peq7QAPGMH2A9R5MSSyzeRLoOQWcRlB7Ba/uY88+ioXoUAAKQV5j
02lJ45tU9uwCeBtMnzlJAr7b5r3F1UvB93WbhTwibRaDAI+SPwPvObKPrTUv6g8Mll15mYZUVD3t
CuBgVa6Hmx7rzCRED3aBfVusWx7ihnQer4SH4cyyljJAbxtmarRxkliogVwbvt2fW0tH9i4ckmHe
TIT/WpKnQg4IKYva3P2p+BRcnZzdYPtXfIDOTtTTjjtL2xC6CXiAJ+WoKq9ebdX08tD/PyD0m3pF
fNMM0rUBVoIXsY4OogZ+inR45vWBXkJ6yv4IRdXCWsRl8wUvPegWr1ZjKclErDAk/7h+np+p1h/h
vg6xIsia/6rk2M4oD4KhqlWeqm93e3WKXCFrhYMbRsywoT/0l/HAKaM1NRXQFnpgHf5lg4WZ+Bpr
ko79Rk0GJHu10za6oz3nlNGYYlButqAmee9/C6HN1ZqhvzlB5Sg2kK4TQ/Z75bb9CVpD95HOdrUq
K1A9YacPXOfGAu1rBT+XV2TDyL9wrgwla857+LVixkzNs753yt1eNWbEekI0XHo9XDaUV2H5Spku
D1ARqoE7iGWaX9BpdZbDLHAdPyRtXvQfxKgT7HehW4MIaOaAjme/hBC96lpA4s07IERuS9SmWvPr
6M4a2z62gw+nS5O0fusyFWC9MCL++IK1OVGp6LeJwf9KjuJumGxCsWpYDFjt8ngFo89RwNUwuq3w
TmMjY6GaKY3fHb5tiUVVfekYjj8w7pTSruQL4GD6o7MbhpM7ABKlrfO4SFlfKlp6zT8bJsH+Yriy
F8+KWC11Xjrw62wnNcy0bTw3DnTKMELBVyrJTCqSlOYwttwg/UHD12WtKv6tMA8zVy5jKBp+wiEc
HB+ucCSSo3T4Pr+AC5CJRkZTZAtjfhiI5K3YIXBouETna8Ly4GXoMl/yShpql62RIaERRtjeV9uv
RFBWyMVEe648t7TozhW0nvP9Wo5kqe6cbI+RsKVcDAnyETvPGXc1wCL6K+nlrf+HPr07ipwatum6
1DsdjWqgOa3oeGG+heFawFtE0NvLvXGC9UMh84PCLeehoXKH722YJMq296tUSn4MbdjKLKMLjFpn
O+yUugW08NGN2HYwka6GHdofnIgoAvMG0SFB2ibR+Bb818dSx/CCxJM91dwAe4+Ryo8H6Dq8ivBv
1KiVRwLpOnL03GfJFHvfa1ip1YEMAXU3ScODPIVwKPQJIE2yzr7AZNO92XuZyd3p9el8L/k+9fDt
cMcXm6/HuQoSCVYNSytjns0GfsJtj2FRNHpXgt4Yidx0ukd3JhXqgjvrDHdJoBlf2KTVVWb5T52C
ybDdD6WiYcoLptcnVUrZ3n8ZWCSLH9J+B25uFwa1MfZpszwsdIJlbbY4kVGYwogq6nq0nSMBuzwu
8nuk9jTQovJ47RobGW7tiUJAfmO99SK494x0uXB+wb8JVdHIZnuZJMzpMLe5MZogdnOT92AYKEs2
TT/+ONJAzlXDxmP5E5VVit+WGebE5uwsBfULAwnwNDINqV3iZEF+mbdruxWMfC9mgVN+WoVCGwps
UnR1kH5wbqYfwYoDHiP5zxJSroCJS2niZmk/orQSatjk4HWGxJZD+DSextLQb702xRxrks1+6/9j
vY/SPKhCqu3Jnj7sdpXTyRKsaNCB3uNj8KO6fxBdBsD8PeLGgRtv9XvDNKRoAgnPZrYWjwwkGDFR
lxTA3oFTVbuGQsdcLxhZUpUpgYal3s0n8n7+qGnkVIxtRxZdWePjnZpq1at8UwcO+0BbtzKefg89
mD5FE/7Myv/rDvMwhMTY412mkgF0avxoPTawIczkuy+sBzoftrPYftRw/5BmfiyN36ul5+Y4YFSe
DxwIKDFnK6G423lkIN8WH+JY/q10HDdAM6SP9ZBwgIzT6GhvKB25n8sRu4QGXKfe9eyn4YtRRq6j
rBtcxZNtQaeqkOWLtngR7jQLDjDypS07z9UF88FXc550VV+SqTcAdLhwqn+uivz2JgzG5XfdzOlJ
syS5vmHLYlq6s3jTd+MfYnQKdsYRtMN6DvLCOvQK+DDVus2LalFhTw6BXr+Jm+JAFrMTyTWZAkKq
wAhtJW1kepPjvCD8LQ/O7Pb/8cDe/504Uo5AHMqm69BeU7iT0tZqDbT5lBOnAYs9WAh2fci8EJTt
R6U21XnaaF4fZJc1DSq1+MWJ1vK7OhWY1kGiPuPJjiOZeW17ecQH2vkeotaGon0bqHdnzYSmu698
MMZXnGmb9Do9diCS4BrR/UopB7OjVq5rqcKd1vTNzakhE7wlNp99LzKzVh9Cf6XZlm4Z+IYTu6/A
w7JcAjlbCKTcBFq42DqAt3kFI72vPPF7fCI5wItYxFMl/3OowSXPiD2SEFriUnJC+QlI2MLBI4hj
witCTtfdnWm6/TH9Hld+HkXY5fxG7PFBTFqI2xe0v8PDLWvLVWu1R2fd9viY1pXaf5IGhVTAJp3z
B9vJW3QZ36E99GfTOnAxtf8pl+E610Ps7HnIk14X9ZUsZyCmAph/kSQaCa/hdyz942ed7BflDmZl
wv1UVCZDWVI9jDs4WCT243MgrJo8TIJAkekbABZDiyAX1SHbzsBkBWWZNv938REgw2Xx6CIkBhb9
1uhXtIP2P8M4sP5IDA5z8Mhkmp+FpcLRtD1TBRc3KPFhYou836cuhF66qz+poso4ra8UKgXO3YCm
yIm8nUCju5vw9Cm9NjsZrwuJ5sZrCCvl7D2yykxf7h3V5dzJuR8ERDNLS2lctnRhrsDzgAxSb/in
P+5Oc3RguE7SRGK7cckn/WECJ0YS6FLoPkf1SuH1SIIzTgRmQT+hEK33Fd/7Jfnifh1TTGgFY63N
XBY47bhV8ynHxOiExDQKgWdbzrrBIN/9ZeO7IXXvi6KfSyg0Vm+aPbGT+SS1DUNjqrKMyXU6pkRe
UR45ObVuhXPtPt3x32o4rOxe1m4OoxrRJrgqrHLos32WKdL/fOjzLTQucScB3iw6XN4TJNS2Y1aY
ubl5OfD7BLEFKgBYy0+HEdUPM9RYtI2TA2Bm5AiSQ0aqvtfbZeOt3AiYjL2N5O+oOviJ/pjhNDag
Wfgt0mTFD2lQ31AL65QIrDxdFbUWfxtLlKDFREjO3mOyRRND88cjiGFzFHN7CmVy3gW4yiR8UkPF
6u6Ruyx21IxCA16IWETZX8Iyd9J/BddRBaqxs3YbeSumI88D0jWPxUsVgMjp1LMuqxms9C5mKDg/
NmUgyZlE0196qwjEfYS+weJxbepfJWXkNor7v6lIQMZOPswcOJ/NzLXm3tDs4TXWjnSleAQdQJKs
NSojswBlER19Eu2sIiUq1JuybYyBTcpe2hWJbR82rkCx1d9/dN0Q7hXTEbI4AgoXUaKpQJxCY+XS
7nIA0yuPVcQeBTqlnC7QR3YGGIODtQgQaNYoqeH3rgfZKHRqlVbZxWQ2pOIk7ia1bfz8FO3rILPi
+f727Lyeho8oN4nPfBtfq2Y6OoxYfBLurlRMTwe/n6YLDD9ZEKbviu6XeyDtXg5/MVgH/DfmwNjA
ftoPrQXAkrdJkgrfU9d26kDuWI72djBu4QqV3pENbDRCmo2lSmF/KtDC7FHgJ0h74RW1He4XemQt
8tEh3NprIFtNSQ97yu+sqkG0ltLV02ZF6a0A8Ez082UDGP1CoZi2IX1NO6ZV9a/a6DrPPOxvXuhe
/gCVbFxgYvjueX5yeJLSx5b/p/MFl25k1xjpnDksthhUhiThzEVIQ9ouOfa32DB2lbLUz1mFmrOd
kjQuj8SXaTdbIebko93EcV0UM056Z9UWRMxMbrVy9z3EN3RrwQmKmuRLbfY98T6iigitEhy+Jo5h
5Cc/mCR+o+1WeMzoocATDllhCd+VYHy68sLQQJvjqd89ibjVjVzyQ1rgez05VAvacvM8+p9cylWz
COutjtmuNulFLIvu+t86T0AQ5oT4z9jdth3S8wum/R0AJrZ3WKgqFypHq6oK90jyo9Vudm2feTM+
lH5tj/TFvjvLCFZfcUhP/sUC05XKHUUjGr9+4a4WT+xruHq4VZ6aQjSb1s+93c1V91d3aa+ek1Qp
jI+bx8LQwwuqp3ew25mOLEzLwt4le9UMioFPP6csh/2k4sK2PzAxM3TC40aa1kCAZhvuzSKCcKaw
cQNwqxpSoihKjyr4DYlH7RLvNwFsI+HdljAlo5OubQgRcQtBl6COt9airqcn1tSQnuVJuGZuzL47
jy0nnMyXMS5HtaE7lFiKI/Su2hZx8AZ9X8jSoqpNvhDL6Z6iFqztGPfXADyhceEiuJv/h+8331LX
EpROCOTv1xxjhY8hMdClxkBrL5gyr9t9P/QRrxj3mqp3jQrWUaypnyFWr6zS/EbgFqhmWVqL7TJX
jclMqnfZi9hXWD+xSUULSCFs6s1/SIr+rh8ZIR4O7x+SheqyMTrTK6tdOlnOaimOSULvtOWPuOCo
B2W74V5wI+m4yjLELTRH0Wiue1zkXx0Qx+JtEB6+hNg84qoTslwMpw3BB+J703OGKCNe/NYl5A3i
1EtQjpM4BWzen0DQSo/5agFLc52Z1e/80BU6iRlNPpWWt0lg75jb59ml4urT8Wuj9q7aDL/nvec/
cPCVk0aJs0WSry+d8UJI2SX5zAkELSxCfd5Ldx7HVA3hgBZeoQpIsbz4riXuPFVwr7eZkDjN3eKI
hmyLbuRAjY8hwn3YArkxEvRjy7RIkK54VjjmjS+Iz1W6PGKf24md1e+bAYo7A98rJoSsTcJ7BnhO
CWPE+1ItNuNdMclNiJaUwd+3o+eXiQ6kF3XBJd+sP3qdRpMeAKi+2fhVTMMRI3j6rcM6OiU341rS
LEvDaPcLUsz8A3YS/0gHS3AsWfEIULeyIxTRrKUOOf2VzIAih/KalyA7Kl6q7Tdfsg5w8V42Vzoo
nuSkobWdLwFKzp1z/tHd5/e8b22KnNuMgwkSm+Seys1v/4bUVA+W9O1E4oWI13fAvT5QJlnzcEhS
zdS2XHXnLOpXVf5QR0n84WoxjgccccF0T9h7K5OlMRl9LWuiaq4FUdbRahJ3yQ8cm93MHYngztog
o6f7WrSzi6DE3pbyHPH/5sx8diDEJaeu13OBYHjaklksb8h+owrPYXzC387vTks+bpUBqzcQpPE6
RE/yyOGxVvdmZCccXp1/4ICd/ZQJeDFce4nexLwBItuzkIVRvW23GHynQgQFYGuLN9Mo0ji4nb9X
BmmybvnFo6ewUvRslmzyH14wb6yGKG7VoeQNT17ePOJYSi6tizE+RhyUUE66RKhAocNLXEDy0HLO
eGDLhbz/D3pQCZXke5+/Q0G8XuXC7ZL90xPUXx11QvpNCBBvw2/5Rvf4zffnFH/O7pFLvWXfiG3c
Rh7v7j2oqkeXK5fk4rpZodXbfWm7oXSQ5Ib9QNOfr/BjKgfAMZh6OReIsfV+x4UEfFs5N7Tlo6YI
ALrV4JpbsZDymNPbQx0rEHVCW4HJF12Ih7JG2NEdrpS5ead9dRO09Ql5AYah7MTfsQdgx6FL9lOe
xlUW2WQvLLTkSgnLS8kcdwyVbkG9v1gv3h6oF1UxdKU3ndrwm5DQ5GyRy0TGqSok5/+pNnA55YIL
QOSxMNOzCkWLFWnmrDEdwhx3dCc89Ucw9zb6XbSnbear10LKHxbi7hmg/+9OQvEaOmTDKqyRCOz7
rvgXMs85hbvSEXk+KrvsYwcWTo443mFCv69sPCb8LcNnznzks69Sc7R7tOCF+fNdX+8EMpeABF4P
4KtTyQQOUogBK+eBtFmp0Dt0LiI8KUKiFtad03aMrS1Kgs0ok/XP7dGT6cU+cWNKP6WTJN1Ao+eB
ZT0MURz6Y0S822qZQNPOAKF+hJcCTYiUBT7zUtCh8RdaDjThGaDTIpMeTh8Ad5iTfqPEWsFr33oC
23gVmpqdj5XoJvOrGccgxfL5k1dQcyYfPlBr/MYBpSAfqLSjwpp33WxQ6zPi3z+cWNgljzhYNKBo
LIIAh4bGinoGIkRjX98z6jUCN+yDENmYGcrfKFOzimpUxKN4tJBUstQes8JtkO8fJWpNpJOgiBA5
IkThxf/I9lc5oqavkyb4hxFZ8iaZY5A+ZFMZ15rln4XN0PuyEJC6r91UpK3gY+CBpSgzG9MI5X/T
lGbnhQOf2JaaBKnnY/Km7E33UREm2On57VE3x9hXe/pguq8adTGM1GNY2ZkEN1v6Wgls8AnVrNp4
UqGjz5UMMgIpClz5aDeQNbCQPdmMd32rgWWtOVaD81YyMQbp+5hu4RoDVNv+7YplijXQm12ZiAoV
LNhr0PWOi32RUNHOJC/qAiqXQo0IMGux5PLGaMWtpfV6UWXUggvvNMrq/jiNK/FElY8rWmVVwsjI
TjIY2txQWcnU0zget/wBFBpWkCz7Q44midEaN7idmcDgiRZ0ECzNOME0Reo9nh5Elm23Yj4W6gs6
ouDE28kXJs+wgvh4t/kQpXc/CBMaRzoGmWT4Q8rRlCJiLdUF0O21+pRjR9J9Mg0PUfFlgP6akLxY
WMycmI81CjNcHcuaZJK3NpC/HziY6qGv48fs2uMmd4zTe1IszP/ncMJW+537GlgaiVawDw5kJNxV
Ft/DIgFYQnnEpL3xVtsXbdUUKS//8IiGQTaX1SNUdXbvnBSTjer6p08UtXjFFLurGdSKA8xGJoiS
ghCmsQoWrgXEoDxP0qnNoLRwQ31VOMbY+ELy9S27TkE0no3XpNhfwTAUxslLYnGqKQLsAmewZKjP
/Lo8QPezWmX/SikpefpXK/F9sCQR4SWIknWxz7EiqTsydksLKpXuA4B43bMuoVSOG6bQTTHwD/g4
2Kj8nbYlA9ZzVHh2ooV9a0pDqGmhHf/WAaPypYgJdQsWK5cQhNzVJ5zxVlQ9KVO0rEj/Y5KgQrj0
jYG6jJ/Bhpn1Qf2GoZFYcVewNtKby3Y/225edgCL0+xT0RgvfGY/BFJhxXktKjJFI4wX8Y85ljY3
YPuMG/wZx6HB4MDeanAxBqQOzmwR2zaRQjiCW83+jODmq7yq/ymrxOBEChpY1lExg0wojkyMx/7e
aS24JuvymWSY00qaG4XeXdugpIG9OIA6Rr7/SU7ekF77S+nYWJVwJATi8nefRn5f6tL6eOvKojp8
LG6LuraicPCYeBhYSJyi7v4pVlRH0mj64qaIGpZoesCV5fmp+69Ez6lKBfZPpE1dGBGFJoYS63Gc
aLZCoqxXENKpdO4CfbBjsnugEtmt0rxorrvceChvIYWK0ZiSZ46wuugg6wHbCAyVpXbwm92mIBWt
J3gpsYDZ2IcM3GquhYbzNFJuRlihOBf4/PlUokyYV0b4kYFv0LXuqSp/wy0J73j9n6ZegVBpks8m
6uexaAEDJGV8mjcB7jzVAnHBTQaZFG3jQ89311ZPU/sYC4ui8N3BJC1rV1bwHb3v/aBX+dJO/5lX
jFsLPn4EUpVfZghPoNL5PYUkZvZcjJcuNUj8XgDqwVZw02twpUJrql2K8XZECBeeqMDxu0pjDjyv
iiZWn+BXvItOS+wTqoHQ7HE/iT7ONSVk78diSIAqOE1wdhM7pHXVkhfGFUbQJCLdfAzxiKo+BfwC
7ZkHitBVLym7kN963ut4wRE7AX5ky/DjpQ9hq6GXlJ9EN3KpROfMxO6PrEyPPiEhjaznm2XyOCan
PXS8YRGN4ErZYZ9dOXIgVLWof93iGlPHbCuL2opHCSPgMNfAyaME8yqUMHOs1i+b+lnGMBzk8uAy
MhzSEkgnmqKlRnx+uS1LR+Y+XcWYUmNeAzb0fTTpOEeCJbFfOBZSwoc9A0epGKItDiC444AUlAFw
YGdf+YSIpss0OZf0n5buehvDJmFo1eVmBMg41I7+XXwJNGGhtRJQahYMVO9Oj9isE3JW2pqq1EMR
PshQTRaskBpv+fR1ZmYrrCHYoD7rZN5KAdNEX9poTO4gb/AYhrmWHgoH/IkpUKtoJaQd+2ZTgQuV
VE8CTndjeTs0UubbPzOAy+uZMKJANTbt979+jeMPn0w9DSXIyPjJK3ysdyXjHVBjRwVKQ9F5lylG
KKk1Sl69n0aSrFqNnvdJVXN09r00NuQsLW9BAlNpwluT5uzM18wRiIxmBBe2O+pP+/Y92e/GKFjo
mwsg1eZtfUmXKpXdgUQEUR24wF06l+akUAf3qjZsoKerOzAJzlDGcgSmGjcTHyC5DBmAd2y6o3co
HeDL6YKqdeGYBSt3Hg9rrF57Whr3ukp52OxmSZh7Z4MG92zbsxoY2/bfae5257lvIecS+ErUUcQe
fNRMVHZqSQT0mH93y/A4pM7hnCo94TNZ9KVYnLzJ8tVERCVgQRafdi+w5heUJFib0tyY0Vu/1tqJ
uY0Se21cZSWKJz9vNFJb2/+bensjy6oM5BKN4iNeY3pBYIGPb8Eyu0Di3sIS6B9PraYM4itqnKbg
KLfZhskt4g4AaMMKnIsjQdmxN8ysSMSL1bPg/asrMQrx2H0pp4UanSgNd0QqxJVZAvD8TpC5gEO3
tpPBssCtXPRv5L++9s676dW3QArbn6LabUBPEvmnLkiBB3Cg1iEIMxb3DTKC13Eq91QT7X9dw/Oj
5VmSqdiZuHuFCw/HyFoPwQMAY3GwsFY9Jnac28VixWkMbAxWupI9tFblNVSk+CV7sAJaXVzZBdYC
ooY6h6o3wxM70/OeNQo4WCfLulrLni5KLrrE6RYH1KAHPidwkFffiGCEgzw5oZjDNXnENvHdK45W
iN4ZTytwyBVBwFiCyzdobj2d28pNz+20jFy4WKytG2M1uPtOS+qIw+EPE0/aKf4Bq6iVGY+o08sQ
8jHPbel5EwhADFtL71cRIOAAHrU1nD8WdQ3rBSBCtaAxdVpfxVtaSKIL7Sz2z3tAdRaPNWOfYYVC
xMill4lp8cAcU68gP1aUpqZMrZYHAAe3VZ5sE8I7DjiylXvrvLEa+K6iYMFMOuhTqOXd1Ou/IeHs
qwr1clbp3M5Z2m0YpIuhvCVD2rDarTd2pRe819uxUSoMiRhUKp9t7BTo04D0oe7tUwBBhbB6exb3
/sqmHbKH5z8k7Ew6f/O1AdD+HPm9nnU6rtWk+OLyTqwBwkbCd1XfEcsyQ+mlNDphfKkCIOFl5T9e
gsAy3aApejHKMjMfrxcV9YJ3hs1RDojX3Zl//x1I9UCVeOLH9q/POYACdudQ73y9/sns+DwNjTmt
8Fh42H9F6FZjLOwoNnKRtKK8/tj0o2/KnvqeDcoGz+DbPhwQ5elyytEs91Iby9gEocF5RdfYsjE0
j8o8mhs4etC6OduvXStbTHW+KhVi3ZbQIad1P+oj/SGsTMRau3qX0YEv0zMbk3IoCbUauun2PYaX
wRIRI5Hj96vFIRk2o5y6RpD1xMePSAfXFzXrAFdiUr8EvcmDKHYNxwtKgLxra9e8PlvNvfqc0iyQ
4MRgQUK1mlHW22hmpx4raoimH2RG/F846uvWXjHSyxdnCxvNafkZdm7Sz2/UQBFyQytb9hPDldWF
vNzp+vnaPj/KgDddvhy+NZNh0UdSe93s2pk3vfZthZdWJRBEk1pKZIF5t8fEOXVsE/R421mrDqqc
B59d9BuH7LVB1PBZpjwwFuBm5Ly0CuLcJjJ1J66C7XUr+VMlHyxkcBwZq+ChuAw0aJkcbR8VNn6n
UPlD8Ny7TkofbqcNotKeaECuoU1k/W90OFiPMpzk3HFGT7kevSAhqCihJciHI0QPnVHySbCN/mRT
DePQQtgoI6thIDCL9IRArZy3DR+NMO9BLxMSjlSj6+Dx1L80VBJMjTLnK4GOiqtzqseWreie/yuW
5AAehlLOjXPowYTeLp0rT2EHeocbNkz2qoiXuzGtyv41YvD3Hjl2cq3w7U61eE6c5eJKiiOXrsAU
m+3OjlduaoeaUWH4Q26nPVAIHIWWbpatSaJ2hXnAlnN6DA1F9X+/grzEvYQoswfMDX7Ry7nkDtr+
BpdOwinLoRJgS8i7FBmBUR7SstFazNR3hMUP1VoBuJ3QzTVsi2clGA9CObCN2tFKntFeQjK3qwm8
xNZj5RDDcNUwrW49iX88UCjnUu3r80R6NBHWS/9bSaxFbVzXDRfBRKJAItSIooofhhK1rAekmkVB
eoPyCy90XdOXQpJ7a2P1oHqbQNX53NXQScP103nH0KD41BzLYkNwKwgPr4nJaNXqD7aLqDOJi4oo
f6WvKSMAzeoYyhc67P3n9vNsilJF/EOsQASjfv90U0Kh9b9xGkNhpgaSxpwRX1s6F0MgZR3hKlKh
aowYBcuwCcmgl2Vdzn9QIvfVWSRCr2aTpYkRHl0kCVe2Kt/+pAKZ8WRz+EWdZyEF2are1ra/ExcA
HR4XG7IzcMes44DYWZjatY+e/TkM5txQUUY7e5sVzWyKLBL6ZGiXrGx2my9uQhhPjWX22+PVhvIS
EKYXVvP6Prp4Se3F80UZQlvc5pMsifZ4k48cnxFtsP4EZVKA4DA+vPRvocxS8NgiBOfFvO0xJMTh
GjhwcMbiKP0iTyzgIuj0J4XblyrWh8oleHNvCNk1CHNvTcVA4MbA7StxPXCHbicy1Ud99kfxznJC
HmXxIRAN0WO0kACx/buS4ru8cx3aIYUe2wGpZXYXuL+NnLM/lB1AT5598xA2d0fAa3cectrCpmev
q28Xeo2R1v/w5ntvMN1i0GW0hbFs491C+MIAi2etSGA3APpnF16YFOez1h+uRCSfy3L3c6Yuzyp5
KOSQ57xN6GJxmaMP5xNgwq/Fehh7hZHSk165VhViPszS9bpHgvye3DVWz//wnbZgry5OUCNVjQEm
/1osN4O4XSZWc8usgLrjuH+3suT0Umk2Wd8fWXnK1VSpTru9Ico/JjewmeQNZ2xOt+sNmiUaUz5b
S8r3KdfsEzNpForEb5uR7gkiLWh60HqAYqbB2OpI1HcO/1lg7dqDUoAYvaTBxiV9uEtbV2oEF1sH
DoaOwJ+FJRiAsAYVNEBEi1gS/1CrdTzjN4tsYWtpp9KNPLWpKGAtZj0/OkVHCL3B6/fc3kz47Q0B
W19EgzbIzVNML2GTLZuzHaprUDvFkaNoHAYX2rNStTX6fW+0dC444OFiImsxyxZFS7KOm7VU2JSC
K4EwsLF1dKX2TB3sMCFUI/7OLTt6gDRyO1PW1suAN1YUSMZJY0OEVsGUAyDljYod1waF4jQ121kS
QrzocCJlOl1NdsXSK47jQJlKwFFIAsrXgB/0uV/XQ+GzcMRcoT6ojLiqx3lAcZxjxv8SUzBtmbBJ
KlPmQmOdSwZYv72TSKw7NEX2POO7WE8rGN2TXi8ZRgej2ciFzeo2dYDcXw7uNPZNRefgc1sty/TG
tugd5JuuU1Ggj3ofYA1F3wbTaZU1me1rALI0+i0nakOyGRbuLRrShnpW+rotVdV6PAjHt7a85qLU
A6TQOsfwsPvi9m5nF5HUb2SR+Yt5GAwDX0Vo2ShEUnp0fHoewX5FCBFlHx/FWhnjV/nwjI0UYGas
BfqPTrECszvZ6vtKc80N9KAt0XYelPHqt/zqL4m75U2jF9ItZhzyGRoXTksMDxNAmPGjr0jEMYpo
Aw3Y2FvTdGCcN+S6QwjsiqxVyTFrXmhwguVKybAXz6BStYwl7Bv455AORpjoPXVjwD6LQVc62wOt
aXobaaYwVsZyt324U8FTQlEYTnNkro61dg+VSTkhZGNqpNajLBvIv7L1Q4CAjzerU7F3pPbcSQvp
bhKhjM7a5JBIVBR+tKCazZCb9FEnqQPWEZ3uw0MWvPGvNgwpMTsJYuCQEEc8Y9l1jzaYmO98IdmB
qlGN5Rl5FI06A51uD2JN31CRwi6Z4m5nYsvZcHXxcw86fTXRrT2lnbXR5cizq+H0sXszV1lR8IhC
tACWCHvxHHvzxSNH4jeufQOOPu8Z+fhWuC9Va/5puhVrEZw2gQUnpolGspaNsy5yzk4pxHpbltwo
kUDE2zjFh4ObkiwRSei5lbyHbyqDl//LWVB5216dJKBLsI+1USNWIn8ujY5odM/z1v75cLQhpCDC
eeJu4vv3WIXJ8ACch2yWumOBUFyB2JYIQ5J8TTh8KOuYUTkvfLmM9NxjYo+ma5TyWhkWnjqryp7D
kUlDRLcK4drB3ErZiPucfFaEpY0Zt2RKI9l5K/CkvuICydaxLGUycmbxLGD3vP3Zf3TPENXExn8C
kiAHDlllqXDZKSv/bredIzRwbEdeF7wtezmKdJmlUjCC3EtJEO1iXOGrUlqevooJ8Y9W0iLVOWWP
/LjSqxLpYxEAkr5f92JNwYN70n2ZvJtn4r16u/B0zbtbGiZwcqWbJzZpwiKbApTMBNV8f+BUw2S+
Ze+UgF/RZdZWjyhqeQfzRGVkjNdUK58odFoA0iNFy8ZU/dUGQ/hvBS3W2iexJU721uqHQDnK5aoO
UDbeQ0mg9OhQ7foJrecrr+wGe/xNiqNlXcjTwePPuiIXHP7QdUCEMSKWeAN33L1FnhdxZkDcf9wu
sIn04Gi4N5d/qRKQj5PqW92MSdImuJD829yL3XPw88dylweaVR/pES22aaon2YEd2GtQ44mLCceL
5YYnwYoE+oz05M6i7CLbHI6cDL8Lama/DSJBDHU6IvDQmhi1paFLkTWlInqERRpnwsAwGKzVyu1i
mhohUEK6d5IQkMdnw0QWdp5lddIPEwxCWdLrUopqZHB4+AGSBwVgCcsaG/yKJBDTNqXvWyle0N7q
9sSSpWPK6fopvPyw6KRh3ZjAJQjgs7uWprNQuQ6Hg4aBIlXvAKuqPIPKC+JT9T+sN920Zl4adYgt
ZhwcRWZCYZNcmnMUVERJGJPba38JvmXp5uktqc+ifpa42yHaJNxoE10hapbHu0f3o96DsP3IljNu
mD+maL3aoClQiIm2oumA601iqpbi3tqAQJ/nYIGyas0yYiYjVVqfnrElFp5O92mzSbVvXpM6Mesc
B6DsY/TA4YSfzPALfREWBHcQhpgfeq378XhoqmK9WadL1awXix6bpeWdxK/T++DszzwRtuNpj+Yj
pIpxnSpWwPNpchzD8NYghLrEQ07YzeojCekiAEtPPwnEWXYpiAUET8rR55qxyHh8mI42OCIkuHhg
n5oF6TmwBh8wAlS4iQgGd6CiQ6FZ4fA3NqntZzroeEkMOQS6srghO9mfX/XptisYr2Bhatu5P+pc
3Q4EJh0UjXZb+ctaZA14Hbu6siPnn2evxxl2k27BcBf9gd0qeNAyFllrgKrucC+p3nS9t5mO9IBp
fThe2wLq7+9Lixqbxj3JIX2g0CXg77i+V7tPYJtYyVekPugiLc4vPP7Y8i0vhsQAO4yqeOn1cYwZ
di5R1+x9o3KPLZMBa8DSyhn7sT5hsQnpwwVhBXxfiubugyift46Pv97O1NGjafl+dNOw2U/FQhng
pjNHEDtwjKq7wza65bYGeYFo25ixQDD9XqWfQfvaM+0WXfgvGZTFTUXKEzNFSXzMq/pAI1iFA4Wu
OeksFNeuYoN9P7ek0jdTjWKX7FXeDEaVMTlObFsQMiqSDKCMQZaMCnY+LdCR0iVlODT2N/IaGd33
LUdchW6oVxyogq4obd+ZoMT865ztZdQEZ/GxbnO2SNGeQX+ySuUghsZ6qnXILCLDrzZqRZIhhdFc
MkUkvaUTlwwlfAx46JjAm7EL9L0eZOw6BKghj16NfvpWsbWbwM0Ha2S/wtyEXW6R3OimNlUuwU5v
QO7aGCzl2+2QXUSUdSo2DWuc6wWvYL5EN53Dtfy0R//GQ8Gpo2VhJVCsiM8WNbrasfSE561bWqyD
pq+hqpoWMkGv5Ri92mM6bn1mVTzszSjdrl59t3ToBNS2efV2ETul10H2XChDoJFa8JZy1SArZqs2
SimmgVwaxHRDIlzQ2W/msWxPEb1lUjbFFyXpjftb0t3KVrsLIFA0//JlcvQk71niWEUMzofg9h30
mcJS2edc47CfwZffml0Pl/fBPrgh7pgeoGKadce9e/bdiQnkWe87tv61XHxW7h9MlVm9j8TK4Y2j
RiLndAfHpcvFSeNKu8c0La4o2+ET5m918tLAI8Bd3hrj99A/KYBmsj8m1nH/YuLE4CDOlDDdj05V
jYUxK5rA3ATV+Na58xqiiKsrxwXR6v8cHoP3p1IgpfHovqwCUdaJcYJIEGwpUpkeyUCEd/j0kf/s
Yv9hWB/XGfLacVhadYKh3JpRsymlviy/ZjXB9X9p98MZ2OQ2HqKW6TdYLc6kVUgo0kM2T9sd65Jr
CKJz8HRqiTXyBVs/ZLOuSnffSj6wRbSrthH045zjBcrL0SpodmEHlMfnar2gBw3hG1VQ8dmoKami
MF5ShHycwtMTyVEoeA8eMoW7sICplTdCYN23SAuyeI/HMhyWhRX4Tc8eD/e8lYuoipGxr5Da0L9x
HEz5utwnrdILjrH/4PTcR6AgMRqeZPZXXVL2VDxyrygXYOA6ros343BqL9PtHRcogYRXGs0znrzf
/fyRcUPz6huvxKi7bD/wxSBvbgO2iriKSHaJ0wo687bAO9d+Dl5MJOpGirmE3thkQ1JLd0Czzegm
SdobU75+MGJ83wfmdZ+7m7vwoMu3YpJJj+KsVk5VhFH+ntIXfCyU9MFDCOop1ZFOZkQW8cIU9L2k
/tWig4CiNGWEj59lyiJs2og0OG9Ek5qT2plh+ZUZQlh3HBRnW2OpLuy4gTtjSIOaqlLv1g/Bfpv6
A2S1x5LlgU3xptwbYbEpwcxTPtvxKdLYyUXNNsubQO++eOGvAPhULvCVBrW9E8wE63kvkKApqdJ7
ZIpSQukgLKSIQFZwBNY1RO1Rir50mawlfwHaKP8fdsyKXe7syfqpmR2csL0LT2zAGmZDOlLHO7Zm
cc66xrlZdwsvtvWFoF8X3OYB5uCt/MllQJWP0fwVTS3nOeQ8dxbCwUODxSdlRZpmbqW2Y9SDCvGn
VmcJ7eQLGAWvmuQWR1IPOYW6z+4IhXsNTpdCg9jNGVRKmYD20lttW2V61AOZiHO1ANx15Yw4bip0
u4V10dob7JlkkE4fAlrn+uP653HVMm/Iz9IwILi44AvTSAEVJsdjQPvElLXg136vwyBoYNodKk6i
xbbxR1K2RzuDdNi1qXqY+8dJA4t2I/PUdXFldfq+s7AhgDKHCwXtMXTvnCxKsVf2yrA8xt4fwPER
Bz2zFCswykPsuSFM4OmJNBGl7aobKDZtytqguyzZwuAAN0IOTT2fQU4ftl+jzvV2rTFzZHhhS9Nl
tEuyBjM0IVRbsuuJd1nPQdro17J8h4Ai58z8iBOcEpNI2f670DjXeg/40UDqaTFniDLhOxoSxX5K
cpQ+Buwc/inG7tZHQpfW8MFdFREpgCIPpnT/Udlg98vs4ZUyDx2pgQBwJU/9PF9zT+D0D0A1NsMn
xLpf5+pzuiuzh+IkxfUmKl8BC4TnFvGfq0iOgEAMa3bO/wOps5JvIc8AM1pPuW0taYK0YQVZvvdo
1lH5PuGGidZWbIxgwtT4rZ5tShpEcmka7l0G/CxWkKJYJJgV+AFq6vkNOY+oJU9f8U4dQwT+G6x2
5ZEtZ9rMR9ip+3yyM9+A6W7olGPIJEn4/J52Kw5hAjPIkl6x+LTUegORzpXGbAybs5OHkWdGo+0a
FYUqCNKZK3z6vKdHaU4wI5/m0wcjS59q+vIsTG6KG1B549omUyO+BqI4ypJgfghHSbqoLraGBnj2
w+cq4Hym2TzRBY5fPnwGOZAn9CHrxPbcuRkW6ZMcZWfQgjmFYkyWll+D67ztGc6ASX6F5YVqBX40
DyVOpC5U95boa+vRaDf0b5ZY5NCyXp+hJUkTNJDzmidTNmLoY7uNTB+ybbOSUW3KomlCCd7DVgYJ
WWIBfgCrnu0mXvW/b8CX4b0X+uZ5eCcG/IKi5TbUzqZkQIB6n7s5R52ql0uXjmNjM1ys9c+CmmBU
SWFjFj/8mvR6rpRl2OvycviKrgiR8oyC6jvpE1lhuetcN3XUaY8zHp1cv4FVfkxHvx8f6NULK7lP
xwJh+XqbNUQ4Pzjoy0ETCQ4S+TMjpTTg2I57tIWOSayduqcP0hx8aXOJqKd9KIdWZHVyInrEyWnq
CgVMc0/GesZ04UOtAp4fVeGoJnqEH9O7Quf8Uy7ke5+dOvq9MmGg+G+xaVoc1SBUcwJj8GlIR95S
rUpDNgT1wzsz1R8VLApxWj95mwjWVYMf6H/oL8Jxwz/l/2eGDMKt4EXnQdQ1Rn9BT+Vu6w4Tx4d2
uPEh1DejfblDWdYcqfhw8Ud1AncH6Gpo8bDTsyvKVF/ivFOVNNuXCAQ9bLieipqQP10Kx9usLvoI
qCGXhNuHdjb9eBXi43VGH1YKECjBbwZITA+f+n2y/bYZCwGdAjPtNq2sqwGtFpiqj8IoAurOhvzA
9N4dsCZ8IPeGybFcyx7vMKLYGw4Pl+ljRfia3bFy/ROkDavSPazPQpIaboiNC8yx9JaPq4LUR6zK
dVDohBVd/cJit6zorKSIl3giri/NdB/EFMbj+w5ogw9fuJ39GhKmjxsXws/Mj3nhsnDDh2MtNNpG
1nKy4SSSw3QxNA0+ot+vPkmvWjJ8iF7IoL78peR3HG5lKYf/LMatOaTTw9CHzgQSjv9WDAC5ofNo
wFYGaJMWYAVd6WkL+ZUh4Dcf3EvbrT6fr8aQjHOAEnlCnempBVXXRqAlAmt/n46mO3s60pct2ZW6
h25AHdQqtWRAcn3tfTj6p6eThoYbCT7Ks+S6Xb3EOLqXWlFTg4WA4PvxBuKzJQ1dzS/GA860/Zhj
31Jqspk6OWXennl0B2UmxQhE0o6xtJ6auX25AaxY8xAds1reDKcB9l/lZEhUw6mXDR0jVCDj074d
QHlPNUWxXSROi1g5+TCK/4mLOqzW7FF91JqCYd4ThcqVE7vb1WNHJloqTAKbJfugGsBR94d90sX0
I6slsxAQ7lCwrjgLEsUfMRdD2ny6N1QCCa8MIWD/dGqIddA98URLSdAeFmw9w42qnaEMoLHxEIiv
gsRfMdnjfZPFR3B8U1sW5v3z/I2m2I+kCDcJDRd6MATm3vXQVDeGuokHpqG0jDw4Ju2W0aNIIykO
S9pVhwz/v6RrdaKqKKlH7/AkQnwPo6mmX/Mh+XbjrT2VJMctBlADpLvdKXUSrry9y1UHIAe2Vtfc
OewduWvnT81CBVSR6RIgZMEYH2LvhYYGc2zaSWwt7/rBiYgnp8MClYkMWf+juYsS2vXcc9cYflJ3
q2KzF/MiyHk/ynYaZEj6t0sBYL9wRpZAgx7uwvpt9tJBJ6xFUkfN8Y20NPAbCj6qXqeRkATY7qnU
6MOCgz4y+NpsLF7shfECaZ4L+NJVP7o6M+p1PLtB1Ou0vcWZ7N0RAKTNx/NqGIaFKCgh//v0WadL
NLcCF/gD6+4GO7kdADMxBrsz5FvD/pCpPaQX0M45TyOEt18+LoJV5ZZnpfjNdjdFX4j9CFwoRRKo
M92xS8K2mkZx7NcsmM9oIPGpVwkZFcQY+nePERVP5Lvf0FGGnjJgtx8fuRbPI5e8H21r84ip8Fbj
CYyLSGZ4Tl7J39MDCIza14+yDptn79o4YQ437gdO3zxD+Icig++XAFkv/D4tPYE2M9ZqqkfvZDov
XAFFx3bKXwKF63re9s6bPV1qvBM1yEFC2iT8nN+fGb+V0ySIGM2IA6NxxLmoJlsTUujepkU7E2Xn
LkJbOwSJxCTYCUPoWUdLM7sg9/L1IgULPuWrMc+NwqDQ67Y3asPN75e6Mshipg2UueM9fQTQMDbL
aELHO4XWvNCjl2ENJ8Ey7RLHFkir6t2De2ip/u+/NiZCTkqP7jSbShota4ZkEC/SMV6ijwsSbNAw
S5Qb1bTSNI/IVPqF9LTm6s3B5VgUpco650SMBTNAd5I/lADTLwbsp1EL7gXmJbXz0giTbD9RdskQ
gx3LdUHQBhdcOVXTi2R0Wj/yy0zWbcRFK9/v8fgbzGtTROCohll4/M6wu+l70DYb4wQtFv21Mjv8
rShNVVoBAoHCdKOy+DQE3KhsQXP132YaFGJatDmaa3HRG5AVZ35j2rViORYF0jy+BkpLLzbZvjt1
2FjIppud+1sJyL4ki0lBbc9/xoSm5w5vdFDRcXEykZflzg4GD4jm5KXz/uCkUjz+1o4gu/MIySO9
9mzZ3TeZ7nNUFN9WidpLJp2c0SgJxWpGpKR5WAGmRDtmSJdJwQDTpS8IHIoh9SXdXAFIycHC+ieA
CtwhHCqBknCDsVR87LCftGBhi+geAt0ckPdYSyq01YCHVY/u9m6k27PWO+7Sr6FlEvuxndCtDnis
nLi0XM/FoIKIOkicR9w7TgrM3G1k/ZOwJ/c+2H31Qt8k4EniHcyOxbArRVDvn2jUaT0z31Y2b1/j
7Xj/RWxMNWMAmoU2j4L+hLBkWNw+6sIvIxzA6RwBe6mPiA7dgYPQZEGZsZ4FdyvCMejN4sZvMpO8
D0vI2xRSBihRTx7KFDfLNORiqtIYRPmpXQQSwf1xKYz7pRqClUmuNJW/rz4EYSaZ+0JEoDeaWRPu
2HnpcmXhrZ20AYBGav6uJRE5MIrUwcDjFZt88SS1KAVsZKSATfpsfbl0Z8kcH3jIJjrv+O4Wo8AJ
0jA6uJ92WuDvfKBoNQhQwtmQuke9rRFlLafHJK1gOdweKrH6Z6q4Dn5Q6FNM1KuxozdVDslBx4Am
RoFQnWAQFhlQEsi5R7pzjkfRn+UCrZmKKzBP68xV5WTBa3R7uRjWMbm9x0YLKnn51yqtzbgmvm3l
GXPnwjXb3K/5ANKzKa7KuqBdz6UdYP6dkOmxRD2d5LHEAgQZ1w2aZdkMzzLPo9IztmUzlLfQI/HE
7uPi/Vc6fz5CybeHuLdH9KWgP7nBIn91p1Ddzea90unz+5J+TAuvN7yhmjmSnErTUDWgOsbEe/bF
qrpCz/hhPyCKDF30gKU+efG09L4O/f4/ZI2Ct1Zyqxk/xEqtKpRj/OvUzkr+VSjOw9aGBICNmesS
LB+n/JSKFTUw+EXa/uMwdysPnFhhievn07YdDEPeNnT/YsQ9p6jdVZrr/1q5HBhNRnHL/q/yH7KE
xfnWq/TGi/hZ8qyM3MoZ2torloSljdxFZD4C90UV218tkybSm/Hi616WesoeudVvaGF26aaYW68H
oFxhk2HMCeTec5XlikIOhqFC7qROke61Xy8e8B5ujrXH1VQLg5zfvThidTihabBbbdneP0UX6xOa
AjFe24gTGaH+nzOVyrrKzKC0/ek7T6l82b7gho8wqh1GA7egK5OXSNRSFKs+Y5A6wtyn7SA4KD+l
eKqL8VZuweHOa3zoBy5MgUSeYB+c2m9qSHAJFfRuBbzEeGtj+eRrjvg575glULPXi9P16ugbt1QZ
PmZ49o+SGqqNijYi66RTV6URxyrFHsRlTE/kxKTxtNqkVbNTFkuxSZppKF0Kvrds3D34A3l1WO2H
RJXpLU68PiTZYnyhV6Ily6c8hvdYRBJlcpKrGhFEVsdMaiLr8aB6XIBgOp9z1iM96i7Vb9T8yy2J
b6tHBpgahQsSJtvfLuWcaRLcDG/tJOb+Ff2JcNALNuItbsx5FZXG/X70qaW/xJgDatFQnxVI+1ma
vlp0tuEWTqQjsVDiHuuCgtjyp/xBV8e0ufXYFAUlYAp0/tjXC4cKp1Sn88mwYiuSRQaXRdE4lFqh
RgLaYRYZr6WdpERsr8zSwXfUr8XCLByIQsC9dumllgIWCp3Lakj2TqZvVmrMRB40jkbaQDxovqrD
wv6SbKw8fouLyRMhH6VPRRgsDJYioj9qdniiGa6ZbgnF34bU2zufldDdND0K8j1xIz/Lor/hHQgM
eGmUhPbc2M7vWVH9dscCehqngnf0Zi4GbOinfLa4yEvjPqTNtdgVPK4juTvQX+5nwf2jbV7EQP76
gMjY6689E2hRGMg7u8c5jjUcGzZjMrO+3clbIX4ffhzdcZS0UWm7rT63SyxEWLK6MAvSTIgTi0ep
AzlbggmloJlzSpI8Jm2rM3BeS9viIlA19/Sus6zVkrp4XttmiBJcMBtZM6CV+zezFDSUYDdN2vbR
NSNNAShPusW9dwWbhJtjl4VoJH6lEfxEDSQe7Z0pWSTrq9ASbo4TOBlIOW73QDx/rNc6UDfPiK5v
gy0IlsEeYAAW6aVQf/bFqtgKE4QywyJQt/jqK2foH1tIHaMA0w90sMaZcnZzSi2cV4e/YYvdmVna
2OV5ue7ZBobivj2+YkkdWGSil110Uu3cZZPucziHaWIPIfTYP07W+I9e5tOQaViCLSZKPCHSJPlL
jdZ9W9SigwEGt2CNoQOI/5UY3fN9v9/AwSTpafxo2QuHV3Ya2P7vxHO2s/6zedwkyIaJwr7NTjFU
2FfnMcrzmBq7zzTk7ItQjIYazM5pZJ/qDM4cN9eeJktgmQzy7DMUhs3t0epuUSJBa6sBFhB7Arte
iHgiVfBC+HTfhDAI7Jhlb+VHI2soAx77jJiloJtkh6PD7OtU2InSRT4CW0W9/e8MHMa9NL44Uk13
QsQAXtX+doQ+o4suzTRWNZWXWhjYWpxXQIQjGD2Zanovdg3JscFBlzfNZw10dbhblwFWxlRZicco
GOJnuZItZSvtzAeYJaFEajL9hOooGzSSM/Yhq2vP3+FaulVA5aMNQrJKqcGUt5JREE7i+uArSs5A
lr2KXQ+8R6mOepH7FtglDW1WV+4wR/XZ2KyLCDZIZXpeVOYsGoMzX6suuGfe1u/yWOYnI5PQs5Ev
ukhShkcm+NaB+2im7Yf5qpHzXzIbNeV1JMLgxRFAv5cnWfls6GxGDqlMAZk2y97d9mDISy4bbEST
M82swB8o5XCmnyLeXZX3wKh5eq0euL0UNnMkFumK9gktgv4YIIoBxwJlvs8WQdURR8wgIYABCkwy
7zTeOQ5h/z6qYDgorZt9BzLrzNzrpbRrHBZ7qLlwUxo9Q3+IZMlT/mId+CVbbCF+Rd2QHRYwW1IH
+dRwnzJw4noRiDbWt3w1ZHsti0l9gD76g4SPm9rkN5YNfiZcWoJLAeTghz8/TbFouFATAZdQ8WIJ
FzcOP0DwWnZcG0VNwV3Sq9h0U7Wi/EGWZkqrhXk2uJLdaqRawruQU+s9c20eCIQ8fxLvulyPfggu
nz131h7ul4fpQUDxHdiqtGmRpN0//OjVgQqd2ds17Szw8yrGzPK3Wduv9nlmX1UJIt3K2MLYfne3
VWuNfvOp8cc86mFkoC2yMj5lAUuOEdY12kYjXZZq84+1Ew5C8z9yR7O3Y1lJ2UkqnYc/tRFy2W37
2Gl9Wi7eCDb7iUnXCD/LWiIWfJf3HLfXQTG6muXnXxnEwRfkBefDjHErFemlc4QPRykTua+fnirK
FgSLLp4WZiZxGUJGHhiKlOjnjKSDeyzwaC3i1aNegDkYrKYxchnUFXWFnUen8lRBPX23Hhd2JA26
kkvs5E1/lfEtx6BO/biNsR7KwItd/m/rsIyMpF8U8dix6NBoSBUxsAcQInMGevNZnOwBgzx8dNe8
MzwASw2iiftsN0HE9xhGBS1nl/wz+/k08NAF2JL+BMMOpclYSsTe2I1xwZBw0iKm2xN20Sm3hFQ+
6kpSGP4c6nZxBKQtWgJcBqJ/gFJXBvH2PKWlK7amWXP4cRY0pofSeTGZ5rngPsMHs3TbqlpCmA0A
2wLHk9VH98UoOjk9DlnOMEfggkpqgFwrm6s3V8M/mYAoMPY2jwn0EbcL9R+6Gt2Pqj7iFqpGZIYL
LnYzV88YpiTTml/Cxqx+QNzpCTyc5EshiufTWB5TR8wG7UL541XU3LNjA6oRXLu98SOhfz0MEFqr
OSgNKZV1DmjvUU05xph32Lf+zlXIAlpmdOOwc3eiD4zlTcUu7tGV58cfJ9hkAV/FwlrG2AgOMDbe
dlL4jCnK2xPJKRK45VbNHnIiRsZf6aoxOeouWvxW/Pxo/Jpl3pYAYS2AsyF6n73d3TnXFn94EBeY
A/FPxP3RsY6DSNOjfXlgJhg3/Z/N9NtzMWsMuHOmkQFkgSWxEeNOKy1AKuojZjjtYaoAZuUpYF+e
/+QkLLvfe1zAkJJJx686HDvWYWPQHxLwqbt8FnJF2JK99QHxbxHBl4pUEA46kOIp9iQKixO24xn0
I9hNZORX6uF7L/xxkTi9tSmlzGV/uQc7MlG8QE2WYmtO6pXrC+lOZxqVdmc+Bsu78Uq7HOVwATOo
rqE8zzUyrs8l31WK7yVS/iQo4Z9E8Bi2kjRmbn+HhJOwBf67i4ShrxXLG03E0mXmcqUo8Aimrbc6
W9XVJhNs55i3u2SRUReKwmGpNhs7C8bYy8pq/wtBbJdyysrPvjGbxFlkdEwvaTV0HlV1yFHApNfo
T1rn7zoEoMQUIYaLVlMee/+4uNCnZExiE2uq04Gvaf7bM4RuY8ygDBPjUUkmwGMhOglOLhcvgtcY
PUe0CIVBTfOWgUkJk0RkG+yDlj9x8Y7cAw4ZfK/L8hS40+dS/XLv7s1XNVBTt9f5o6hHU69yq7d6
atqv5hvAqZsn+D6uHvOQXBAU1lkUuGNIK/9qwlxwn3ip3619MseuqWNey5RtY+ftMy7liaCmPOmm
I3f0mlFKCyqF6f84HHVWG+b7/mvZVfF8dcxNn0A+Wc5wLR0TgPgS9qLG5sDcRhILpMITw1Xk16Cp
pndNQJlFGbdbkLVDan4L7sXZuNx+/trMlaMDn6ffzTp7DoYZ4NPuozx4UGkYbkH3lp7Z+NM9bRot
j3DLna/J+/9rRV7XYgfC7Ck0tLF8NlZ9ERabH7errcwy2DZG2o/TQHp5gNEhG1XU9pbw7AaRgmZG
3OZr8NpvhqpQW6qH4CxmtiQACEBc2ycVY0q0OYLZtLSRyU0SA2K6WNbE52aaglWP7VCKF61puNHt
WGoo5pJy7eVY9ivn1ZekzDzfZnYOMcEYkUS1p92Re2sxLw7Q/8P4uKC508jRhRcx+P+xQxpiBtv5
hXcHOycffkjC0BxXkCRNySXjJofPU+apkYT0wpIMnXIa6DnHHaK62SM237xdA9wGHulWDcjM2NWA
+/8TG1H2Nny1x1OcM+OQ5bjCV5G0q7pzWEvE0RHKDutw/1Ebc5U707WgqOAeeQtToJh6qRcK9uGp
ews4gEZ4vchAWnX5DMMPofpRgYqxYLdFZy9/UDWnYpowXjKiiInZVxht55W3kXUbFZrAOX+zX9Eh
atQLMJbQDjFRcFThws06SFRhM7vSlO6m5VpQYBS3a5Bg4iSDFI4zKrrPj9q48jSMOn6fsQkWhQim
X22v6vkjI6Li5xbBiAK06LsTW2uWluVLfz8itSGDgznMXB7FngYy5TxvVu9xPtA8S7bmWBLKxtaw
NTgwcxpKgOkR2/JUL1JgqlBri3zwlEZKNu5iO8BHo5puWKYJ4/e1ZhsoEb/bQuk8H3ui61LkgI6b
b+gV36unEwTOwZW98vs4KKx5E4D7Rc5wIgZWSG/KbZUXbITF0Wi8Rrp582zVpxjcB07e3gUWbR3M
kCNMaicIowqz8PrIuXa6Y7HPFobz6qn9TyobKAbDwm4zHSoxFMurR761qQcef0tdTPBVp5ED97s9
+rMtLryvPs4mBT9OuepkRhltGRFq8K9FljtplaPCFLxkoI6dEJoogLvZm4A+ErAnfjhrCiq1rtcv
qf2zQPh4WjYm77db19IwPsxdXJ9FyTFNRD0qnG2Nm4i7Yggkc/YTGNNxjw5DtouMDQszQ6eb+DkE
WLlR+npNO/6Xv5Q9ZV9kD/sbohP0IqKzL/qRK9+UM8QtF/CfT4TZ3a4au0bQbLtdjH/UhBiCT39v
qE3d/GQQyiHi59b5Yg0hLUtfLYsSRrTD3H/Rn1/Mm+CjvgRC1Om2cK5i9IwO0gIY57uXwJVZojeZ
JqfmHcg1GZ0uDyAfxalAEef8quttSNZWcdZsXMCioSJECJUWRdvgli/Iy4ONAN3WEQGuxaJ6atOt
R1i5spADu6/aM0FIIGyElNsrg3P5bpLQX4jLZr3tOFgjzzX8XomqiiYX6t2n7TyeQovlzy7Xj0yb
9tHwRp4t/KxcMIwx85Awn9A8SeW5h0yxwjtjpUuHNKDmNEnZkH5gYEuP4apsjNhkDviGQ/k1S8Vf
gv11spHQkefMToUWeq6GOQzYXHvXBGn6TF2Jos13rBuTneT6QtZ/vVwLuPTwp+LfiSq8tC+vJbO2
P+JC1hSxyikd3mtaUKAsSaKyX+CxclY2SvsVAzXH/Nz2tjF/YJEU4+zGdCRorbiylZ/u5Kd7Mmqp
iU+Mp7+7dTU+FCQmp8yFYef4mw5f1HCuSyRQHKyK+ZygsgRRtRclkeNX0XQTXJWLWHca2oDJtUf+
F5CIOXnL8XggKwyFemjAS6I0+iWkJofumDxAMmzUGZLT8HMpGQ12wCX8Mf3WpztbOE8zuq9Q/OFV
QsvYXQ5zzfyeiTMAv/tcHJQjdbmO94v5kN/lUmznOmDmz+NbbRhtyL8pDpMjbIml6xHXa2TAPesi
r6UOMYCRaO3kQpn49ing3peWF3JGPoFqQVANZh3KlvXJ6UHZHdDNYWtO2T/uKe4SFNa/rWECPxmg
WDEbaAHNY/f0W5AFF7cZixays1q5M9nrusBs0s0i7RaATh6XVB7hBzyNrWkXo+NsxfevFeAunq+W
95uSEceG8pkMhAdJDQta4V1kPRHvQTXxuDAPlVLrVDoA2zML9+gGhp56fmYxLgdw6cI9/ZI3ItCO
vXUDFYanVJUDYS8lURehT9mRySHgOSU9JZJl3XU2bPI/Sn3MA4yZ/kvbhu2YIpkfFQoIYlf9AVcA
tHxT434taIP5d0pt+eUQhV4tLuZNVFvT+FIg/VpN/PZYg3UYNyn/R0m/TjKEzBY2OzH2ZUPUoN++
jFYIz/yhfsfYq5FKdvZ6Jqbp7WySPawuIfeGGYEuc9HVTn+ciTkwV7xH0uLccrWfTNiqdu48roXs
pOi4gtBtJ+zA3O9R16DYLP+X1q849o51l8CkPl+U3h+Y/ksPvVYrgHeHyxUcdVcUtwx/67S1EDF4
0lZzD2VXb+dchKK6GF9pV6kv8hGRq45W7j0TWnPHHPUVYoY/Y+vkmKnJjAVFq2jtWOE5T2SrWxev
+CRBR1M0DWrcw2Yow74Xf85FiHUPWExRmlN0m2wFSlwbtO60PBBdwlqyRcERSmoHM9SrrJ5iU7bP
lN0c3YdIcjSFWFb/zI1GMQAvYd0rfJA9B2RqznhWXbN8m8WmLK8qUWMf+JoK421OOARf7YE9U66E
dmZSGrrrQTf2xTK2C4XZf+ZGBQnsueiDPEcnuD6hQ+Cg6P3s6BCRikYqtZ3xY2sFVcYTpSn9ewZm
9H0m812yn5YRYRETwVs+oY1ZKOqXO0D8h+xYnVttTEa25b5T98MUKIMfAQVtFwGSi+QRvAlw5dcG
D9RLQd9mmDEDRFvMUWv0oS57NjoAipulxswNGSdZiX2oBBYs3vTAyh5hYG0f83uuDsv6zwKEtF/r
c8k6bZedB371rZuVOzDjP/R3cqR9GXhRACC+5k6kYhzxtlgL9LL/5fdo0YHfbJzSBZPaz0STrMaA
6P2K/kpFha0+kMh2jCAdkgDudKxOjvNZ9agg7iHikammHj816jAZt7f22Q3HGJUzgsnqiVxExHO5
vqe6I7elx/u9DEdRqbtkQRUKIikOL5MeEHeXzw381PV1P72m/fsIcwpgVTrLQxjJPMF3L54+Ny9y
1g0lPbKSdju27yJrwCuSWjsQHWCZoTMJjZIoiS7ohRGfRQGgmQ5p4DtK5TB7jG4VJFww3ADYzIhT
U93tBkddiQkhTvh36ruTxmpMHZ0NHyxjZO3OwHyzk3jHjUMOb7cKXEhW8LzbR5PrPPq4z0ekNmTT
pAhTvv90mbIXGM/08+qp9ooMyb7JtXBH1hrNeUdvsdBDJLHL9IkLF3+cZSBmODl1MFTeG1yb08Li
GWYMnxkN9I2Pgar+lEyJOV4Z3wzkN27h849yuf9CeTwDZGb8t2gquE04B2Qqg1ZAfJJwY1y5K1IH
tZ0JbYLkCN//phc9J+6L/76gc3uIlAUZJMWIzjn962TL6756jt71p10jyvHwdEtrBOEvF5mhgmWP
Y+j1Q5QWRKbx6W1OoqSOgILTfCd0b51MJYDg8XdMavVUTtyy/Doyda51uGUtunkshk/Raq7Ye+DW
hXowJsiEaMe0rYCIgk6ls/Jrw5XU2MRZpCESuP/mToMyQdR3go7ZC2bE9KlZlNSjBun/1m/7r7Kb
6Fv8h8XBXA6trT8HJth8Fr4Y8rB5Y3qwE2Qtv1jCJGsnKaCefRWE5pC3VLiMIKyu79oE8YsPkmWG
yul/gVPjOQZa6txxRNVXW+DifD8S4NbdHfleA2sSF/tKev7RPZ5P+zf8xAj+FpQwWyCfHd+Y4Gr4
0M8g1p6wWW3H1v4/BJqqIS/go2O0Gtpz3jwxbKcu/8I3tdWY+V6c6PMphQwY8lmCo3KxEg8J8VQg
ZPntlTZTF4XwJrXNvH2ILQnyhHQxY5NwhVXmD8+RgjaXZpH6AiiYrKaJ8UxSf+mgY2HPnsarukhA
gMCpOvothWsLBzU91zktE44GoRppZFxcygozAFtD0qHz/Vd4mXWglm2PEKkNx6rb6Nr7Fl1oQddW
yO7IO1XaBEKrqByjrS9ca6ss0Znj4zN1QZNSjIVuV2wMkpmoA4ETlYs/o9cf/pIusg1l9GAw4WAs
K6aOey5zUM44T56I4IGQEagwDxxXPjsQgX7FU/MuxDYenHEw+jkicur+DfQMayOFsMEGqDOMmikS
QAiIVluhgXxt/M5hRr0OedQZoyaStDC76pdkCTSZJHc5rIrNtwvRmeBBry5HJjZ+X7urQ7c3rZjv
DJA9HbYL9RKimOxkXM5T3qB8woBINzMGISFNph5615ue8FvE+vN/sS50847KJ74F2G7TcwjkGB2o
xIxxz/eOny1mzCeSbTzrcPaPaw602KsuwDDqUK0f1YP0Swm48Nw36QTg+ah91FEAaLXZzs9JufA0
Ukc/WjilpENfxIGd2OxETb0+SV0YhasJoSRq4W8qufDvXLxNdWDUcI5rMbSklSzxQ5mSQvXzt9tw
wOnD3oYg6OSnYrSy2o3AW8318+6mpUCORfGPp7dTXt4T2eQtyc62flbEMt8i/9fepGxNpdAa5hAZ
T4L2rRTeAdSTNVOdiHrhz4nSUyGy6ufaW1YTNSkY0MtUDUdCtuVdj1KgKqmISUbEFpyoei4t6IbJ
NRvn5gfE0JwEZyBZBuvg6//XxVsyMtWClDA0+16J7r8B6Aa4QFmzNVSwRnyIAk/TWkDXfGS1tadQ
l/XNvqPmOuqBraItkD5ZhNrab2HNL8SUZHuKznbnp3q8yR9r6gvGAM28HrqVmQuaVfr9enbLsqly
uRtBQ4+x291tkX5sZ9DeODAiIqWqGSNXcpigz+5DC0oQAPlRlxT4hP6lB2c+JDH2Au0YGkwOXCxx
t4odWQnp1HEBjxQx2d+1qd1pwreqRpIO1AuHVkQpZn6Q6kayS0cvA3VaV2C0K6n1mvHWN2K0cL65
9tmLUkAoCwcM4Yf8LSMZRUUoCV0pDjdUuBESYkZXz/41HETUO/3pwyaZisv/BlbRCzmleSGc6wd9
gr3yQT4B7nrB0dj3j3qEgUU5scIavgJDiKkErI7mFf+MwODyqOUaAxopMkCl7pviNvZVg/wXzadW
zNh7th5FRAQmujDwagxuL3yAoaztLwvChf/8ghzncortvfT8omuvdMDk+h3AbT2qM9/0Hz4XUnmz
AEPgqdWSf3aKBFFWs2TcRFi3s+Hgo0Qyc+gH70VV2kVBCm+hvh4UY8PpfgQypfT4f21jD6R8oMGM
pURBcIIs5kgS0beve3k9wzF6vmbITeLnGJ32SRke3gCTy6jCmWi0vYPrBIluDqU0DWIh9Q85Q7lF
humxvrxf4M0LmQ78+MX/Z3ueTFOJHdKOYwgdCV0mbJzaV+GpCaF2OoVWu01bQQ5GaHGOHBWK0w+e
/o9Sk5pQ+FirvaNsLKBQ8N5o3EgJfSjaMyoZWwCn7rhd6/HZZGIIgcMQJlFh615QOJ/9/arBmEdZ
otXulxTPd4MQTXnG0ZQ/74FHi7DU9MDdvAkpfCxYQnBE+L/ZbvpLQX7uYiMbO0/DDPkYR1y4OA+L
bpHvXG0jdrdJt887CGp85dAV8CiSmhx8qYkn1TimhC7b4OjS9+6gFYBTzAZTKo5tgghY8Exs72Bm
d2JpWgg9GOpV+P6wuOsFJZFwCQevj8G+MWqkFX/mb08F3WUjdf7fI5nZWzFjNi6oPtxKUGl86f5O
4ohaABb/gPxRBqVDuVy54ifua4zRTh2MJtR/5pSrJBueiVX3vSgcb7dUfFJ3HOnhTakRlhDQtsqa
UkOtpy8Ie0OEQUKVxqO3IYes2sH3v6mVB8laFB8jcT5UFMM6qYZ/9aoLZ3lc41YX107ks0LgnDeb
jENdZmy/7No7qo9BBa1eLNXTfrHLor48IiCt0CWy6rWVo2e9t8rXlUjqSlThO39LKOSS/AuyrWcV
rfPUcacA5O/6N9Mf4Jfoo8D//fZEzgUuH9lMCc6hqjJ6QcHT+fXJD3UiFJHzsWI8Z9B8p95GbGg7
gvrNz8+afmYfXQvgNRWmLUxPlNR4ZjrGPW3/6PkWpTXbxflZ2w1jQb0rr2VDwXP+fPIRWJpTygW5
0g8sJ1AoWPRYo4dR32TY8y0WAei35YUACMQQfCMMNWww+mKm0vMeg5EL7wDTTqmzZNLrXdb3wHzX
N5TtKHne5On0Oz7ZQPVBI5I2lcidK1cSJSsStvsDv3P9ht2auAD5liwHJ0TV/LnwJ6f0zX8RStkX
mz+H63FrTk+0Ml6+43jD8OhGFkC+TpW/YcJX1o+CTC/D/HDjGS+FoNa7vpzypWknUTs29XZZEEFB
KNMwPOxW4Uhlo7si5eWdFnP3HVdTxdxYlmqXZm29WAuKoWlGWtKPG6PUH5xdozKTfb+8Kx/r+Ipy
MDURaXmqpbn4puftMEgcD/I0pinQHI6U8RjxFM0qFf/qOE2drzlySXlpuVGOqIzeIqiDan6UiGrh
ol9RlZrJ1R4TmDgHx57WU12Vm0k8wulXpDZTT+JeRtmZF8xRW3z4/GBnx6xgzS+HtAlvBG3/EQP8
Wp6IVegas9L9wUZX9742Q1jv/CZKg676Mq1c8JM/ZWvHYIMcCQn80+TVdIg0MPUMwHid48hMhUjd
P2btYzzhW9pYLTkGn8pZUXC5CInkuZcXfDi0gSSyvYAozcX/eYJ1Oo7n1G+KDTCEXKMwDbABHm2z
sftCl5uGP9yTSCRqqYHCjoPwxPy2YtCEdgcLZktJuYcItqdssZww5ZnevLWn0Fl8I11Qm3Z+C4Ra
65Bzy2xndYBqb99FYiUldjaE74melKzQfyAocMUqovm79tMjJpy8mGRpU1JX3B7UT2FpibuZ4cP5
4UI9K7qEjOYjzjgdP84uoi5RipHM4ZSVHHrl4ldXL2e8g6EpnsAp7y/pRVMgSiWjB+kLUnsZWLr7
kF6/FdCbblgeMF1x9M1ZDWp348V6WiQ8+ff4qADDPihjPxA6jaFG8GNkd3nmow21XQtmA74b0J90
mwGOFcRTfMz9hSQRyo4p5LFY/y76HOjEqIpVEZ7zYtV1mSvhFDYxxT8Q7P256fkD4c34mzt78vhQ
DWFDWHzJWlip//DWLelK+tF7qXBYLr7n1FjA4A5e5YW3CRoaJ4J0TtY27riRusXxGZys3ehfSo2A
0eY8UiNX4iBF8D9jSyvDIIm8Mm+Zy6sxRFbJPcFsnMcCEUR7yatZJo8iaEOH30LVxYGNJfQ16SXR
tYSczkReG2kB4uwsg76N88mWRfPRAvHL2fDcxG+fIrHwr4KDv3UAxmoJ3ZvhTVCDp8wHQ23iENOu
CulAeHc9NS7UQv30BXx7WhnC84B/wyw4v/3rMVbslzBgXZGjdxcYA6+/c4t4doLGl0P0ledHD/bs
gYi/CiPW12uDmJBbGTay3dD+7nhdWllvUev7cQqPr4r0m8ZWtVQVT/RgPsZz9OPf/zwqbd2DLJ2T
QXKbv5Jx6DO4RfTdtvJ+OKBGQ50mc036jYWRRHzFpjy/hR1b7NIUwhlbOd+z2lJZ6vN30Vu31Jac
4gT83YqeoQS3UCyxOlQnRXwDUhk3vRxsj5QpVWdk7OIPmzkceWvYmLPlrr/tj4LaESU4D9vqLazf
iYT8PvQTzQigB38ibgq0KShEn8kMA6LCeZ1Y3nzR1M3/t+5CylhrVKufxRxQDFrhC/oqZeS5oGM7
MhIPSxhbDprT7yqtafgL+TGUhZTW4j+eIjcWaULomR70B68mryCK2hAJfvh2vliD4othMSjx/yfk
mjidoAPIzfLt942x7i3yEcB217QVpYTyEG1J/HgrOq/JozmRYqutniwFTA8xQZeBLqGbtZZmTxfu
xbWSZf3mGlG/Rd2LdSAjoFXPjcZqXOWid+aERjgbw04FXAWGC383nGl5xnE6oy2EJquPDEzHNOrK
EM7+9wM14tDYTaVrXHh00QTsd+QB9VjJ9axZMRyrW5Z85rHMMQyFFAaVDLnjFYj1Jyo42k5MyPPd
ODPS0yV+rPjzsXb3oXR9ny+g1kTyR6xKkjSv71YnBdrD4s0b/sytCzIdDXdjPXu7Nhu6j7epXwfT
563KJDWgQOkIR+tRZd+2ZHxf7Kv9TEhRiljHXv6HRCa28IU5jyrfUQVBZyF44IYXqKxHtfCq2SHe
8q31Q7rBCPRiHQm2tqi6fMyWx3aXclAKLyCwbhQzc5ixL7xjruwL56tL3dQEO0Heses3Wq8YEvB7
v2IA6Ius1VJ54Xyc23VbIGpoMhJXZv5rwVzyJ29V4NA45F6ICgXQwvP+YLID4Uy4IWH4qY040Vb5
VaCjqguzWnr9Aqz0jI1dOi3hoTKNVGGYwie4CiRgSYVkb8MViNqo/dyC7YTgJF3MwMm5LYxQC+es
oShLVQy4NKoAqLhB82LciEopeMHCBdRlWOx8u/sMRmjD8P8Sq84nwZICp/Kwj9W+HPBorMBHVBJh
j0yiLg7yG4AqumQVbEOKvAS2QKE3zwNoxFyyIjT+07IXJ76NyihbxqBpJig9f+wjy+tbKf2DBHDz
BE0An8evXWe2C5AcxDPq3WP+3+CASbeboPPqmVxlW34c+jrYrw/Yd6jlBQspEpG/uppzY4HWGGWe
CcCA+1oSRJB9bVQcamgTt98Cxv/wGR9+8qAyHcHhE8Pjp3N8hwJnLLDh6Ri5ZUs0biEvvP4nacvA
VBRe3IEJ00/mwEOPgkMa+R3P3BkB6mPatACyakpArtI1XYuZeVe5KjcC6jyDDU+dTBfElRM3ImVX
D35cOKuA5TpOc9z1f4qikuU/2qXejkxq6bAEjy+31hAVqa5Hcltz8rBAVg74QM3XXmIviFhxh8tg
oRqS2QyiQvjrIoE40Wd++B+aISJWgozVcn1VE1d2nfvU3uKTPNNR3LkK6ytFM40j13aFqc0GH3Jr
mTa8DapYgNyeNdCwYldncLNk8lUXrUbSk/yhLGe60FhhpKfwpEZRdrgm6n+wssq428uFIIYwXhJq
EqLAUkRBQzTvyhc84IuUc5qqXu/yKLC9Phv589MVtrDRqO+/8gLd08jg6Vn85JKNM8XVX5htH3EN
q4L1KTipmDEZICaDID6LgbTyuY3zhmbABAYW+6Glaj18GKiiz+ZcSvvtomZiyChi+RVeMtho3byA
6ji4iXs0uMe1W1THwUs4IxBTjLMsL1CENpO/YZD37vr4QZEy8KcIhY/ll7gf3Bcx+yGvH08OcvBy
wOrygsgLhBbnoZKDOywnVYntkBSpzWarDViV+xJhYJqKp/WRX9tNhyUD4oLSv+W+J00Wn/HmvPee
PfnSP8weJs7RySbiD1ee6RsFvYwwrHst+7yNfGy9YnkRGxu0+oZVqoSYLmovNnzt7sZ+IWMSabHA
OpI60+u8/8NlYCYzrzPA7vptklQkyIStmLPT0yO6lkSbV2MEuzA2G+CfAptqDYKEgpmQ2AurtAQL
OeOjk3NECB3tAoVkOIskUDPKW9yA8Mx73E470ndhPMw0xPRS2SOU172hcTHWkJjKYUFpjrxNvFdB
/owmnqH0VCL2SExAA3zZ7yM4/lN3+ZgLAQsI9qz1xHfmmfgEmRExXJZpwmmMjvjFfcKS//NR2LYh
8UvV9D1WW2bDWRM6ZBHsin5FAacAXeoqloEQCN1ar1k9qQKjlIpRKxgqUGskP86wcrOw9NYvGcvT
KQUbaEBpqYzTgJ2m3QvU8FUCtrTtucGBv0UXTukF9aG12lQv8Ay2LMMYrgVjqwC8Hv1fNVkJjWfs
7zRxnfHGLXfyC+C8AUt4fmJ9Y4Yo/BpTiUTVSw2wIXgYIOGKEeI8bi/f4o8qJNPoR4yOlFsVC70y
j+QsX2YbPjh5koAYze24SGAFQtGw+yvytEdo+6oTqK/NvQMeHoBse4qfBuJWSXYBeKGCafAb+fQd
FAwGrdoU+rs9c8s6FgxfKaUfZAioCntllWo6H/iRE1D6lxBDpJBZNUvjrt3tQuLsbqf3yCycX/Sk
lghoQlQXj7KHLqJYTTi8imZY5+mcleWbZeEmDS6VBUP8JKWgaC30h1hn8qNfoENiIPJtjKxEvHbR
doKprbl0zHStpj9E+las0O//NbxlUuDlDi3M0efpbiemcUBZB0BuUyC7/gBoAw9nBeeH/Lj39CMI
Kv3/u8zFLZmTnaLoOeTZ1/qu8uyH7hbgwqvPy7POidSfvce9fTfH5LOwkKiZ058cyzNdKxAz93oy
LMvuKVnXUE03DlgxKfV/k9JnuKz4Hsxt9qamKy+kUmOZ5HCPG1bnBmxUkIKXTgGOb8rR0v2Lke2A
rUhg7IbyRILRBe7KGkcXs+1NUSmqNWqjbLXKBVFSjofbkualUib9XfqDnR5gKtgFRoU52Zv5fCj4
cusl1OZDF8/RDs3gTM3s4vUTRRdUFROmsaG+av2jy67HxL/6aeqGX05JwNRZdrwYvFqNFdeNEhSO
H85oMmuu7TVLT9y6JKGpngbl56OIsgALOfJBYjW1Ds8VTOzvS7OPe/rgQhiHP4Q40eyAdXTovsWM
fI9/jRwZ3PdQxhWiCM2e/KyQMr7hgGR6EOkFyNn5mftJo7VjBcuqWLmLPWu6f7O/R6qgWOJwCeCf
rjPwdA5ZeeGLZxoMFdAQuho8+uhvIFG1dedMr6O4YQD6p/hL7xUDFO4MqaIIkbjuHLDAMShoqvqn
YhZwZPaQLp5o2PjuG5M8cy9M01vebZG+ukLS2YziL1KPZ+tcvbjt02+sGCslyyWjzLzrODiNhgoD
PO7Y6PPW09KNVu50GuEfDf6Fe+6JuKXF5pB+n5r/qLTdjDeYDZUzvbdRJRxjmxj5u0+x6peRMLQt
EitokL+8+K4+sSRSNU3I1n7pbsw5gHm+d02JaKWM0jynBA1E9V//e4dq69ZoQm+5eSYgyjYFC7uL
0S6jda8cubsmrpQ7yYmzYuwaPaZJ+kucl8o1zqEErnJpf0KQOCOLm8PFnoE1pyHDHgGyhvIBurN2
f52OSPN2BblBasAfT27dq8/znnc2UujaEBz/UfO2c/RK5J5duP5aJvXod08iV68/KPPIU8PbPE1H
JnOrUYLxljUZzpTEWK0w4G44O07oX2OmMQmcqvB9gdFCkxPsCOxSQwJ+SeoVlfU2Z0rMsHDg+pD3
gLAJ8zeKV0FjoeZmhIYd7IaoVlByRvjKrn4DLiTNtTU4Eq5T0LS8pm2tu0L6jlTIoMeCmD/NKziD
/EywIuC4sRtnED/A3wEvroBCYc6e0GV5ni3rMg+TwG6cgT0yNon/Co1d4oun1ALe4+vtSmGPToCe
znvo0W02MLCkUz0CyCLlGWg5bbdz/ZARtaXeGteUmqGqOpGIT8DcBw5JM0Xn0nSunJCI2yvVM1j7
qnHh6CdVpwny4uO3BZr7++2X0aBxJxZuayi7yAx+lFa1LYoHV4HCu+XUDOVSFw/MJWxTpxfYB2oT
pWm/1OL/kZmTjq159hItwEVtu+XUzD9aPKk2caVHVNmBQUgTei9q/5Rh0QgAOqcTXLeYEQqZz3fa
C002hSOZy2FU3l7ysxBHrh5XWbUPThVAm6CCtBQatWRcStwaIE056lKfr3i3LTAlBrERVMtORNgh
OD5N6tPJ8nyjOE3wpiAyZATG8k7vc8NryCmuo6dUWpL+VH/XPcjRNzG8aWwhuH4zBOVDLK7jBFhU
YvmO1btJQMD2SJato1H7ZLwryhwokO33ThqOl41HxZdpJwU1OKB7jUf7kh3eZkiiy8SyggxKMlo9
RSYsXMEuxf6vFLIfPWgeqZY3v6Sug6wlT8fSFfuiEpFs6vFuwn7FFiItwASTwK5D4xHuumwVaiFU
vpsPkcwyVjiznWeZdt6lkhy93aEbK61SyAVkxm874sCExZEDCP0tA0OM8YfX/o4nrMMv5aN9XErM
XNuWvND0L+8kPxpNdYhzqA+qiHFaFuYgmioaYASMFqBeuBYDxr7dezr+zL514WXJ5QN66Jzd59T9
PZqaqUo/ZOnpEs5RwHHuxX3goOQY8oHInPembk/A6h+OhXcWe4EK3rH01rOIS7ag0h5QI/4Awln8
s5eQlYv0OhLpCZlQyq5HDXt1sY9yXDSxFHCXOq8+xs+EF9yOz4ffVPpH8RCRGT6HP+klCFmpwsSy
e/rXWxWwHIyjNXv3eZRCnUdI+WHdguPYaBxPgd4LqurS/CtLY5mpUe3Y8sr4ocrEYWWJCheR2XaR
tLRVIOqJcURmXUxv4qc8FuLNReTwnWDXf8dRgtIg/ET5444ypGMIgmOH56P8ekmxRqOeGBCJuJsy
4v0o7XkBe8qiiq9msOAXuL9h2Xba/Y07iw9erJDRFVtLDrRwnlhA28hS4xUss8oqvJMI/xyG99YZ
IIloGNKcUW5wHyIJYeZuBpl0PaebyqbMCLpuKoPhx3frUfE9pWKPve+ZfN1FCQrrSd+P0d2Ua2FH
MqjqqLyAndh7Yzga8VtpTl+p3FGtw184iErqVKBDwTKsGKCAWbs5Scp58tNR5C5PREtKJHFTTgYp
56UN2GqZ9kC/Z5jjAeusMmv75eLe0ewiI1mnIN0ZKajMWOGH+df2Um69QzuVnVpe2LsBRFb85RFL
95NI9754NB8/m2v+vuLS5VDdgi605fDQ38CpWqJ1o56ki6ULpmmUOhTbUbl1+dHMUbB9jKt2O3/s
mbebd9v5MQFoukqJzj7WfEXAPLx2b6qEBI3jdPVSxUafKNfulyJdY1tgKaXfb6IODasohSY+6y6z
ioD4E96fnOA7EgcT9CnhYUtLPNRNUc3xU6Nx3Wos1lQz74QBSYuhIASQAnqIqzpJTXIMhOlG4L88
qZr3/CuIXscEhEJOdtQ12AQ06URbWE18aES3tWBSbIKJMhRK6G6xX426c85d+n6gwPmPSG9qfCtP
I34iRBDaz1hwJATAm4FXEXjgy1siyhxF/GxoFScJRucyTOK4yzAl7lbUaZYTQ3C+5e/duVNM1wXq
v5FtuNOLsfV0dkl56cz+htqEuIZWPI/14NZzQYF2jfr3GtACjC/Ig80431yL5LbFGkVF6aURlzZ7
GneAyR1VjlEPlaaT3FriecnnQsjeMggj8W81o5mVIGvOrzNDss8TBVbtqHt+xaG5Iybboo35lZXK
jNUKlNhlqiP2w24eYzi42UnwHkCl4baWrk/uell2qTJ8JFgB6uAb2GWvZrHKKHiv84OxQfr7+Ytv
2W5cGEKoK+JrY5b1TNDIHTq4S34zgJ9qLRsZ4VjGE82ofQTj+2GIMimRjvzWKC8V9GKUgmk+kFOl
+QDqzOu5uMntkKKBxv3+UHqLoyptlwm3LOtRWePin4ESxpw1DGvNSno2fdx6qsx2cTeRWlzhDUQX
uzxOshJxAdFM7nw2hop0kQlhXScn60vp+tpuSIPW8L7yEendt983r3MyOEoWGNVwTc5ohtOTUZBg
kljHTi9PIbyTHNa/tWzhD7UYqTxOQV8EAiuobl1FLQb7OBkP/ObIOHH6DgtvXlSHpVFTlwu86cB1
UgBjPixct9ORRXCq2/2ZatSVkBW9jKWiPGSfj0SFxpUJJuiVC4jQaDBxeaNQp44711E21Xh92bTk
8RZP7D19vwEMT4per/pXQ4FIMu/MtKbiEdEUODTicv/Ymoa4dJ7aCP1vvp3Mup6c3nKLjQZ3v1p7
EedQV9rwAhwDBjrU+ur4yFJEKFXM4B790fN6a3ShJy/n9GnqFwQ+yXWdhAowJizSFZncSgSnFGqS
XQPnXngsPFw5Zcar7hv3lAu69a3tq2Zxln7CAvnIBh+UVK27LEx5tlonv4MZr6NiHp5oNWVHojb3
+08tsyTKhhk6L2tPasn+BstNaj/qsFlcxZvnPY/WcyKkiQxWd0ZJW7sSi510jOG8ahr7z6toATZV
COyOHquzqkiyZbN/5OeJ1jkUjSIvQIeYR5/5GHp2xHTeoYm74QovRn0/I5u+tHsZz0adVONjLkyZ
xJjPzPSk6IfcoYYZpMDAcj3qHs//d2aftL5kXERk+md0uQPu7oR/22D9HzrP+BDq9YJnQurjoIFn
KoSnep+WQK3DZXz0GoWy0Aixwko+d/eH6ZUNgzBiKsEEtpuP2C8DPXUT/++HatIIdEfi9jqGv0Rw
/uTFafEP8kBpy9sSrGhDn8S7cG1RebAX4YMEppsHiCwMD+dSAz9m9RmUoRIUaJY0CpagSzF3S1jK
KTb4eAjmxhU5HH7BBUsPrbv8Ax2gNZp5x9Gha8kKZmCdI8oJG1J7ZvdJoKuJ5HEUgoJHTR/7LWqZ
iUo3hSIJB0oIYg52fOQSgAdfLuqaq8KytluKY9rsI8Nnzrmc+tFydZKuyTI1Q73nonZd0oyrOWnt
YdpzEIytDSLPuDI2PXPG52wPGmbJUREeKl5aheM22HVUkKCafE685Swnoe/JtHg1TXSXAf1CCnRj
NKPxwgR2p/ankRHRlrSqUQUkpNKC5z6OMQCbENW7x6v6ieTniCV1T4AgUIg5wld4M6ZM+0Fsmf/p
eRL1wvCXlTVN6O+gMZoLS41onMFgeQuvCqkdYJhLUTp+Pz9GsZ0AgLNty/v9Hq0nC+BvRYxxRdoE
jAkuzZ9AUOa6jGCqH2WF8qDPd9lWjUfu5OFwPGYcv7R5PxN2y8M7p/RoRd0kRjR91iC6xKYg4Zgs
NE4cFcMoTjYhoL3izxREyawGu/+6M2iJWyGtUEIz22NzVYDjSnUYo7LDUWY4FaOyQFA2E1LOViOh
zXhSxocJkxQk9w819Xc24AtTx1ZGuthb/Z+frH98Uex+vkUJVqLUSggXIf6u+ErCWmPnJcHXS9xI
kpuOLpJR3Zw0t4WL2Cj8UkxPzEl7YHmxKjTBL322T20VVNYTUu6OjKFrhEdhgsAnbkWkrPCkuzkf
XV5fReJO5CHjEx8IrqgK1THX49VTqTxJ64Ve6xpOYokrPCkhDQcS19fc+8cWtiLCwgZ7rFwb744f
qcNKOkBl6SzMZKPCg5kn2dXvyJLiwgWS+0Lb8gu6FLGjxezj3ub1Bvi4oGKWlidImnFeid5RH+sN
hheX4xtjnbCqN8wNNB5kg7a3rjC/iN11xenMto6U/1pdHoAwgehKXhT4An9Zy1N4lRIeUIJEIDRX
Yfbf1DrlHIqrOrBINyoWoVXKz2wbTJ/joiVRFZ28ne9YIxRGxWVUgLuk6qhLz53Dk1HDV07EgKhs
qEnDnjVJX/LaZbkmcT6X8oGVpq/9M1Xv0NGSgfB1cPUemEAZ7vdNk/ZF+H2ohgrJY65qwl7FQzLf
vwlzagODKsZ5R5II3bJfm9GDUkQJvKSiAL/ukV3W+kQ+rH8ozTpoW7rSJ+vCLqay3neOjLBqaYIM
zIlD0lv7SrwvlUs9c6PD8jgs+G+Aq3iUlz1gjAsAUQrlPysRqRMRAfWueLmKXKbYuurJHjrjmu6r
WE3hWqws4dh4M3lBMdObyuWPMFtKpJmusD/h4f7+zb+AUg0Fm3CZpUQnGxqy8WCKmSSHE//cbiIA
cAEdyN4DhOIHY3x7Tuo1IFRitVeuVmoENqZCT5430tOTSv5mUcjy+DRji64RUWT5o8ALPmJ2cXF5
ZOVLooKiZADGD1tBVTrhwnpRc4kJSw9T2UiZNIG+zhmGW9x+XXn6YfJhh8S18FhTr+4K7tfoieuc
IEnR+KiH/Ga2btfrPBSy6KZyZa98PWUrJBB1j5pxNafQoT7KRXLiz4QIUh3NHAKAYWJmLsiN+UnU
eCIKVhR4wP3ODp4B0NryVkw1zXM2MTjeRfYKnm5Ptcyq9m2RNu3dfU4nuJFuT6tlF+ENl3GZVVBX
ls9nwp8/wWcR0sa2KQexbOknmrgp2YXxF+PPpUO6u+Na9XO1UoMxbITk3a7uIjQNN2T3m9y81nIb
p7KLPvxmUHoPzlJElvc2qE3DMzItwzwsKr0CTdPm1VsTSRdaeDY/BVnM73zZjUO6NQcjl+hqlXZ7
yL6TMOrbhhjmAHDvng9R1/Njzhh8fMrl7mcJC8UkYjFt73qv7U/Cjjab1t9O1sxGfW5w6MKrFokg
MT43LdYgdk/0JRjHtqSW2YYA05XLCvAc9HOJ8odao9oEV8SkRMcyDrHkE30R7SN+E8jrt1bwxGDs
jn6Tg3RqKdUhzr8SBSTpWzDNE2xUzrjY7BaPzgbVeeJueWWKw7wLdINfirV6lHMDkLv8Q9fLGZJM
lQnjl5WDhAaTeG5KiADA5lbtK+tm4MYoUZeCbhZKFoSN3TWaM6gn+BqraOaNapMGfaiH4SBtfPyQ
/J6S0ifFWEIuyvm8zGcBb4NrYlJKlkJ/5sroIEgJCwiHQ2T6veF2pff96nW6WOktO2IrOqRvwnex
wE+xibR4veU7Edr9UIB52NraVsTjQV54z+MoBMg1Kmaqm3fOQKgIuhPl0/MDnPSLZiRo8TO92YM4
ofAtndPnMicGOdDu9vmaAFdwBx0XLd5zqTNP2yR+90RXdOC6vA5+1bfbzd6bv9S36fQz70XQRrHR
755cXC6pVbNJbEXVPTtDJ9HoaKFMmQCZBmv27/h25Lx3AS5WCySUQptDlp7L92vamgr5cwvVHlj5
Z2PzAeXlDNKHb7C2t67W3kZ/xFx6SZIwYByxJ2/MWvPMuDsOsb3GO+b3VsjrEuwmFm8lAsUJQpfI
yQ1V5YlHsTBo+NhJDC7+4OEn1ecS755ReooZwaNuiNvM/k9kIQ+z6YZ/PzoacsZziy+scF6pUNC6
3cq8kTlmcz/8s48jCBiwMw7xyvlcuX5MsSa5kTIVh1Pqk3/tuBOO1cXaURgHYZ7S5YCor40FG5WT
/ITwQPsDImmpqa50XkJcwr686L2p6dFOBz7f2fE92z/zRL23RYbb5PmPUa0I4bUEMaQdUVhxDrPS
LySKYoEGbdiHaCXYp+c1Cp8SXbw6SwtgRnuAc9D0Iab6Bvb7vcuKiM59TBdnTIpkolbi5WG3MJgC
td2fUsS9Y8qVWeFCRDVFKMvOadIRRHyglNRR2tZuBJubCxJxKG8rUDH+PXGBVO9W8Cd1cZ5Xaak6
zXZnxdOEp6W2ir//3r3KPh6mah4kBIeeUoqKAhFfuRftshHK0iTjkRFvUIhKcQ3isHxYAK7nVR7v
KNd6t+FBRL0+a05lTTnYJxpUvJI03fuBS2f/EPF+oCbfv6yVTevBcF5urGoM9/wW/dJZjsEy8M5S
+aPmdo3jrXnfQOZcMd78oPlmFe5xpiDf8/eW9Lsjn94e2TebOz6KzKHQ8gAbrYUQSI6OVy5MPE4y
smR2Gv4nGhS8RytPVR2mjHkeMgA4AODl+aVikmchK50qidJOYQevUUmTI4lhKFWht+Rda3acncrM
qPwvaUUGeBuyAfCXA10nWFX+oUWRVGmRdqyerJOGrCcCQrr3CdRvsqptpaeTklJH10x8v8bQ3xoQ
48K0uXaHn3N3uQG01lp7crX+Xz/mW/HO3+imtOtthxSXa30abFYaF3WIJZPP+M/uxTzk6/yVi9J6
aJQqhkqYqUrRBqpRXPM9mvumC+18BG6x1sC5/2BJmrg0PYHIfzezB+shk8ypWdizksSU6JZxxkKI
XzMc78sgPkfaudSkZA8U3519gDKr1PfmjiTFM/91yKohWxcETQCmJeoo59hVJc5CSwMe+CG2rZlc
cp2fC4kzcvRycuU19mDY3c7EYiSEH5amyl2QlfnKFn8dj+UpoDGWzWKFU7WOa6JcsuVb+V4I/bTy
Sx91VmanbHF+zZ2Svy+6Fj/vA/ziue+Mr4zg3VZv4fxpUwhRc67tLlIPuG0OIPbfSly0Q3WMqQou
UhJnWbeyETA4O8aVUXX16WtLuIr6ftIlrWRPimlpin2Ggfeq2iyy6Yt7Tu/aQkwsvIDeIFhflB45
QqjiRQtRy/2YnfMnfUcba0OeKPCnHVAdpMpQXRAg0V6D9Wbbeok6a8nyd6TOaFlXd7H7AST6ziGf
vCqOsF2SBw3EfAE5hHHG/5w52aa/gNjbAG5ov+yfih1bZ7yJ7rIwHxN9+D8fLLUE2qvdACw3dfsB
2bZoTMNXmlDR9PCgvulKa3L/w2cYxHYB8T9vrxuy8w4zCeVN7AS2nUMZRHoV7XPUabqt/itIuxJo
wQrbA4+VaGHVSlnQbULtNQffqT0D2HSzaFSIDBWQDLviSjK7msmpAFk+w1+NLg6NR4YPv0psz7OT
hg7MIF7z76PFrD4gWf1X2Z272GJEMpPNpI1zBVgNL2KBnHj3hWx/Qs2V++OADlgdMBVzJe6pBon0
Bd5aRBNIVtCSM0h0+1QQ9qeXGckXiKwkQYC12d6cfztUpmFlACn6wZRH/wuy1rqWqJURSJ3dMJ+e
A8o5x8UGj7Yf2dRlTCuKFLQ2JxceI5OMLLdrM4QPdUQ0geCnk1P1K9y7Evg/fuhNh6gaBuTo3F6h
SoUpPdQ//QmDynXh5e03FNd0KnsFQgi7+numZNfOtTSkusOGFhu5GZDePhD4ZucmjsOopDp1NVXi
hdLKBVx5oeQzo+iHD+uFg79x9Q6mmS0Klw+WecJrzaGc4inoCZW6NBJq2rx2mBF+WgM0l9TejnXW
goiqVSd1zsyIjnSa5FjoJLkYQJfLPYuI1TqMtaioJT527lMHiwvgfyLWmj8rf+Yc8Q91EbBIQaox
HivE6JHmQHFb5GVN92amqnR2x6BoUy12NHNejex2VpMZA4GQwWN/q3fjCltpWLbfvfsYXA6HnGdG
bFtzT9QY4W6aX+Ir3NzD+vCuio+zMdSJXn0rrHZ/q6ZqjGbsiQlkLPV6M+WlGdgduc6J2GfSwuDw
Ea+M/n75qFBIVqJcxVyM1ZYydzv/KldQV5nKcqwhR6f/PEWCMC6z6ic7RPiAPm+dvbBu9AdKMVi4
+EuiUlT2oN0IGKUEE0e5P3PA9quxTF35kKbuZFoM4jVsyijPICgkeIPYlq5BJMN3NRJRlH6n2YGF
uEHUHt7rzqrEqRGzcpO5leUYfnp3BjTi6zDPuRUUPjc6CfWAY1lSSm4/DDf6+TV5UWWXcUt9EH65
6q7UbTqctKvwwmt3+XpSSSy6GExLQSvp5gQg4JECIcOSkoYjd97fjxftqmUeWrlKoNNuHo5g7Bvt
iY+F4Dvi1xzA33pCYatxheEBhIruXsPlrwFepySNl2nSb4RFmOkJ1vGvxh8bY/poygi4n5dLzKGi
A1Lp5JyroKtr+YL9b1UT/hNh8tZf3HPhelV/p4zHwsMwgTmDohdDC+Cp3R0dBo65NEJtWp5ElXXC
K4as3MyeukYBLPIp6s4uhCg44yFYf0kxzfARo/+jOogHKJJabnRKJqID4oong2aCeLpLvEC9NMKB
oYn9SjGRB4XKp8s12Nv6Of3gme/5H6NKuICl728HqSHeYb5WWWNK211tmun9q1fFA0NwuHHGAWC3
3hoEaswMNQyFeH0+izyf1eiLEpVvKCeBt3eq8zvKfjbg8EHDEbLH+Yw0LpwcpFO6umCoxp5gq0DT
shSgkfzyikHiFviUjKRIWSgKypOk8gQAVobbnVHb3KvcJC8miWlv1IHU3MrNZNgcz4s7RHXe/cD5
NE3iCiA53dn+5Rya/QiS3GLnVN4y/MDxztf6zbUM2tsReNcoNr0cY04B7L3fDdjLzLZzVHwmp9cY
or8HeGyW6oa0O2r3LY411Az2+Qnldw+MmPWMMrxfBNn5iHG1Jp9jkcCR0J1Dj8e8aTg5FnBlnVvN
JKEGsZkqG0lj3niL1/G/VBkL1vyTDxdVQqNHl9+r/LdsAVXjjTLvzxUYP3mbuP/67r/VZ4NnUq2q
ARtz8v/71oFwK+XN/yY0rd9Bfc5BipOCqo4qbtfswhhLktGdkpnKygji8FXBzkMhC8kk2+Jt8K54
L2zSlv7pwVIh8oijHQ5QPy6s45aBNvPpWEQksSGYxVR6A5ceG/xFDUR9RhFi2c/Uatl3LNFMDtX/
w+V+9NqdzCfOAP9g33JuIldVpnSi/gCwyQ9IPia11iPPKSPO+9wrsao0CJj51kPmE6AtPQXuebq9
ttUo3YOxTtNLLr9HgTTfqREPNec/ocfgGxxGOGR4RDaHEGYKBTGHLrzCvkDs6KlU56jKK+osdUDI
bbKfPikdSKhNbMN2j3hoFgDs8jSoQKSYbZKPgliK65oC7/wnkt9EbFu9dIlAuXyu5j6U+F9H2tn+
62w5XddIHCxCSMS8YSZcW20EJZKQ89mGg8IGLnS2HgV9ex+C4Lv5Jp8JWEzVw2DbdtwH5o++uDKO
kZ1QsMeGS7AWN8VM1Baqtim71bxYguG1PJ+E+5bkR3PDM0mNcZ7J1qJAd3eMmUmuu0WZJGQezA9N
pEdcAW4oKaJvFZr1uAGeyDfY7k2sLL0QBwioQpVAdxVHL2YsEP7/VT1jYSiSMYfr12TEvbovnB8D
z7Ee0B2Kqjnf4osQx6qav7vdCymzawIvpq288iowaGerZKEV9AjVxX/dvtZ3mR42Ekk4Kh2K9y0r
KAz0jgBmn6LoI0+KQtDg1k/4iOWWXkPxd9xTDBgW7NpPwupqblw+muy3malfiX5qDo0pFosYO2oZ
8LHh0VUDQW04G026XMKbgGX/KoQdrKmADJwgYEldn6FJct6dtCBZp7qjbfuSpj7qqz/17+07cl0h
Mk3bWOCZBNyfqUYywwJwD5nJ47AmNsoGMfDv8WoVo137/GhgFv/LQpXkZTMq8ZZ3s9lBNVgP+zuL
iZp2Ewc4EdZpX5ifvONt8LJf45mr0YmC90rfbCRobqkZaURUa1t5qCUCEBfTmjkLpc9b1tUe4i9z
XrYoxnpm99gBShAqM89tka2XuOYbJRLYWDruDgyS3bQy6NeVvy9FxlDrB1s4p7iXWzEIk1N29R5J
TzvSw7BF/6RNGAEEtynmGHWn+t1VuwKaS0S+S2dv+vV2XYk2QRj+rDM3CcJBPgOQLZlSlTMiPCAU
EKe4qYTv3Xjj4T7ldGan6TM4m23L3ZRjRllUDBHlHfhVIrjeNVBUsc1Hy+Is1uoJb3zz3yRtmfPa
r9dfLH28I/LDhhwO7Tlm+eK6dyYkiZiNAk2ojLmU9lLEI4xmYM/O5Enm/8E9CxVoT2+74vJxMSPm
lAASVA0amGKDGzxiXPtd+F60I/qxap4C0gctZ6QRlMCjjbTLEYcK8QwC0cGou3AnfFV7uakPW9HI
ueGnUfmDtdJjaPpV4j4oy+RLB7nECjWzjNDNXpHpbpM5PbH6xeo4S5jkI+3c4ooLo/n7LPnpXPfp
rQis79D6i3pMbvWU3QCuVO+WMBaezYpAMCMOtdoG10a4bfffInvujsLpI9+HbEkMvyta+g55SvlM
KJfSF451WrOFES5Kcqj+rdyMihhNEg/r4Ydgx1U/9813YCTEyvW8UyHtk48IhQa5z/vJw/f6GPJk
OqR7TVFBjtZm6fyiGwsVH0All+yK86mx8wOewg3RBV2uREVHyBxgMtZV1+M1Tw9bslvTcF4YMpHO
NyAHzN4C3NMAvGm8gjl64l4T34T/jkHCazGhmVniM6NVBMYPP57cbRAvwzS19CbQXLw2Z++KpKuA
p24tP5PU2026aezaHkPjlHHlskt60U0rbG5Yih4NvuvhiyZnmfEstwzsOQJ8/xSbZcsiLMX3gDpP
BnC2qPQHt3muaiyA38eNYkhPqGwJba8THhvP8lkcYcg9lkh0scNh/KM5YeNpoa5Bdv0FDxp3HnPH
vTuUt/OpnjYw36Ct3D/X8SAjZGtsGMlkduDX2CXaoOrYVaHt2jCK/iza+1So0CLs6YlmCu+35Byo
6NZAjVSNZ5GydS43tFv8y6TEbHnS+mP886Y/D6YXBlszzKKmzIeUwAP7ozvQwCgHF0nk0wrcKJHy
1UMRJCF2GSVmR7lIEs//lMCOmeCnvKHRBYwuAZLETHqD8+yO84CL3Pgq+lvdXIlNN6iuzU3umMP7
eJtCT/jKX553603iwGD3miAldjg7bHjSqv/S1+O2b5IFlOKbgY7bgbi7TklgDJo7U/fFWZXTv1mo
IEXncNMtg7b20BmVjMCRkPNg1GFh7YGGv0yM3F7W1hW6/BdMWezjUJqHWiNV5K5QDrgyTJbvkqIb
tGX+d4unoL1Dh3zvlcumc98kS8ilCYzUdwpKrf+Dl409Vh7Vg3fOcJp5VqPXPJvZ/mh0LLewCRBY
Dnk3SfQ3ldXLiS7XY7O7zRmwn951ltzch7R780OgrBadNknu3IfUGSU5vPzQZ3JXuuP4GrR+hHyW
Z0TCRmVk3CEisIamGXvBS1fv6wpesTKm7peJnV4DH+VyqqI9VirByP/xUoD4pmyUgN0tJ9HGESr3
6kGYGxsqsPQvTRdBLjjtvRIf4PgUkAjRtJL3a6Po9yotux46M4u0lSg9yOTtQz7343VakDTD9986
aOgnUzXGjsziDRTkdL1m9AaniXpLnvZbeLbcl8RPiLIRJElwgf2ysceql/QxW6E/FPP/egrPu2DD
c4wKinbyOciotrxd9fXc9sxEUMEF10y78HmCcbIhFTKJXwlO5m65wSy3svlXSrlFRaePYeydm4Yr
yC+o6HQqZEH69TUaPJ6PKa/UXyk5NAWJ+2aVCfFcQoFIZ6BXCdHReMeL13DzvhyWdA+i5ukinFpX
wpgw9I84MXhnBVFzaGlo5JVrHr33cLQ/j9aa35rwHtFIRV6GX2A0Ny9W59Wz4oHSK1D1kpectDw9
LRge8L6mAqvPiMBTVh7UFRMfMmt1ttZz+d3eJmB5gggpZ6hhvnF9T/RnGgG0ojL3U5MV6DIS/yUJ
MZAs6G4qGc+rx1F0qD/W1kdlNDsNLv//tBI3iJFZ4A9lkL7dOEjjeg7Gnpbiw4MKt1z6T18cIwcu
+WfL668z/lrjv5oS2uTrb3Q/UiUJsPt+QH+JNWcSf52NzMZylf+x4gvEFOsKZBl+7R51MuSlF4Ri
WIisaQ1E4v6v9Xq5bt/KL4FJFYvGoHlVozCL1KHeapcGPz6Wim0sByT/fpMBY4QOJMevRX2JTSbM
F8FvYcXRYWMe4Iqiq8przvFYDye3TRJf6NtmhxVnO0f72Kybtvc/u7DSnMTBpdfem1q0hRdsuX1y
4qAIaMJNCSzsbJ4WdFiMzsmK/nXTtliw2mYFRRpB7Y+6cwzwPTDdDR9g4gZR567p1RWT4woj4HNv
gdo2ttvzac/QB5JhC0LVlWSB4rb9a9N04vfbBPT37/IMSWpNfUE65a9KKRy0Jon+mikmYpKBmwJp
U5uJPKd/rYpEL4QVqxojTgqStf24Rxx7N17RQqN7VtIoOnUVqXx3TZKQEM3TC3G7OW+3nRDfcOT3
e1dVfbTEF+q+2QS1mTNBDswBcS6qsEUc3GquYpfJc7ed6pZAGc9gsCU1HduQefcRCpk4GmTA8stD
c8dTj1VXS1QhmXeP2NMAWwiyVOAwdP9r5zydB9bkXOba8L9ymsbLr90lY17sagtdRFE4Nt65YWy1
g8qC3vyKMZ6uJ+wk0qFdZEcRCjRZ6JnR7AlHN4MUdadGU+ijsuWCZNapDmF1GyBQtWx0G6S1ycuv
6ewdv414/KtHChACKew6fUBCtw0XGMFxTwcdt+D1VzR95QUW58WVPopcuvVxwWtF31+YykpULPGK
niiqW+WvXK1rsffwXugdRUca62OwBH2svKbeXEnJNLgSjB8EglcvowoqyIl8h21NOHe7lnXWIwp2
ISVEEHqRjoELHOsQbuTT1XEQn9DTXmGj+5P1iWnZbQxkTTZ99NQ8mlzRP+JIxjK+PrcN9/C8Gfjt
dRt2M6B/90fiZ2tR2ZR/4J8caten6bMK5iAvkLUWDYKa+zaqaB73KuKh6dwIIYVPxVDa7By+F8Fi
gw6Z9jDSiGL+xM2pVaNnVSkgss4nMvpngPV+57/YMtZMfn+qiHaafb+R4JwdgoO1DixiW4dx+OfC
ArythNz43HLEWR2x+V3MepNvgQxLJRKUnbU/yXC0v9jUQfDqpzm+ar44w1OnX/Bs4qGcQF3JHemS
bJuokPjGiPz2LLgWZAloPS+a22yL/umIned7VMnxPv39WVy3vYQ2vvUjiyfSJw1xLjtG5lkxz/S7
O1CkJOFmTKvCdYqiRtuPgifMp7N8lpRGjepCVRpyfiBR4tychXQnlvvy/PMl2RSn4n9cIhi4Wucu
8K59gg7Bu3VwLa54m90s8AcJB52dro3Qu6Ch7cpG5zg+Oa2zm6L+NPaxIfnCWY6yQ9xaijP3FjJW
CHdUwBnAZe7En29cqOhrAxROZodfX85lnLKWOnRdBHVGqK/Z7c/T9XGfa0MiZrkPamFE5nJ/X7q/
e39KNuspT9Fm0PJopa2Vv99Rtel4TnZWEThBYM5Gypck4Wh7v+KEC6jwLHVFc1W8d3sbSrz0ogmz
nlQAIvzILhtOOI31qV7ASTtAcX0+IW7FwjDT1VPsIuGOAyS4m9Qb1XHhr5n7UT5K8fZY8xhkYF4N
znVuXHmxjLNRIog2O2vu6pbGF8IBN2EfTt7aJm1ilm6/0Aa1HWEgbFyF2Ysw3QlrsCjs9SQEpk2G
8l1qSi9rdLsidCU1MXtBSXAv5Tb7i51ioeNvyW5WpQrvZJR5a4JUdo6EjcoLDByYhu45tW3e/ISJ
FVRMC0hh/m3ttKylS0VUHuhNDewuazzJtWdlQrW3tRe2G+sK10iSUdtS2zIoagl+NPg9B4SaeSHL
KWvETuq4Db8Lr537Gdvx9/JJObLT4XYvCUF9TDg7FWLQYuB/EB6p0Jo87NWklZik485/ir1yVNUU
3rU24/Zo+Jrf1U35K4hsYeF60NSHVbpX6ab2Y5YNkr+qK+DAmYPEWBoIGA+4ovBCFqLx2xrDsuar
FB7P7rzcRswAzsbEfOvt8SgsikOiTJywqkrlRb58kdLzew+d4jkZh6XyLhYk1UC+flvcKBTS88oY
jUYOXaGWg2+e8GocA85vgXDro+pAxzWLZzeuQgLHiP7YUjDrQ95rP6u01gEmJBbMivEIgHtraamo
5nwIfQ0RvPtEXuWboc4K1z3/FbIjZsD+aXc8LPgm2Lt3fkGNDM844e1jkf+Pe7WGSWgMIPTPMeCj
XSAuKDDuW7bDgUTYZJFFHtxa/6lUSDldTsnDl0CRBrl2hpBrhVokq+DV29JajuSiP1BnpzV7AGlk
c7W/CYlbksK41x2761LfTgae86xQI31Dn3bzln4A0iy2ITyQ9e9glVSHL6gXCWiin0tHWoi7JgsC
SxUHU2e/PNUfb/ZxhAjnhi6Qfq1aibn6zKkCU7jbn9vKAX1L1xPlUfA0DiNKuRn3NBOkCrYFnxh1
9nA5l58c7bFSsFIUfEptxEcA9dFjUv68fvw7UDGqoI/psCeAJmW2Qg903Opu/OR4feYmZeSE8x64
ORuVagKFi1ijYR7KNhwWHVIW5vSW/nP45lvRHyBWztjCnYMtywa1hF5ur5Wb9pl1kgaR/Z9erAnO
FIZQQZdHIRkAhO66ZftaCGH3dAzOK9UQ3tNfPUIbuEwsRqjuHdhLYNHM/XVmxQMqRNHJk09KOJWT
4NA6EGemZxjHgwgfcfWR/q/IhsC4T6qtwbqqj9XmRFIhfDoxRTDCI/+d25l/tkrEoBUTAQ6AnZVq
1aN1KxUke31gV+0IC+4+CTrtKKMQ10olopnxmrKZEoCUPMPJSg/tLaZvHHo13VI3QVOcBHLfa0I+
O9NzGlM3yvfS1mR8vdLI3P1GTSpGVmqjdMTYztkg1kLPHlTpOdscuJaitReBiVs5V0c5vHq0zk/h
Icvjhs9ujLlRqc1dw+z/KHBy1ltDgrNe09gj2Y6qvgGGz+3PVjg0G/+6A6TZr9e8PRCk3dewmPuX
Owty8uZ7StZeB7zT5euJOXNl6ZHtWo/wFn8PDALYbGjmObUOTUlWGNwBCk7MD7Fi5zgb7R69oz1b
eua3HDhpVGCRsFVzaHCUj4TaZdOYe2vA1t6EPGShjN/KkBKPWa473nELolAtHIulsmNO9xjpaXyE
m0Fvsliy57OWvGSxTMYF67h9HpGrrwuGRv4hnYftBnpCYYiJdYlJx+R2DA3BFGhamdxlKZRdxxNY
XCpSFj6hqkE7nNOYoJ12YdHlW4ZqG/v+3tHYPzoUOcn8yifV0+ehn3q4qnNLdyBTRCASn+o0rwzk
1UtyfC/TtSgjR7nwveaaOkY1jErHq/9qy1p8dSy5QvzbzBGMIPx9iRSONMWm1l6HkYEdwdjTXU+J
oELiqKRDTW4Je14f989YwVWmR6VwJRWuxnDFXyPPJoSLYBFywr/GKBPBkTSzYSYBJNRCTkRzZva1
cbyNS7e6miWegPiUij3QaXhbXN7oFnFfVjFZsSHyfZUZoxkTRCrUqtMMIReTAcwqVLYGrfK9URky
mxEfeTg+ZwBnDaMghGpXIqjw+yj2lFNsXw3NmDgcNFUc4BGQJzAXnZLWbRS0y0L0dmTJUllf2SJg
hnYsMDxnw+LFnvH6ulm97NPABaGrKau/PHrrFvQwvNSd1tACyEdw7zvMOMEeBYy1G/HJjBiJXlLu
WEkMMbM93vCaf2MvlfYpGKUD8oEfFrDrW5y77vSfYnOlORtfsq3GzE3fCsrlea6VaaCNyMP/qzhp
Rf8C2I+iUQrF+ERFwThJBg3VZsldjIenXrRQAkQvpv+T22FK9ytaWApfHIFgN+cjcu/pLBMcTUYp
I3HywRp1SGOLN/BeDQQxCwRrq56yXuYjUCwpqbmN6+/zD6yrTHGu31NfaOrqgmksSd+gaKzquDI/
p/DRgiDhKUZsbaGQVzPiT6u26fSNZQG4fNnu3mKr3KAgrhPEXyJSU0Itwfb+6dO0MpJ3Oi/g/ADb
Sy4hYtKYufhZWOtNdZrfEv4ZZiOPfPfg0eozv195Ao1KPDZH6aHjluZZec+BU1QvKnJaFsH7KBar
xCmFGL8ofo8vSpBC0vEDMEABKifuXGgJD3R1dIqpxFbVdZpnnF+EkRYLk7/5l4rOxTadRypzavmI
k0mOVsWaZRyyYXyrWO58UoskH+9jlnNC2wnO0GhDYjRqzD02ILVhqD4R2pY3w45MaBRkaTGfCTLN
hgEONjnkOezXk0e9gtIIenK9mb/M9ISmBX+JCAXWOIOrLvsAmJ8Eq36Md7sPStiCWz5k5Q5HuOFB
nLqSUE8EjK/b4qWtHdxq8j8EUrEGaXSpjKJsYsDKTUTp9vs9c9IxYxWgv61lSLKQ33AomyLpO8rc
OVIl4pVNuW+4ewgW93olJ1haZKKA0QMi2Zkl6liUASFk1zxurogSJiDzeCePxt6EUSg4W2uqPzfF
d8+NCDm9qp3AyZjWN1ljg7T5vPPDUD9nuWhYu8bwbAL7onAVgJ5HuejcZpwB78gWgYaWJj3UfH1Y
i0l9rOJoYm+wkhmNmNJuBBHiWozf/ir9sLXzevKr/hlAmufjPnbXtqCCWHsmbPsmsnWBVqjwzaWF
1R8MFpegzDHHFhErU+yOmvDzEilD1BXtY5opnM+H0i2wKLf3v5TktByrkliKDB32POcvUDCPGrR7
r5bIWeSP5VFbAiP1VIetW4UHN9T2M4Z04qVqYXXWKvZ6olZDvCVHliq85g21TsfH5M02gqXvqVHP
wyepq1Xp3Wxgt6mVg/9p3PBD43tdFKDjWFrp0wrIPxmf/7x1Wfd28nDG1bFZ5isjAOls6AScOf7i
LEDUxxg7CEa0Ovlonv7PJ6k01oFvT3UTw4yhaCauYIxasugCNkTD4PZpbaf7jkAmWQbyDsJRjhvO
FPPSAb0pNBxcFIG9v1+lOcHMZX+TWJN8ADPsAg33snvHJy3u+7ZgmXayorXxmVML2mCbF/mgdz9e
MKjHI1zPlVYIEfpThDwZ9D6EMFJ3meecRiKlUTZ48XbesV4ukyDBG5Yco596mEyjWiuLI4SbIPGY
63SyOfqHLyG8wz423IbZR1QiLXABzFyDceFvgswO25DdcXj5S0lrw7wSHNftDttJU5OPP1ZhrA5P
6MVWv226O33PpaozIyU3bcRC6WiCs3fw2poGKy/cqNTNO1fOPoKXDgXWOko/ORII4FYSmCOd9Qmv
2FgUgyzCN5YZhp5kujFEWh67m5rI4qeBdD8BtA6IrLtRHmjMbchm8qHn8oSqtBXscrXYxVMFXx04
YIJa+3hpwdjNW1hWLhMhidwxSV0Ezf4h48FxJVcOSIS5uoHHgFJRz7WAD4rWCgbZVc6OWhDaEj68
tDdi67h4jowJxBiQAFBUvWnER6VEhJFNXprXVXkDJtV5igxzdPQHi+C0K32Sfnxu3yCyB5hMVbZp
satYVoOtqz5FxgqrL0kJhGL/rMlKsphKjeQ8L64KJahz7fac0f2U6RFCaQEfL6Lc+qKjwM2hWkL5
fw1h3m0826tFQCeOs3/MqJ4wPudB0iBp1No6V5RVki7to7p7yeKcQZYSFucGQgD3sEawZCsFi0da
wD5nEDpmXnXY/RLAo8fqGrE/C42Pwzij/cGqHu0O/WNkG747pfIRRgCC5iqWoNDNGg5WTB3Vinz+
SXqQQMvnl6g9OkKa3JCXuDD9wkfAyLOamqDXW7qxOrq86zeQdljsDtBTLACr3uHO6qd/BBn1Sy32
I+PU1hZTK88WNhQL4+0DTPaI1jgLWYheObPQ7DrFRCtmYhmShIB4VV/lc1zP9C22binJs6ZJfgvR
mLxBKjEy5ytc5mSw/Cb0OuJ2CpMeVcc3aDl8Ghn+XA1p3iwd4SLhLJ7EU95x/J26vLR+8Hd2LSD6
DwX9pXXo48CODOAO26EQDos9tttYdMLJZMiyzRhAeS+84LosHOUfJhgmsfyiNKD9nq7CLM0LpUpy
ixkfzqwX/zMsaCWBd4bz/Yl9Wvoa7o3br1DQ6sm6EojEzQZkEwLA84vCqoxE6513f/65WGpuxRNR
B56uKw9rKuiEesIIpjk3FeZHe+BpkZN1t6rDtwMGdcjzipF6n1hW9RMy8i+QGDNj7wI9vVRK4hjl
RtsQf+yxhedBm5SOvLbct1nx/PW+5ldHS7QC44IG3I1gQqEFoxJFMqTYNEyRSv3xvWu9fBeMbad0
aV1UEIfguTS6JFPoBcXxTM8hWAVbCwts751Dh0EL/yEm5CI9s8zCJQvhaeBbND9U5qfP5cjy9cfJ
x5LJtCK/6BoXyZ53jCMfwIKQyMzkcUNfo2Rkn+MJL4Dl5QzMup9P4Z9PuFzIgunuEMQ4XerpEVbu
qRgFlWLNzer8Q7QBeHRPeH1J5KXj3t8YC4jqrO4dh4zpOeWIup0eavrhW8OewuB3MQH+iU1ZTtT0
IUE985xvMKuG2mll8ykHnmsHG7MjX+MS2kkuf0EtNrqDT2nRAume7mCWofOECeo+oYmMCXyBN/7U
zzFws3IX0pD7olBc16sbkRP68nyOwaek3tU5kF3T0OF/xshZxfLhMW41sVN/ZO1SyQK2TyQWDiNp
m7W7Vj8XgEC5Yhb6/74FXs+yDBgMNkerd2WqP0HlyR/N0iklI8mpS44MyiRzy9r0aviWY6CNBK2+
y2PSVg17X6bPLCp9iOop1XNDlk03wkiDNvnoxPC52ymFxw/7I2V25evWcsfuBZbGu6FpwaJsBRt4
Z0EoVsPd2MHVVVvJdD8DObrf/XIJzIjaGnwx9kjbEzIsxhgaUp4h+qV1SvN+BukrznAndbCdQi8z
fteYTJucMR5WYMFtPZvWSSmBFjB7BDhtMeV0ZzZmyr37VKUr/7QOiHN3mI5bIT8z24+OBeKEFhTM
VX6drkI3xycXuhHngYaucSKyzxUogTrzOlqVCGijo6AiTSWoUMU2tnGuI385vT+EF0kno7aHZK6+
rbN2qgxEZMT3dukB24hPeYkID5fszkqoJocGKHPtrYKEWJV46wt1+yaMq/PuwysMVctsShh7+URO
jc7ez8d2MvD+STPg/fi43kpRVakbOgm3ofglFie9UkCFnXSbtVJOiA5ekCKNsnnRA7iQAZKTKzYL
PwVJt+QvAp18aSYJ+GferuI/EiK7s4XmsX+QZGq0DoSXmEUUctRTfMij8gqvof94pAwb6POdTLuH
HxG46qY+EIvIvE19yOIH7pSXfOL/mCI0I5AQ1f/8HIPYSnhBbdyzi7F5qUDIsms37hZQxLiyAqCD
h1fWi4rZ4L6iVnvAHIivLXNAS4E2mSs91VreT+sPhTEDe8HvilIIvJDyzHK6nh+pKHaqxdzylnMH
bPrO8MX47EwWhFLF07+eFu2o9pLGe7URa4p05XLrKmFDlXPOKuEJLG1shVewojx0gqcoBv+hZgj3
R/89Qm+rHyHXg78dLuKWbKKLmEPEcjQtNsD2mEE6CO7ZTmfvYYFmBQ2t2rFYNgmY7ndNIsdVpDX1
aJym006xKCFTd3DCNDG7khzxIki6tPBVrXLGnpsXSlx6h5GbGFSHVQ7blH13hBspMsSCej8LeUM+
NAfJFKRPVwXyg5fA7XHIgtce6pKvHm2spRWZllCCL3g/M0/9uGC1T0lzcgxvMN9u/Q36wS4HA/+3
BtmAcyOzsHLs2eVPkPAnUuyDz5SqALsphCTQJGft/z3ChzT0X5h48bPXPDeX5OGA6T/KDp8857cK
P5htzVk2L3fUpL1/JHy1PaEDJ36OWdYW0TGIHsWJoMqeW6qVBznFImWounEsIeeiswPTB/LY288D
CTgRUiGG68efwqW058M5FPmRGcxrSBXQCsBP5V0L7w3IHlBsZHvjFWiJNyJY7RbRILPWAsoByz4d
m/Ny/EbsPPiY9oAKPWIs9vR4TrkuwyF+JnZDiSHwdn4fWuwbzu+wz27aLuCbpMqXNM8u6M7xEvNq
QA3HN2tU3ncJKSOJi9GAw5g9lLFLIMvKEhVlIppYIgmuvco5ypWRhvsNUCdOofOQS4rvQp6Aq8mA
udXpvf2C5GN14c2qrOOU1OEtvCfE7m0XIUONruV6GYcf7JrlT6a+paDbTyTRGU5A81lyu33dQBi/
CkmYomcyaTJD2utQSb8YfmYkJBJSPUZneGx3N9xLV4cLGkgUrEqz2ghg/hAWnn+PnhlZFwruOwUF
MWHC8UYuX50gXHWApHLlOWL8xqNXCGOCz8Q54zK7cjmcSBQz9cap0v6z99Mwc+iDnuJ368bTgo5Q
thW6y9h4wZ6EmBboRTEM6KUCUrz2+/C19/lLQbbhxgT5j6k28u5Bz0QScpmBrM1KtNLH59/xvJrt
3YiG1RzDgVwESFzE1ibGIr4cIeYDzT5KQEUAWoZmNRDulO6oS9mpeHdkLffMUJxFGdlB5Ew5iJf6
rAcBeLQ1T0+v3AZs5YSXmxOEkGHzzQPQDSfe4lTEU15Z/wwFnHTOcjVZldnznRtHdHj6zOjyXNtX
f0+SlO575pc85ZQDFJP/l+bHl1TwreDXz1112Xo79Z3CCLT+ijkXEVHhEM5212wKVk2dJQ2ywaRb
SGb7d9JUTjGTN3GkFZzSOQ/AQo2T5GwB8vV1oWgKk5Zu8Eks6PMrhKbUs/VLwPzBKW1T1DxmQ5O+
m75WsuH0CdP3LCgjRNk6aGK4du7AZ2LtwQWlYse/3m6JatHlsKWune2uFQ3A0zL0rcuI43W/9g/d
lkhUiB/G5Yleaqyq3b67RiOsZeEUdFZp0zrB0H7JkBqEi7mvIz/6e6iRTgGPcrJtd06KcpWXW68x
ZV2xKb14yN66Rjd4WM4D2p0apboYBZavWoODAVg2xBcyE6FZBxtCBwW0lAmB47XO0YdfWhZrlTKX
HefYOop9AE7g9W5ef+hrF29RQ1dAukk4rgzVAJKx7hxVCuU1oqtf3GEXT9/jezwLjQF5O1JavBDG
b4ouciKVVMx8SDcWjDKdMfzJRz6lADAcK4ixa2QftAW/3KiGjJx8JwCmxF0gtQHA84/8zv1KpHaX
FWQGV8iiLmx+HKjEodM2YcbWtolzV7UAf/S6DHOlLpS10kdiufWnwkNaZ3azeQaeszVHnJpZgIdC
xeKV1VoBE2isVthv9/FYstH5Yo1HbOh684KjFiSftq9+YstFptqKUvwLSaFlSpDcDOPMFgLgLMm1
J5Ao0ZOyarHVbdBiNvcjzm4rcoR1iRDrbOVF1fbt5Qj0aqxWKWbON5ZdUxDSoswbX12Mepgop4bk
A2b0C/ty4fLHSGRsjRIOAWg3MAAGvzwhSwt8Ea4EyAlg1p8udkjtAOimP8gAJ9lEkvt+wNC/fYFh
p5g887xge/CvLUkrZDEoiSNZkSrSihCL28VGKFne7tqvFBJHtspgv8Q+bsI3ihpkV7Sw0NO3JALL
V7dXpGSd7E5gTY7CqDuSYpGkal5cGdMHcGQqfK5Vbk0IWkrZK2qx2Fm9TsnEBQqLCvUSWw7wFiTw
dvZvO9/Mi4ofCC2n39ombmbNM9OywnpSj3EbVrfYFA33lTHR4VyLiTVedASbaoIylyGLLIiZqWGx
tJMYBROncv1XJx9VU8RvKhEVZqa6KvkHHPhVdSWrqHPjYpNrHvS9tmy4GxMLqEEsVizpWJXwQQnC
OGIY7XAtM3w5W9swkhNCFCojJtyODtE+MUCd5xPdf3VF/19KJOkLicDXb8lwyC0tTM3SvbXkAoVL
Xmc8biK1E9aK/8QFIfMVfj2/fwdNtwoxRfX0hHMe2tOUkQY6jJN+qU1kqxhy8KQcoTeyWhVrGGRG
WZbdE3P2mo6U3kMwq7hQkLQQiWE6SEPnJZ14Otdl8s0tk14x0XisaPfoUqXjY8PN14w7+ozzO4HU
/qwc8U8VOdRHMo1GdvK+MCQtomH783oJxRiiWhMRIPIkkpkiAoWE93iAss2PlR7xGtySaaGuPbsL
sQjg9Y9z7a7SOfaNoXugIqcgkml71HUHSGoyJcs2LgL+Xh7sH3lNfADpLsk5T+njYadb/hgHYsKH
FbZ2v90WjtMJGm5Id4t8kh0JsgaKhVxiNn19n+T0PwsrxP5SD67mrTGWshEmBU3dgqD3ZbKHCSvr
vke7mKlBFW+i67wwS+KnWL6jmPnb5tvjljc4l84UZyBtdINoVa95Qw3CSvSLoWE7O9Y+TaeQV7er
rz4LsdgX0UkhcbmjTTsRLeyBXXQp0dKF6aNR+GZDA1wLQLP7XZDwenHzJnc56uXeEErulAl7y26i
PT8GFfbdVaSYB5IfpFV/t6GNAi603M6RQ/RcSQIa63/kXt6L0FZazy4TZBANYmNiSwp7p3J0Ud2/
Qkd6JxvLULOLXfNHLxKVYOJMfCw9Vl/6SXUmwwHc1IdxWnPh0QgB6gGqtKZkWpfSZGuoSji30SA2
W+tPCAi1z6R9QP+FGuVu/+ctfPtYxoJdrsOO2YWCXNNMqzC4HFP4jmH9TrwEXaBRwGMjjlKxhmcp
Mddobs3sqNeq53CLGkpm5dWO9jVxa8XN0COWs4sph1NlnYwQrr4q8OHq87qP6b5L1jAfEVndsnts
WM22Wd+yFXb9x0nTVq/s+errGChH9AU6g6eiqmlwTQRx3PdQr5WDw5NMyK2am/afYIwtFzi6Kd+/
auRrnQrHSpTHVEPtA2i80iOUPZ8lkAXCtQQc9hidbMBM0MzzPZFaKxPviSMz5yhEaAD1wjrs5BpP
wqsomGr5c7P3bMEo/ve9SZaL+C8WNK6QZLn7UkTpqpsRpIFqgOaIAaLl5JHJTih7DS34SzUghBAu
Wd251KFqSu8SdHZTPHEwXh8pihiqH+DrMrDEW5TH8FOJmsewdMYULZW+C7YFcwIeWXxAd4QnH7RB
FeG35FJIHd8tzr49Wxf284vi/8ZjDvKTqkjHxIgyyJSHY6zhFnhC0G1TqN38juVIn91A2ouptocE
Y0USmijPddual8VjW8TNVxTkw8FtzijlJT7D3Q9vpl9IkR8R9sPRbSfS0Kj3HnIh3VEni923Qa/Q
N7jdcvjNwzG1ivErCXpRdNshkRJ+TZaIwIXtIq/hCoCfokV50RpHpNthw7qOGMBkzk5Bste6S0gt
+mQ24onvhnt7l8zakwc4yTbZwdmnyVeWL0TUxIyhmFol1Y8FqEqcevnRubxIl/MlkTPEmDGucQtP
G54erI/ISym+l8P2LpHhzWhwEJqYW1xwtF6SS5X5m8b5YGhhruEBr7kDq2vxq/3Yl5FF/TfZyRX/
66A3GtxICfVJ4wLZdBr+3Snt2pq19bPXZRTrRK380MGgWLkiLtSYQfUt/6n6WksrzXT5OViwbeje
CKcNfKKif+RKSHAIkeQEIsccdQbFNvy+4YdQIJCGwrJiiq6Xqf4d93z94lmtldBplT2VP4H6PR1m
5y2b4SFbfdaHavAMTUUNfRnP64A7Lx0vB6BvXhv912bI2NVz7FAatyrDKinspgLBMnZfMMS1P+vo
kL0c6AOM8JToAEZPK8bKeV73wi9sD6Fck3KwUfNMbLPTZqa4Qp4w4dOizdHPbXe3oFFZtQZz2pYU
mM5OLY+W8NZBG6QGXpbIXdzMtjPHj3tS/PG5ad5aEYzdinALSLctp/PPHxRRw/cOBxft5CoHVBxQ
X7nIPzVFAzPw0QW2POGtmRxPhWJTbL1uVrCC9vCfVsCAbEKmaz/seNpO2YLl5QxjZZXmZz77o2K4
jbLE72M5MOPBNxNfy+HKxjnlzN469YmkxWRjS/i8ofKBXCcB8ABRLeQr3p8ely2V22eC6uemYPU0
mdYt4UpIHLvye3KRmsI19cphVJi5g+CPzvG8xL2uL6oPTHO/9nTpsNFFww3Tqx3aOkDN7dnI8xdp
C7VPUV54x2rQDVk+erpJnk58sofFeJ62Ri92KnY1MYdBzh+M13pPeCx6AlZxRmPN9TzJ6jcq0SEO
gyorbFp/6vnbrgFupKXDMJH47eUOmQdEv/LGdnxxNQrrB5o7II7a/hk4z+DsnFbH+ugthoAqHvM0
C1t6DiMar1bVs/fXotGq1FbLXcvpYmAlpKw8vkLqoR0XDaP/YLzWVTU39WGT2ac1o/NnCLb0jxX4
VreWvH/lfBC3SfXw159Ch8Qcs+GMxM5oX5oB6VSovd6TDua3HDCNspPmNNJmsDnN1lANnu8t7VID
x6b3WhqA9ZU9aivQe4O/oHyRZq14xQTLtc9gVwKzI5hJV6MKV9JPXVXnE8Bt+HpMLP0TksyqDZCK
EAL2TLb2ZpBZlOh9AcCmTpMQU2YPiEtmfW+qVStBeRu2OQtmNR20YlSGCYY1ybcRXaNUbkhxidjR
vsLtjb7kcoHantU2veSBVT/lmXSIKAvFe6n7BFaz/1lc1wYBcDAiVjsGj4VGjmRunPyy5dsN4kS0
zuOPJ0ScyfwNPaD3HWMD7GHXMj61o7v8GeMyxW3zPD+UySzonvbTTnSNJvwSOV+8/0Hx3SsZ765R
jPwQZ2OfiAU/Lfwn+cR4+l72PopG+4ECuUdOhMirJA3UqnX7R6RKCaAT91sVbq4+QIyJimjGdlCS
iLsymjh4tdecO1W0Cueu+/Bd4Gz11XrMQrWKxMP4SSYDewyFonMK+a1D9pfYpDM/G5UyPB9eEQ6K
3l3Xg0LNecTIDfhBbiVkhFIYSZAXFy79IPMvqXEOACh+nJ/mUUTeqbiyiNtSiXuRFyy+nxHEhpZU
IhIvzMQSkAqcWroi+qzqoCYSq0izIj/3RfrvnXU3ZczwndqAwLEuIOtW+dKF2Wo0+aNGwg4slgmF
DMCmSs8/W2TCvo8+KcBwobZrWhNVKqnUhy58unBSZvznCsWAdGcueYz4ug9lYoq+S+8o1RmlxYH7
q1EvHuU51QzHq/L13DqIIaMwn4Tdb3/19LMaY30ZkrodE90FSQBFJwA3WWXJuJj496c3V2uJTyXI
nuYh8em3o2TmsjwJOim2lm32aQn60tYbGBge7orDxAfFFRUvfJJVT3NdY3MuQQ1t13S+RKA4ReHE
OJNsRbZr0UP6HOsGIm+VSU7CK/Dm1GP6xQk+LWdYbUggmZUDZ5THPDtup4ZsdVpaX/lIMy5oRNoD
iAkp269Sha3zxsp34E2osycXQZnBeldUt9GKzD2hLfjsylyQj4u5r19G03CgIAVBApANvdYbfRPX
fQPi96Kel5q8P07PHqMN0agZiWRR0cpLx0aDWyXZkA+DgSRxRf/fOeDOKzrINJ4R2vEpIEuj+O+b
NuOu5U2t6obE4+qq3oOsMSksF74CjiA+gU5PgTIf4vrsLH1sLXn5eh4pdG/7s7Xxm3FdyIfOmLw5
JssyPXVwUy6/TiwJL4xkBcFygz0d9DcWWdx/rS9iWrylQBttAKaRgfzYinG/xK3TLBJxfiHfcyJK
bQzK7TNYkZm2Fuz4rhVxS1k5d4nvOa7ZWvmliezzlXLN73mkzs7pK1a3U8k62KAGlNSATZ67TY+2
xK0+8BQK6GEPaneJ2LsQM/MugvEsU3FmJ80FgvKBoWXS5EvYEgkfR2/pbFviIYRTl/h2NU+l59OO
XXuwnwhTvg6JINES69SavUhhZBmU1H+0RmM5rEZTLkKHYAyfxmssTT1nE/kp+SQ/1FhJPrQDdR9i
iaNeX7sLw3CXqOJwV0gsZMY2ftMRqvsnEgl7BmAI85I11SpeodZqNq19EQupKP1TjMWEL7WSoGHp
Esx2bZkoA6TuNKAmVgOWkfCkkmdLLEMAh/NYRr034bdkICmnToUZFd1Nrnw2hS9Sp1ETMjXpoZ0k
gfu6oEq6xUf7fyoQP1lh8ZbSZiktSBj4uWYj+Q2qZ4vjUMnKpmJkJi24GJZSe+hRqSpHdLBAGKf1
smRF1xiCSGFky1+Du0sF9wSIticvFA1EeSJE/HRUGNyAYWN+DkBacqNNqsj5vTurecn3Tj0FgsPj
g2jtaxARd3qOnBrLYs0C9z4IfbLf3eMO4VIsuwJZ5FtcVmYJ83E4Vw0cFA57YZE0nyL7bkmj3ZSi
mRIMhKC+oPd4Pd4UJmcNa6h5/KImiKPJkE70kl6psh0ZWqZAtgU0z3geeL2xjnfZk3t4n2ueBdqV
8k+l7w7pSoyu7DFmkGYYuAKUUsydleUm5Fmrmce8+or7h2DBFUcYN1a4ozI6T0SopgNtm6P8FpI6
Hja2Ai43U3mKEfpO2JG/RKvZSIhgLUL+olbNDzAyfImAIhYLoLn9M7X0Q4MaXfy5CdTP4d/tKJlz
lC6+5SlnMvxWjlxrEqqZdpwon63OWMVKZHo59FUA9X6qQxpR2NBo90n6S5kKBIGnooIdH5/dIrUn
5vhue0/03xBlwXUaZbS5WSo0s5I9R2v2OPzzTtAPuRr64NDHPEf98wzvLJcSoy+ZgAzu/wh6U7Eh
qj4HPFAxX8iRmTc2CCAV9PFmEVixZ7yZ4LHS/9Z9P4u171h+ReHNYpTcbiK3uKPxnAGjbr6zibay
zwsAm9GzP3kuMhmhCrlxef9g3SCZyodwbtDaTOhkpnKCbZIJp1rWcfA7Jtqm4dp++9FMpyalBlo5
6yMnuWGIUFSk8pBZayr+phphu3V0HRNWBywYbmjibhSbU8nD+AkhD/LAa6Yl5l72GLZlxYgerS2K
0u854SzPtzfZg9hjnlD97RaH6XgN6pdxsGzzfpIMWrA7Ipi2ygldJYgws5ufxqnzUV+iAx80mcHH
LaEQ3pwdbmW1Zo1ucPd0KSOUoJS7VpLhxfpaTKYAs2Ye2vnGTsfjokT5V1F5CQjcs2VTMZNBATP7
VOpiyrGcV9QZFAjC68vzi78r4RDbl1oVD+uMCE56nAnLMLp8hDlK2xpgu06tTNE1fLKqPMQvXz7N
CQ4i0DkyN4i+nS5rixqsf4ZAHYQkX+kGQrdzRReSY4X8iL9o4Ljps0IXy05kDTHhv8HnqiwCDFOg
Fb/RxB/VBKiOg31asVmnPtzmfXuTGdVHqzyuxX3UON2w8XjyrbZjje705iTWhHIFr7dq+BMtECeG
YvCECyQfX2IW+2NQnzLQFHNX4GOtcSRNeJhJj8AZAHvrGyyWwMBV41HfguSMARr/zLYJjfMWh9pd
KSm6mND7OlKbaZDmSGczNO7jryurR+ze3v18ZpZ2V3Tp5fP0RVvSDCvbrhVUiVPDKMQIyqsiUDaB
DVJYLOoIxQbGA0g0UNTRsXWFSV2lQZP3HRf4XKOh2hcxWQfJZ82NH3e4NvYAW46yz/c7Ypwu/7x0
8/pc2bZrceo8f0b3B02zys3ceLV17vRsqqt7IbZZkBwly/7DqrU94jB9ldyAEcJ8pxmvLHiUowP0
ns06KxfdNxq7ZT+nOPrm4IhxfNnUta4UBoaihSkE5ToNikmNysiezGh15DdyoBLenTgcIqzyUJPA
xu/bZskR63U9Zp/cDfCPKBuHT+zefgxuFmXpJdgwjrwqhgykNAF6JqMctECYAhxWAbTlC0+zYJPW
EBDe2tJE0G++kjSFQ1jSfCFH9MDebOyxD4O9jaG86iWj4jezAPlK5qCWbdxcTBV9YTPN9jZU6209
y8iT2odHwBIsMPrAiGweely5pKqeA8qtepKBfbi1JLd4Fo33LwZnJTX7MIb++QmAGfEUYWmF7xND
XylGYQUrEjXyWUSisobPEfHr7AH/2/zvoem1jbo8tqiQwUu5nlN/MU8ojmGg1jKD0x04qd3SQq3z
+SlU14A07K+50TCSDjKKd3pxVoavF6zVuu6wWou7gbIzI2eKSfxdFWeoH3NQT8uJo8S5D3bQpNQE
isJyVUxz6+JnbAdx6mZd3yfpfN1Y/fwFp407ifUJSDpqgzbApI7OxtdEbwYXbvKbfM2HbZr7cP5N
/1CXxf7vbJ1djAf7OTigiodaQ9kPZQoaOUT8ykx435ddhigA2tK8OWvCOsMK7ssdLL7C+4e1b/js
WVO+PEj+C+KrB1FFc0w6MrM4c20KkgJ8xxbzzjlOIM23yx5wsfXgWR+Yn0dxVHUQThbofcWH8dqw
Lfjb6y2bgJKKQCYW9C/eL/YrW45yXs8I5yCLarL1RhXB4sY5pIjy3xcQbFRe5bnNvYgNoxDo2gD8
wK6lq5fsnIA+mO5f/0O6GHKbC6Q8xHxOIi2h9Q8QTraGm+Y5MTsLqcqgNioPP0HUU1j271c1eW/k
f6ruU74VebMqAo91GWXuWQ9zGWaQi+i1kPn0OEBeVzRuU8zkVG789z1WBlpVXbxP3stTTVFrkHto
WkGY5HuRm/r6BhbWV2GPkiLwytPJ5evGr2Vtwehe87DK5hMCb0RspYeOiCdgrs5sMnvR4oIE3+1T
14KOwtloiQnrEOjT5IW/c3WVVNvDEenSDvV8RDJxbBpvvVDkgUAENz6qC/gT8PghOapdY4cUjiQp
RQ16n3nvGX2x1/Ld7HLhm8wR0n8UzZ3UDoIUsZUKfLfI9jDyhs52pRaPVM9QtoLiG1Xoas1poP1t
Wq3KqKRbJQ+PlypB+VvGkw6TVG1aoESp+sQ+yYjAqy13iC9cOK1Y5nGF+iTNufeEPL5lDT46QdUu
le9dm8mPyLl14AvNgg26gScQrUxvAUXcvbilkcaRuoBKSuZMLKeKPx/mjdk0u9Xh3raNW216yDWq
eVBm/wQIwUgdlnpPcN+deZXtfvK4shvNnvgqh6uo2A/WAc7SedcHafVrBiYC/20Lla8hbL4aV1lF
ptQj8KDOlIb5iBlFVctEZKDiuHWZgxJeea5EKsCFQtBXrHIaJyfEKiMlapIpn96apEl7kmaPOYUu
vuLmDY54vO5F3V6v7uadDXY1JteG4T5avlb2SGxrVJU36phKX8BHvvtWVnMyRY/r81bXYQcsZjKW
0Ji9BpcMgrIVOAT33TJT/ug27monRsFZu4PiKVWAP5W+dNfvjiyfNP7a9F1HU6EqzAjwfGwJJUPB
xSZR5YRKWFKKevWeqcv+dId/zdgBnoqzR0tWQ2oKIPHKX4YSBEBH6wJIigOI6IvQYET629LryUaK
POtTzTCvYODn37WpY6uBdOHbBy50XqBah4nIJrmHdtGDJcB/6NqlT6zX1pE6CdJpqv4nntZjh6yw
fwugNc9UiNs62T2E8j9wHOHwwzzvefR94ttdsVipXAGOA+I0vGWkclE8NYCPPacd87AC9S/GFdYH
t+RIAkVX+OFCoA8By2HyxU2Wm8JRPUbuXnzGlb9TklUJBMQsgj+KUtIOtrvnLqKxbomd0P7Znf7n
dZv2bNaSHIQROb3OyKrwMKfwR7P6wr+f0LptwFEMKfcV+KmwmdKp9qklsVzJDqQsFz3HNCL0Qnh5
pXrnEOu+EDJFMU3/yszxbviwI2ie3LodcERmrYTx4l19OkcvjIPzUeTUjSP+prnnhhlBaS/FmCM7
X6w13jjpVdF2j+IpWGiFffgn9IPniSwZhFV82kpVByNT8vt0IbDQFG35DRo/OMSgrIsuSjR7l0lA
tlTQ7nTywuSAkCqXrYU33lycqVF5YSXeb5pX0dSp81tI8du2GIz9DH+R5ZTOh2cxfaWDiN1Ji4Sw
OlW8xQBMyqk+qrEKcTbcMc6kyaUi5ahvpId3cXwFsbXaDcxLw//yD0oogleS6k2MoKkeItC6Y/7F
erAm5m1Gz+uzWRuW2rP/E8B0iQBaW+a3SOvHttPsXdErrrnnPKNqA1jacn8wkXmINxOnsxJ8EBVs
6xylAJPcfR/jA0UlzubczJoOtejubwsuJvNA8wTn2kxfEDqOjo+UpRMhyrZObFeOcFsF7afR1uv3
SsrD6X/Ntb2k2+2PvC7wI5kQN+TNvXDn0Fi6kdgwxMSGay/9qSb3RgG5oMjicjAhraH8XaNit/aR
RVagyHYv7Hpb8zVHcKW07oOcKS7GaDOOG6n5KMMCdW7D0l1g8or4QQZY/egO+X2i359Pt/CktoA7
yFk/GTArbkWIjmUOJbFx7Eg3xBVGnT1gc49iHCVwPEd4bkJa95vzvOKCAqhapLtnI2OWyG9rD3HK
r9TgxaHwefCfxFAaOL3QYzOhYiAR7yWhVE0B79ZuOL9dMVv6Igb4CWVx2CFXV0PwnSnvrgCrYrSa
49EZPaANVLDNUY/wIFjk2zNy0u8ssDSQUzkcgVh5atYwwu2CnISADaAu7QyvKDkmkM9/FsoMAPwu
KEGo+dcUIVYBpisJl1nZyw+6vIknxJQZqQ9jOXziaI+g9AQmLQFenjlEkyiafoKiK6rBJPM3YZUV
kv1S7EJd6agQh9LyrJaej3NYlWgISfba8QuGadCxJpl6r9nmM5ALzdW0TgOesnRxSX9jZ8eEqD9M
wZGL5C/mecIIB9Y2DIF2GfEw8q6REic+4h/zornDvoW8bvgY+aEXBbM7XoKxjHo0wUGiH6X2XCVq
Nn1opGPR3PP6qC/ilCTRL369RQV8Tcmy9G6/kmiMLVAJYu28ulhpX7P3+DQmlu8XvnJm9O2L3rJP
VgRpsGezRpyyb2n1EIzyMm7FGkw4P0Ox1oR1YGWjEMUJdmcNvPOkLXlhBPt1BTf2qnmhIOCK4Q+r
BqnoZ3RhX/utNmjjuzLOHB4nYUsK5K2iXfoaezClmRjlluGoh2uUIiiHTD1c7DLG/GWbdN1QDvfs
bbAR6sJgJ8NFdmmW50pNuBp9cUpJhURKWuqYojd2NRogO8TepwGkXY8Nk61moOuTlBxJqJMDlEmM
12MO9bj7OL63rkzP71vxTm3Opgkb3NEKBpxf7qpz17NytopxkpgHwyIU1kiOVLWqM3IWrjjLhQYU
B1gkCnkm45k7j/Wv9vLWYzm4WvG7CZjQ1WRysn8bjboK64qeWKk417lYStAbN/viWjfGkftFlARz
9JGYL8Umav+ukj0oWn/9HrdzUixJ53rpm3MTf8BXKuo/9umUdEBFzam+28Vic6QMyl4jjL5EMMUs
6AXP/8F8GFhAF5EVL1QOpQ8ygOyztVJZKC1WgxgtAz2ggfLtVzGt7XvT6ITbq2Ej0eST2VEUvJRe
2fJTmkBLxvPi8hAE8iUiENEn5PGfQlp+oDW0cCPc2moOjHMN75vHdDIbnbJBkCCNnNVogGPtudA2
9fNo++rM1FQJhPTLrWFhNMuLdU0F1TW2YZi9JJPczxvBbSsBkBMUpBak8+pqdEIQ4drYJEr3cAA/
+oBjE1ywrD2DX2wBOcL41i8E4Zcf7+YrzFRNvnnD6M321hygJgS33LWdyxj/ounfCDeNr4SKgv6Z
IIjZZqC6n8LnloNZdH2ZQTzRFqnbvb9ljIdFRcpAw5GjZ3zKN2dA53ygVigFCXaljQnx/1GczYSa
Zv554kpDI0/XzgtsOthWI85LjfGk/IFkurG74eOymrsEB8hhKaJy3RKwBGXTcECjwN+y93GlpA2o
HlkMmqH7Cve7GJ2opWwsVX5F2KZd2C+sT9+Mvc+d00T3b1aJR9nD3xksSdc/lmzFQOq8vb8x0s0O
YELyaFYNTsHqIwYjxFhkAiyZk8ZN2Kx7a6RBtksNA+mdAEzqPvzi7At1M5OK2NFYAheOWBonpmWZ
yjlJ5CvNYBA+zOm3hm5rJLQrt2lAbV2IStVbu6KIhimuYddjNQxlOk1SDhqEXwlkVEFEAjv0OCyY
aupOek4muRkWr32fVDld5I3x/27QR5HPO4s4Hoxef+ECLQ8YBZp3Jlxnvni+FnQ4DxlXPjbDHXGi
9ZKsaDn6VbAdQADu9L2HdMxxwGOK49jKP2jeb5fwrUJCBV1Dht0f4Ws1uUe+xuJYgsadmEqeD5G6
alHOm8MN5Pz71Y+TUlXfWkFI0ah/X6d0k3IkM5eHk+QD1FMpnLHvWGYFlfTQ3KDyQcMYrUPUIz9m
IKQcAOl9vAQ4h4Xdi5Wdw5AEC4WpGcbxj8h2m9QyPfmA4xlevBrN+q/QaOZRAa/JuwkReL+Gyset
xt8t2vOcTL6HoVnH/svSTYBAR0NrAUFcoxUbSyF+Brz0HEsS8pb/09hUR2UO1RfuX4qmdQd2bhF3
UcVSq6ajISeh2sDlji7hsBH3rDXHclpfTidKYvwwo0AqkPuDFWC/d3T6CK2Rq0mVj7W3n5u58HXA
yXJTBskKA7NheYZT9EX0bwBxJfMAJd6uXu0LgrqvuJyLdXhAOPlTTXTwEBoEQzFTVusFS9ryMGF1
u4RtX5NmCrkofHCMxbADP05wJw/kNqfiTozn8l2jl5/mmySsMG96U6/xebCWfnGHk7qoBRYxywIm
37Vk2DdFyNt/jwGMGe/Xu3ChA/KAi/sHbpTpmLGfXhcqomCKTJi3MPZrUgyDr2romkM3HQ2BeiSD
cAoshFmuSpuXuo9kqT7AMS/3DRIcdFhrwdkCD7Sy/Qsw/Nok0Z1qmmcWufetx/06r2skpoE2XwlT
JA5rF7PlL6XCH4HOu6uPoyMLO68W80DK5uVNUrTawVD5VziUffFFK68zcUWAxTWOit5inY7iPGqN
XJnyZ9JGkO+MTr1hfdI9Aqs9l2ELiM3tiaS/k6To6p3QMOHjXPXuc8C8Dpuc5dSH3PqgOiROzc+e
cdzANTmIHKvmMdwjTiLMi2RtQQdJSjPpYs4vDHtUd0J7o3hJmCwsEXZoJdL9xV0rthb2PoxCDCCw
zN8V0EYdHdNk1OgcBHsJdRoNB6QyFqWw1g1toFXFda9c/dpuiB5BptDPsRDGrkymAHnjtdF4HkGz
1E+CUYWRcwreU8ueYg3ZNou4VJ+k0EgOJaxyL4QvblRRCUp2HJj3pP1zYZF6lNabRtvA+4aCFixZ
NtwbpxM2h8BgM3BsDwm/7c2pKTrIQN/UvthwetDi7sGSNL4BlGhxnIangeIC1kZVKzHrJFstIqXp
G+INmkhZkz6vmPqv8hf5jHUXsvRRccFwR1+vVAi4HNJzz8XMP27lNpgGRb1U64wkjN5nYEphoynb
b4eB1QSFn/w4GyAHndNCZan9MAJbhuwqoSJPmjhU+iPkMhlNCBbIQL5bz/xw9TUyKSMmKzZWs+Q0
OEXVLGrHDgF1+56HYdtTyaw0j9wK7l/yhxCpzM0JyHdPBmf8sNea7msHnRXv78ySvEe58hh6XZ+f
iBIN1MDX01kCqum4Z/gjJo5GkLpIMJALcY16vTxTZdxqC190Rx0zFgMvwszMFaniVAX5TtAojcj2
4mVVY/eAJSk0n+OMGP8mJwPpRIqrpWzU3rx6zrT6C/Z04KBQxrlhSAndvvJiGt313TLlgmEjuBhS
jpY2tgmER6Ba+9B8v2eA0v3zgQlrlTS0b5RxU/upGjVvEo5NE2l9W1xCKyCJX8fVl6gQTSN1rnw0
po0G4FzyVm7gl+XNoF8HWzENY6K/Cl7L2ZTfh71utOKujnvMFs+IT3PjgLanm43CZvQ+AG4nnagH
L228xpBSESS/WYGWOUkduzq2tB0a98XtcrjGnppvryTHw8ffzIl26NKdaQPqAYzEYNUZrHMJwz/u
kZmojtMVNJnrHAoxNGRpi06HrL5PlxUmBtvE+eiRn+/o2q9Cjlb8YcOdNM+3pbM8DACbGcVT0r+b
ecqCtESUOxSScwbiuNiv6o/oozphCKaKElf6aYCUOF8ef4GDywQgXLcmqGSCvRXgcF+zV0hYNQaq
g50yYUFxpEAIRD0Bs949sXWI0taMKcijI5PT+FPz7IBoz/hj5CMBNKLXi8Fh6eZfYVUCpn1rFsv7
KQbunqce/zFg18aIpkWnBbBzNPhwlKqL/C1TP5W3iApDGPiZITtmSWcj+S6CPWK7mDu+RaqwWsz1
VCtdMtKoBGAiZW3bVzx07NeUaDskjUx6Mcbq07ZimReEUjcbO1qaHNH4HXIiY76EHtrk9YLLgcli
a0udF7GNpUIF4bYP0zkHkAoDQ2sk3MqZHYdaHWcn6zjvrVK0mfPq8vAQHXi9f04XKT7mC9eFfJMB
ML39E3H5rSWijw+7yTAPQrNvxRqobYRKIQWWCaMVdbhA/Ic2O2TIlm82z8n3R3sN82WimhNliZ6Q
xKgBf+35LkeJA0fpoK65UNWk3BV0n/R7Gq3ZReqGL7rPzW9quEZwjLCFyMaQQD7RcNgoPDZYBVS1
lrzEqQQTl3PzZTRhoLZmRYvKnr20yr73AkNbVrVCGV2cFhidOu3H9VP6mVnHoyQV9N8K+y5RWqt0
6EuaiHq/rTqjKJHdmChG7bPQlngfW9KcpoQAwrd06qWmykCyvY8n+F/L2/CnRKrTWBB2o1Y2LBv6
RQUIQHh4Uirqv4Bd0v/Vyd4dCQf5/ufHElzlvRFSyBM8TryJIxlVfkEwi1icbIqrSr2EpzvpNt1s
jLQJXTfJ6/D66opl8VKLLpj6B8HZTr0Z/QTKPN0GNe9SDufeOFuPkuN9zboPQUzypXyYdgq+J6/i
y4GtnSl19vpJY1VdpEw11xoAl6IYY1qpeOVlJuHxhqiz3oPqf+8jSaiH+opLscQ4t1+NSBhE1WdB
jl30k7zforn2XtFnv9Fse2H6+rhKueLzPDHi6DFMcSJ/lp9F7s6R5O9FkHmzJI8P3ZK5qAF/7HM3
/2L8pa6zeoZGoL0KhHJ+ZCcUyUR/9EfzNlgGGdTT6iJvw/FWZvEJyuiH1h3+BfFQnW7Ndo+Hof3X
tfmtl0xEkkux54aa+cH+eVHtV36yFK4d4FjHKtxApkzJksPzNxJt0+9+Jp9fWC/Ahhv7vSG+2E+x
G4CE50Xqt9aqIE1ZzAjWICjn0zumaOS/dsLlMIlQe8AwPBgZuF4QW0zm0VO+zg2N9IAzkTDkxjLb
J4GTqIJRtqZlwU+/fUHoOxfGgK328sK4Ye9eqgiPipc0Nc7dWq2FBxNdK+L+xrDgS/q1ZToGTxOj
HLIyZH1eanmStuhshB/ICI8eQXsxFFnTNbAV5YFsYSbwj9+CmYdpPcuPLJdK9rWdpsijKY17wT8C
m0HfTjfClU8Ph8BP8lCxsx6uxPkIsZ0WlCIuDH75zESMyDEHDw3yzhPU9C6/SucQjdcKC4/lnAwH
GI9O12m7R6z0XSTNrrDuBlxZc32hdanMtOGQUYHBM/g9Yt7KmD71G1HwFuL0l5Jq+LKFk2fabAgZ
D6BClksglkwWlllJIb6U3wdHinoZKiUELQEkUVxBxYWci2NkNkuMcWWbafITO9Buf77JIih/M61O
IMa3TqjgM9ROnzW7zxZPpOwCiim072VS0vnltMC2jYhwohXVTpzTm6aWNmzyB+bbFrIK4Ccm7GNc
kwRc+20aUL8oKKI6NWZ2p3Zrkd2X6J2iUr8CVqm9VV2JOoSZUFoKJSib6N5cKHt3/ILhyH/o2BYs
VgMKWVgwXNektH2cz8TmuNjvrFydt69BQfwKJT+WunDHj9AqGyZQEnoa8Bf3QBInUbHlqXzlQYVR
+T5SFkqmbRbELhIV9s553g/OhZGEKNajpWWw+7J01fAdOhAETMTDt6gC5f+hKZoFhJMZHXZ+RXyC
T/UWSHQY6qfqy+M6OljvjflZ4tvHKzSHKkdvvRQ9VX3J2eBt+SoskIAHSvmmRyumofVMMgy09d1a
bEp3gPnpJGmjJeErgowbpx8l79xp1X+7aSqbCH0jjjOEAR0s+PLW+gD0KP6W36MV/QPApMbCHWqr
fkY9OJIPw2dANe3/dhyM3lNGGNjJ+Xve44DbgQG8SYas3FNDSNRmRc7F4/SgZ+U9+pJtZ2zVLrzy
9JtDqct3r+AsxXNHDWmsD2nuf4aXTm8e2tfyNETlcSDN0HxOzhef806NXKnggtwrorH0YwX+v8j+
/FeDBkOXJzOzgBPfAeU89BxLm+MRoJM2iKM02QmFxry4SR2oILH1btOzu642/ZK+Y+4U1p+vkyHl
H2NqI87RPHFFdJJeAmZU7+OMw5vPBF55fYKVgezAXeGuOY7FF5ivMGqak3D+Yqc0YVNHFmlF8jqu
O5FZZiIO5N/0CNgEehZtKLlA9TSI6Vo0625CupgB1e6PkuS7a9xOj5hYt5F8UMwSSGdYQYAm8u4E
ryMpnMpmvdFCIO+6At1riq+btSsj9DrW5SC3qFDyySXf+4745AhgbhvtT9cmNhu2z2yFoDRog8tF
EpdIk2tIW8gOpqzAdPeP0ySaOPpECeYLoIQXY0NTlfhRkuR02KvspBazWWNg125naYJxv90Rqpzl
Pi80sl88Y/7zAv4sOcN5lingX4OchA00RXxpvq2KgsOr3Jvx1z2zT7yJqF/m7M9JU53GZwL6VQR3
becK6ZxjbkrG8pDizpEPKogGaXlXARaxOHEeGwM0t7FfZtZmJj/gEu2skNqZfuzE0wtHaC0xPCrT
3YeR3HaIRXKIr0PHGtFQJF9k7EulP7yYDkBtwRxeO2Y9/3g5kky86rq1q1OJDG0W1H/zdAwjydcA
xsp5DZKVFy6LMxE15SjL8kxEh/uTQ9koYtxAaGE2hVas6SLMFtdm/ppNM2WdwkcGiUjdISKduBAP
MuI0jJSOvIAzttEJ3Xx2DRNwoGBmQkg6e3bgRADONHhPcqRChWImHHd0tH47a9voF871fLDFoJ7+
xPsA7k1oVIPU940xOsBXX01/bCqta32iDihgHRimll8CSiz3Y5ohup9sOWSx0zwtCRw8nl9r2baT
s71RYjYQDGiD9s/1fKCKd3ch/WxwVTY0gTW+DoDpdYTOlB1LgGkT368qfRV1JiYWm+NWFyteyRuU
B9epnf1ZQO1gZU9LgKr6cR1o0ik1zKvoZrEhf1t5ze/+FelL3LWisxxNibWrFkDQAU5XCs2d0fsy
NBz7B53WUOqaM0JyoVrNJf6jGmjS80+paRu+s45GKGydkY3Uitx2R6+LCvjzWxucGxyDm7CNLw2k
jvX1aprosOW9tpAZpN1Kf7Hj3HQZjW0nr1NOI0LRiNH+YnUCmAgQnGqDCKc/wSWWzEa8+xL44S9i
wyXmq49BKkvcz5BdUYTp0esGzJQGva+hPqotcRx0RV2GK5fuO9QuF9t3WMhw8GAjBMb7Q5xpoM5C
5cm+uUBX9LiGL0ryFX1I+rnhU/+9lZwCLUpPJFC3VQjd3t3K90yEsaK5UlwgAzUx05tmeI/Y+Q7e
DmJlTMQ+TS/esR2pBxOROH9/8+UR0TNzKwMtNhZ4oJTbKlTKeHKazT9onBgxZz6zbui69Pqovh1T
3QcejFhcW7Rzm9NdaCpilJ/qT2dlyAqwgGsfD/pFw013GOqmyqN7LBk9eoExmKeQmMX78S07VWY7
o4LwbrcSC0He2eU6O43OTuh4h8qKfIkHL3LwZJXnaAJ9HOLjJynBZUM709/Y161ZAgFP4piyUjhT
dm+IZzvIJEFvxApvcdV8M48Tu5YnV2l6OTSTrDh1DZqcMQn761jiwpGI+pVnaZzehCijmeBMGHcJ
Cb+qD+sjlPyNBo9d6LjjKKkHuagwEFTqGSDIWNnDYzt1ugfAJRLALe9qme/EHl+aLba71ksh35X4
Q0lmEQx1C99jfhDEieWD3pC+AmswoyBG6qk/vJ0pboknN8geXa0ydahaz6/Hi8V1+RhJDuCgZrow
QiHTKcGdyAZX2ZbUSsd5dKWkdSGif7Giw7TT252d4dHrSGcic7KiHh55pyE6ekRfbILsZi5RJQVg
oj274K7BdzsXSj0S2JEVw4eya59AaijWzqu4oN4bfJFPLWlkZOXNMp6JRRgeIBwUL9V14VBBHS3v
CwwNGsrAVFoRV+iT0Y4Zz4AeNJjodjAmjh9On66OtWJysR58jxPpznwVDXhBKb1KcLamydzrXA5e
3GoXkP5jXWaqnBx3TPAGaqSvzyUPGq9UgkucOz4nbco8yjJwRS82PgImdzoC+BqXFtEBuV/+G4fZ
nc/x3aJ5Je/wl4RYykPLOyXml8NNwmMdmrpQPuipY4VQMezQZi60pMnpbd7LY2gC+fsFInu1Mb7Q
51EvJiPIanGP0Q6PfXzIHM6TU2TWGBK/vLK5l1nDQ9xZYoQj8ULyqeQAM+mRggpE931Mlrsn1j6f
wMTAs/yOTmW1eXM8I9txg+zBrWMJYrDPYn91bOXZU9XFAO0jvI6zxw5MMIehER/8zPYLEExN7YBi
q7ErJyDgQD9rnVCQaCaohf7l7FKFMsBp+wduVjRBKvOZUwwFtW0BvkziURSQtkqyNw2Wm8IYPzNM
X/lbZzEjC3Af1HdZg+XV87NBILJZvEpj6SWiTij1zBPjgzEkH4wuTB3RC/JShIEAZcGeLk/nfzTU
0XB3RduYpD0jNGJpBRLy9Rxo8y93Ova9EaMG1eolLx619h28ZiAh9fC1qE67dm0Vr+9eCAgA9KJZ
txgN9XJn1Y+6y19h6Asi6OOSUqZDvtjubEFaX/f/YUeBdqoDpKmuW4S+Bdodi7AgH77Pe6d6HdVU
BhqRa5jDPvbuKan/OzU+8QdJwn6vDMYm+WtncxgKA66J++OxwrV4vAT4FkWUfeMiCxn/5DnyS/T4
BSZRR6Qf5ZvMnxOCmkCL17xdVykE+gGSNtZlJKM835TvInYzvGavEPoHvkGPvboI3UcrsNp9RH4C
lTKZPdHWJRWjbd0KfL45vjoqXTCrBhbWWwhhZtSurYpvdqSiXOzxR1zzTMfZlc1mu21sGuSq1Rlg
piQ606GUFqKSq6XynI32fnkbzHb9QokWUFQBqgELbes9FBHsvAs8sOLxZe2mevHdaR1xI7+BqDIx
cF61ntv4Rc/Sm3jA70juDWdwfLXsl20Qr2gEjMb1WM0GthL1zfunMiX5+pqppttRc2R5NtCc8uM5
E7FvIoxE1hRTsbRuqIIFBbDvAlNuZvaLuFW3OHaxm3Qn7Sjx1kfWarZvdximC67TxHkIHTUzdXyK
IQqS8Pf8Sdgkn07wG84VcBdvXETBwhwC4dPd3JpDluLP0p2lN2+/rnEwcbFVqWzVszfN0JGzQ6fJ
dkXs6nHnYh77lyiPo96RcZNShXg1A9hPFtNLtknWYa74a2s/pPfGfH58fxOxBVOhwr3k2gBotOXD
D3t5OHdNBpFqW3PjEnWcsOgUkzu6bm9hLDWA0VxEzMhmb7fCG4+xpY1kHTZxCVZGuCIpyo9CeRVk
jQPyhO343GJTdabrC0337DliXxROeOYzgnlGk4s9dYvJX/yJkJgDXycWQhNkFuQ8MZkEvfIwatTZ
kL9G6KGLZ8lB7y8EihZR0R5NKri9lx1A7SfNmyl0MwiAre9dFtaWHD9Feg/vT7ERQGD0twkhEBke
2sBN1+84VIL4BW1Y355U+RzN24ViTQ14LEB76uLHGcsfO2WB5cK4nIIauhOypRNa5rg8d0KYyqtv
ie5wqvy4RtmYU8OacdJu/nu7L+JFQjHEu6e49jMS7wGJ5R+Vic4symRnpgvbtjGZdRXqfk4ihgzc
wCxULs5cwv7z7pscfgcyi1VdmvJNmGlj5NbRtNJ0LyvgXKukhmQqQn1BqDrA7UYr7mW+cbvH6FKr
GsdDkBr9dhVIV753svVrFXqPuvNimtZ3yDsu2JRiMLuR5rPVcWv6+ijpT8J7vrLmGpbR8pWe2ab0
wk3TWy3YiMnkzhwwsP1e2XLWG+d+Acwug2/e3pkiGkkH9rC8N6hKxQqcYdte7IZSDhII+7mtCw6N
Ipa9rQcJnW0IOF6wg2rI/TbvPW929JVedW26/z99VcYS6tGUv7xPx4QO3uSQfPH0OhtMGMSsxM8U
QAeuiCp5VzkWOtWDbvz14aIg0HDQOi9orx8psLTHwNbkfDBkZv/qDomKFj1xy4XcYuwQNoN6jryO
cr23rbHRe1+5f1FGPst83kR1K33xBL1PRsC2SixdNFJBANS6Sswhm7QDBiIvCIiHlfWN7iOzEt/N
st5RhGNR3+PDdhlLhD8Fbz/QanJAAyMx7CuTTlLLo9N08HY97A1j5YF1+TtD+xTBew7zaM1cmDGr
WJ281v1hNYG8m56Kw+ZnONySEQVBYrQduQ4u3FEjGnEFyfHsvEIvNOn5Xgbvt1gigd8Ucsqp3Zvp
2GMkh9v5cmKSSd803GLPyJ5HtB1yJZjqSF4oPlvbq0OtS5x62AsJ2Z7/MjuBRzIijiKnsePfWECJ
LZxWv4WE7pDYI5EByb+lefEL6SyRtGRPPlyUYzWO8E0wn8K0xqmp07O6gADcqL3blN7ZPxjt7pBt
EyOHBARmcNkHJCDOAzUOUr6uV+71K08/WAKmTPm1bOR8vAq6v2AfCMsQP0q2eq9pd23aT0YYsMjm
75w9E18rAAema6EmEtabvM2G4JAMjEiDqNjV/OQz23Hj8SOytdWd3uFVKaKgF8tnkLB2f09I/y72
O7lI98/QsV1Pdn99RKqTSAVNKiA4PGopIXsC9QKu31F1RXWAY3sHc3rEB1/T76ejhjM8RQYCxj8J
bro7l4Fkjx8UKnzYHSX6G2cIPmC/PJkb0ChcfJrVVXOQ1sd5awQRW43MO1eiANWtqORqfW2tbN3z
m1jG5epZjvcgAt7Uq/UogP/8wvGZR224VjZyaa9f46Spyk+et76+i+imWPuTte4Uj99O8NIytNRG
WHa5JIeAgh9GuKe6uPIfzLxQLlDdaV1t3sQt0IXIQqJ0VgPdh/CdYJoQvXhBmCvcgOLrSAQfnYVF
RCLBqWDFqUQ4Ol+KjV51KHv3nYxFj7eC3p3MRPj5S/9cy92wOppu10rSEYbtGU3apQkAenbXH+ak
OBTInSQ6pfur9mpA59H1BuVXZfwW/UzXJlIqS12Sg5koXcqNJRzRAB64ZU4u80NjU9Y5sMpMhI2m
U8GnNoso0jBg/XOa8iEQPENvBFpkX8sXjSPwt58fkfPmK+qPFtt9fEwR3gMgvDkMzz9/god/zbz9
iUIt8/gThxE7cGP9N7Ds+1IAyVLY1nM9eAz1moUI5/KJXHWeNfcMYkm4UTBMqqJwdoaPg3QsLkp/
etIF6TZ3xME57d5Objma4OgHPVlWoVyFi3wF1T330TD0tPGxyi8yWRl4MirzV/bxUhEyj9AF57M1
yzJeA9GP2J6YCzvksWGjcqbi0y8v++RyNWvT17gblDbSa/SwP5z63KKitzYHpR58oVK4yAvLu4XT
TCSK/fRCv0IyrjFESxx2W4Ug/8DWvEzi/+ISPUYNjvU1W5ljiQVQO51GvMrqzFKx8slUdhSAjGyD
0nzTK/RyTrAellYfE0vNP++pfzMjj8PD80znWnVkNeZc2cvKOHDaV6OBZIxHXBbKPQHRq2OFLLPg
8gN6HhFazZd1f0XYHJ3tL/LiFo/S7OWTOKZwFJOqwX95m78dbAwAj0jbRHDNXTLTTxXLjiIWmfuH
6t7A24ynzkNgsKCYxVzrcp2Ij8caNVN+QRiMFlibeZPi8jHiDyoBlfzIKmtQACtmtoxbLPZHRkYa
F5/3aVYY386gHf7DdoIN8gwnLh6jmdFNWonoM0egv1MTWi4c54n5mCYtXgevub1THW3lNNGVh5LF
Q0P64bDWg5G93jbdRlvUNa8VwevYO9ROVuPH697FdBVtrbt8eMl5IPLSpQRRXgeAZlHdoi615SZw
3Pvr+Ngu2VtsKgkCwMhUzRaTi3de/5ny6ZB8Ttqq6GQqthD/hZ50NwhH/+yZge3sRiHsjgwFslas
HLtVBn6xS4qG0/faBL4EPshHyK4v8gPfDWynaXoIIeN0gYudLEnE0JtIDZV3EWkVXbURO+yqQcWG
mKfmUUDk3ui3j+IP7Y/UO6nvm7scL3fFOwMTsYFQxGcER+iTv1YTqZuaSPCYL1V3nctr8UM7UAk3
4GL/2mvFM/cBocsIYHGzafRFgxAnMsBAPl9bBHgYcli/xQ/fu0lHqiTGp/gtZggPddJ4o4BXimfq
e6yEmy6Gkd1pgNXO6Tz/iFE0jGtccTqgiwopr5dG5k0rO3+S1UmG5nANFwbu6CKAddActmrx1Ig6
icZKUHseoDmPTXftPpa7M7W+heVGnrH/nB/KsIzw9jApXrJEt04xkVyG/G2AOiJvlec3thIlpxBA
+6qatkuZbrR2JuXo8zJJTZ1OTmjs1uadB9LmnOSGRaAZXPHeDR1YURDHQWzHQAvqQWkcN6EiyALs
zGtGZutSRUG/4Tcm9X9pG8F8v+3m8S8Xuao8J5vgA6ofZyY22MXj+anYGDQHTAU24jKRIy6QSIZO
z/1YUXB0dy6esmO1Ew4uhMj66oiNbIJBdWsPsnurYtxRv1BywDsdR2ZYMRMOhqFcaecwszaRt0E+
YJJIxCW6IGYTSUDQYmPqmqc60IMfIurEVZIAXlY6S6nv7O7GVAJSeIXoH0kYe4GqpqTlDmv6H+Q0
xlNUMrtgFWWlG4K+ujG/LzxJLhxtjqXuIHLGqrA9kodHhjlVb5a5/PyCZk7htPOTRhV4m9p30Fyc
Rxzkd0Thsud1wHMsv/6VuyQ/0OCGR7MgEPQd00jinwVE50oQuzjKfmj2FjQIjSnDlpPvcW3QgWoN
DI+FgJPsvCndqti7TCASn452X3zfb4gfyyHUVqM2pLnNojC3Ibhrb3zZCgwpxNfwxg+MQEk3TqyI
85MRUe78/uoBJYhJHRk9hsakD3Z2KGhtPZNyFbAXMD+WcfOO9TCjGbf9MWKvMhQaKpL9dcJ59lz5
AhxK0Mki/3iY838rY2XOxwMQlDJWr2Betu/w/zZS8FWVOHc6qVAmwLcajDNg4Y6DzJl0hJ1MQVR9
Zalf26X6moA74uqjeveb4EUySCLiu/flJvz4gVGtVCBq+MVh7pos6xNhx+zCMzUBQXW9rCbmUKYA
pjnJBHQaHd5ScNvNVdUNgo7vD/AINSTuEKWdDhp+/T9jy62+VerArp5HGcbwV7s2ScRClFs2ID/w
TyNW1Umw+3sxEybscMRX0PFZqRm0yCJNhdJul+U1jM0gOJIUeKBYgOGRqujXThFgXFH5+SVxRsi4
CVZIsl1HtoKlbsBp091JxB9/Lbbu1ATm2MnVbrnuraWP3KCA2f3sSnFbT7e0pHlHQHNpRwQeuL8o
Xs9g0PFPnZ8BDEEJMt+giWEUFUogHX3gg/2Tw2uHpE9MeAwKQ0M59ctQXyAAx/V8YqJmW+DEHZYl
r+MFuGVWvEufOG/Ifp0BeMjcY1708243NL6Jz3nku8iizVZz9gCLVDNUDNo/9Wf8c4xIMw7G0TC+
FdYQ/BPP1w4Q1eiJ3zWvnsnXtwCkFkqa36hjjeDXOH3uGlsptJ7eA4nHhqLPG6jvls8Az//yOQcq
dfNkz8VisjsdZH8DjEVVs8ZvfRssx5JsU8YgTE0j9HMdkv4egGO4Bd/PxLlM7XrzGRPhynr7fhA1
z9PVfqDZAwwUZAPXRztVlEY1Zcp94hqwzR8eO1lA7LwMM7vuYlXZK5W7hbY7NU/leZmuZNZmpbki
1kJbHuw4irf+WkgNFLjtDBeD/G8RwFKfFB7eBnzIx+wR75ioR9Y3MlIli6yDG5zfHM6NlMGSEU+O
fYbvrW+ssfKu8KnkuMGunIPnGjb6yKquPlBsdTRan27T0Dl9bOoxfaITKjV5103O1ToapZxCL1Ge
OAbMLYrMpjTjT9G+gPwB8V2e1v283JDIIjonqfE8kkoJX6cKn6pzC5Owzb2QUcGvUdXu2vY/ocT1
2RmBI1o9oqBeGI/BWp/dRgYy9AoZzxS3sErOIKwACyB85AaMsoBD/c7N5UNAsRe5QQEz98B936Dt
FBtWJEKQtf4VgogB2Y3uxXdU8eQyCkauxnCuVGBKPfAdtC9XkGsfcmznID9y7WB7qLC1J4Y17uU2
0ZA1FsHl0oKAcRqg52Il1VcSXBbtmKJJc5OZKm8cDc5NoofkVYo1I6nvBxAGSNAPvrcmy1l5aKzx
IY6LwLXsOmuw1JBMyc10ooS66gMvTeUm1HEuXgLJzvSNa6sYJbx1zRd44Fx1ni0g4pjxOhALh5Ly
5/YjU2BKTiJuZ0vFnngt9bFKlRD0M+qXBP1yYwhwCQEfJ3vGkdBliC+ZbcKv6vRKvx1AOLbTZSMD
k7+6fxUv9ATod54S47Wamy5DMubEUV3j4BNKlOfDvivYQavwWZzwcxgbCiezvVfenwAdaz2CwE1i
XYEBniAxo9vN69yMiIYeVtE4kVPSEKxUE8xOp7huyQd7LQECz2D+ikvM/CvrOnv/Vbgz+6sT1GnN
c+qwNjceehzOIxYEXL6c51b7e2vl8pB1Lb8bhW4C4KUN/CJxooO02/SCR4tQkPR/KPQPw+R2wMtI
YSYkqtrJAfBGCf/GxNn+C+RHEB2vJmrwT78LusOxWHGRQvBpiZyZlZKS82QHjUBFX1z/CIw2kS+7
gkSLzTb+fnLqKfmSRmOofVhTTo7NQ9+qyNO02edrAwuMsvCCuKheX3YRLv4giGczp8Nerm4qVahb
JqwpXHI/QEJ7eoNZ18qq2cmRGxAWQm8Nqt1ixmD5daCGNuKpnwUb1wQzTSD+PV926DiyOPi+Y6Yd
OYgLhVsZgKOf9u3yLzY0mgGZ+74YrD8knerSpoQJ64B76QqHA3+JMZA/sGBYrkZZ5uaokLdnMxQb
mW6/NtcGbWhLFLLYKv1ixuiyO327Iz0+j4+3A97aNBwROeA2hWxrMvcpfdarcDGFuIACjrclUXOc
H0t0a/Fu7B8ftoxVO6rHKwHhSZibB7MHmOM/MKksoN74DvJm3c69rb00NheGkp0toKfZ/5kCmS5L
P7RUsonhqn0TJUiUSNuCKxjJ/1PVVLaGLDjZw3AByzfXlFsnNLkqLF+tF5LG9jj9SNLZcuNShfKA
KVziYwRK5YeHeF1YR/K7yBee9Mq2hrkLnCugai13Au1kS0oIYzBKf7Zq6z50OY25CWMUQg/n9tD1
1I7NQgJRoNhAmYxrrYZm0w0pyk78WT4AgO9qf3yVrZxcFrGGXXHHQEnhUoI/dShDIsC2RCFL9tM4
wnVWW9bNTw5mO7Ty6EIJc54x8AiOnp2DNs4EDjwstfFgwIZ2pt09ei0NZqLWj898Qu3O8ipD00M8
6+hhZLb/lyUF/kVFCR3LfdqjMyA7IrQ8hmH0VlYgu6BPcFKteIXtrFHls6QnxzGjgbiBsGiP1c12
GiljO5oo8S4j4N4fdGcuPvNMrdO7cR0BC82sVf4iOTFZaCMKmkvWAVwalEMhFL1auN2INT1nBQca
OhkfjZ2AZF3n97tzCHLiazHu0tp9vf+hAGWd33ceOurQNIIZzpOoxHWVQ6kBF3+kpW7hrE4cXY0c
GZ9Sdwsho0vd2ATNhb03Esai4FCI/BrI0QF713e6CO8xoT0GKxjNbOtwfXr+iRIstNMIcUYMR6il
cwzE/gEdbtyajUCKyHTnoeJxpmPyRBZFyXKjoi+zJkBTHQ54mH/tHmlOcfMQmkHSDPy1+p+7KNno
R4WdU2eDtaqUoklZHMKjrMEwCp3dDJxOeeGhxluauYXMDQjpPXn1SnnKNiXauwGSNpFeMASslXUt
PWqN+1ox8u9Mq4HgA269m6cvuzSD1HxRYB7OB2+LXzhwtNKxLwvyRBgXMpuNcVyvIWBSYTtzYEgH
8BVXnLXM7XN5kW69pSC+kRWNqCleTSGpb3oBk7tSVXNU9JdIOF6tW+fA+0VQyMDalcYPTPBUZ74R
E9nMDwSNHyle9B5j+lL7RR3p25dHE5T0zMxf5NwG8AZpA3/YWXl4xGK2xGg0RM3hm/S2olcqXLE9
Lat1rEnysFz86Mpu7dXuWFCNv2N+XL5LdNFjp2+I9wl7+Or8o8VEjIrZkCLsEyqUVzJmGVUOm273
bGbkwLLkRgyezshQd5PQ67jmBEx/XXtcm3KIkTYj36QsMlQ8YcjrvcUhSxtH/RB38XP/SaK54amK
XaGFdnNBFC1PkGbyGWODPOxLImfMlfmJj0f9aSx1Pi7q/xwxLNCBqKSMqEc02vU0h4PYcYDNUV3l
G4J3n5jYCJThZXCMeJHiCtT8LSVDiq3H7ensZ6BjCkDpm4oNaHUMl0N7fIL5inY3OVo+gkEGJyMp
9tyEJpZZNzn1T93JWpjRUsKCHpcPYqbxP64lgQcmM1hSvS0ndAu05KtXNge4I5kGQJREoyj/Ru1J
6LuRTvgerN7U/1bRa/eOsRTDhwauswnrKH4uf1Ud3WQPaSrkTw83u44g5+nDhHWVXFtH5Y1NR2g5
JsmZaG39J+11nRJhOkx11AWkgI8y8nHMibWjTatB/qlN4OtIpNbfczutatC8yShLYsqWwSXbyFLK
2h+pEIcys4++moHtJ6V35pS4bJbN+WsuGv03LXegTZfxZgIRiWZmkKkAD8AA8kjY9KFMX1VIUU0q
C45Psn6dn3GCv3EK0suLrK0RresxVznlji6nCcnDVjMQFHXTUHjxRDFLStdby7HwWguEvAdUFQMR
6K81quWHKu0Eqc+CxG/OH/Fr+JI8SvaOx+ZyO+yqi+6qR9z3feMBR0vgr5LCIOAe6h6xocU4AdNY
qeO1hUhu7cYJx1ihFIXpGNKFbF4sP5DimJUnbWYalNcNhFgMUts+j3fmhtHN/Tn/McNJdhUpewBa
g+XE/doCLUu8gJqC4yNGwKKpwBoaKY7DaoOpn8H66zGlJGD7uTJmtvvy3f7XSKS5kdntUdozTB0V
GtMn2XSVqZB+xTVriD5YEjB+3XKpNUIZYFZAsiP/b4zg5bum4TnuEBaUEMpiyoGEnmpYBbk42jwd
VjEdFTQPOUyvWKuXP7zzd0NqaRU+iOeuvPCuyOOpH6yGXdnXkt1p6/lKpbjAultAM141vlcZoQmz
EqqFq/qXW5xhCNLhYbsvgTfAJS76t9sosIC7b7jwc3EbDShg6H+JKMySl+h/JJO0UGaGF5zNjuaA
pIhSiUMySQ59g1sFUYO5YnTBsKjaaoOqS341Ucr4z6x4sPUfWQvx4CBWOditsbCM4cs43I4Erq7O
pMXFvFAwcyY85VcQzFh+4CTmF1eOmttXpsDz1VlVq25UTwjkWO0t/K+lE7RG9+9bSdJSUevF8X/q
r7cgceQCe/JCEg1wlixLyDCFnF5IfwjYKZ5hekh22GHnB+5j/2qzaNQ+5fzFEewj9bZ2rfjbKNG8
5dRa5a0coK2myBIL7M3EydymSXR8h3apItIvHzojH5kWEgD8YM+P3R9Kq0b76+CBIMpFXkzzONHr
zULqp/NmGM50tEap2qdDB3gI6hrWAXcU+ser7PuysD9zyQ2BZEhLUlh9nmf7zRlaoh0hOaQsRl81
3ns+Y85+UDnUFrMlVtnNB6nKTleVSWZse4hogiftiYWm44iSpuo0pzSg/ZHEsdwzGzwNgwyFH3IQ
Go60fns2eQqlhCkpSA1sjtnVN38RHSNwS2tkcLUXOTQAhjstPhxZDYGxFgeN0mnJlMOetjr9QoGl
OaskFwnMVnrBsoXUnSys/llRtLlVKYucTa3wXKpv4cIuQVpnHkWwd0zKrGiigfeN4+i8gN4d9SgS
T/id3i0S55SFGYorZ0xPGs0sMgwV6XeGazbY4C3lkG/zK2CIsKmGv0E6rkFFbdVpyps4P4Ek8SVU
pdKBKRF2+sVq1lEs4TxbJ2YSZitVJbe4OFFhcauNw220luZY86Syj0JADN0UcOahVSVqfVWbg9xv
Je0jyzq2JyL5HpBgX29Oemb4XP3XdnMPpNpeGuqIngAcaHfnE79ErlAXAdEGHCVPu8x0//sTbsIx
DDJDuOkbKrAKz3yNYRi7cDL4yUNrrp8+fuU4aw4m5D277TM3O3ReAcnkRWtga7GtHq4dkJzkGnax
HD9r0POv1VHRGteUmt3kE/nznfxVlxWlOU/tw5vbwZfyx//Qu5M0kRVt6q0A4OYMzSUNAdB8jPEB
TAnFb8TfL8EmyN86ex7s3ENeP1EotHJPdQNH9PzEq+0o5KvlqhbZlXjFH+BypJjgSjRR8Q/+eICm
cKX6bkJGcJDweM4KRSMC3OhEo8dGVlrNWpvQaAwpaFYkmyNxFnwaq3kfYiLU3d0Jxe7nDdoYSh4u
MxykPpG+dZL47KKH6WOh+i27X+csIoMRWLgR4ZqcivbtG+/CqMvXypxZ2LXbAl7lyVTaA2i0WtBT
br0gAaSpKQw3uxxy76oQo/WqWJ0ulMCSV/S9HQIMEkedG4qP1x0GOSOSckutNB9OqHrzMO2ig5+e
BPoQ3a8UI50IVcsWdxQg1/NM9iisscuu4wA2rcN9hdg055Cy6ocpOCIVqzD8NPF/w1tIBDCUJq4Z
fWoAqwkEsXj9lfD8uLa8hKsJ7t0LD1NmMVHPxmgdTdQBfiBfdcbOFJxTySO8qPXTWCLiNw7JukKn
u9jADOJJXXP+ECVQZMPjdFrSX+kMxjeSzNHqkiss5QTFTIzsxJl92VSC3TL14fjGgLol87ar4Eqg
xiNBnc3z8YDbs/RDYnWEirDUWOxS9QNIoMUz31VNpQK4qDLxTvQCS9+ZitOE9jYMwHp61Ojvuczf
bakbAjKbRrOtaqRLlAd7x/qSV7sksk26SG8pQSTPEhbJiSYZjd6a4b6jx8foaDG7yvf/HBCBwHOP
ye8m1B93mjSeAhEGk4/2HxdlHH0Fv2i2b0mJFCWxgUDG+L2QNzaIWjCCKMBPUNSdPcFmNFiqVDcJ
NDRG8DQ8En3fymtraCLksGtZDX7u5om+pSRNc5/cK7QB+wyev3E5qeEN7KV/wbSHuwZ1gs2HuFzn
LBCxqrwRCukK4sFxYyyUUr+UdSoVp8dvRl+egwnBs8efRfayQfk0lzUrM4UM7G546r2HsQuGTzn7
pvhmSckb4funEArjg02iO8gblA9RXgCxmM9JQb5/KGUuWVo2H4yGV7WQ54UxunXjMmqA6bMOhxBb
aC+oAY1Li94HrCISWxEEJqAwaTzHCLzFsLH6AGrbwuoR8iKzeHPjlnEZVWNx6BF5BrdNmXjPkdSZ
u/Taugmvr2p3tQky7KKloBjrscfrXv0JWRv8VWDrWQbQvfWzh1vPtLOEk/0ULu1ieyEVpIUi48NM
FqrfnkPFlHKtDymIx9xpN9gAmV2fWfriw7UVrs5Wq0NUTtKGXktLo0dgjHZP7KT8fzOI2gINnrGd
7q2nenf9wfKza9Q4dEV7Y9STU+i4c8kPJyuVIgFLVOmzkvz7q+CLMZ/iiWm/DRvJOnWoCteJsS/s
naSZmxveQJai8IWS0FEFJdQIsA0jcrbZJFRPYP7isZPnpYCDgPhtkQyiXv54dRtJnkPG80NJEvlV
6L5mFzYVuplN5Q4+Day9S2lJ2QVtoS/d6Lsn1Jjzn4VmjBKXkXFR8t5EKy8exrgEDFUJETrUw/KT
Encsa9TPAJXb1IESmx9VlqKg6/8jwO09cTPRtc+J31UrAUrHdcNncNpjjydK5vMLbkgGsjiZaY0t
GEvzyYksTphwnSLAdg8/GlbDYAK4EmbxYrihgrvNYS5yMKkhu/zjBC31wvuHG/ua2+HLyya64MrE
hoKS6uwDIIIe2uV0C+vXcNsunkzdbSLbMlYAE++PvG1hrSyx2M7PliLOspON8TyzOqz13lz7yMAu
xU66Vbt9BzST+QQ1s85A6tpB0PVjITr3ZQPiiJuQkUJ2U1dBYyj9GUOsbCan6IRaAnjHyM/3oKwH
L7vu5xs8viwC7W3rpKtcD62T6Hv7fXfRqc5QtrQrbmy1Lh+B2p14Ovtnr+c3Al+0RfM2VOCw60kD
KJEUQEDrSPNWpuO8R4YO+fql5q32hZznIsVL5l6W6GkHmp0NnpdAfyO2o8llD+576RbRYicOykxO
gTa2Nq3wF6z21huDnAqywAbhBp50gtPxgOg08/y14CSob3leEjP7cPVhRrXeScSTbNq+s7iv468l
lKJQNgZBCAcmC1Jasqc4GT0dilPWgmG3d6pejpsjJrA/edBOj/yQA2vRpSWDkXfFRmSppvbRbRiw
xR0r9xExFC5Kr8Ivw2Y9eAMsbw2m/ollLQel05oSAJmZHhiQk+n+3/ggiB/C6wgyAMdmS76M8a4W
9gasjcsu7NRan7hduItcv4Vwhpg08W/pfCoYWl0eJJS/lNEef5HvybmkNfQKcKmKlHByuoQInDSi
rFl/Oq1bvPyNlllBboPmYufDl2rDXQ87mEWT9ViDRB+eLofZPhOwxGR4zKTHYuCoCEg286xTs+Xv
ZQ1O1lsMdwgqS7nmZRNaTfx+Tuj9pjs3Bd8UJQg1ozjJWJC9bTw4aHodd8+JwBE9KNMjp2Z3dEfx
8ls38baA8JUlKV5BVHnPamI3fA/EmVAG1Qo/JBS2eZg5sgdQk6MW2uWzNZAcIfXhdqiqeBKGR/hZ
pd1u4yw6slBIR6AQoQOG6AOpYWiqt8vrOyF2JiRc3l+MBrSFHNVG6Y7XArk8zT8faLe24davZ9kl
BplLk6A21MsByH5+PyTJOuSVZafKOEOqtwhsWQb962HOUKTRQTDd13QP7fBGTmEBEvW7WWBl/2bx
onB7bHc62rINNM92G1NlaGqstX2FuKs0f0ycwPN+VgB3LF+/WDoTeR0PUAHu7IPaT4X+QwvsQN8N
Qo65kS9dPxlWwYg5OYgcHmOP6u9yV1F/m60bSKqm2rOezDAR/JfFwOKLjH+Vpv4SXtxIEBN87MbY
5gOFf9sJe/27D0tnb1fNgy7FuYR3uj8i3wNCOj1HesT8tS9E4Nlf5Scl2PAzXX/NQrS8XQahrj1M
YCPao/VjZhydKNpb710SAV0jR+AxZl19dqsF0iBLbX0IHOPFfZyUSCRQ4kYKWklqbq//MjJADOmp
zsGaIBsoIrWoLgsCUewtroypxLHd8lGMdOB6Hg11U3mHBXnDx7NI17z6SfpV1jkm4XQJmylUiPJj
EIv7JwOJNqkZuDP9+z1bQS6HNUMrAFiS/7UyIbfhJiR08h+w0TC500YPJ8ve4F0EYLeBaU8Gv1Wg
KTiK/pS3PFafPJX4Uw2QgwCGMRgrEynR9HrDDJuAxSxGnSFXdRA64Wb5vQh4rIKRsSyn61/FU9XS
tILDXijVCweqDQRgOEzU8oII3AArregh94nvPF813KiWkywvyhCmhtVxBAk2206h10vV2cdVgJg9
qrRXqnJKsOdmxt/jTHjpP6FybG7816E/UKP0cVbVT/3KvtApBpuglpzEeBMIfAaYVcz9KUKVdZ8r
xb4KE3ulF/0EDSSpLgpKeSdsjVvTWaWsZu+Lg96arvemhBGa8pqBOjS9uSyQx7kA5quOhdxQHBDU
bE+SmYMK4ZnIXH10EXAaaaEn16W+oTxRbcVl6M5wssqH1HuswCha9f1qHgeOjeIwKq/C2UpID2W+
yVh/fMLeTyrCKgkh8OVxE4ADBdmUZjjrtvo3uL2qcwGTvL/eDG3NsJ5Pvl7AJdrU04vWeFm8FpaU
wHmSONgDT6VuYMPh4k8StNgUqe4+i4fp4qZ3XDjVpiwOYzrUDxFwcb+9XCCjmRuqxYZokRnmZdiy
CNU/Uc59PYgG0Dzn+LQBTSSNeFHuSRGGwdtL8pMhzZ7faFSK72e361VZ4TA1NomZi0lmL2M7Vzpa
6Be898PCf9GgUMzYUPEfd6S9LszAdgsdAoB3bMKmzJqBLTsgS1HQJGSohAddMReGUiLmOCOaWbJr
LYQrxryyYLZl0JO7dzvNZ+RXJr7uNDk/N7I8jQ8pVxrlNsDmxbXJcud5WYJOECGWIirlYzt/0WiG
BxYXoIO2BbXXTfXeOsLbgOiyfopjFwGe/QQQ6Q8L76vUHhmxAOEcaGvv5tUFSHYRciRibTA+GG6M
o63wdHRY08pVzEqoxyNSMDNenxGyy+WmrsTKcjNupsZNjHjaXMhUTZM8lLaawifrQ2F0vd6BSSk3
+sZTfywywOQ9/2tana2zW86yweRQ1CF0FfGQsYnKu2gjlh1Wq1z2U5ule8U3HVPunJJrGVVKv9GV
bpP3SSIDyZAvl5mM5XlvloPC/YpHn8ccYToUdi6js4mJERhpIzfU2KwIhaaKeml+CYWTy8xdh1pW
myeaMqb6gvPkMHRgV/DCHNPrPtwLG1LFhWIgYl1Dz0OsiVgl+EhPB7MPsbgaflmEgBS5jToz3ZPy
BrmNQ5fRRvOo5jpY/W4DPvxEAnRowugPUbWOL5Z1NtOcfFnFWCtmyGgrzfOSCqPtqB5vg25m+gbp
kaFDH4+xjCczp4931/LnKBkHqqbKJqIyUcZCceDrUv2FL36JCOffPWWqa6SzSDp1P5+yWKP0PWgL
RMgNThH8w3uC3+azkGVe69G1662CGuazTtymPBuT3MJPNku0rIXRRzHHKz/n73ZFQQgKyH/1Iz2x
JkS2Who2ROMBxcx2xhYewa149tPjt8Kieh2uzwF9/SBnZCcIlfpyMxRQd8mmtgrteWd9iDmW30l5
gujIB7mP4a1ALEMzxEtUcGNJc64qfzf/sxokykDeDe+I3VgwzNhb+V6iy/e5pHvznUdxyq89HxSI
Kc0pcldbQYQTt5OkZc41jqqF9fB3VTLcWhHKcHT1TTaW7PWO8z/bCBqsO3x8gDD0sT9WMVS9S3tu
DZpb/OGQW3PyKYjdXqX4Q4mnCNCQ1f2g6BgMxl/TjU8nrzx9Ridh3S1zUJM0NNwuy9SYSbPJmLXK
u3qc6kjL1QW2KBXERkPbE1HjvArb1MfMgW429CR1Bcumz/9onSdVvL5KoNTQ1Ocqs8W/Go0Wkq35
QHnb1+QQkJZibNHB3Z0GyvbIH1MLfgQBsvCdlhm0b1Q2X/9zhoVyuAHryWZmvmZrsRkmXDzrdSFP
nKJhERuRYvfbmBNR0mxKCK3rfRqERKwr5GKYTlPFrMjfZOtSoNE9u51YWlxhRStH9Jj09g3yd0pp
hAH22pH/Ym4MK5bWBzz9qFsRw+e9UbIV4J7VgYUgJzrhpuyRkcWl5S1b20qrF4CQBmaMWWURiaJr
3wLs1M9VDyd4mfMqogHVWA1ljW/F6SHwdRw7kqw+QGsZuvSUehehf7PtJ7+RxdIIbsOnWNtrTUdU
tGPrZB29n0ckauY14JvuDzc8+CxA4OzZiZ5Zr2Qaak5uMKdYKmSZ4PWXSUUI625Ajz8sd92EjLK1
GuuMYJBfq0oeUGa8OdW9qh+Q4PxLL1FJUCqPlPBctE99Iw/zhJiqpNfsTmNRtmT/wKRwzBhlKknI
gDIVrPewpofkKnmoK78BFz0/qfshcn86yWozswTDJHLhs+bnqiKHIgmXiFmnKP8ij1hPZmoDfqCh
WUszPVmvhY01hX8tb6oUHtAANlsPRnIVJqjQl5vH7nDibLBcrhYcnAbrIemob7OIgGmLpLOdodyV
vUl2uOvftOtH3to6XfEAja5o4AjB+lzMtt1+c7tLfw3PBiyZdeyiULWoKkNcV5UZ01ODzicgTG83
9ZNK+QKRLBa6rfABBNYh1EPtNeqaxiKgtcmMKJSwtaTHsg1bejEQJ4M664/2jmi/yw3lCQtZm+oR
VzwIuJpMVI6lgj0mKW7ZX2AkiglRvj/wO12gcH2btEPIgvGQm1BsRlGZfbjtfXc2yCGc71ZD9Wqm
kCU84wq0v09VifNE98VzJeGkcLq4OkbbgYLVqNVsfvZzPYCEfmmGTGqbv0auJkpqFUa/RxNQYnAV
aB0E6A28Khzb5FXYs8Z27AfMAE15yUUKQeNOtg8nr6jbf0Ye53gz6bjuXsTwV2odv8w/FfRvqkkS
BBf4OUYXdKstAYK6f+I64j+oyS+7q+6LF4m59AcybPUUi1eO4VuJGDWM0fXtQiZGS93W8mLZy2rB
ET8AXX9o7TYSxsTkuOJrZyaakeFC1RPEERTut/R6v3I+OJBsHwOflBn62YdAvg6fbrm2m1H4TXpn
zS3lcE7PPB6O6KQI0YADdZXU2rGm7L+1FrgmR/0sr9Ou8vdaBwfTTLdhiqMC7qadm4VWnBChs+z7
rrcnuTBDiyMrvHHfQ/0R6/oHyLFLrnQoNxK4X8veR6ZH0j+Khv13KZHFL8a46Oz9gvEIzAadLOvq
trcSDM3/NwbT/Hn6GjTok+2+EN8bBcCZV44dAMs6W67cVkgdpnFFEpTdgQp5UxQLrC3lfNKDpJyO
4L98kSDvzyPCthzUe4E/el1qXyNFJArW/f7IpNRjmkXZQp9+v39gXqqArtjXbPaZtmZ8KQ/qS576
I2Q1BOttFroGfXREcn8tNs34TmiCgdB7B48W48cerudoolt2UTAA3cWTT4xE3Cior01mHgfhBvC1
9STCIP58pXEo4e0QL6LaWT7TPux4ixGwaKNo+Lb/yQCdXJ/VPr76mBfY2BV7p/bCwWd6ndoYmmju
CSfwq13ViZoCsuNFdilioQg1tLGtUMmOlgLigvDJIoWmI7kV+s1+olqOe/7RAMlNdIW/3yriqs3x
PL1FwgR78QL7x/TQ/aNRgKohZSU+gO1h//VlPHaeKTG8YEBWpB7PzpyylM9e33viky0ZQTskSXsN
QNX0F1NvTGhCGIxYDv415jq92FRbQ9l1OPt0EYbE/KYULRI26yIk5xn28+fJ/fGJQK0tQ6MLoeiT
Orl9KJQ99DqgXcQfsf2It+aWdNW/+xu/f8j2DnmnCxSQh0XvKYAv9xjZVjtlDuiqevBP8Hl7tyzI
CBThuvNpeTjAE8O/BE7IMRUfbyb/zypYAMSWlU9fe2V5YVpYB4bgm8Vz9zKXbqmSpEiYLzEMkpga
NinCM944pik7BhNnRRWHnSG318gHXZTUkhAawU5Uv4QwHx5RI1XVTw3d90hWRi/lVLUo93D2AWrE
Eh05lUf1w0ADvEhSeXj8qpYE7Gs1SlSKeGnhZrQ5m6faE/Y9MHGLjnEoH9euPZfbh2SVV/ZODuVO
8mlYWh47fq3dA3ilpAACW6B9XFxi/oa4alFozNWrFBKWRd3UZ/sJ1I0V2cKMb0lPk9nkpmHlu7iS
KJBQjsXEn6/z9sawtF8CFtm086OOgLI4iYu/6jzZz53EWxKkApAPbpejYSTJinyHvs8GJ+TrwZT8
SOrLzLjnUvrj2ydXeQc172y72Mw2Z7auKDRi4/FqAm2CoR2vHi+Eeym6ZjZkzPFgOfL6/kU61zpP
ZmhAhXyMENl1dqo7ZMnGeuzP/Uu2jHEAIuJrxY4Dn9kiii4meQdmIPo6OB2o6Lw6snBSFMwo7HRc
a10fFoEhj2tGJ+MbPFcDD16FLsKW1EGOT3XDYQg7ePY5eOB4hTHugfkzEzDL9jT2ajctbGT+pUgu
/gOoZgedmBaU4Zb0i+42OZrNLTfXFVc5kURqrjb7211p55QKnwQ8MlUMAr/f6dhr5t1WxTXf7wHf
rf6fTt2ZYGJzF5xgXcQ8sTNFFvNlKdOMf/01QI045Sv7w5t6s9MYv1Of9UT7z29czFXd8F2daWUb
WI5umWVPDiUPyL5iCSe4JXHE9s3mfpxQCqqhMtqOmkMiY0uVo5yIBhvYxo0YGmvBORhXAk6qNU8W
djg1ZDV209dMXbrEZgeGich+0xddm+qurpDiCewXq8B5Atm10SD1FxY3sGWAraacv3u3nZ/dpAFv
7XSzJNuLNZtD6xbgBj0mIMN5HQ/o9sVmibD43VvrZLov6K03NF36kzJYgUcamlEhRlxlXuKTNiSL
BP57czRURNUo6afX6NBs4K91bgiPdwnN2S3pBhL/+GUo2bW5NpdwBjPP1M1Jyvt4N5satmOXBWzQ
8XCvrnK8y3Kk74IA5lPYwHKZIDzA168zT2FIFfrsa6anA0J5+BjjpGcqh0m7ZXqFXCfyfjEP/Yco
kkUSXQJZMyzqWEC1x0iv3FnMBJ0uwwT900FyIHiz+TpEcv7Nzb51xB/mpCgH+AP8EjZvAM0k90hC
9FeJhwP4d4ErSAUz2L8nloeTqu9i8vAdA32JEFeg3rGXCxAjraF8AleVgy9S/m1CM864k6hkiBCy
V6s0+LH1ME4mbX4NG96vja7um20zYWZlhqVvqHZdt8vzMcKpq6i9jwYjmMDtDbJgvdc0CiAz1woM
e1FW83q5YDH/6IjY3JNrsoZN6o9s07CwftlEaBbQ//dUXA2fc1ha6cb/oSUsslPjNkVVkO1CQqq3
rSpllb4cZ3KSj1zrWCOIm9U1eTQ8IRPxVTlySIwT4X3TZk0AKaYdoSj2CDamv6NbLNCUqVKxWn4u
Nzhg+2FNdT5GNN2PWP6QBVtqlf8vsrjmLeM01qUkSc87JdCDNs2ry0Z+l1DZchmLDLFSSSfnSaHc
NZ6sHTtdgTQz8eKlYd/GPVxjwAs3VhjmZBYu/XUyMNpGlDbAgF90sJLxD1aSJNTjBoPfMCwshLiK
qD9cEvwDjfsFKJz2BwiqNgzZTiJyoIeAqgXjSnGqDnol4otN4ViMhxMdTTwvh4ty0nlrAIJsAx3h
C8UsrZ9IaJ3rSBmUJch7C4v7vEe5SxWMIGTbINeN5tlyVbKnLb9STL14r9JAKGGKRkJIiDT+1bE1
iVIYa173ybsnBPYI3ZH/7A5D3fm/tgkplsLweQsGz+FBUHdLmFQ/AbWUqacZLfYjumSfL0F5P8om
Ks6odjTNr796cnJPBVa+enk/83une4I+iENOo42tTsuKFp7VHzUo+oWzAUWBl0kH5Q7rYI4IN+Gv
OkLbSLHorQeVMZSddT3bJB4t/EQOTfVgsTFpeKtrtfCiydc1ZAaemL8KzmK14YUa0D+1QVvE7pQ9
7EYod9l5y82GxdVjhbZZftaobRYGwRssJlSI+AGeGO3VLEkQmHQBvPM+OLJOUmO3MY/0P5Zi6p0h
kVTpkIcXaqg3shCrCuebuLnsfyJYKGXAekWwaKCCY36s27lIOE0rKt3p1ByMEJ95KEsfmKvnZmV1
ZdFgjiQe10Ojxi6RL5WApJiYMXl6EV+DOlBe9LWyX2ms67xfU+cy41vL2r7ZP6YBAclEGdlRJmhV
VO3eK4h/qS3TBgB+EHt3+7n/C9BaMfHUUDtjQmekyiHDphdyIhff2b7CywsYpTu2TJpdHG7r8tNq
4hQ1ZoJ1mCBoPjVA5T5a2D36N4cniYkpVZHoWZ+HpvsGwARKgo82Zmp5pZv/wJGoKa8HC4No2gF3
oEjlh6uTxcvqtgNPMHVxkezkiVFFWtZYenwVp9w0uVEnPfCuSQJTNgEWU2CZUNAU6uB+lEupnWYb
Ntboo4K69WZoYxOyNCzqxHWzA00nq0ZeuwACYEA0jrIo6+S7rrLbgaCPdkI+ke9M86Lch/nL5Y4q
01IhuevP9D9PnP4Tgs5XcnWJcp6pE8oYiT5QiLrILQM7KZQ3t1FxtNNRt2cMjfgRQvfi8PI8pbWX
C3nlGwGmyjSJ/8xAmBu8a6tnfo9SvomqQLQRA2Sir6GPi2ilfM6DyG1tAiSBmP+kjXrojIbyW/Gh
wuLW3sg3w60NvtvyelAC3+l/wepO+9Z5XEsOY91CBM5UO6KnNc5GZAS32l/FK+DlrOAccQqxZ4kJ
wfiWPOncpssUnMrNI0DXPY0lWtdf1h37PFrKwdn4lK2OHy0TwMdPVPIjFfPg85OWqhCnmMOu/BMd
u1XXv3gNQDnxv31PKatO4ZBUqdIo+UFVbxBKgP2fy3hOu73vn5xnuL/ctD6BPRqQ1eRUnqxunFLE
KBaghpz2mLjY2uXpTglf2WnXoCmYtZpxbhhhZjpEhiGKbLG+OMY02jTyy+LhomqdLWkej4AQvkPr
iOBpqD6MEraHQOim+bIsAHIEj53kFwpvpIRZOa0Vnng03fxvRZSgG4csxS7NE7QrSET/pQHo/waY
EdZVE/DgoWS21HDH9CA/7tU74r5fCjD7+JcJzYGjKL6YWYLXQ30v4xiaAMZm2vuFjUEAyDkONR3Y
FL3Iet3hbwns1Znur6bD/h5uKbsVAd8a9sWGHJZIVM/mJzgknBH6k6zU4kLFisJV1Kdzhu/5B6Wp
Xfez74x+Ec8TNxUntWCgdCAhI6F0CE7Oav+bUULypetLMfvPDehkddB0FUz+a+/DldxjLHA34E0e
oIYwiMnupv58K3MOEGuU1RwHCgxZisMw+YFNaOIN1xgSc3z+IlUpj9hJsOAIz1KyJyzUSkDhdJAp
KKFfiCUoO6n+u07a+ZoBZdl+jhkiub7Wsji52ISQvOy01QFr+ICY0So87KZ4tKkLbYlkwApY+1wT
x3jRHUvPpmbmyY56GpvxdNyWdmA1aiDvjN6xYZ6DHNBxenAN/3660UQZIDlk7jpzB2KvG1GXY+Lr
4YxGXRAUcInbxG1O6JlV00X6QMLTFBX+fzytGmJBQpsJ/O4efrySpGYUn3dhB18q2KO1EAdhUcpQ
WEeIhL93J1syS52qHQXUyn6dI8rJ7HXnAik+Ifx3cFoqy631VFAkXMwx/qMHg8moDvmkJMt7dYI5
8/Fuwz1Y9wjTYHlgDwzeyU+fQ4kJ+Zc2v/eX6MSHcxN6p6LNLygMHAqp0yHv2Iej0dH8szHNKJu/
4e10iCCYX5ENBSfi0h6+JpIqPJ9gVYsuMy8+3yVH3IRe3KGljDffgyGQRU1tTEZmQj6tcOGDWJ0p
5R7tul3eQhyeu5JMDE5TlnaALGhTAN3EAh4TpLwxzsVgBYrFjI69iObr6yNZHJ6xb5QcCcZod3u7
xUMoRcKKM9SHZ/0iATkVpf5+cjsuInDeXOX9E8gef7NKfuuVEHU9GWZH08bevZdZfnVBvzPeL7Qf
jZ83yN/xeKWCvQZC6Ao/XgZ4+R0EoD0+ztprGdwG/9PuPm59gHbyPX66dDB+DH22qd43fSsMec7w
+C4eMs89KtASJQH8IlmIWJZpS2zsCthvYtoh9Q8XoH3YTNKXmbH8uH+TQAYvPUxpjveuftHgqdIs
/a4nL/hClZgpYFtV/P46PVjJsJfGTf6N4ut4qizcMEi5rDGNHcarRQ8KT1fdButtXqr1HWSWl81H
3pQ48cYfzDJifh2us6nKTTVhGUCu0f8SqYGEwzZizgCXDxyMTX3I0nP76X00I9u99pqyVQZQnB5l
4SRkj7IHo/iGhd8ClFLW0rRLkcJmc25EqKLtvQhAflzFnH8ynG72kmfOqnru3bFNVlR8e+xVZRRD
NnJTTv8m9Gx34Pb3/1SvahlzWGkDoayBslnLi3Qa47VCvKgSlD3bpk9WMCNRzkABDNRAza5UJKNd
ZZU58uofAufEVWXLAtZV01807kKBeZa/B5fpXKAA/ey/hWW0pWv5RGh78Hy7Eb0ReUO7WKF0xJ5S
HQVEL/9JNPO6EynziJEAbKS6EOoY/847j84/x3E+QVlC1bxc4vxrX1plml5k+zdUEIqhX6ZczPc1
ZbVKFmKl4pY9Pn7//K2RvVosdfcX/Trkv2m97Q6eBMsVp+ycXwgsD49f2tYIqdYrukVxzy2SpHFS
fezWZXyk9slWr0VEm6HhFutdMuIleNffZvKEN61EvxscjhYAlhkCknyakLrBqIAWSbTcOBmvBmFi
nHqS3NZvr2U+JK7hbFPh1ngqXoe9V/gfNfOW8T2AGPCzHMZkcQ/Uw01ftQ6tXvciKzRpLQT1K9Vr
27vZBjEzcsHQLaGtL4OiRyBsHXTQZkaWixVDNqYM36ydg1MGnqMLKia+BrthCf7PXL/nDaZdRf9v
vOOdkJlSEMRP31lX656SRPixWR4jjdfqfPX4ifrSzJYe14f2ykZIv0Ne/aTpra/DVfdjoxq+vg+5
z6Mei+ahmkmo6veOJpoEh1VzAzd6xCu+ch7h9wRR1InHWt1v8skStYfkRZ2YlMUrz2SMYPVXwiGm
NEeLszlCUGZ5i6fK/HWTAx8WEY2V39beF9GRe54oqXoktfhb/BihZ4O8MvKfO582aNOKV53FtN2q
lG9sTmax5AwEr8JnnG2cRj+1BBHPIB/4pVzucuncTr72ZTutkgtoqCVUsFtFzNDGhs1jkhVGG+3m
G4pubU9c576z0aNZs9+BhzI1IX6iL3/jt4FIhNhoWrTt1mlaat4O0B4hJ8P5jO8CDnbSGINY1aXI
CYN42a7tNuTskpetL1ndZ4dwsufcXZoUK/3YuthvQKkD6OUEbuvrVEZx/kMN2jMCOJQZG3x8njkr
QCBtdNeBdkolbUcIHPYBlEKgAD+K4bLw3YMQRur26mWGw3dGFMWQjZtFnqqWQgaEzmgcWFaRJx4u
9tCniaLvAVoFDtliTmB4EYPa5nkbaOlqBfU4xbmv8ht7OvrGbb9ZMRbB7WJ0ru43FXKi/pfRLhF5
0yEKUn7b3uPa7PfgQ2I/gk7JA12fAFaRqnmLSovw/RNWIkch9PGZ3mjcCAB3XeK7tYzr2X81hoOS
54Od+VEAJrfoc1UcsGzHtF/NLBE8cINqK3Wdccfb2b9oG7sHqUCeQ/F3qFE5NB0M2Vh9HkYOwkPA
kmcSxIzQdZjIkRl8ykgh5bw6772TnhbGyMvTcSCGcHBS0Ag1r4OrHagowN8w7AwBc+bO0YyxxG6R
3hmhy6NWGJGsGvmFuOGj7xp0eRjawLvhRjVPYtU8zAW2dRwnDLikXF4pFev5NFmpYmsEl6jkuSrL
4MCW48PQthk3gb5qziyZ4nG1cYoTpkl8TWkzmGLYWnhmqudE3sSWumv/fnfg6rv0rCrp9JcJO+xK
ixgywlQ0xgCF72uxlJjNKW89kv0CNW1GrF3ySVYuJVDUFcaSFbO8PEaU/bExK/gbiRZ1iaGqb3nu
HCoD78SbGk0CB5XfFsNJErF60HeSM66AQM9wOXlzlPLrLNO12YQ4YfhEkWN1ISZ8feJBhUmbynET
uVejeRoO/DUFcPD4//qq+gFlCi2wQWi8WWj0EWZvW1JW+fnSvTSPPoe0RMd+JCejHqRsBUXWz5en
tCy1gHHc/KEpWU4r71xGy7fY/An0PX+WgTHDQzvJdvyRO7QhZ5Vx6nRhAKhNnLkSWsJwQbn8hxG0
emllcReCGGCe8xGgAA0y+A5MBCfCJT4IVOKJHZyh1bFKdiml/gA6nV9c7IHM5Cp0M1oO0+rxZ+yY
seyvvyhxRHcsNhcxD1o/Qtn2daaX4yOzxT05CW5Ekq8TxuksCNDFkEAvumpMHbp1SE4mY5YlSifs
8Jbe4DsQckuykrrCF82wAFiwHb6RJ7+pQiEKg+ULeJQ4HOEdGhz4f/7ghjZ6nUizk+w+a+pYX0zO
vtsSkHeKLFhK/61O23v3tL40nXlDaA2IKXiShY0RzJoQdRqcZnQyZec5rLVvL8xBi5nJ7nou7VfY
w3AC6vgmwZcuXBmIGYZKzamos+N0c8FVpV4lwuQtylQSoEINWdY6TDGgFAYSgxC3fRfk2bH+ma1W
at6mUmqrlBsMEPdOjzQZLDpiDy2C0qOYn0GefyS0liUIxqR8CG5hji06GbOEYnDXLcEPo2nfdbLn
Hn75H4wBxxYLmqzvM5MvcIdFrsQdqnlzoNK6Qpt39UqXskZBikGlPBV3MPGbcIsNyFH3CvvrNXgB
EAik2xsCdmB0DIuaQ2vnMHyOXSPFsk3NNm3ZdRECnSPKuMMR+hkKEulFxmTUCWeeGxtT/3g9GSnK
/55tinoyb/x5UTEKSNUSu219TJGV/2Cfu0UZlpwdF/sxZ4wZiRbkYQhXqENivihN7FE1ZO96F787
x5lC55y0uJkhe78Q2VrQiWny1HJDps2mO/eId13qOOsWqLx9agiL0Y33MNe9yAG64C6ZJPm40Ii6
EyUC8azWX3h0pFmS9ilmdN2NDuKfWrY4GszjT7rgFHrznt0zeBrNUSDK0VGc0H/OqUHWXfUOZHBE
n22T4PsG6mM8VlhpOUJsHtJZeS8oYtyLjZPPVmuZIG2Mn48e/5GMkjrdnC26By8R09lzepZjmMXl
dtaeIAEqy9E+XHec/MGCd2fYYg/Cns5j4msBLmtyhuP1yBOEDPBtIwh2chnEtD84wJ060aQDD00Y
k3Bm4PHHucnrQNNDucPmFFo3RHxJwzIxOViHWWtseKTHePzIZ9vk9SratDkMb7ASWvZ7Ag9j+CoR
ighpZq4fFZiVTPe4d+oiHCQ+T6XFhxtO2aMIGbwxVPznlEih1RUhuC9h4RnneOYQJugQDwSkmqPp
u+h92vr00yS7jrnsGlQ8V/bzxfcf/iGXzZyFwGIDAPuGbfgxwv3i0hmwYMSDJqDEW1RpqkSZ3jBz
nXEkoyJMO0iGhTw2Qs3pFrNhkWhjvOPhlB0dsFORlbXTsf2K43rVvKxxWrXsfIJ707zMABtDDCYP
AVFyshaUASeMflTdNGSMcI7YO6lG4XlyShCd8bynT62MEQRvPFQ6xYytzr2kTpUz55YbcNfy0rca
sYrqKx2Gm5k8wQ3P36RZ0rG9WxhuOt/X0hpllEBTtWJ87UlrbNeCN6FjkzIXQvsoAeSjYFXuvjXW
OR3Yx5Q50ailKeCQDqmslsAuV7iwyGvoRzJMsj7Zi41PT2gJRZ3Em9Bqdd/K3UBHOVYZhgXU0lQh
YzC1CRVTJwubB7UuASaIcOlmL6e2FC+QXHs4S2BH0uhZHz7sC2upzS1Q9Jj5FEUuQa9PVIaeIcJ4
hd+9zZDp21G57xMa3VPB/hsGv3VnVDte7E+2aOEOg/yhNtqd3ruj9Zv5Bne35Nj1n2o/uMvAYQfX
Dh6lfcCXgIq73/5jRgpCnYkmWsOFjPP6FvAtBUWlcL4GZxZpOh/jQUJWjzZDx3xoWFpwBf9HSMD+
qs8EdWl4fN4Z9QsqasL3MDa2rBWAGZp+t9RQdORbwVYt+4N9cLjfVIwpKZ9mGk7ullJgguTUfHdZ
6R4Xlt+IGNLDrv581zUGCTl3GHnA9Sfah993YzxL37FDmCieCWDU/8YwnDCRhRpN+CLx/NL3s8Wi
wArYK4mbddiFHrxapl21pPsoeEeTIZjsPP0Rz9WcKA1jctR2WLizjGWIcAoLK4iMnr8UREc9HxPc
UJik+G3vRA/uHsfqlWPKAZSydnbk1KWGJA2nM4tEcSsTkDVAgmwZ8SuQA+frDzH3QhZTSr6UkJeA
4cSq++JljJnwbOsCiOppGuJCWISBT7bLe+XAnA3WJF4DkwgpDDy3eDV0mw6eQdxzgXe81yoWv44B
PcxMFyXShQG6cBJiRrv19RK1hhprNEFlUh6ycQSuUZf9L903lmQftaOE1ZS4I3Pd3rvW2zzwBJlR
4uYNzCYy2n9hgz7t+xpu5p+1jf7w+1OtM1w2+8zwr2kv4mkCt/7/Jc67irhwzPDCNJzSyXrmBHV4
ckvj19xbr7pRv0nyvgwKeEZ/4S+thZWhbKr7Bso8szChXWGZfKGV3EcnFWhtI0NEFXbRF8Y7jTLa
6lAgaK5lv33heK4m5msbVmw7v7bHNHnhqziaH8oX3tRtyd5aOAYwr1nO+Xh7Ru6yoSP2KGiDLVXG
yIfJ6gbiAscYwvaU+wyxJmsrnkiUXt12uce8XFxQYkTexPxVzRYOZ2Muulocph2pukmn1rl9sbjM
x5wkaCbRBoxD5Fnd/B/KJjhbDLk48WPaBTFRHeDHJ8hnh19hXhuXHZwr8lX6smE12vEJx7Wt/fMC
jLjRT2yReH29vWkAWH1hhTzlKNV5LyWFcjAu9bRaRfImsjVM3HzAkMf3U+jXaHKj/WY/BL1pleMK
pTTCvnuQldW6XWno/VIAwUBjzPiPtDoK0CnKnRgfLwJO5HAy0EEs5OkW+vama5cEaGkBvKYPLxSu
1Ud1sfoWGe2Nj7VbgGR9mk7WY+UY6hQACC8BEMPZLyiFAghPuDNRLlgSHIo8YKmc6f3bZJlyIZvk
laioBild94KhqJDs9bB2qiAXz7HwiM4PFtAHbHIBJbMjrIDO9EksfrnOzenbGluP/W3GLqLpykPT
GXVm65M2p9wQB9ha9g4eZ87W8X5A4GOusN+Fmzeu9cAVhP0Y3RZRK+tk0PwKIPTAaYXtSOMModew
u5uyGgRVbSzhwRkmvmCV8UTsOvX9DSyWORIy9aV8wp71xUaeJCeO4KTuAOZDdOQpnF9RyiDljTe0
heiDFN7b4s/x814GqQKljxYpY4DvJqEj1fL6ayGYi2F7ozeMRxPZAfs3niBqNBFTHIjCzWhDSPA5
2UFAGjfvkdk8nHGelJur4uCx7ZYnJMpF6dbNjx/YhaMvV0/F6n4is/KR1a+mqpgmR8uTHstFLVG7
nqAzyqhQVV6JkDjYjRhYcW8haw0r8B9RPVvMwVGMHugNvsF6uy6k8ayaRclVAcXxi6XNBHWUDqad
AbAfX2JBCUKpNN+V0glFE6P3MAoqzrNlEmExtVZtgamrtI1UzfbxG/Hha4/mLdV5Vg6VQCFoGg91
ZfpTo53MCEp4/0/cZ5pRIB9l0wFwLOyh4ejnN7J4GuIKlw2t3vzJgG7A0ypoU1a2JTZO/+G5qOUP
mfKooJoE0+ocluzQ61rWhAMtiZpq19dzH1PBq3XcY6HHLqJvk64iGLhwBQxzvEsCpj+vvt9CnyZp
csQ0ReaCFtKJKG2KSuf/o6qLSLGVcN155EV9MD7fuXhTcoVM9njz8iXTNbm3B7jFSzze3jHttza4
/h0TxM794OovGxg0luWlasVTBDtfImlcxST+ZUNhuhKiCIozU3WCKwBs1Yl++1siQn5IceNw/phN
oU2ZwufH81hsq1VIedwuLM2h+I/AUvQ1Nf+FebkJgLpV3hWAp3zDPAfYmf+lPSZNRuxF8JyTlk/L
HET8LbKdZNY0e7vqMnhRy4yAYUXKZaVaqIht34p/5jCHJKSaERKPvAskXJiNCuV2xCpwgSqFHifM
TdLLXeqBKoOXm89TyX0icDY4AdFHPmRQ7wTVu7FwRzxXhaH7WMH05aEwtwj/mZ6Ck4UQqabDVdcu
QHjgVfKRxLVU3RwPfSRS344dYxg2DsvPAGFqIx+EpFGR5y9uloRO20j1yTiJF2EIjjPros/JK62i
W2hG0fNqNQO5N+K5m5v1E4B7tzV34CSDBoHY9S4ANTzrfsHun3Pd7l8nq40wkJ0PQAeA66QDZ8JP
oNMxtJkBssI/gEIKLmuXRINEbA0zLSEmdpNUpbCFsGCXhfvchh50OTwXIunGDXPz2v+WjVahWBQA
/jQGJTB4lxBWhOYhlHJU+cWL01ljGCEic665QG3kP+irjFEPba31j1FG0FMwgNQkY2CQ85zjyuUD
PcMYOKZaHpX7526OBl4Jig+KLkAVNvPb7C1gi4AiDD4GLNkoVy/HH7+1sbu698LDtBBsGMffhXtp
zVLoeRZ3QgGUMyvzdXxlob3oePm+q1M2HVZPkJWO6O1BvB+3EGNYHftaNCONhGPmiadr8hT+wuqT
xe6DY2kuBk73nnDZut0x1YRO0cqzIBojBq7Aq58VSx5vXPdbfsnzVnq1ibx7BpMibcNaWUGhRbmy
GoXE8TReD8Zklv+OSqis25ubpLbQa6Z3mWpQJsjuHov1HSO5eGw8sbhLWZwly6pUatWk4qzkpqfG
UXYhhLx0C57IDOTpGnJDSSmaMI3djU2CaugTQ26p2+s7KO3lACkHV3FpzTxJ4FgVAi+IjJQh0IVg
ABYYCcd/VT6nwCbmtQjIrmMJK5PMN1bkVjnQkftV29vFbcrEy23W64UTsQeGvvZRG+DgqghHH3yy
CLeI54SsNFJ+3ptQs/XMXMbmQZuPG1iKRyyYAii/d9pSBDZzoRcx5EqJjaQLIouDKtFETrZgxKNx
Zj12+ZBdjF6y8URUkKNzVwy21FN4/6JdriTwUPzfipfns33HvcEeWt7/OVvt2FzKSfBxLo2vQuyi
dxG+Y2cr418RYhI5OATgC6Gy+72ZfpNz6IG9FO31TlRuSauZtGrOuc2l6Yv7s66Ny+d3w+lB9wWC
x7MqrYpKffl5vI/LjQG2kW6JHeiY7+mM7DY6TYbjyredPYRqRM+1XZ87GyGfq0HsCubHNoneOM5c
eBQAlJZmZM9ezgBtx+0V3d0rO6ZlcbsgRxq3femyCYKZBTGR5rN2gNgSR6kdNiVf2WD7CiBeyarO
n8oczVLuhayv/axVJ2Mhz4C1E3+vtqZWgYVB3S2lzyhtcSCw32bQVFW2YiSz9sPrAL2D1fBKjFAf
006khz7Fc9rJ8i5BbsRfx4/JDnf6vMbUYMuySvw9w5+b9iskdNgzsjdouU0IOb55UOVXbcjBT21o
E8pSSFmoKVdsDO73F2jFKq5db8pwMogfqpsUmgFRJMfUJ5o3yf2f3qJ3CgpxZPb7nkW8ULBqgkWE
FALUIb9MQtLntUh576l514ff7AAAfra1ktFCmCjNP3in/MTb1AqIJ4ZozydunKpHpFeRi/m5QsTC
acUmGdp6fBMbaM2aneZvPlmBgtpNchuVcPiSwLwNP8Zx8W/XfIvHNSqS5udQkmxd65BPzKRyX1dQ
YlxYa3eZWau1GxxW9uq1pNot3hYMogTnP+gVJyMSBX08xgPOcnNjhyceCTGyJSBq0MI/KodYUTeW
1r8cCEiFwr887dlbYRFNjDtovq2KiA1tlzB1YJLI5VO4GyM5WSprKlKhJaXLUJaqU92S0zFu5lnM
+rBYV3ZgAutPtCBUU2hrgEqLBw22nCMOobJxvdX+9aG2Lt2879O8LAa+X0wjzZ1+Tjixi48IMy57
RPb67nHq6I7Ca4CUYPuKSu6vZVGok7VHX6PgOjsNK522XoBbTNrE7G3oHDdhaebuNqR8uPG9TNvo
umKZWCfJvxcTV+b+jwt5iQsk+ygu5jqhqzJU8W7XkZ0f+0yLGuEuvezL4/LKudq82/Dnwp8lRVFs
CRxq2HUYPfLkiLcfhTVnTR+PKcufLyWfqkJHR/HWEh3/6hpifCMKD2ee2ElaNC528YCRy3LT4tAz
l5oIRChHQR5QpMU5OQmh0l0KS0LMIBxLU6CNEgci63XgFgIuJMIxMYZpVPswWG1SQOkgUiJagnwY
u/SUzCdh0OXWIz8C/wZT2q/iDwj2PdQ0iPB6vbacxaB7JOUYmjl46cK8s5kFmiubfhrOu32vs6JQ
XlZmg1b1we9DmmmshKQvfX8ep6YG/0KjttjcYnV+4vBar760N1t5p7bbw0eL2trTTN1TGOacy90h
7a2V3P8nQVH9QpLfT99CN6OCuUBGOPiRNf4j7U9jCPmAdrhaF/wzlGtnaSgQR0E13Izi8TQeAmBD
xedKwPimacyrkGA4EPDUnBl8nMFG0UllGq8gsOeLKJxSu9VIsPE/FOfTrNU24n+iwLGT6Axh9kus
ddULkVpu+//8zz5kzp4DjoQzgz2QxLKLBAmPLETF/mMEYJkK19tvlhquJypGI1u9VK3jySdiS+aJ
+xsCnmNv8UvoDHt4CXIaAn4Lhtvm6WHWrMjJhy2GSK226MYcf0S40tod4LRAT8N1SsApBY1JF1sY
rufKGtSRfjjIGTiDpGDgxbnp/De4mEiiSoa/Pgcc3OyMj4JF8qe3GGwVK5EHUlP1bRWvZ71fYFSB
CpWOPOgINg2+w6bmr7228xT9DIwNFn+gqzyw0yN+FdsJ1D06NH8Fhf+kWWHsaFq+DIPgCN+nesCb
XuE35WQ7+AoODxscOhy1PQCEHQR24oNWqCpUTJrqeFTS+KuSH3cRV0beB1mx0a2ks7RhaH5LR5iP
AcWUSdVF7ez1s3Pe6pzpTIQrCOo6wQoXDGn7wpXZqWWbKxD03/utg8kyIUBlWbH9TFrD/qQXSFSy
9Rlyj4HFD9RZTAlwk2BvYL8K3wJchHeOIPqO1N9MAD4MuqYHL8fi/sjJ868L7ft1PKCNZnzEoG3o
KFtTfbP6VGzKyiP4RTj3zSf+7JzvvYPuUNUxLbNmBuvO5jj8OGZ2lOLhGQy6dab69l77Ba8qHGEm
wLSmjlGz/Sw7zCBcCUzYT3RMTe7HajKb/E7HGawyDU6nbEXS/lOtDreuFZnooR3z83fGH+d6IKcL
6fQqaCMQo+BC2697FMTOhuEmUYwH3HmV1S+Os2z+a/3wY62G1zvSZHDJG+PKSaCP6QELhp4sN0H2
dmuJpWoE6roMvAu4pmUabK9ta2hZy+IPCYCnWSXq4EG5V4+avL4fFZq+1IfThNv7cFh7MqXGTAuz
8iwINeWZUdlKD8a/1EQqEMaUd4dhH81t7J/TVeOQX07e1zM5NJ5CaXI/g/hQytjsQgJGCEPeOhb2
JboVzVBnzzhjdb2bCcEb6VUazUCr23RmTkCDHltC5W16khL1+M5VPg56KmoYIxHT12Dvy3Fd387a
IqTjuoc7JVOizg6AKvklftPuLBPzBTjMc9rkcLV8DzZ+s1ZEUbUhQSQfkQbhUopoSRvShxRuYtrl
gnqca7frAFMKiOkhA5HJLSzv49RAaN4SbFLdDAzuboWxN75ZILdSVF180O5wBfMoQgfQwWL/1O2t
bRc2/zBzTNeSxNxodgeKBwDT3YXJCuZ5jaAU6Tbck1R1dpO91PaQ4X3lKhoT6BFLEL685KEdzq37
I5SG/4bpGXrzk13tHhyi8JaTuFEOk+VBg0xjAz295LtngI+vudnD6zhR/C7lcsUmE6zDjg1kFiQk
yPv9tmcuqEJDOHTYhiRwziSkYT8jMHztgdQl9DmUosStmZARMASd4YdpWEogOHeR7za68Lm9daDQ
jIRtp03es9+7mRoKUpRGXSGgCpCmm/rOp7cgY4WvYle91oF0pQpDD7DT9TW2hktJbJb1glXC7EYs
xhKAzPQRl0IdTTFeXxc+kwN4nA/gMxzNFl0xmvZkkF262zu5ufVcGzpe8ZjlvoSArXJ5jBIgc2vJ
qPGeQgUADxaGoq14aV2LFnofLe/L0WQXbT/39kJ3FMuR8uFKMQJE4aY1upPKd+UpXg4IigrFeyMK
602SvN7uGB8msLVvbifGUcQ3Hr/CGEVjknz05waYQhKarqF86byZelCw0jK+cs6ZSW9y9FFFC/8o
TPVSguDKX1eGgd4zG1wZ5PKBTTAMXdc/Ku19QYMW9Cx6J6OaadRAFdg1h6gmcm7fCjaba7X9i66+
FnHZUBugedj84k4Py34lsGD7kHeAKRAlxCXJ3nKjnEmXA4d0aOhfFjANi4JnydCaDFhkXIMXMDa0
Dvp6nEpHzgukf+HIwnH6I5qBXCIrwHc6VbHOebtBriW8+LoL1Z0IITA9j1vdLk8aOHLT6Xo8Kr+T
4oNYgrcoBkuMgtdJv+ii6cTMiHfR6xhQWKKCDSnSbvdRur0BYVtRamLwVWMOG47NxaZS3amwgOrX
KnJgn/tm8We8dt8uVi5OPb0ScLSTUNVQJJjJL0yUeRCY9xO9SMbOGGb2LlQmetuht+r2PZHGcNSW
oKWRohR5Ej5O0FJgRAOWNLQg8aVtPQaVQ8GpCVw+vOsC65zOcsL7COrKed/KukB+eb11wrKMA17f
hAZL0LR20YfnVvAAa4NVsBLdtq7ivyU/fYQ6MuIdZpQYwhxgw89S4rCQd0OtPz8lhQbgkmLm7RrQ
0uGYtDunZsPZxE4MWpcQsHMDi5a/Sc02HgclK+m/SgvmfUzwnIpmb+TIKUFtH8y37QrlAPQdIQLr
vK5H8w++cJi1CI5J+pV+m/rNxJ010TSL+8wHUABTfkZBkR9CJWw3G2/yjs9FfZcSeR8VZsyO/FlU
8DRwpAO37fj0wS8gXSqhi7+TcGgZXBjOAsJOtkIBVFQ1xcjsMHE0DwjxSn0nnVTiPw72j/brO/9A
PHv2ttIIqJGSEoZo4UuXsMVxssITP2rtDEvn81CVDEJ4cy6pQ0pZw3WqdbQhfZI5Yft3gmdezdKz
okv+w4zJ3XySk1Sg1AiO+X4PMdGzmZdPqbPsSDDA2Ar6EkmWpDwFeOzOb3BsWEU6PwbX65Q97+bu
SPs509VtofXG7d5cbXeRjKGPUPxccZMoCMDYMRPlGVbyWTmexVac/akW45biAw73Lvt3XSgoGZMg
ufuidZtgw66o3unc1/nmsN4t5IiueSlR/5fntbVKDUtkVJZfvemLdaToH61+zXABVHzZotHXwN36
XyqdnGhuCuORhwmSvfNABXeZ/L7zu3lKG5FJvUtUlngorvi4ph0sQpQL7W04jpNV5YWAuvyQ5iIW
vL1nyIAg2doao+ja6J9JE8WaHMc3XFHFJCODLZ5koqfktWN5Fr48WfASnN/ptimdyx7PWTvHzKOc
1MRpr3CJGJzTwnxnnn/qHH8UmXG40WJ3bEIq9I5phS2sQ22ZN8rl7FYIYr8/xqnAgsk46snc5SU5
XrNdP0/g9LhimcdC3E7r4EfHdTP9QrAX2R3KPcSm1tJoTzvxVDP43CiDrJbJsdze90sP36QTZnm5
kVh3mcEawwivGTq5eK10npsO4NwpDdomhjaWnNSU0HRT8Z/qnpOG33I8RJfs5/EoN3wHiyywjRlA
Gr9IHdsJQJn7/WlpVrj0i2N0femdoINXHjAQlIzgg5YBxcnObL7tmyNqzDvbxMjKr3gJkdQjU1z1
bnC4qSG9Mph7XtsSnp9O3UEf3hn8fCgBOokizsZOQ3qKs/oIwEb1xQ0rVV6nUUYu3VylJ5LNxrhy
cIMx1HbARUYUmW6hRTPlUSvVB/JdSBxN/pLbzPFA3rZlyPqd06AednuL9fpd8jYBqSAJ4TkezXwX
p+JWmJ36pnTX/K3SqyYXIKo1sb/gf4t8b7EQG9M0ghM37Ys4cTKzDk3Jvk7sRTx4gkb02UlB36aH
Xd/b3qTXHSyvUeR7yOUF7zTlXxHsR6ZX2/AtNrkZhTbNFvAy0PFIrb7LrmunuoP/0ZejD212AkH2
pa0rxxzBqXhi0VkmqoVrOy/VSomv5a4GmMS+wSqdJcpYdfmmb89pmULQGJx9kn5ZlnfgjeeKnMNw
Js8guoC4xAOFoEb01J6tplGSJd1aMIuel8iu7PbVIhsH/rzbpevNcuDdlJkhRDvpcoKoTp/FmRe4
1qG9BaEmoH2lJydSObdTDQWPw2OYuSoVS/xwEKwjzEjng9Uh8VkusAICOIFvlaQiehb44FDxBsw8
jfcFaM3hB3o7YGhuIaevBFI2WfAKHGpqgPCUo3Q6JMZAidYBkWonj97OkWd1Ywu5qznIcNXN1GWr
owi9VUu0R0CgtmXvhG3BLj9mHlQsz1C/08Yo0uoyrKoznFWKilI6S+a5kmuQ1AUGt2AFeEtHgCf5
jKdRRCTXkv8OcaYnvOCe0fvjydho6dYmdAgvlFof00CPxleNOyUhEqbVu2XNPuFcWBv3AN1+Z/ce
GtlJO2nb8uX74PHLaDu+BCsvqUbs5HAr7gFG0hLDjTxde8quVsIsrh9Z8Ge49jEbNUX3WLO7iIgh
FHI6HfZKaBWstu+NLIo3Vo+NwAAOPPg3UovqMQxV3mCUiouuCgUKkPwnXNoVtKTRJ+KQNqX/pJ+A
EDhKVspZSyN6fy9BAlmjqX1fjfrc2k95fBI5xivHBteqxsqVyp7ZvPZa1fX7gGZo5aKzvfk8MY+x
p4FzZ2iWKoBCqPwmiEjNCAsltxhPg5uOMN6g+9HTlFGDBJn3pkqTfQ+bp7hKrhAJgcQdXN+sCGQV
A8L8SoRIY+puAqzQ/9nTKscINO/ATpe6cjJszy+uRxQyMN/fec3AhjHUCF9ZH/Iz8tJRBmLlkxGt
MDJ2ImoYvBgVqBBcxEyTCWkjZgGFtFG7irqEUce362zu0dLy6tZ8XICetsyu+DKHw4GaU/FjGY7X
74uCpPktosWthO2mHuhc9fVn155YkZnKY7WnRES+BdG+LwpPPnvpZljIz4YZjSb1qpIKywWJ8sJi
VOcA82rF9o+9a2NFB5HWsEMb6HqZDT+uFc0IKiOfH4ioFenmIoiwCyqp7fIXDpZBdbBGSbYs2MVR
f6zJqtK0/n4AM3LWL4+EpbQPL+d/74Om2lbKJbM0NBxV0NPsIlJj9GzxdNEwED9KaiuWMhkQUQqr
o4KafkQLy29bLh9ql2VRVQ7rItJNIabdlnXoid3mQsjDsRZrxljszuc1aLpZWMXWbyslVjDxfkPM
2aaqaXNh8J30jq+sfkB4mT+sNGDP8XYjeXNmmBXi8479p691QqhipIPwygGI9B7eWO/MmVXgfLcy
976x4PybGJOXLE4bCWEU37UvwE/I6tgM/tZvHLIgTclFUtMXzRaFgvft8SHum70ep7B6ygi9oPXN
1KSWn4IYWviYvCwailDVjfmS7hpRmJUKPel7CTdUyA7CbAdxtqPjyeSqF8ke6t6LiJ1LDlc4s203
xvUsPH8E+KQkaPWHGlGug4sQGld2qo8Wi7yrq6f+heG2FB5tpYZ3Cbd4ULDnAVuq7qyR4iPCyny+
YP8ygygsWxarm/ZavJnzC/78m2uSiHFZCwh4yz647VublmxmpwAzSNd7JbOyM1tvzpBAjneGDbSk
sbZhDq8qOynDOPp0/LozgRUkwmBMBMEpcLS2m/lMWGerd6KQfWRwHHH0hWNMffNI0I7JvBZg+oYZ
x15PAdjU8+wnoBJp2qy544t9/SqR8P/CLa8EIKWDwXyFa96QUvcO4n4BQ0L0f9ia2ApzTNeql7KC
BAj/yT3lTkJhh7N29cPQtTLaltv7lnsQUxE43c5EbyfvQ4tIWhJFikdhwF6PSaTLLla4dhjaemHR
rnvfoxE1xlbbabkaSbwlWuzZO4cXsfbMIxK3EQiO218dBZy6osjWFifNO/l1HfssTHVVlHT/QWEa
2gxuKtc9K+ff00/8FLKiFRuyy2AvPzqdl4nsnpjgv7dViXVBQm1vlwuYtRCLv43Py9kRIGbNErYZ
VG1sR9MdgJSZps+FTbpDJ3YlFFrSAaeZKi8q9CB45jIt5eTBYNS9D02ZfeGX32ki9Ae3qWlV+HM5
6Ib2WcoJtl3gPUwzmoYN8mIYg9FIjQqglTRMXOXIxnpW1HZtVQOsi0uQkGQi30rx46JHiKQtxDbz
6/b2cdqD1jMV9Nw5VaVniMb0+eYy7VSVtfFySnn0aDv2OdmYr2ViWIvyShgtVET6VIAwPtr/fgwa
VNDtEH3QsqYYq1k/zy4bnbVf3hL41fv9fl8tbJ96ZlTZVt2x1tVIXHCnGPL0tj/Ka1BOYeSbSd3/
C4c1eP5OxVDap4kKyoPlLnyJBm3Rm/Y9fi8ZTyy/5PI/dCTKtK5s8ZSPi7WDEI9SsxnnaJUIRzA2
8lU7ahcVs1oMZxwBseJx40n37qSwtZ+2fOghQPnvcx7LrBj8MKFOFoLrhOdvroaiOi0sZkKcEGjp
wuFsVyHWvCXd9Jch7ki4LCp5pHL8AtBVS8od4ZafD+MR10qBgqryN1G001+T6G16jdEaekJF34Fj
ZJNGXtc0eiC7WYEvMxb2d9MLBAvIpZ5CqiRm5C4DUlgh8UdhZU95XnYKUsmmmWwGqQhggZx2lCMj
RWrBGaPPhwjz9v6BZ+5YSaggXAOHhIGCxd1bKvsOSLbFY+ftdrwtt/MwYLioCnE+D7cvYix92S1N
159Zrku2nYfIeyQggkZPPvlYWIagZsmxKPgVBQLpVnmNMI21wDNve6APjRWGWHbtgWnTcdqPNChV
jS1MW8UJ16RbrL3TfiX5nXbbQhQooI0F2zd8U2ppgmDzkZBJ3QuanwlYbiIOrUjJk1wZFg1fbmBF
P/CXHLW628LlsC2eHKNHNYoLvcvUrtG3nDotMwANVZcaKx4XyIAQm4lmHDHZyQ1TTDRYvK7NThhH
keuxX50ziHrrXfiCtHSUsEAMQBEpl+Amiu84h6zsaqbq1vGckql7RRUkV0oIGeMoHqUb8ko/+EdD
HRYe9HXEmhb9W6Z92DmGoFfw+ELt1P2FBE/4FeG5GfSz4BK5WhvxOeW+MBPpIAj8miZluBl9Fqva
dxQYLVgij4oL2Jwhrqp/6/A9F/ZcmM8bPJwTLmJkxM3u6KVR1+41t1F2VwlWb0RHbFsAV9mlqi22
2Ku4b3h259f0OncOAdVmg/Tt/ACYpf7phnhmiu53l+rl8ryfqQzVUH88208plQi3qAYd3ol8CjPP
QWklFAdiWHerBooakTFzCHRjZia89Q4JcI5ARALSLVrTtyi5HaNpGyCcadYnc2dFM6gGE3DlvPTo
a5SzrsLfg4EuSW001iQASMZUG3rKJ4OPFQBd+0953pwiZ6XcRPOd5s9fpuzZH2Ic2P1UVp04exfV
BlkD4qEaDAklFar27cFkJtL1pT9yDAWRElcufl5SJ+2NSWAhEp/nqWS2JjusYelHPB/h8jHGOga/
TETOKVj0h01PH1emo0bJZCYiSR/Hp1uSNrHUcQ9L9GDnnXIJtAZFu1WdI6Pl3h1axrRUP35hAoft
u99ZK+Mjq+1t1xcE9q0LyGKOxe/4epHDALxQlH6DF3kwnHK0VAAT0kvkX7CGQIz06/0no64XOLK3
WjEkATB48mj3SgJgi6D3Wm7CNeGKMv8Ibtn9s8ehzTfMuUGidHkVegKsy7INKGsYbzxFbVjJ2mge
cEa1dMvigHvPD6xjxDN/kL/oMHfPNw0cc+iDPVMbB1lGZ9Lw/GGYYcGY7AQSVAbQ1KYXLHMUaKHe
SY3S78mhO1pHvL9pWwwLuMAR3KFFDNUxYgjN2l9Ip0yBQCfpcaJZh4ZqePy3keMZtwVxSoNYh9H5
4cxG/VTGY9vbGovxqnpC2r0JADIIbD2hDbUzMkrG1E7nUQ98wUiRTJLrQnaM4VGAqE9Tjr6zDOts
jn55A3KPZWTfEWI14PrDBOyYlA67jy8uOajGqHbNfBJeQYXK+RfW4igfHsxpC6aLOPK3zWVJ7yAb
wn85U/n9Zxy/Qbc82IfLQHwB8Mh5Avdse++S7iyWY+TgNeKRiRk+a9E0VoLa1AfE8g6tc3QZNbOl
AogBOZ72Rj07iLPe0lh3Gb8jbAPVaeN/iGSK8SQ0peRR0W+2ncSrFVhWi/FzMSxi/SwGaCUTEkSC
ynb3AfOydfPecoPOGytzEtN4m3m+dbGmJa/2N8v9Lf14GJ3zrSIr9bn4LebNp1CBLD8l9zLiufiO
U/EmL5cSaeZu2K5vPp2TGTotTXkh2NT7TC3XxMDgjkXA5g+Fugn1o2rbPMPiDxiZkoW9OlnoDmIe
cWWjcdoGtxnNus8lqATNswoYWSMLdQdSB1fnH96+hB8PFLTBV7esnoWttMIeIB5RECSQmMzj7fqf
RbaXX8vsQAw5YBy3qBUdqHKHuS95p5KU5eth6JEfI2XlSas7OCfA4idWmlMTNxYJVR6Hp9Uq6mX8
12s0OCLLHhmj5/BZhaVFolPqxPaP/+5sMOPadJ400/7FDyqbDWkF2y1a9GtFCzlkAatPsitkdNke
+ZMnqp/4puS5NeJwqs7XUC7lmWBwG1TqvGiMKqvXdH4Mb2h4ioOknUEHrCgmtpqrVy2evRR8xTWd
PN6RnUMFGTr2n2Yjf0AE+BYXSMYsUx8kSyVs36dwdy4gpuxS3XQUpwztu/F6QQuRKP5pnPK3pcxf
15Rmv3ywqKdKeqXIel+rCV/I2bfcveUuSyfjciHDg+9fVlKRJILRGSSrSPJXX+4RAEhFHh/6WPce
1e026WkWXgA+WfPgzhCS3TqJE29mVYB0VK9L7+aLO530ClOxjGb747KHepO/A5UuUWvBmLUh8hPp
1rgMFXa27GkHGgTXmrKcR2Ruvwm0ow/RSFZM2lbLqhKTJBCWXtvh53aNFFgrx9exMFvUcJeW+mkY
kVfdMwNdRW1v8ADXd5W6/pQYIMgUs/rSkJXh6AgbtZQ2ErZQexZGaPNjjL5qdvw9Dcq9QtBqy9i4
Nte/tZtfuj118HOyKCo62ax9I+sdCQVo9ysmCnKC/wsR9pjcBJ0cDVinTfe3gLdR2UM6XswF6ndJ
Xx48ph8rzra4lG6EgktHl3NdAWWoaR/8ZTWHGp1tIA0CuORqAhZQaXxPwomC281u+lmkRRHqywb2
OCyi/XqvWZqjOCgkJnSyNnkDTd/bhb0qTf36666s3opvraK0twzCl3D061LoN79ovmjh9cvrO7SA
8e6VIKKuBRaSwOTA5QNmGifR0DXi4Qp9IzwQmfCZL39Q+qrFTi1Fc41tQjRLQNNc1J4U/32e+JVV
horCVRPyIfKF8blHOZeTq2l9DiUSZ5VwMfd1SlH8u2TSJHe5BHG3F8CeJ/etUPOEkk7mqq5TyVuX
bliRbOGPsNZVKAYoEYhjsigFkaXH/IkVxBeeV3b5D9qVxk1+EZpM65jqmGxO+i61F8vmxPi6tWxx
/BJuS/1m06/lmx76JYd7D+7HO0gNZmQsFiMzVnPTCMpmfSSl8Ttn0y7nBQvQwNI8WjMvuH+X38uh
QYuoDDT2LROX0NCmB5Q+KMqmliaHiuzy14/SGi3uR63Lw7wV+O40HM0lSfkfQz/96Jsu6t7ZM41l
4OcB7muimdTH5oJ00uedV5OoiQrD/n+wvbZv2POPY+AfEEELDm2QkkB8yid+zejSmMUgILigdty/
HY/U2aH5/SBg2wkV5L3wkhfInJ30PP9yCkUhAZbd7+FJEhbKch/E5pozn2spVqhzRGGrGos8UzDO
kdlwSvu710UW698khJKluH3Rc0z5UWm/vSo1yxFJfSz0OaNh8MjsRhaq1D62foN3czetXDtip6oY
1HfkRna6BmMuC4jgT+oa00m2cWBqx/8RtRexiCpzeAopoE0NeHn/qUO0/+2PfKoNWGe7IqgNuuZw
9bK+AoePfvbO7weh2/beALqCXqYectsPvBGAh4FiiI5gJ6wCIgxPdSIwRWRrzlf1Cusy3iaUMyqj
kAQK/pKn6G4+NIYwG53Xa3h5LMCL2P3p+q22YgNlTkmrkXb5fSJpMz/672I9ky33xPfbX1Lf4Hz1
XfTqbZceOsFNcXkFR3SJlb2o+qsVDJC/Oah6t7D0y8zxGlwevmJ+emrDSTPwc8llEZAz3t3wo623
AU0a1MS2NV7n05EOj65FumQ4ADnQtoGKYLgyCfXRGZyIuexx8lTYH95kf455y4lXbcXRzQuRh0Fy
yoqH7lqAyZ6ViwMRg8qAQFW+pS/fFc2A6j5dWOnS3zsNuaSLYqYfeGjzPsex7ZWJSx5wAc+u+MbY
YGjGtyel+Q/n3aAmj6u/vve9eXJVtFCD7W3fGHFaqcPryHLuiW09y8loEnuTsnUgxplNsJpA7HTW
oLt1fLRUTyV3rGFVxRmea4vjFFXuCLn+99wWCoYkgvRBdLQl/xdFUlaNFDLnVEq4A12UC+bAW8Ik
O61f7O2VeQHgROFHQM7CCT6sAtd4HSKm/rHOgd786iOnhFq2glM9OKUBUpTTaCgXI5H1GOWNvQ5T
yjy+t51/L4UDTizfOHBPfxTZ7FTbJ45lzPwuWHvbIXo2KMeg4HxtzHjQMxKk6VVO7TEztGZexS2L
jBM6yocEKZQ0fviO142PPMqx/MhnLw1NglaQVHykfpiFzWx+59GTFffR24/SfQQGuJL5mC8dCaZG
Y0mNvePpsWJA3kIAoER3JvYmYE9+ZLAamuW6aXkKhIxfDSJOlOUIby4AVqM9AdmfQXp3/Nriqyko
a15Evr6C4sl/1bIelPav88Mr/Uc3161p1gyRsiGgCSGk/Bnst3WgWSGlL/rb6NqPrGEJv++DbKh+
kJnlDRwOb1i1q+g9PHP5uQ/Ut3gfu9WPHFZioyt47wni9zML+R25xEG2YyDzLzx1qTUIFfNY9H4j
zaCFEJ1/iz/FqinFxqsKw9KeHkA09MGwt1ZkQL632s42bmOyJQmSc5H9GxnQGYcKWTklMofC+Xk+
grdTpswqbpM9FoVFQvLZSRVZ4mgwtuVpMUMJ0fhqfys5gM+bxIKNe9v84ob3s/otiITTh2O4TBmM
1omcjJOJSOkPD/oqNSxqpwd+xqjIvoO8oXRNnbonsE1K4aC65zHEsWmqcusH/AQWp6yJqAKaXu//
P5YeiDf2N8K8ByuEE96tteTgbnnFc7miQflKzqpCwCKATPp6E6EELBfkkWQytIcJTRfhwVhFviwV
dEuD6UolJzUgJO2zjgdegna6ws+esk2hy6Hu/S//0Sz9nOwaoonWIvfAbfzm9t9z2Xn0uVag+tcf
5MUo7odsoYfNKE6pd5nBDJY4HWJcWJMs2OpcaZ8E3ubD/kaPayooPGV5meMIzN27XhxxYvMaWYQE
B/hhP5qIiSGyVTpEXvGt3+q+cplPrl8mbTrML8ulVnxieMJr+JvAOCjLcM7abUc+sJko0F8WhRar
r9jPc1DzzaXhRuwhWKyxed/1MgZQ/mraZmH5KkQfTlhJgyxNZ7DJLUmFBfYpeIz0+1rsKgNOq8hX
o6+xi+EXq7cj+dUxqyh8SZqpkDfOVRkDq9Cqlt2diOT1TsaZhsgUJCHgHLc0c8qx59ET9pHypQQF
rB1qrj6IYoPzMv50JjQUDC3daAX8F/KUGLOw0ZsFiYBO6983Tz19T2C0Bm/arQf8SBT6GjiQwDie
jZyC8ioFIDoPrbz+tk7topOXzUNi08fqWJkPiJwRitVeyvq9iiV5nsppbZhplIosACU4p6akKhER
i23ikMebGkFTzbbHojJyNbWDZo9PqR/1YA7BcNYBlKyWH3jwnFhuuN87BunZKnQ55M2v6D6G1Jad
Axe7QkttK796xEH+0H3vl+CzpvcKoS0cTFtd842JmG/Fw2khiWpuPfEuOBNAWVQDKb8WVKSRXpoT
4TmfZfrT801l4leFD+DlBdpQCo/6MFvi7YmO7rQl+JLNKRIJNwPgYBVmRfwXaxGgWRvTIsEDOHl6
2BN4SjsBLCiiJuzr7JvdNq9ILZT1CfaULJngDsgu0i9CXaOrxqMiXEyjxQ6ZVdFBsDACx0fjbiyx
5ovO2OktDi6hN6+CFYFMtLpLI2shaGssUSAVhRYUqthtmeKXPP8W0MgW/RSxIsttW0ZuaKtppHZV
oW9T4emSnJYkiwI8T1Z5OBgUJ6A68zgd1FMUeqc2RqqcYYNOBDfQca3lN+dotAVbuOeQcOi0ioUk
xWwHzl6ds/7d0jD9VXyYuo/6cfRb/u6KmgGMMnQELyT31TKAYXodH1fOBR7DoamGJEb9FZ+xn7kr
TSw2TXNWCGa8x3xShjFLCMopQ0Aydn5SdEsLsHZkDL5bvwz/NqOJogjjYw3xuSyPjRaGUWpltK8Y
S3CnRhPeR0Q2LD9wFmEiIh9F1omFZWf2DsBpFcA7ugCoZDEIzJoIiiFVaER8dsgqMVFTaAWaW9TT
hehHTINoz708X8t0gH7JqM53uWntWdvk/fCjivmDlfqB4tU2w2IPOF6J4RifTwC6MsiK1F6Bf6Nj
R8K++27hAPfIftUs02XDyjdHrWM3kNda2zG7h624Ui6/5AY6ay4wUIr8HCXjDQ+LiXgXfV1CUcua
8L5GrGl6YDMW5DSy56kfASYx/sWMWg7e/UKHKRnusFJa02zL0GZqiFoGLktbFaWqir/2HilxqZyr
PWzOxBqkgwXyEKBcGn6hGprDoVWGoWz6JXIG6qwiOp8N1F8wn6rkc+DPM4M8FMBfqSAhieqqHO6V
Ewp1y7IxJoKudXKhPqRJ5g7dsOf9XP3q5C15KXJ9NJ0Ify4yP5KcnJXTsR7z1k8D8GBxG7BgSWe8
ZDDpfZByhy2b9pY+TTKq/cxQ8C9j1PGYM70T+BEUvmXJPo3CfXtMWyYBeycldeJDgOYCOY0vQ5uS
1ebWVIE0HyhFIEeRT3/opNsFNVr+MQv0CrKZbN07pOLJp5PbtMw4R8tZg+dG1TS5k9abSunsw43k
iRkY/75Mb8zQIk0XuGBHv6ZVg8VCUS6uout42V2qBV0YYpeJ59/3o6Mx7I39jAVv5SxjfPv+/4m9
aWBCWB57GTgJO2lMOfDuDohhiP6avl4A95bs37Qxk82UZVcrU5YmoS7zt6Fgxge6sOs+ZEf4HGm/
TZjx/byK0gYUjWrYki4uBnPajYM18FseO1regBQ7IS/DJXsdGga37Ya40etOSaHLyoWEzxj6JeUQ
cQXB15AVINtwSbOuxLziHB/VtcclA0+jEfm5x7bf91gw/N6PplLNp3urh3WgFDeewsw82WFLNayS
dGiXNcz4imnfQR0yGUjSHTc8Ah4/g5xUA9g+di8J9Ya30zEPiKPDHJVOIw8+iUOLTdhiQGROIolX
3vSOD534YywU5l06SaSlcWoE6x+gOP6p8RhPrJHc0sJH3pGWI1iZhj+9ovrxo5LITdOzLQZjKMkn
hnT6HIPSpYvaFmeoi7JElIae+pkrxHKmFP6CjG3yOvKDcbjMEpgCNBTtw53BTjqTqfCBBprkSlAz
w1wAHKYCQ59SWivVJmprIRWh6id78MsnpfQETe0qemSDsGddEUR+4z++EdDRt43XlMhMKhliYYFa
klJqfwiqdA5ff4tN5WEQjPxwVznbTp2U1JHdEClK+n9CpwSorwg20zTIJZePk6+FaFI77kocDcwr
Bdp8+ngzvR04nvXA7GirIk7W/fEryAUzko/vuzG1N1fU10J9z6JBTBskIolykGmoYpKnf9SDFjB8
AiuN7wpurNfmAtHAJeWwDJjWovNflNbBdaFlzjOohs0NXXeC8WWIttEtgMBxIjxF5vAtBRTMVHms
FqrRM7qI1hXPvCjJ2k2IrJ6IQu6Kaf7Ew2u8L12aq1BHq9aS2v9yLgq2/qq/9z/OWDVgCzMBk3YU
aMgiAsNfmx0xC5Le6tnj4ldL3qkaMHum0zXvGmt0MzED2muhXA+a26MZdMZF0szoCbv2xaqiDHBZ
ijsMliw16bezj5RlBMV7bIU86w0TW6N2NP4Ek4R+knwped/HhlGRL9w6WYvhzlkcDY4SOc/30GyH
ZDZT5d5N/EdrWFifkgrazgoi1nQuZVgOtmx7/36TmnJVkR3KJ/JpRLmdToAauQQ9GyCW7V9DFzFc
A4udjk4O66KU33o9pbszxS+elEFwfLWmLXr7dfWtmmqjO1DMr2qH8K6ys5wy3hl0h1DLzh0DFBQL
kGuZIk2oY1H/BkWOPQZoorGBaXz/Cg1zNAvppuD3QQpiSSLGhcxlXZ6LTzlIJBeSfwX8lC/A+/Qx
rvoq3/0zaUk7Y5FaL5OezJizQ5vb5axxOFyUDht8v3tZd31cUeJrpDLFKtweA6wVq04ILJeNNXe9
YOkniNTqDHHR4cd1flQqlxPTsdVkE4ZQ72MNMaZ8D84ROMvQctjmFw9j2LT+IYp5BaCg75cp8i2m
R5BnVB1S+uJ8Z6kyl1mbLFRvBB0dzsLpHGbHJQTpJYV66i50wS5pllXaR0pCDTo4vDo3OfM7aft3
VJ0FcHbcAjdSV9snioUO8Mh5Gf9Bet2EO8g+dT76qE/Mlu5Sd8K38QW/5GUl2Ae+LgEY16fRUegH
VUVTRDarrGqEejYfGmeJHIbXIGP10d3mkkCI5SZ4bd+rSIY0sMNBtBSbmyP+zd1ysqjpFze0dulJ
qmv0ejjgfgQCtJB9XHcUMsNqByIzUxlYBgB9kD3X5ueddoFueqmHvFcNB8spLaBgDF+wBUTSkm7O
pKDiEvzJboL76NHKEpI+L1/GDJ7q3K8JM9Uz4/MgrR1aosUVA0/YdX6l6A6Wr4ZN6uUvCOZsmeYu
+VCJg4Ddsg3jl63tLU9t5jxU+2qns8MpfuDQAp43t1+zW4GEeZlZm524GXReqgK/rZtaSZdp+o9w
q/UY85/ZUN99bMh6aPi0chNcPPCKY/h5Z2lzclvyoXgJaoDcVHOdaxhlM9SB9DjgeaZDCHbW5gct
y+apuS8TlOQjz4E6HstqiW0dnfND8Je1b4mwRunC9bPSbwsLtiVvjCCtDab2q2ISjyHDYQgfg/j0
kl6xbW6e+3vuXEvOSW02aE3P18usxulqtmUphD8FHKsN8uoocGbfwoPH5jmjJL5JteJkcnGhAWvB
/Puyc1O9HMjRgY6jt8crGnvbGTSLxVBcgzJPjKNTCwqR4mNthdgPhP/5UqkVHM8UQUd/HzzNpRhK
Z7b1f7o0KDq+qzUcCU4Hn2Wko8yu6AFVZwT0Em+KUSEimIpav2p9h62kEekQT5fzgqITPcqp7RA+
dbwG7N+8MQFOoOPFa2FTn93z9xfNcQVHCJSzUJqBU36x6x3p4DaJv+VoJzDy59c/Z+23m++2YQN1
enTkARKsqtGrbpKTb8eeamZ1cg+Q3KqfpdtqM6x+cJG2lcQMxCZ3wtm299vZ2leG+KNrfIOUocZp
9BGrxr4oqhsWUQ2UCuz7UrVp2J/qdYZwvbGXgTmeP5cK6fQAMsRG0Y3PL6tSsxK5GcnxJ9w0MEdp
mHLk8Rw3BZwq0GIFBFCfSUXTy/atnzpRNhZ3TSbXL8P6QxuR7H7LD11cGH5s8tlY+a2xkIuxvZbh
2n3utQqL7AtZSR0f1CZ2ZDrw3mROV7/2NiFbMPd9B3wU1gZzff2frK3wfRzoH37GdkErl5IFPXhX
Zc+ZHijk1Kk5DHJ9tvk/zFYU83IN4XcTrHpHR/pIAEaN563ViiZzR8UcGYEKKcBe6zF70vqz6f5L
I3lC/D7OZMHPPnOzi90vaYzG/ei7WdS/a1FTUaD8D0vsB71ugv6D1vo3+sESs9gMYkAlDCn5wIxg
IVYsk9xmMG1UvSR5gtDG+qlLvW9GyzizzWmoGk1dbzstUbmaZXjazLFoogvgpRh9XT5a+7Z4od5H
Qf4QmXmYPpsPRBBS6e4aN/O3D1N65NiK7SgVB0KNYzKxE8a55vCiKAld/p25ejaK0++XC3/gDPSk
s/iemj1PvOv8J8hoz3PLLEVmuaIJ2BGNJ1gQh5Xwk4x41nSaTLFeei45Qqhq0vcpzUt40fhVaOap
zwLJvXagZJSlY2aePGLpjI9zDMIzacNauHuusKqzafX7EgzyvyPmGSxk0/USqkKIzAtcRCCqu/x9
VBtJ8ehDHHb1ka/aCWjz27oSIiuBcZzoN+K/9Vc2COVH/UJnWyRnFTSDGlIaPIkmOuX94bZzlJb2
rc734GeKXEoHbBYGcVlFBUDmSNtFS5UCfpkbWijIQCv+FojTlKNKmJcX0oNZpOfZM37xwGFnivYL
GA48EpnakX6ritQqviwNAqd7zJxizRFuLk3Rxoa3QEs6i4WQ4GGV60Lsk+/KnaCb23qeQc+9BS1F
yYGIeZBW448rtDGvSty5rEmO6DaBH+OYAoZFkPLxi/vB+zXJYYPAqaa3MrVRPj4gcSSyppoZWUaB
ZbKS21yktV0Ka9GiAJHexm508iqwJ8ceMI9gGcs5XK8BCzHTjz8n75NuLQjiZ498wTxGMgx2St3h
AVA1PMCBwiqwA1qMSo21WrGvzHwGc2NqaW/1A5jmRPVtVxWTNFZyS3f0QabVBFPSSGBDTB5cZ1sD
SF8jz4Z6u2Xpwaap5EiguVNAYQ+8WAi2xFmFxP9wNgl09CFWU2r8lTS8f5bOZUMq9lI8VOgjCwaf
7oKleLmHpHRwOXB2xuCaysBmKXkJCX3eRYhSewqyGJS4DbYLnz0CKHehy0aCo79mZkgXLCTotROr
AtDB4jPKddANhNfq68wFiK9N/tq5h5oIdYAmg/olFfJRJdc4l9kmmpdcnwsnsQsH7eDhX593nNN+
Q4X1ebSZOgE4rxmPqXf7JvTy6jbWnJpretMHzqPbbGyM+8UpmlrWPI5XKWx3VzmAUrTNAXPBj/Vl
rtV5PKLfv3NusIIe+js0IgEJyOGVc0QTaz+/DccMu1oPdR31i/zXpFbc8l/rg04ApXZhB3dxcoJF
EaKxJqmAWzC9Di+IF/QE7ivJRIVJnftJ7Xu3f15xsGr/aJNfYb73J300qw3qSnb8X52eyaFt208a
XpsiNIkD0fYfVGogUIMOyoNXI4Qzks+OW8kyjIvq0WS8aK8zJDpYXg0I+/TSZQvYPj/yQO8IPzIJ
lEAMHZ5kel9TTXP6Kwo0reANFOXPCbyAFAx4gh3wBPErYaftRhYAOPkbGp+J1D7K+SZrK5cux+u0
5sgu7EzHxyQ9JzVMCm3xTKHvN5tD/qio6vg514SLKwY4Pmp80sox8+ilLCYvtYxDseLx1iTpUgrQ
vEWk8Ue35x7S9/lqD7EbTi3DFSSNpLrV4Ai1e2rjS721enYACf8x+zuabzdnnK2gaaWQenCFZzR9
co7oTx/JqO5YBTaFRW0WS5qyFz5D7/Llwo7QDBl2Q4Cd6tzJ3FnSFFpJMkDSfCcu0kaq3oFBBe9L
0ZExP8ZJhSpNQaJGJPwFNdJx0WJS7CWxIUm6OUgwY2DGtkcwtgvhhyJyTEW67zJPOZ/XHgCpWdAO
Tjs9ibAeI3zZeI2AAyBb8NrsfQph+SemZC3085BdDpcdG62nS1yN7G9NEVZ0HxLLm8lLtV2Tf7v4
jQo8Ij3+aRMsNEo3+kLLG4pgCI28lCsqJh3cQRDF0KNqb6Rqi7ONaq3/ho9SWTyzCJq+cTefUb3U
G7ss9wGcXG8TxiBirKkSP7poYiQ+VBYDo/4vwzc+DTQxV3QzsxgVrje+e/Wx8NJmPtmrj7VfXunM
faYw0y4BkExGq1GvSQKGdfNCcagzDh2AMDvTG2RIWF3RQU6CUt3juZQ00nIwqTbqUhvLtG/yItr7
eK76WuYvyeQYUt+0uj5HScwWz68S+CaraNBuG4DsfrnE9Ox8fwjQfYm+wjKWkUysfz4cDRM4Bo9H
igvvE69WkDRozBIp+t1bqDi6btEfK8790NOsDbe6QGsrIuVUsHNPEMyfIzLzXvpdPpwl4djNYwPY
jbKF20Ux11wc28hIlW6pNg7IreLOjLMnZyY/4bJGQNtDkWGlC31wslBgQ6QEFL/nhYnw22gzGG9F
CiBeFb9oZWGK6MQK13KFx3anOHUmStmPmBaPUgl+69o3OTjI09RbBHaQQDSIQbNhZTruKVbPHKoX
YB2JIgFH7+h7xvinMuDTWqMfyqFAuhlYBkm6P/TKX56uGsiCYXi7AWjSB6K0AcM7iAjc+u9S78oW
x6yeRyci0ZEvP50UCzSGDGmaCW2xebkRQ6XGx6+2IsVxbEiqw+CmGjgBfl9jsb7sTfoEAp/wDujt
qAVM0OCcb85tIiJUwTCojlpBrGn7QNjJmc2huyzR82w75pAf9EZ5jeLHRIFO/vd5BgxgDJAzFbJC
86zHMFlV9QYh7SFjmWKA9qDpkIK4AtxfzQiS8h2x6sJf/bgZhbxxv3scPq+wg6bMLHhpLRsvV2lN
G1Yor0nv5OzTSJCY8FlVz/6tBa3yOaKp9xT3lboMf+nYVuXm+mj1MYiGxBNULF5XLqk+dfTJK+Gk
xTW44B11rXG4waB9bUH3wFITVssG8/XIznBDNym0uvJ7d4+r36tVx+PudnspDYbCuUVTT41KPSor
OJUWq7iNnIdtef7UXFS5zD71AKxTGFLRFTeTwB3Zi29Qduza/DhnWjKg5IIk8R8DnBGdkAj+xjM+
CHWFrdovq88Ve4Y6AGhKDJGzbeUVfBfw5+hrcLM0nRQOoH6EQZvXRf5PHvsEmiPviZ/2M3KEPynt
fiJlfeXq3A2yu/wiSUxTZqovFTX+B3eZo0wxqO9OAUpWrnIoGBbKjCfFEq1oXuq07pIzwxWJHDu2
iEfxEzUit8jLN1w7n4JGKHInGQaeUgEO1pjzWmAJ6li2wkp+Pr8BEsK03MGOSElnMG1F2ByRm3XY
k+sBrgIbrbqXRHHAvIteFmlDvSL5/E4BDQH5QKHWa8I21JYnpxq9PZ5npYHPk/TfwCbibGjRP28g
mkdIlvLZ4lBKFpdIovL8aywLV1u13vAqMj2xHiG7ubyuT2DVen8OidnGUPP45K1tFKAymv64r6fL
JMogWHhabiAqzakPJPMrPE7JVVhxWqVFJQeKfDAEGhsFtg8r/BmRd6/BeRf5vDL+wq0c6ehjVMqk
kg8uYqgTWMYpYAUksyeTQZOxfg6GP/3y82Xg8ixyiv+iAeMztGFM+dsou/MnJFOmgPRZ0bPQ7qVP
pYk6Cwj5KayYdREGnakeuaZHQz9C8Ct9qhK9/Ei/e6gG2+u3eIrxf30b0OmgHNvoyZr35VXMMIma
Hf5KvNahUpdlGgKTv9UiK4uivhHJAbCYzAhdgwkVMG76d5kafXlJD3BNEo+VJ/4KCIuLdI+dVMae
FcUNDoPqGrGp/0CT0x9cUqoHTbQy+0Qadl0oivPKPgFSLCXVLW0xYvc0U36OBbXcIzKfcmGJjjyM
PRXTixfVsgYDZfpvKugXZCaRi79jZuFuX/DgRGgMuhBr3YEuJQEW7rr08XyhpdYFRWZYjccKSYg+
xE1VLqkurRrfc7D+aV++VGD01o4cSopTGHhbEUZDbnmryk1XvuzF4w8lewMcMMOYzYhtSTCYchE3
Tam6udjEfFjg+5Fon/41ztCPaIqqWRFsKqqmC6OFR5/VPZcYZA9ySDBuRMR+mAPicDCNSNCJMRqw
GHAEsrMxNiaVmSDtbXrkVemy6brVs3a/VzNqj2d3OyW8Q+K+eJrgLtlV1JiV0lmLDCxFCZbDndxy
3Fn95JY9ILzaK9IQYRc1RPlTyCm9i6GhBcJLmDhRN9Oorw4fIUWKcmBZiCxUB0OdlMRcSZVCsiIy
b/jYlOoK6P+GKocTQls4LbClUG+lDVArimZ1JUeWkZowq0/VLyNzH+KtwZGuqTV+LdaHcJKF07iE
3t9iUM+vFKoZwPjqOxLGjpUYQGSb/bIEB2kbB5TC7uokA6qjViVTdh0INJCVXUZj8M6/h4oKE+/h
NDGGh6axQfSmlI1CRtCm90+NPRJwLF5DkrHBhPPyQ//1LK/5fUx7kdWE3SzPNhuqNpuV1sp7vEkM
pB4P+pDinSPu0qUA0FY3Raz+90OE2C/Gc4gFEKWjX6uHw1CjtQbH0ts+ml894NNRceziZ2xBw/bt
QIHp9YNFLEubY8wRN9BubaCtMgUSebNsI/1XZPW9Oy3vzVNf3Y5uguszbCjbr4AQjotYxe0DFjYk
RLSZ1dqMUl2wIm+Dlle9q8JswONnBiFp5OluWwwspqIvTwGJQLPa+Po+lTWp5Q+najQdZkTWd1uE
UQHWlYGtlRzT1LYJXE/Awx4EXGBiN6JNVhCskc8D3vaKuN6vhBsBhQ1xGymmZN6V72CFBuLC8CMF
ShOo3yoG6f+t1H51Zq6qrwqaSsf3p/DX/0wxHn7t8dwO6CRF6gCB4vw0feam5XbKA2/7KLKFmA4h
QoPeQMLUfllu7yywdh/Ypk3FyZsSoJPkE+DJXomOj2XCpXRrUV0uDQweUIUOtWTCEVr3L2WFhjYW
ELmIUt7feuL/5dVRwouGOv40PMXwY6vOrqmJ8fsD17P5/CXRD/xbJ60jPZnLSQm+W5HZeNLS9oWd
O1KXV4fhZ5cnS7z39IHJFpWJJjmVLtL+s0EY8D1ynpr91dOy8MMT10vxOX1H6YY47UxHrtfLqaT0
VluiD4rYq/ZRx5l+6N84yfzjAp65Ug9LzTRKgO++YZp7LubirXLeNqwvekoQxxLKO3mKfgh6JVmy
thOZjD8bsz3Mu+EZblZfiu4wLt7R3UrFtmBRL7fJdXOg/gkNihwl4nEvi3g9VgxIWXBe+bmtxbdN
5AWtNSKjS984zs1S9ggr6nztXUPVUCan8vISk0lkl40sURuOxVryXSuhN+xMjzOoSJ/E2S0IIVNI
f2m7E4hUTfBswCYm40caL0o4VwPZ0uJ7CeNqVaaOSMLVbYENpscKILpWq1sLoggrBVDuer0WZO50
ZJuct6A6+7XJyGMB42l0RQEnKZE14Rgn3stgJ9Wk0e9dTPGItYvuZmvFxBBtAYEOqPAU1wxQD9sU
c+fS17OiAVDuV6ECpEp1tncn1GlrCP6XyhN9OXfqLdmQ9E4StTdnYCeCRkJwgi6C8cPOaWHvUNtZ
DQ92s1SpzCvExpGGLCalRLq1SGS27YlkYmanbRVFw05pG18l9bOIVHVdvih9oLyuVpFc48y9BIof
l+iocCZqucqVkKTgg9yzH+A4uGbq4XcsWzG4hiEcG8MtVkmkCmPFv8hB4AINoEC8k55Ig627Oh1x
G9qFt8zw/jrtgGmOqhRsJmhzb/sKj09znBF6KM45EBODgXfrUP3pJScpWUBPDYuTA2c4tlg6RnWs
fP7ddZzJ+YqmPfu0Xr1eNBE6NEji6aVhaJ4enFKDIuuzg0YLejc2LhQjdUArClMXLfAmhy99GEDt
nlOhH/pIgkknKPShtf25ZSufgugdt/r8w2qc269x2gbq2QHhjI3hc42/AJS6/AIURsAWvgV7AiKR
zYHFGjyLRdcJU2XMikBRk9apr2Eieciem6aZI+1j2dx6XUPuhTVInIaMyhhPXlL6c597B47IAJnN
U67OHy0vhixaXVe4fVvy3AQ8n1LErL5cFg5wjGzsOsCag+FPrz2rtNRedDJGpvVgNHGutJCGd7bd
QFpHtZ5uqoFANrnVdcbu11T294cLKj1q1U9+P6lRAW3NxV707K+T3HYIsSrFn9bwARQxd9GKrv2r
X+30CA8Mi15SQITLc46ON+sVOgfjekcpE5OE0TmF+pf1U41ToZPw6yx1X62N96caTO3MlOSeqUVz
UyM/8r2IGC+PNxdMErYNbvgh6U8qj5dI5uN9XK+mVdM7QG6GUicnGx1ciQcfDjWjkqd7jKOqCXO3
jpi4+zM7+fa6R4KuESFURJ9hhQP9b9xDY7c0OQI6Ass/U9SKleOsbqgEs03jAC/8cP2PIeCi4JSI
63YDtqhkeJcJBxu4iW0MhS5FuujItL0PeZgyHIFkYpSDQseeJDx9sk6d0MGrHhIXJK/ijlIrFDqq
UqhMhRFeFJeZfu57Jb0vVIHNdz80ce66GCAhpyOMl9fTSzrgsHp7SY1k15yf4qFCqDNrOmhG/Tmc
BTuK8Ky6X+4a20q32zhjzZ9YAFe0yaiFKCgHNUJ6vWQsEX4nB6BgUCQAxCmKiXHxSBm3vcjEbMRk
yB/H812GORJUiZyqzeb+rBIB6HAZlVj48GtS6J4qpYwdaUzp7dAitxJtLZPGouikBrkdBm5dXD9/
66ngMK+uVetaOJ9CWyQW+6QxaqLNft7XDGzOMnRkZlevNdF0tIrEbU7Y0qJl7s+4X6Bn88EtzJyj
rH4Cm2lwP31aO86WkQ+uGZGooaZiVBgSZB4jhljAEtaKO+m5TDG593FfW2X8qgtRWwuw0FAH3SFh
SsGH/ji44S9A5a+AKwwZOJ9OULLD2zheLo6KM1uVTHYA/FZ9etJosfhMoA+zbgJaNgfokjKVqzBl
Nm9dhJswDrbZfidfl9R69FQutKwdKuoy3ve0QD5yWW8ZJyxeOiZZk8VXa4SAGfZlcrAv6NBtilic
g2Qh6oHwHHmVPFcnO5MEvrvSFuGGNI7jQWqyLo0byWRmZEDEM3F2BeSzVSUuZUSJOCTl8dcGrj/7
7bEiHNWqyvcqgyB6MtC92vg8MnUf7xqkpkj5M1ovyUaFlazulqw7+L0R6T6EjAAudaj/Psvl2eEa
TmoqzTTFLRiDlyFsUh/CVrVNx1bI5MPnPe6eMjIrk7i2E6G21d446OTXvqxxb2iCffkRS7n36i36
xDpAZ+emTBHm7zH8dD56K0BEGChR2a6P12l0Mx3HZzIHRBbH4mBEJ3+AoDSxAVGgsi0pV4Oe+0iG
CZesoi8OHCx781JYeVlFJb4iMnwbkuqv7Ph7RMcM/XJvqjyF/W8vadzaohWVQZf/gUZWeMlWhIq0
X1PRA5wtFXBB3q7XEe8WIADqep6XV+GPAAPHToKPXLYjFm+yHPV2IWwaYk4ljRHBuhno+J7m22px
30+dFjs4ZhWlhhH+Ezbk3LXl2O2k7BmQ3tLbu7425+0f7OrqCjOkOwmD9714yLtuWHmXQZc0HqJW
3/KrxNbq7h3E0r9mLXQCR5YRsMP8IdE3mb89D2bx1ahFrPXaTVjM9WnSsx76gAgM30B6HlAmsDyX
nXltHjcw4huHPSaXOVJ3jWDrw2IBhlXaMIqKUWViiZOu3A/lK9BKmVGJC8khAH7jGqy9HKDdgWVO
qz4Wfd7m0Xnjw/jHuHSrlYi/8McXxPXcMNgxtogf3b5ugsjrmcXE/M2eKQ5q9ZSxAyiGP+XkJ5Kg
GG1lBNCLEf4+ff40eK9d+cXYbQx3KwXq6e9XBaLwWZwv23FtVUOvrP5Ftzb7hRdjo/11vykoFd42
5yIO9DY5Xk8UDReDZZ3+/5FRhmv9kVWD1fLVmMQfWmJF2Hk6v6RnIoA03kKZPXYVvfIL/yRCGTcJ
8CcL/DB/DBkOPjDpRbd3gF54zxL6KcmbQBhlsoMk9SPzdHT3NHIkUp7kBocSJVyQySsXlDKylsks
JwF2nYxNASQaiv5iWuibG8j36c96LUBxOMdjhBZoJIY0T/quvF0fJg1GZOmr+EaLFxWqlKFPmyFA
gP+wT5ZZtdgcFn9Gm9OYfbMEAquOFa1FPVmwn2tAYBMr1uy/MdOzYa1ibxWdCZZy/aNJ63s9VVdn
z+BVinXnlEwKTa3IRmIYWHCMQCTR+LkKmWS3pVbO/GHLnedD1kJzHo1y9XrGzDatIxbxVfYe4+J1
W+bJrwdxVTZG+uglQ7X9d4lCpd311NF0ZySvx/KNcqb/z4HdUGFcBy1dpqINQxyCbn/xw9X6b9nf
/sRnXdAnnOXVU30OJBv9hNMzTyvboSe4hI96uvnA8anTWK6Z4PPHuxa/civtc6xGMl0DHm3MX0KM
ujdGwuhVxM6XrgwwMgIGT9xQgcGvXjwBN67CF9FSm8qKhZ55mj9dVb2YaxpwhoA530sQ+Hy+aqQZ
ShyS9mcGD2put7ceiQomNgM9U6TbdOuEe5PQu6WQJX0KpoLz3z61QPCJQ4tLiXY0lKdbe3CM3nGZ
3m+zBTjjVmrYNOZZdDXGd0uHgf2x6f7pxP5Ps3LA/BBwL9hAjmWG2Wmf4Odb3tJWDpK7vUFx6Kiz
xignGCxZpCX0uMrnZp53RWJ4djFxIiPIYUntvYpsLPZeth+SVtIxqw4ByQYmj8RWGBKzX+iHcHbN
twYHQA1VaEhWk1BFyD9rvZ86DVH5gT+TZKkGshrI5Z/ioo4In2Yt8tPjV0VXVdJ1ZEGziQ4hASt8
cnXuno0EIN7M9VOTWI5OHw98D1KlqqTRGo9h50hpLPglhw8iW7MgF3cyJsMbHp2jZU7a+KyF3di2
0KRqWj6uEOBwOXKYaDoN56svQ7LNcZSpp2YYb2Pc7q6V/o6RkPttNN11RHX7jXRM9Kj1K4tJBMmM
ubRcqkDMSFOfHiWVlP8BpN7APSaXRieLZRibLA3w/rbK6EA/4Ma72t3uHjj6C4jyYUAakNXvtMi8
D0UzGFDgzukPLMmJ0FnC75013XPO9/mXnsqwGujQ3fmTvNq+AJPruJ7hzx1XKPBPmrEqQWQJbODF
xyjLjVPFqEbXtEvoHmXWKwvviAWfeGszrfyHtqFHSIQQJ6yqCisZlj78hVERpyCJ/2NkIjeBUFVk
Kcaf573XwSgOqm2k1LKLPtigoz9Vpdo/BO0Am2h8GJOFLGDwJCVLI5CTA7yXqV/7HHX2itYiSjTx
U/x4+AKaXDkbe8jxtlCuiFnLjvKgY2Du/ssQRlix17ZH1YXemoXNe1/s2JD8LcSK/BFv0ZQdmtiq
fvMe/Zc05TdybZaFq9T5wRC2XWVaeeS3r9zCvco7ySG3nOgedsZTKdjkflQ5vVnsBsvMDlp0AFRz
iFykxjblOKcW0gBPRSFSefpw40ezgxcs2G7+030z6DQGCkVtPF575LUpOqsbCMJ7BaaKE3fTcziR
IpO+hmQKMCgzc8W/nVigOVBVm4y+e3bk04dZ5qhysDI8VCnnOnWIgSNYoU87DFU0/P5297fENNaP
RLkhl/XY/LPRyLT73ySdpcT33uU8IkfpW7FkL/GyolPwzfPaHcPq7ouWKBVgmMY74gT9oINZlxWW
BfgGvm6H5riZGUsiABq8ZLFwx2w7OkggH+8kzSIHVr00oRDN/ynSpnpZOXZkf7tRMw5FIQo8mGw/
Dl9G5icBLBEMz5xHFp3xQ80tNKc+2axueyVv+yaPUlPlAcIYPvP6GXEKfrgiqvlzqAeRNOhlkT/8
Kg6bOAXKU6Z0ADkyzkxJsK59XToLBD/Sd8saenCD9ocvm2D3jHbE/Alb3RZhD1fERIzALgkFyf4P
U5RFvY6MmbSqeU+CKvFsHJU6altpsX49qbmo4MeOkqC+OIPU0OIs2MkHzDwwwG1Y2JMyJjDYsT+2
pKnw9LTXpJHfIwLqy9K3av03ZtmOSi9NtZkZFUxaW6rFuxSZX8Fy3TsyDMoHXHckgtIh0oRPPLLc
4lQvZw1foHZXg6FjdBb7PVuk7iS6TTFfkGluP4sGxtdo6k3EjVP+VElXwlMiSRbHsdTPzabfx+jX
/DgX3PYMdsaAOvFZ3k9wXp0CFajppzL+X9dLhCjvgxxNgciZm2i2hpXlrZbGPSX7U40kTb3v8B6O
chyPRYJjJ1wgSmadCWgWB+nHWUinjOZouoHTzj9bbzn9NsN6Ziwj48ZTO3qbDJyWw98R1vjhSq1D
74cBH/oW6inhNP5LajACJG0oN9Nx0UWvr6wcW9HYMGmBH4OdMZGSrNk1hYGO1uN3DaY8f/JXTrys
7cNCY94HR81Ii0g1qOrOGZdqIfNDtCACxdU6CsYmgFY64NSjJimOjhtFSFXBS41EjheUENoEmf27
1tJBHFssrQSJcsGpyytNGwUiq6q0q4Ofe9QSlESZxjZ/XDtSdNgRmhD7tMO1JrCTlX3OcKODAXd5
PJZqRWvn4NsVKNDcNCltOBDKTlQksHcFU0OWEEgHvshmeUD8YLhLMON9LIDa6b7w6Dugq2IlOUH3
MyMwYx+QqDJlIloTINR3GrT2iQg/Ks7/pZNcmkj2c7LhspytbPo/iVF4U4xEQ2GtQi7E8VtMQylq
M2mBM8whIdw3J8nxgyzJoS4Qfj5Eb264O8UUMzvpG8QwPhAQt5tR7WBx2iH/BmO9OCbv9xW3ghZi
16OJzyYPvKIQrUO5oklpA8lyYlwOL5ZI/Igp7e7nZneDCpyaPFVieRieBIe/pYc3ggaDNZUz2mAD
1jrm5iIOOELo+hCLh+cZRwb9gDsxTSF00+XXVEaCcGoLT6pIA3f2OjlLwd2srdSDnptO3sdRkoms
8BKYrp040eqG2R5ywikpJFVaCB+nIiwwMc94izHck1etV8yNQ2vWdjT53VjqteZpl7wNmIcNENd3
22lF1tayD0e3MTo5le3RAGIOKRMC8xd7YvoH3ibB8idKrt/3aKMpLq59Tyd07R1dfHOx+6x/Lrfx
1pocAmrZhkamKrbq1T2IyYQgzLBmyDOt6Fm/IJEY6QWCBbw2bvm25lBVnKNlo8gN3E00eWmeTz3o
XK0asaSU3T7FWoOdJlpUw6Aodh1Twvae1J0lKdQjLioexC5wOsRTQPAzSbp+IFPJdXehEmkV9hYU
bEzvtpd1p6RspxM4TcqwX6AcekqHRWGckEzlQGyGrjmQf2lp6YWyIacbDfPzBGU19zDrJucD2Hs4
hdEXve+LElvufIO66n26uhljgBy0Lr9gs1rXbmi4peWjcYg7tEaJLHRhoApYzYVxeFUQLyHUqw0G
x8Sm6A40v+CuuOat3g8xyeURmJt0sg9AhdtqneMifyvPU5VEqQAv73XNPK/jB+p+qNBNWGdalPLK
lSGxZuk+m5RUn4EQ5loSCZSAI3LcrmhD87ph4m2w2ZvHmY8+RS5h5HUgrTpeWl/WtM/2U/TUTvCY
UWtToIiLTO1ZJts008xCRO1UqVSd++1zZ/N+UNdOJrh0p4B+LzAQpsidqyNVvnvIAv8Ef7UyaFj4
39wkcj8I4XY0Md7Fu4iP9hMYwqfCP5Wj5Nhj8CYBVjLyEX8JZPesmngvLpd2I0TiSluy5OjYMWri
gz6RmlSCUhkSbkzaCtdPeAdfC0w9cJBquZiB+htQglIkOMXXTIGTyVb5oXkdR4rbSlVpcnDG5mqH
aX9U3HhwyrKMFVwXaMw5EtpgHue82b6IT8lrgm3qkosDIUC55pBvMS+j8nf//HBEKtgQFJHQoIhZ
3bXy3kWjkHuiedBgiuLogPQwUDEiIqMVihPINzcCEZjLJyQJ6rsJECb431tqORrQ7NwZdg0KsiPB
w9trD5WPqOrzn9wjrNBonUZwN37lRBrk2Livdlv59x8r7aismH0a+8bgr+HKzSGlZNou+zZh41g9
9bLDbDdtH6ubP7gKQsU5WQnz5bXOoS2m0KmjoAtWTs403E4FvH+dOleIdqavpoVzSu4ancIp3pa0
iFUdyJ3dCkTfdCruVoowN6oTSR2Z3zJmcQertzrd0S8owG4bf/9pIS44A50icXwYXik6qNLIpoIT
o4vWT8pcd1ynlvy4z+XQopsBCFyAWV2F/7FLEf30QKMVGKxS38OuLG+1ypHvnj+lE0BKaAJXjfg9
nkU9rIxUG06MVx0ONL/hVmROWKOy56y/l6Y497bENpXUweaGgBhbPzIoxafFhpDgYVmhWNFwhu8a
pSEpn8wDvKIBImcRf/IvkkOh8q8onoz50r69PN0InjE98O3oK64gNPQd7vc5TSokPJYNsq5j4LE+
/zGUGq1QXtNCgIW2pX8K8ARQXJVdPmUmriFGb/caEpW/hmmpEV7syxy579MiqObWlSQuqtJD/ntw
VQZcN+3ozYJ3lcJavChINDI9xjGesZG33PETCa8fjMuqXTduXac0wTuxljE1//QavWAjmrFhvWg1
P8oZENLPGsE4O4wPcHaeYlSNXqchXjy4NmKRmQfaFLVHx6Lc4Nw/SMEH+LhLpxBSeTUmoM+7zWdy
kzhdihHcSjtaeDpeWIeVhi7l8UaiOPXgeKzKzGacrVxRk+LN2PPHjbmOPEjltjqQQtmr1/Be/zF1
3ONZ+ymBVUHF9g7gPX9wRdAX2pas2P58MqI3dUhxMHmt14KyPosGZDjtvOcZGDFKDoLqHG3QcnKe
nqshPr5BEiftz+iYPcRZOCjqbvQOuj6JyaECxGnfbHaZ1lt2g3OXOS6xZIZXrdF4AbeEJp8oXMdt
xwufR6GM25J4LXg1DRpMvmPec2cORjW5+LLg0mS98+HeehY37MNEUeCkHxKoiQ6f9CkFExgI7sss
xAIwcFb8RqytmTJfhaDgJzHXuMWLtKjsQJbI0AbLeCGziCP3bS0gXMwRKMpRmv2SWC/xlewInzFg
o4Pl2Q/RMbpbtQJ6A5BndANyMBBqDThGloNYLQRCq9kY6CkH7U0rOH+XuhNTpOXxVSlWEYrhEgno
AcsgmefueYO76nKoW5ADKV0jEfWvN0RNq7c8aTJFEAJbwA4E5/SQOV+XPLoPVEXspRhCgqQ/+wjL
Ui9LDy80odglGKkYvP7zQJWURsdSuDgy9k75NWU48r1lXNxkUkoj3kYrmWaN8KTjUEYNjSpzIqzw
i/zm/W/UKxU60XM9ijrsGMblPq1I3qftO4I8tQ9npp38wH2QZbtVGcKxEot4sBtxBV88PpbvcM/C
RRYRDkpxlQdTl+cR/stbmKr67EXXGqx5qatd1vuOJEG3D9wYBnbeFhBIsiM1aX2U7G/bfusc5hhX
9t9LB2zk1+A1AZV5OeXo8vjY3y1Aa5edumW5hOkZd91GOvCFPp8HPuYZmN7YQaRA8yy+WEk1/azZ
RxC5A6aEADXitvu6erBGvGHhx72Q95774AGGV9qGOqVhedI3X4zLKUmMnr3qfvHarl+8A+0xaHV6
mqoq+XUIm7Umwo1elzOvZaBqilGWZU+MJ7lEmgnwJvzMckF48+flcwXGNa7FgdlXcB4HN2/ljoa+
50Q/VVPM28dgOYs1QahGU+snizFg2L6BKIBrTB7p4sru+9tUQ35ga/TYMxFrHX046pL468Q8NDaS
hJBI/iG5yxSy8kR+sdaGVPA3vGjfCpGfrUekkSyKvG58Vn/yavSLjRSytw/MK7I5ek2/2o6+hsXF
/SGgwub73aGfQhd7srb3PeEw+aBsjR4JK/y7dxwSrLzTOstgIvhAqLCmgvYuK1CGHbItQWkeYEyl
orAY2foGIXZXCCAAB3Rm1TtblUTqY28w9dTY1+a1dDHbpw+gmkjlG0fIhxnhtorbOcg0r2AGOJhR
s5tvyh9+m/3XEksBJa573CVznksUmkViiwD8qU9d/A7l1cYGm55JlvLesDCMFPQBfrifnmS7uWH5
bKYFfVxKwD6TSc0EQILjgoQJLRB35GStW4ZNpvlJ+LJlT+qsAOK8cx3gILPbO+6HzD8kx6J2WYUe
AHK/qPz7F4vIkNLUhWQYwKo9qFamPVWPT2v9uK2BJxm4/oMLC907nhm4L8fZ0WNqr/ouQ9ndRLvx
nwmJOpafCzw6ejb6xF4/qycWNC/duzCvZNvUjBwR8/1FYBruxVzwDaQDQBzshqtiIG3nrIL8fpnq
nwqVOHgADCqWrh6pCzfLatToLQUNAXW7KS69Ktx1eZ9RapKQc6UefLsSVsm5ni40eIxfZ8u4CiDn
C8GvLWZMKGSH8VXokP48M25BOn9cLVTvh/j2cGGrF91kat8IrvIBW/i+iRjqy/4tleUm3YWt+maY
5GjGdy5CcqJrNc8nJZU5j0SGjjrMOjD8dyfF9LHFYyN6doEUxOCvECcJWFLmXQXJUWPwkbyuM4X5
8p9XCnEsYc1uFAB3uV25IN1DcIg1dgYK1vs9oL8mhmRhfSOTYNoViVSKZ0Xbl9oJ1THsAUWFWOdD
TAhrGgedI+matFZ6IzHHTKb0/5uLv+2Mgk+3pLmvcq2gSJXPIj2y6uH0KNFSe8SW1Z/6YyRDvKPN
TAxlMM2iOS/ziPsrYBgmcX0+yr7RllgkFjhiDMIKYnJ/zSa0eIILPrRPuNr3hcZLzAqvw878F2ye
7wQLrHOjaviizx4eMsMInf9MnQPgS0yzmGcffcC4F7sR6D9Iu27SKAUAx/pxXbRvpMKaEWXnya6z
Vm/R5IlkvNQgYn3KMwd0/qQIatwqCCayaIk3o4gpWZ4wjRu4/nfTzhgLCJyYiVjXNaTIjn6YmahC
x1iuV09ydjfsNBFsEU7lNazwPEtHqOO6DgHpi17NaHQU4HQHNT+/rHjvBUS7TU+tlN4LuyvGWrsS
VJEWzscimtYqdRcSteBElzgjWpBPhZoLgRfHEsDEYRT5g/cGo/ukY5835c6s5DELM9LwmL09FzZU
mtgSF6iIyUutkE/iC7fmzmWz3pvriZU3HhkED7NVOUAfJO60FLVGKbsU5UzCPT3Qsx95g215zf2/
7OWUH3vsdsFxe7sH7hSIlvhUdMIw0Kfre+y9Qe5bSFhLu/Kto3LnkqD7i2PfGWtwLicQzdZG0O2w
yZ/qQCpOtr8Zz4q+DsbG9DUOfPQ6L+n6gOQFvv5kt5+S6eNw2pInpF3YrPOifLBaUxgEORBG7Wjw
zzsXZLUEC2Ebg7GMY/09B6qBvxlhGWUWZMrd4AJzYnDTHzXUOtGeFQrL4GT1fOuk7uqE78EoWFmJ
byRbtjyv3Z3UyYZ4gI9YnqRtK1vhD3EnXeZWUeg+UbG0lbAQwA2lNPpZMK4tU6z8ZMcQ+QDHFmF2
fMBmncWJdUhUD8w2+cc/2NQvhE4A3FriheDyHV25juZbiIOGHq6l/sYAvpX/FeNVetIjWKCqPU+1
h61yopWvt/eyGSgi4wMLbwDkAcBko4CTFjOLlej3inHwxJ7aBhII99ys/LwRamV2Rqb/e0QhaQOR
TrdfPph+LckFSpUH+Cr3k8U559ELNBnG9RQN21jfZJifueVcDwZpjm6jVfT/Npx/jBBuvREw+JCE
+sc6+v6b8ChozJwXjDXylOS60WrGkc2BeQy3cwhTYqV8YNcNvnsBXiHEmdWWxK7WhdHJPHAtC7KZ
oM79afpxhUopA1tMmEj6VK6esJ1lxCurNSNbmtnIyslnStnJajCvOBNT6QopQZ82fvQ+Pi2SB4dn
fr67Zvy8aEkzYgfUUkeMjn3tHucnjjZuqlrfqW4RtfaOWSLnF73ex+Evj1aN8uOyn+Z33vliUMYG
I33LGWwXUSolHlj1jGBJDnIqZSHy21dPh75BRWttqwhfOa9Psuvl4iwRY7QH9gPWz4W5Dcd79lLz
hqfCIYEJPnQ2j2SLN+lIhBuBS6PPssr/susZkGM8o5bWZLTeO4x1kKcEf6oilgKPFoM4KD95IAPk
gi5ADhZxIdktzOQb/xVqoHrnkQGOyQGRUZDMV6WmTR/mAxVNoQK/MJ2y+bxOX8grtmC0CBVxez86
0QW5vCli0l0lRZEEBunGV10IHAhrXbiYKIihd8chjk6IWi2ELpgIPcuPjvvFFr0HpSccTb004+3k
pf+yYOBUQzxeQ6zmRu3T+sPCZzJ88TZdKGqJ7mpzpmvsFwRQOK7IUYKWoE1Gt0P9QJWtnZwh+7p7
1mNaUKw+vcLLdnKqktcfOLdbOUow96Gx91K0JGZQs6/lzQi7Qt1iHGUFEPRdUb+UA4KFHecwTh1Z
jwEXjuFtpwNgGVvcI/uzWy0GkrBMMz+llLn7dWf30ykh1y6NYj48gEvaCnIQxTqZKiwCIC8cZbq4
zEhZ6NQP1mR0akWtHXtGeNf4g6sTqx1035mLLNkIJOzMwH/I57u8xZnLLtocKgPfi+vO7r65tMJR
tn6aOnBJ+hiKlFNb4sKofV48aakGovjRO1hO+fvvtFogY9DZUj21z5Ya/8Izf4MPy7vwL3Az30fL
RiJfKuGcxicbLKzUKatteLt3HDA49m4TZn6J2BiNWUzx4C7qGOl0IFz8ushk/56dLo9+20Usa+UV
bJ8mTKnq+J2QdgwfsC6PCIixZ2TWPqW7Akx76VClXZCJySrrRhue8K8IIIT7ljIm7E8buMqkQBCl
Gcis5MRaIK7CHzCylTj/+3eFs4Og1FTi3Zs+8f4FsTOVVRQ5r1h9cqxe+ziZkHlh3zDOqeWs84+w
jHs0SWzzcwzgnMtN5cc80P1Fj2XIixEp/YWCV2qoI09IfiL0fVPg7GpVe9VBgNqdTYAoNE0fLNaE
gWXdiIIELDdLFJdi+k5JLS3UiX6Q0lSbWutKJJpCTDLMk8TRhATTE0cmxp9B9q8kkIs1OeVRYgjD
4OjEH8PtcdFK3EFuZchkleZ/PrcDnT2RzhfiXak/zHoPsh6ZujYC9R7FiVb6eo03kOg6pSEg3XsR
rJgq79IEs234U7ypbBCP4ymq+cNdQNtN89G/4SSly5im13GljtK1ZDb0K25KSNpK8RNU/rrwwv6s
aQXN4bBZ3LKfSu9NkMHEDNQO1jGb49U3fkbNkelMDuTpFOz+CZiLuaXcFras27BbhWEG1zFtPkiK
JyBiFz7bDH9dhigzilJIcf0g84lCruK3XAlWPvABqe6RBWPUI2O+wejcqRGUPwxpkFRCSK7/RsbQ
/eq7VacehyIxPSPb4VzVUEnjo1BHTXqduGasfRthgS2MlUhoVTZe7iIyJFm92yn+L6SHGn1Wcyj0
XBculOHO5Fymw6iH7U19HliFxZODjeprSA4u9i4Kk9kGRr1pydSee2oLSlSPGK0NIGNJbHyWO2Wq
4nh9BBpaKTyZKdil8yKTxp7oLuu2Rq48D6ZU8cYDXwHWAMIyRIRoXL1f10tOcp0eCOFcRQOwYkb1
9EBw6rhySB1hF+uGeuKhhquC++BvI6grKHlOdwGJ0CzRKqJwkEc8iTUfgIxGrUzyR2lKu8rk+coT
g80KDNDLPzTWpkY/9WY80WWwSamKRPfKSJrdSmmUZ+4MkAUGsUD5Eb6UIKnH5e+UTQO9Hs277cmy
smWprHtOrV+qsOyv6oK4lERAoEY2T4ui3y+ZXWwlBs3cSvNmipZKEG4YVzevsCOkNlojYElb1T9o
G55uEh/1pnA2ndFzO3ymz5XX7BCwRwEjRSoXMVkXSO9BZ8uWQ1wZinueOVFppePhHcdtrE3jQo+B
8wFi3yWaVdAgBP68QWseSlA8Bt/rLuzM5CEW4om1twnIWX2tE4hCBsi4e764xBCyx8hEZ2DvyRbA
3p5wkgUDFSGg/SgcBnjNvVKYal+XqzWZRMdYE6MExFp/NeWfWLECb2gwo1rVCgYkxlOrCDHpbZA1
j0ypjtJRwy0xATUIQjHvKAKAsFWlAWWw4Aw4OWWY/ubX3qqo9Gens1jUjc0f2Dhyog5R6RiJFnCW
f2h8aSVRX8ZoPEmF++hXpVV8jcI3DPgwPZmKTONUYz8kvntDX6OUpg3ClynaN5WJLVRpTMsUo0rC
nhX+PcfUwA4zM+DXh8Ybde4kkS4fqhJRX3U21P6c0c8KfeN4V6iqxwhmvVL2/qw7uFzo+VHi3qw9
RqP3mxWa85zLQ+yjm2gaFhrki9jXt0aQdbjwemBiN8togq6Q47gxT4S2/+ENERDy4TI14ZfQovh1
4KVKnHg9ZcuNNKJAK554el3kNjKQX+2msLN/dJUINa6G2Qwl2cRQ42eC5NyiR0vAkRA4hU7g4nr4
TG4tm0E8w8y8LQ3clDJ8vuWmU/Na5i+N/fvJSW/ZNiLASjcEJo+UnCNahDMeVvBCTiDbvsH63+lb
iah+kO5IXAuPNM8+5UA3CavkcyWZUliZvNnnhD/F/+uynQxQY+dLqlMXeyA4k8Ex8A6VZP1x99gB
sVsK3HlfuJ26TYbcY7x9pedBG8W+BqSPBPMU45rrvLublZI1xw+GsscmHhhSN3P9VdsKayTK7bBq
TOEh4odtWt0bz1UT9zIbZIgBqdLnt4qFk0/Yas91nxcNCAptOudG0jAnFiD4jFRRRoX5dFD8eO24
ptzaCylQmXkl+VyA0Pk9J99CzslDJn9GeB9VxODTul/8/YmUULliY3T0DaM0/1h0L59BiF3mhDAa
Q/LvU2w7Q0/dPcyxRsitIBgDzBvBsGCBT7pfbyJ5BJ+YQ2dDyJ+tkRs/XNLfDs6mbS2n7c5NZrdA
UvSsMCXupvmBTZp/Z+4Z5T3O42Dutsrwix5ygTJmBGXvD1M+C9KWSI2niY1AfL0vLl890oyKUMeX
s8ktrDvD4yd8IITaYBiQAfTqmfCtbgO0Cw7ScoI3sFAikXB8Ez95FPmjit13Z2wS0EDPQ7VfAJXy
WIIsbi4TiB4iEStqMCFjOC3dyxm9+QkGEdejbOxWcPQSTOGp8wiJgwFDeH9EQU+lZ62c90syLAkY
ljS9Y7pxuQhixDEDYVPuVeY+SwmVBm+L8mbnwnYH8Vis+aeLBf5Zm1A9xOjz/BiV69OY71Aiesgn
2vlOoYEswTbWQvaY14w4a9GmuILFehxti1dPcyViRixzK0ovdFX7sP14VAmWr1zt6mc2aLrI5++p
e2/gB5bWbL3gPLAohZTNZcaOWXPtLB8wd9oF1ub9R+YfHk5hBvaAPzTTNkHYJb0YKT2eOn+ieUub
olQvQy1wzEDhWZ1hseO6PoSmqPtBsh0Ce9bS8AIc0dgINFc6RO44TJQeMtK30qgE1BP3zwMPlHW7
lQf87Uqy09G9XkYXrXtKeIuIyc4MBHHm71TrijpLtYgGErYKwWaa39V9nq0sB7lXAVHerjqKZXQ5
p8IC2TVz7hwc1Y3sg0d9dDGNjZNcxwDHHYmFfpUX9vFEpEsYmbqzNtCe1NWb1cdLOM8BHsE1NS/d
0v0Rf1dOUkm3yZ9SWfna4iNP34A6bb5rj1eURtwg9dr9pmlKCyslFY7LZ6fIY9n52mtCTbG67w07
P7cIbE2lIskdMwG8etlsazw6yARMfNjBVXrht1EeN+HNlPzyvzGZV06yHgDXRPniDWYkoVL0W42R
Hp765Uce64VXQMrNEP+5bfmLtsHN7d9jdqTbRV+/01CkAcVdeKw+oED3qSsq7SCFfS63k3hRkoHt
8kop1/eRIULxeZkQPZmM2n+fHrUtCLoqlcb6+xmR6txfKSto6RqJpUzOGM0u8VOIooVBFcRxmMmL
VUn+q1WeE11lbQ/e8ZRZibi77CCtjf15G/WOLzHSmyDXNZX8+3Uz7J8ZKbBhQCX8gVRxaX7BVEc9
mYjblnTr5TB+5B56ZpEzfKnmOzQslgmpLN4XIgazrZkK1WsS2mU337hqts1ZzghOPs5nuFxBkgGw
z6dzb1cGuAokZmtEd+oF2HsVa+CwDhc1slilq3bUJYPvUDso2mvKqWK8K8si41EbGlVvs+AJgtT3
rfbYKKcw0uy/E0qcv2/rOokd8M1E8XbX4ntjiTCN3ub8anFzrJCBLi/Qz1f+ULoWq5RaAHvbNadz
91ptuPXfNVJss/DEfRgz05abW59w2jd/92h9aBBYCPIGaeFCoAP4Dof4agtY8S8KT1Spce6JaI6I
SFx7A9jIVPq3s3W5z2DzpZRnfuXc/I6SZ9MTEGruuOIrlvde0la03CxauxJ87sLf/nCKwop7VQPD
3bT9aEP6tWuU1ZD7xC7Z7HkE3kSLfjhiwcTH1wXpz+JjrqSgv/+ytWaFie0K0361+M7fMTo3uQuF
hkqdrXMlUnnHGAFvSu4a2kscjHw3zwXPeNiseJkIzpmjBDrgJjEzBl6PG2K/pRwQdcMttgbiJcno
cB96vuFBhBmwb0jCUn7Ju2Nfi5idqAvMonp5QmnEC+ce4aWqe7d2h9RqxR3m7BHXXzUOOYrvZcTd
UrA8g1aqOtcQ2vioaBgLuFXxDR+G5Acr4DSykws7PYLFW5oxeLyDWZTD1+aCZpcq2CTwBkvDMXcj
d+++89gwptbjgpoc3aUCYPKfXqiemjhPdG3y9fToGt27WbV8l12KysK0BmE/ubgi47SabbTtIr/s
bDxZjHOH+rlVzYw0bRXbCsLpwNsqBrahXI1mpCPodIIqtinkwPb0lINf4NfFFujXFJ71TtVIjAYa
FjOEqAwFKyMP+CuBGqiIWuuzTT4OWlvgfk0CA6C25cGxWvBtx4F4RQ5ipEM7lv+XmIDmwCqB4Q+u
xiAuhezWwHnIpXE+bBMw45fYGUAwykf+NtYFYWTgZfvDaDn71gfSeEoFNS6YkRIDyELA5BkvkblU
BANA4qw5TX6QnbvMF+pE++JgnskLBQ/e2+r2jecizR1BEgy04S+GCBGusKJ/L2/NCJVpLRKbo4Fe
DfI7fLMqxZwzfZKyaP7kP9OnklVq5c5h2I91MVp19LNBQF4CjVurzvLeSm2BXVOzdQBOR4uY/BB3
R+mYkehyeJgrbQHXguNMRwI3//k776R4b/BtxCA+XoJzUT0O+/SO05T27ef5IqezIiEX6VpTqWZt
EUwsMdHlUCjzWq1d/5FLD51ZK/KU1QUnkmeZY2NJafHTn/YP3+/Zi40qdM6ShwSpN+zlypAet4tc
EigLZkOg4bHzU3aHek/PT1asmrNMNH1LH2GW1lVa1Kw28ThZHYSfopK8gc87R/bS5urC2QT1bBQx
V+ziJjIqquBocKB9JEdSZlPq9CsKvnLJIzfvXU/o+41YF42XEX95Raxyou0jRH7ezJ39bbz0jR4i
UToLkE3/IUX7+rGAwqlvroimXxaAUs5BQYNyzMq81BkuC1TxIQmCWNG24yViA7Ldt7gqTAOXISUS
KuHANrCfoIsPXYCUiVFDwXdDE7oEXyyKsRjVWFK8csO2+BnQKnknp57hQQRVrZroTn7+C4FsFOho
FZgQNLwB2lr1xqhSH72Yg4+eK16DByVTSu3gp4s/B7NBEej0JXQOCbWpmLSrmTMH7ejumMWO/XrB
/lJE3ig6Hl4Ik3fp8rNZ5K1fjp6OEt2UxOPJf+JbZWYfzm75c4j5u+VQL1CiOAgak+HqC6KT90TW
rPsn3nn1kJO9plgcdzylose12bm6fYe26Ipcb1gziyIcG4JLdzX7DI+bqcV0g5ieRW0usO9XNJxd
tS7hm6kPNOANxM796UkmcvzEWAwqiNQIqs5m9bGylH260JkyeBQTw8L+S85kQd0YTUHEeMIax94p
WhxKqyZwGLDce9QfTu8LnQRxEs+KJFmMQW+XiGlGLcBIZ1dgq3hDh8nie/rfnHEaLLUAT+S8FRA0
p2d9Fn9GyyQLIKr8ZK1gnYVb/KU8jTlLvNqI+fXAp7nANgDBVmXpdxYevY3P9uR7jrmsOsnXAS/t
eoYWRy889HCrkkrvUjq3wc5WdakkEVzOesQ2KIYBn/1VvclXrXgDpNFXUshr79gw5czgnYWuiE55
Apo7kJ2EQohPLijgzUT+g9rEAvtIEiYIjNn6YD9IX5hB3O2jHxyPepFkxvZXpzVykZRCFZVkQKuZ
y4ekiDCNRb4SXgcZ1N17zQt+hMWWWYMk/AMDwNyNenf8vnJlfsmOwK0fyrwqlCqwmzipVqPrzihZ
kpt8XZ55T3ckllsR6Zb81dkzUUClAQAypweatDb2zkjVJyiSAymdcp5YwiGGJ/REZ8d1Jjw0rQxr
1eB+iswgvD40NAFBoIgOLGgH0/FTKo/ckEu1qzxn7o8y99u1Lp4z5TkLJMsXmo9XxoMKTWmKB76h
mGN7OgB1Se3jABKYhwaq6rBdmiskjhv+c8PbwBpasI4kEI2CSHWu3fcxb/3iSYrJpAK3qwTlumun
SQjpgAtffMBL+WmIghSg07D/MsuQeJJV0uSmS3/kSeC2Rh/uFqFuvRSRDoBihklaJOb0b0VJG2Na
77o/uawX+cXvjCNGaQ1zQ2RNvPfkFB1wWdjLEWykUo7DApHvt0vRkRoRgu2n1LRKpHd1HZun3f3a
0dn0GhQncdNApjuPucK3UIam6DcQhYnYQnTET+N1deU0flO9QTCb+QB1Wc19KduuxnZoHvWDqyWK
/Cw2QCZverDO9pwxJrUDeqgzo1sq+i46sexH7WHyEKGAQQDNIG9NDWSIYgy6afaprMII0psS6VJ3
hntd7hSO3v4+6ImSf2btvbo5MXw3VG8waY/tBEvaNtXlTXIGgnWZTTuz5HpKaLQFB3eLPSSpvDs+
U3vOxT3zitTwnVaXh8WE7zRg8dY8ERjjbOnNF5k2JffDOwgAXf9sl2FDqkze+xPqMxNFLeoyiYai
WTFfdwcGZ3hfwAqPvrpYutb9kUNJr1VCLsGHxmZgv5qgoI4iJIssvEv1E7NZsPmMMzTSDySaxXtd
Ax2VRn5k9L/onjnhgv3CGI52BUBsFmjBqS3ylVYHFv+xRb57c0arn9YZHH57SBeQKZ+eDQ47eEtf
nNfJVCXczs2dpCA3VXH9xDsb0Fo1TBiOUR0mhEcVPvkPFj6wC1vYuLsc1m0oAR5PpngR5T7i+Z+N
6zdGPiqcxBgLuc2mMnpB5LRBTlI3pZRq0bZE4XEayodp+rsBrBLDHlEVBClyLHRN/gqwY4GZSpFg
x2NWLtOgPdoI/3vlSoL2Jd1sfWOs8Wbv+lP1Wn3OmEaE0PWrhLRGTy3RaHJgdjBvDbdCLgsOr7o2
SiF8xdb+291OHWsocYLT83jGYraPOLI/vsXL847c79o1mv+JFaqsUL0cQqIdqF7XHqJ9IW9qzWRj
hxDWrbezNaUQSe3aiEfYdScDuCG0H2UWe0n+CIz8iZErxi5tv5b2insrERpj8RQJ40ed1PjOJus6
PATN2CDC3karSWlKkhEuSBH0tr9CAgceRJEMcEr7GZpPbBEj1WqqAL6OYUa9pKTELc7Exwl7G2QI
05etLz9jMAhDt+s0cMitlE9Q6gTqP1lbada/Mpg1/ma8ReOLFrrzrI1e1aU7uDgpaAiGGnWUnSj8
3ek9nIz2v1TkA2cDrlYU59eg5zdKCQ0TCvYETTgXAJtVuS7d2keCqnA5MrAIZk9AIk2WWDg6dDTt
ICjPR838kCfEkSTHhg+vTYWF0Xl9hq+wZe3oRsZ3z5SRNyTNMCRuiD/qKtQmLCsaf7KH4UTWnC9w
J63uDP/FIifw1UvXGK67ZXAUs9BBkVb0qn9ST3hu7b4UuiivkqQZidC6j88pKUG2DwwgYqjAwErK
O8zeT0ofC5kWZS6VVogOnlMEnHZNp5B2I3ACh2sxbxC/imSpPxDRGFZPCwKpBb7f8SsMdcL2sTAk
sj6Up/+yA8fTJg9r+23HOaRkPeclgWdTVLg+nWraxMTbItiFuWDyEBODVEs9Jt8IQYr3uIIzm422
RTJCe6a+sZHd+8p4obf3CSd6QNWvMKkyxV3j0PC3nLp0t4duaFmKJkkO/o8HRXKlVwRmwUohIjUt
jmbo+gdOnPOBHu+TrR5Vk001rgv+EZNwRFld2FWhVD+reakY7jsWpvFv1uZ9VJ1yn/1vCRoUXMrl
SGB8si3YvUQgJnmYDpqVVvwG4vIWM9QBwtq0Cj6RqUBMuD9Q5fg50GqqaHMYoE0MVCypiR1o8zkD
XK8vxIkD5Ef7s6+zs+JeTGwMivYreNoMwOF/MU0wn0Yw3nZf+Rd6OzO9sY6isEOIUkz+uaXizWEI
SX9mDMv0+T7txTzz3jcH7FFi7I2MJOCs/r4CJZAFdLipqgU4AKrVrstnf9Yc91NmWtvAYk0vcc0c
LhgZgXYwAbJ/+suBSQFqT0DQny0Tm8DHn5Vpmf+USkp+Jo3dLERZPWRJwNH/rmPKWVbneazE+x1D
nLtRKQqYCOgHPDdJvjnTF5K+zJTB1qps2NYzD5oTVu7M5NpV18EpPI4xLdKYF+l15odJnBb63uME
Og5dG8Qk7Bx8ntBQu5scA01lhx6UEa0f1yLh+YSTa4nfWIECS/jTNsa+TSpsIDTitljn88DSVGaf
2WqsYtD0D4Yl7xqr1NWJt8+K7S+GQ0+9m2em0jvjE2bgLfS8ywSRcYim9fnFmYQpyERz8C1LF3Jl
xsc47H9sJffP+RjS/FYwrTpYBl8WVF80OCPboElpQT1gj7k37pBD4NHzHRP0lN0MC56nj+cjDw5A
reysdB9h9mQKXqAXdyLV/YXiodL9pP6etdjB2R7EiTuD2w872Lir+EnDtGU+j2HG/QbrNv1kTGL8
cuj46oyS2bi+a5iu7hCXcGLlGgd2fma2bo7C7nJlzlAWyT4NyrSt3pZvIXdrdG6S5RTSW79ALi8s
uIJ0Ww5dnfK7YUqNwhGhXP7hiXautUT6/Y8aO60HvLjjwfZZiRvQ3dAk+VO61xsW0Wyb6z6DRTh1
lOKxPS7yjOdw6oZhc7vL2RCHm/tG53bHJPA8PgWg0BlHajH5fD6r1CBZqIMAXUgcPitG4J54a+33
xHdYuO8oW/Z9YNneB//xWrjk5lmmwRdTnhvwZmIh6qNX8cijaSWbrWj2gPx35l9FUlkkfITg9ysB
2Lz9sCLq3d39OFj4CoG750qFCWESvgKhqgP98tULn659m4OQtITYvZ4uZVtK7A6htoKSVdtLvjZ5
voMvUw7pIeNC4NjpjuUNnWXfcGW12v/DLrwXd8A7oWIzWwrufey/aM4CnPwHBUMn7BxsEkmaptIK
rL7d3BXFw0abduwN+EbqU0sQw/Fv5xXKswvrda9OTdyhAlhwu6d3AEmWWqCn3K9cj/PNwi7SH3je
BRwmzSmhTNI6ajf3ResIruuCDThdvTcavqsqrIFSJrTfgDhIED6jPBCu0dnVtUcM5Ff+Fe6QgLMn
SfVY0oTwxe66u+3QF8rtPgq6v0CrR0oL2+zFr+m4PTfcBvNcEIqGRhDxMwwKRi9fRWAodYpPJzAm
anx3YMgPhswTjL4J9dqrB2cmkRFm/0Cz6bqHwNWrh48PgOmjpbTSIKQVficRAbuEZS2Oz6WsLkxt
F2zvQMh1IjS/Zg/VA4RsLcJWxI552SCmHQgFakAWihfqQfZYyzHAYS7+EF8BsMm1KNxor+5EmCSS
BjnFLJwkbkHoo5n5dUYjS3T24hMG6o/KDsXrUlJZ6lUooWvDOIVvGFPNibDEb6hl80WEEO5dMbuH
/1XOp9UsLzYVBJSQ1torLWB425Ns79CaJ3wjEb5S5sGjYdkkOIP1Mlhg2kNPS5Fzu8Ct0Bfb2cqs
0xBvh0gjnFP16llL2IVsuLDUHtukR5mbdBRl2Qwd97N16BgPPtHv81ORRIQDFqdpaBWy7bhj7xu5
OrhGCwVOhImvSBLylI0N86lmk3Kn/4rFaz5NmdYCHpOsR4rgZ5GFtKMsKNqpLmTeY2A9nCex7m+F
oYljNl4ys4mQ0p3aurngN40gHRRdKI00a8RsT5lRvz+ODhzERXlV+KHvugcgcPXeAZ75DQVsSysm
e5klWo3tvCy9VMHlllslaVGCB5wH4y5c/3sklfeog9jbsKQ5Rl6FvykaiLBnxtzgzZi4hPdWPK5h
PiruoZ1y52Zs/XkxDafvS/6RrADI1Go2X9Sqhp+COzXEsYY/rwZzogCQb8Abn/AkEAW2PlXq8ngm
8BvnsD4sx4lyy6htdsvOfbu+VhAPL7bgf2TCDTcrwtiKTs6AegKh44r2D9NV7bKl4ncu8N8WKM6J
wVDaeIQQ0PctH0blVFshVpsDXCCwGsmwGP6s0DmREGd+jUqFDSQkVjwpeYLsMCLMosIqb80np42h
VG62qVhn38MufbxOB1pQI7RAWdXkDeIyGHnXK6ZLltuJXVNzcE1TZCXHsiiO/qIJ76cD/zMUAyDY
0yxzpGPsPouOgknJxN9hy+vW6t7gSe52ChCyzThI9nx/fLTmdg6AL6batNoqNjB0/vQeqwrTaL0a
hYlgt3FIgRfTvFepwwSvEQiA2hj07OHKUKUkqagjW1l9gYvXtS7r2HcXNyUQh4CCfRyY4V+4x2KX
v7oq2GDmPLjpZ1fyATQEwUWRNNGQcKOSr3qGqDyuT8oBUTsPIpPx6vfvPgCtjy7nvna+EXEzBE8x
Kv0wCiEJjHivJU1eVeK4g8OC6skMXFNW54fhtYUh+47pIhU6fZ4xuhtn/RNY908sk0X/XHPbLp4N
ctXk1Fp0Vhb25IPSVEs1J+vwk4VOdcoNRMU0mOQxsSZHoTb59U1/Dox7LhP7Pb4HC61YZhnVaRNS
gvixrwKhmFrxmvgrzA+S4XrGmcuQWK37diMJVVUpQyjQYF/0f42SlFCzlS16i7p1t1KSbWCutZCp
EyBRZTY5FHnvHeXQ3Mm1LRQ5tL6RDbSmBkUPfvjAW7SFhQ/bIl8ZK7wpD2Ke2oiJ7E9dodtQ4W5u
VsxAph8WKHWqZ12C7yyOzvjhNHtMH90m1C4qUApPHfxVaSBNnj5xYu2CDm1YTDbDxPZe3uqANCil
Ki5BtyOAc6Ae2It9HPQdfncVJlnb/PRvxi+PgmlEvcAFFBo1EMWA3SVoxMzuC8ZZXmrH0dyXHZ3s
Ry1qZIxhTGXAchqV05D7ONDNhsQ+oHNZYKs/OyyDSsxERiV4Z6IOzcga67rAtyXvfKjSEZ0nfjO0
OL2nDDKoGNuYBlkqo2HA0HwMkIfc2fWBtoXCTNGhX6IsyR7cyf1GO7+FGjVHcJQlTtt7i05icQl6
PlPFX4ZsVJGgSxplnkKNIkiZtZMUZqDlgOiH4AUeNyPxPz32ozWfv8nkfjzZZRy/LKmekEhAUwT8
9azkzVyOWzkLnQovnjan12fPocgYLSJKSCTZyWL+GgRGqqXWhNzPO5X9TkgWH8KySBiuesQpohbC
YF+K2y6Low05KbPjxLTKkmPfUSqSuDe485/DcMxxFQMj8RTKqbmjiHqRWiIfb4JprpUyXyPqyUCi
xSlTgew/58ELd8+/jYxD7EFI44Eit6LzQPyihg0MQVNXqtk2zLJ0uXhUwEn4EhGEZp+7kp59mJgI
lz2VGlXh+JWWL3Qkc33k0+hHR30O8cJdHaHGU0lq/vGlA8NWvkQipkLzox4zozW522zgd1VQDx6y
fi6426QFttk873Q4eJS2nqoNPHIQKQc6IEznDmdxbIobn9+JqdhVXxhX/31xKR1/sBy694L0TxF4
a5/Z1Cm+XgmmxdTvdB9HNRYEroQvtujoBQammuChXvn8XWhmDTUN8gvQTdDy38yzH3Nep29aCVkQ
TGq4LpDh69ynR7obHW0Pq2+tI2cnBMkqJcjOhcea3/IvWqr7xFXYk6SVyBo2kit8N8WBG7bnN65z
oVcYTH7M2oNdhbiQeao8slk2+27kbuxCsdILQqZHyDF5ZGd7CG38d0MO51vwx4XqEm5N8lWd6NXm
mrRQTVGN25ZCupL2CEQzCG1SJVrLnIalrEdFktsqvtEy7ZAyRF1YgteI7+K2fb1sRbiJXUZG8mvV
9THMNStd3UbC1DCsVgAjFihQZ4jg3yrEgQ59Sc4mqRgrhox5SMNrZdcju3uD251iiOiR5m+l6qiS
w9TGUHHUCPaxPXQP821pkQpo7wJIyFBa1iU47Gva3SQW0Xm+jfbXlGjwFDbKLAkpb0HxQpm/GyeX
s4VjdVQCWXCeEnyMNGcMtjKNj0ol/nMy14xYPUTgOVGLdL1jTCK+WB1vVHZqM+wDQSd0nl+2xvsl
Of4o6Hs8xbqgcArbM4l9YFQjwgtE3tN/ATJT3aybzKaTDscuRiZwYXEMURhTU9x20mWxwh528aZb
eiRZf9LPWHHdxhBE8gEWjgsj3cMSFUjflTPhBsH6LbllNKnvtVOpTgbyFuMSZxqbJmNk1AWen6hW
6RN7oD6w3Tp4LETAjF9VoFdoRku9o6BZ8RR6q/WX1wAEvyxxzfJWAtf19RrsDecdBg1Wl82i+368
X7/tDW3Q/lKNW4MOcUZkLK0fIw0Ga6SxyHj1ctV2965n53AF2PVAxLzSqVUhGq74uDBaeImwFNnu
dkQbeThoKqIC2BNo5rOIOGtdq8uai3vPn1udgtxLxCwi8FsuJQvDRdKbehUkehPtJLzaHzhJOP0F
WyfeREBpV/pcx2Nvtf+Byc9lfBmxoJgCoOlhEZVg8gaVnRBJcw/tEE7YfrixoAiens5dHeCV60VK
hA/nseEi7rKpjOP4Lsj2dnzgysAc09QQJGIgr6qDj6/tp9KRCtLcpmaU1WtoXh0vBYjZ6fGf2uKp
fynkAjPo5YUm3o9s+n8kGn8NXbYesQeJF7TCxgvP3fMIl0UoAvSol8rNJrIvDVi4k7xPFQr0h5Y0
i9GjYvyj+AF4fUr/1ozdSoqkV7yJtmwv6budd/0iUsXxXdz3cPQh8GGxAQceJq+LdZc6GNP1D4GW
ww5Alq4HFK0wqy/fvki1SqgDbrQBtvk57ABHWQ3I/Gd5LKutAZyq/yyVAdA46+r1fK6yh/XjOHGr
ch2aXOybTdCVQeiIbNoQXY4A1i8IPHsBoPJ9r3ga5OpzOURZJxi5aXLm8Da09aKxo+Ig3WPDCl96
oNlwFPSMaxgb+EiRcB86XwHpIHiEwnrnIwfcbZhg+kIh0+T51mOl1Z9bNcRlFLMtV/qTRT77HbVz
YW/YLZm/SEucgN1JWgcZCkI09dzfSuqfKpOFfqX1G7krlYXmNvh2TLdwK3xGfLsYNjDvFsiOvuW/
IWSkfbfh0HFea3v1mVOZtGOp+Uq2oA/+Rs7OTWRNtaAm36BlT0RqG404+vP9kssikr0PWPe3+sXd
2hFsKrPykTOtWi2OUWMIXp1lJlAqqhfLgF/xVcFXD7L7HVXFSBRdVRiBwNfCYgUNYlU51hWnyqOj
lCP+/SkoRT64WC+K8cKk7GH8B6V+0JztR7bQBjG0/0jiX4ivfX3U+JXCPxcpBVCSv/C2vnVBSXOk
FAGR0wlOAiBsvACVaX4lkZROgqksJRTTSvC75UmW866ZGWCl55inzUvv9A+esJLtzfG7s17OQvNU
lrnpWx3hvQrU/FreRnyWC5RIQO1jDkIuSi8mdCeJ8eMHkUqeV0yZEYtANK6KpQztlN1pGKKNs9b6
Qv+lQge5Nlaw12CdfIs6ZOrQPShBnZK1NmBCBf2JMXByWixYun8TO3+DY4jywWxJS7exr6MqB21B
Qi99BQ74k+HOGrOhrYFcLjHIzX2/Xd1nnotvyhWSLVh6lj31cOCbAQKAgXE5x1hwsJugZurZPjVa
8VuDSiZSDJGtL6W1tCFYf6sqlIDLhMGYyG6mIiSLZAnX5HHO+v73OU2amHnDJJyijrclkkhzV8JJ
ZHe0E5vg/G+GRp0U0OGXbvwJRHi+U/EWYHSDdHkh0FBpdeHqXHWB9TmdP/DFWNF8GSRohlGAAO19
6iUBDmsO4jiNKkbFRQnrNXU5jkUhQkTt2WTmCdvpllUCiEgB7gIomMjSJaRxC9/ymr4VRfRuCPV/
tPROwnZqgD6G2Wc/wtl58yKsYzlGxASPSOV0auc0snkLV0JrfdpfclUfKtaw4uAxqoP5XQDydaMn
L43T2uEpPhDTKFrD1W5Ot7/N3z+8MNzIb5m8iuoxaGBWMHUZeCMl3rXIb68AjUtSSCZrJeYxXWIO
VlqHi35uUNGiZA0+5G56R89mne2BMNJFqi4ypfObfYMZe/8y8WYSH9A7XPR77FZW/fFzBVBdpxR+
xBwBRvnlzk3mAXa2xmA9jWbz0TtlcK8p73W3X2VpP9g39SCGafWtLXuO4xMlR7BcEwb9GDyJIG5V
Ng9U4fBWQ9g+0kmL3l2iy9ULUGdhzhA45ZbCjwKoMXD7zmDpLi6UBFkEtI/mMSQV07Guuc2EYe0V
vhxYz2xxwm4ndw8jSg4NzG+loclY+7noz9gwqy+yvWXMWyOv5CGnbh3dihL1LiFwVuxI3t4PX08a
LCgMFejEnkjaFZCfOvzvFfixk1I4NGduzvTL2tmdKiio3b2GmOTEcjXjlzt1ZT21Ci0W6cSw7sPa
YHIc7S5owS5O/WZhCTSpZX/7h/6E6zAIG45g7SH4odgq+8x0jXAHCNSRkOLZMf5VUXkIJdQ6DMAX
XHngFQe+WNwEgzhaZ67DTm/QT5sR3Mz+hxN0t/L3/QFZEMcEzypw1G/qzXlsKZ3qcFn/3jgdq4D8
NC5/GEwdBnAH0+6V34jOg9QcgCzVYVaz1IM8PjWSc/gKvKhCRIBHjRnAdVYLqwtNwU+w+TRDIN9i
7KGVVyYd+gj3vbx7rXNyHoCQ300v2QZ7h05dbBII/V5krOXiyGvqxxw7wKO3ZYhk3USOkt8r315K
wzEQ9TcG3OVOd2x1GmwL/KKB8uvAX08TueI+yllRFYbWirV/9aUim6OpdQIwABaA1g021x+ezfol
xdIJKQwUVRoenj1ovOFYk9q/dLojeATjjKMG9I74VgJMxS30HKArOJmg4Cd1T4Uj4BCd4N9/mb0B
1fF4pi9nrGlBPXWsuhdHdWt0767WPDd/ZBYYbJpqFAKo7A4TGoeoq87Abni6AKS3aoI5TTp0CjQs
Y9sTBSPXsyPqVVLDW0+M79g5JH/LRm4K/Y+DmVTp/prgsOKl2Xzf+0uT7uOAruZk5MjGtqqSQi/s
sObain2/tn08tiIFrMytDUOroeobc2iIClqlwGm+KbJ67KVTyx0h+KOiomTnELfVgIsFfoXsEMy4
az3b00bZ1Pa3PZcGbThJnmdQd9rUxu3RFGkf6xi43dfd81BP3htnY0HYpxpcTvS6YFBcq6pc/ffz
BFB0MRwk3WSQ+Hxq6+anVGqEJ8Lsk4+SieHezySgApx4hF1Ypsz4fnj6hSYRMoLqW4VQdCJ7TUmN
I9ToWcgT4Z3r2Yr0bZIcQn7qyoS2ad6olI4eudJeD20MhYAre6JfCfH2CQsLKqcIZdg4xiycLVXm
rfcKoTabsVosfBACnGMNVN9sb5CUHnLFjTkt2NQRUTrIzcCRwj0xUURhjMFoZ7mfrehHE6+ySbkb
3jB5KmRjAyiDcRtU9T3sM589hzJZ3TMVUSg5892xGjFWK8ikLZNIajLQZqh5Ccs0Oh5HWn1cAfZr
hYisocn72RMiuMGUHF5rsSkz+zOz8ddqG8lLxE+HHbUTA6j3DPHMSf/edLLSfHNAKjiloQBpl0SX
liqKupyjFWURROXE4W3Q9pk8+7iPVbx10mjWGu6PUp71q6B6pGZEPtOBUgBeK7ezPtvEIKEehsha
7fN9pZH90pn+h69GazU5FLyY9LxEWtgYeObnVdOIwll7oxvD981DNm3w5mA0Xf2Go5X3znMMNNgH
NrIBDyrFzaYoE5miF9dFpzS9daOdMMf6lS7EJ8E5euzCy7t1rOuJzV4ismCEQqNteRvYykItjshM
1iG7BUhYtbTpiZwaWsFqUaUrf0nm6CSq13lUyvOv6lukT1akA7rT0OzwdbYfeULz7fo3kT+En6sm
VJG1kLq/MJiKj5UgNY1KO09tSzC+1/WvjZHYXm7dHq8+5WZZsnpiMqPs3cQ/Jhsb2iP5Go8JpWh2
u+Zh0lwwVn1LeCwkw9VkkTfVB1VreWTidGX0XDBRioqGYJGm1YFMfLZiJwzESfx2ifrxzfGw1T6o
+72m/pHiTwpueZa9HMEWQr0VNGCnRyIO85ZMIvehsri29Ikcf5e4eRqTu0y9Ir1TZplqXHVJ7B6P
Ybb9uZvMy1XR0dhcGoaMbZXhfTlUzw8o3+36h/xd/ChZBTXC6ORveeMVuTXjVAaNTMd5DoQnQWIL
4aI8rGgdcx01RyViFeFTctQtDbdXNhzTafNgmGVoXrEECoAEAHEsn9AKbVd+kPaTAk8bu5eUvtmy
w81DZHmd1PaH2wcpMwuSVvv60jwZF8tg1gJlpPWG65SF+l4qBlZ68/fGKynF++KRElnpHwGXIzL4
NW18HK+dutrK6vOepDjPiBKopcAVtLbutcsvRN8Wrq1UKHXekVjRbUk6ndXuSkDlU9CbgCabcIew
i8jKtYrwdPNgmJyJ1FSM47OlCLJO1CsXf+jd5oyQAeGKKPW45BG/28tO6xa7SVzEBoSn9G0+0FFu
qDSkjVG7SsAlu3nP7P/B4/WnGs0HsrmOeWVIUO7pg7CwD0VJxMouaiU9KOCwiU1XkQz+3O0mRarC
lkIgGmZtP42Lr//gPlOURG+hVO3DPRWQdIKcMImJWwpnWGj0vBdzdUyR0e7goAryAssHsdod5T/l
DbFhfYByB3sSi8XbWqBney/YFVp5XTHfKAO50vdZ5EEZw9XQljk4dqk/1MRXwuznuWarG2G13aVN
6w5fGWVWqMgDNrEzj5KX+bzmURQg5fRkLQ9Pzr/obrn+wCqNukNl1piGnve9sMe1ZMTb2YvO0piM
tJyWywABx5bR5GQjLm2ffB5Q3i7tMDMkOWMM1IWasfFCybYCnBhIi1AERzIhsB+N2o+2bIzs90Lc
lMXqfXweEwxBNfyfZVhvmbs4FDi2B+WtyejBqQ32OQl6yMs1rKf7CWUfJoVcFwkpsKgBNsmEd4mW
Xf8RchxtCcc9Ke5VGSN0l0Rr6U4DqQib4I3DV/7Hhi3AeLDO0RCNMEOqhNxfubyOhM+z6PgqpVPD
ju2yoxMvCfP31gYGSPYjY7+kdz3lTp0uf5LWq1gEZmh7vaE3GA9YaI4SnwXrTXX84penecfVnhJE
VDppPPM4cFMbQInhAj3RUrDvqX5hWwrpn8GWdevlqXBUVdVqO33guzuzTFnpS3+JX4NCdDbwJiK6
5YlYABxBYm2Xwri4F6T0V5mJy/CG6wssWGlT+OII49E4lrLAf0dQMZtmn9X7Q9l5+MDF8P/bBJ0k
C63398dgQ0aASx34UmDXBzwDENPsMakHgaH17FNGXQi5WyQG6dcOlih9bmM1hZMdkvtBk9jHCcpA
p3Sjke2pdbvQyMJGUZXBLW8GeTcaTmram6sltqbLnj5K4yLpsZuP08PfKLVFnD55Zpxz0Zm0apkB
G0J9jFWC5jryPcPRyt9x/IpQO+j8V1kIZ+aqaTj9TJItSWmW07zipEWbcUH+7Wj9zTP32f6Z+5zo
aDMW5Fv7MlFEqZIl8B/nr+AGGWZDKI4rOC8cZsi4wf4yl/hBV3c3cq53f4wCcs/mzs8w+tPGo+BF
8scB0UUTLtknuSabQswEsG6m/bL+jt4fmTnh2UQtk0l8vTtov5rCGS8tKYXKTjskbBpvmojS4lfo
dcYJXthBD4vn3MnvYU8bSuONiSZE36N8bZu2jEs8WhfPfKRx64Sm+iNzScCyWitkbnixI/DDRRey
Aj+eLuXYRErfRE9HH2ENXjuC7XtGOFCXlCKzVrp0IIZ3j6G+hInDCytDmsZ4Le6lyRMD7knjs/8X
9qAxECaYPXpu3IuVHR7yKEKxGYT15ey0GEUU8iq8r3/ybmT66KaXXMM8GRXcEberGegDKpGeNEou
fB01+mxA7ot3BjE7hFmMoapl1JXB6Ya+aLoXyXEO9qAGtQ1GYnqmaJB3GXspBMC02fL3pZBrhCxM
pLdvxPO9YI/hnPmuc2FpOUzDMF3/mY4PaHpHgsk8E2YN74bYDaRgNrjWUxnGuwGSEmm+IWMoG984
ODrANsU6S41LE3CI5VYlQDfrMFOPNOq54plDIve/QXdmYrrnzC4UXYE3yR5RiN1vwN+F2y7lq1Qc
VCN83vnx0/qdH2C6+SY6JW5iF9GoK2O5Nai4e4vCUZz+3bwigkr88+Fqsu28j5lydioxb8FU8uwq
Z22TPj4MxPcueEWEdEoo6JEDFb8PEonMn6/53Xl2So9PeU4+XEjx0aF8ftlcH2R3FVMWs9Rca7pN
bGxWhQcaFfrGjKeTzQFd7Bf5pbJbi/mqNnWa5tTlNNh23dGBdcKR3GlT57dN7zvzgBg5J/tqPeX4
dPFO+SbrvW9mrfEItdN4IiYX3Jh+0k1BZcJslOtpfBnSbyR6YrN4NO+HI+UYVM86aCD1+LMlN7a7
F7IzHo1QV0UlK5iiz/Swa+uMED27BmAukk+pL3QhV+8nXBa/vJSC4VF86VKJ8jqVZy9fIpi1jnSa
hwaouVDJBLKTNj7F0JfSSPJ7JLfo4t/j1dOVEpn8/tTgRIBhmrEVnqqZ/SUbOD6ShDKatzXD6oqe
vzVnxkEWjXQIjRnX9/BOkg37Jf9QndSpkV3bjuQSAj96/gCEyxIarooeLt/t/Pr3f5YUL/dgodNg
GOacCVIuuEUlcUqn6J0PTxF16Q9HIBVJlyBl5bwV2tET83Ur7iRhPHLMmsWq7eqvWRtlkPhePD32
apht2VhTa0RAXsUoPhHXbllqEq5UEfNKw4n2yliNn+R/QmmpcERx3ZUdyIKVadh4bvgL9kjO8VX3
Va75wM659xbfvkBe068Vm4ml+dwW0TDwWEAVTbyIA7xZB2kl0iOI/VZpzHThMEuLZme7Cyshh/Pp
1hLEoE/hAjQOSoeiM1xWd/qvCEV6DzNT+gbtpVanb9eQOAF1cO10xnVsZfbMZ8U3nhTM6+zPlO65
xBAuOnqnk3QjfOizD36hICIie3zCTB/IxRUC5AQou1ysRqGh2Rq92BohTCiccqeuNmqrreCrGE0e
uGqD6+QbAmysj64Gt3pOybXsLal24TVMXOEghDn6g2UH0gfGyvaWgSkvv3CJfdj+DNV0YOJ9ki/v
WsKRlLTHcRRoVxtpuKcvL2y7mTi5azTCbUtWNEdG7wAM4fRGPo9lNFWp0iHRECBjXavVWkYEWXQa
awIdKtKdmulHAQ6oFpgOeO7+iIb0OhOFCuSTIQNlZv+mEhKLKa3XsfvMZzvOr1uU4oI2comXg5nL
0Ac1BodY6350MbycHhG0t/njVJJyf889sOWcUOvYbujUE7zaVNoDJqel/kb7wh9Z3NayxyiRZYMk
sJs8ZtVIdPnE6WD+OQz+6Q5LAUqg+jUs9Sr2S54cctmhzGOlsGO4xxIGUQINx4lFyB0fql77OgzQ
+jbbyajRnlBpQTv/i7BVHJqiDP7uC7SAbMhHQPiItuKAudxrO4lGXBVFMq7TglIHrfNyAi4TjjWm
nTiTtSWuBqsRfPPKiXNbTCe2sqKJTaAyTC+9MOYn26gd8fJnCS8ZBD/4/FPIkKkjMuwXjviETKVA
UJoOflwICAnc/RGF0Z5m7VXo90sDvdngDzYjT3DGVs3Xsmk/SCH2BqbMsQvM+lEU/ERfJct00WOT
8pkAGvgzG00eBDsa3zOZCgzcp19Kljhq82K9pw78QefSlo26tPTp0yq6gEk8gO8zU6nE9sKpxxub
GC8uaSzqxLp/T62eed1G2OWjJIek7w2aOU6YrP3GzZlUFe0GE1rrq4JVtkwqlYbuMPZtuTEaYcEU
e1+0KStn8mINqJUQayc1HxkT4f4KKzvLJ0i1nq3LEl595ZQfeUnui75rCkN60LXyTIiev6Xf4zsl
OT9CXSTtu+9FILNmQ7zlcpckLEX9KmWiH5Vvoj2Nw0TSDK+n4zEmTqyohPV75tdpJhv8mtvt4B0o
58Q7Gr52vaJ6pmjKv2zpLb2Jl0pwLr2vdsBguZoCX2tz9Zdx+YJPGIdT5HWCKvkuMUutSLehzPQZ
1K32KQ9LJF72XtNF+68W+mZX64zYIKAPcxFUaMlZRGDjvTOOf+7PHRsh0PC7zkDBbsnCW/5xfMyh
Ae6XBAuFpBUrbRy0R6H9aFv4jgxJPXpG0uK9LAOn7DspeAGHyLmqQ48zsQ3hwFb/5lq4yuMcsLhm
7BvpwWyk1psO0o4ayl36+b1QSTQckc8JMyUA79OxuZBpuYeXZCtlEj4PiFpnq7R2wkV7RTrY82CQ
8eTdy/uUDuo9LqxUXZsSM+pMOT2OCdw9Thc4wxJaCxcxqMEv1MZL/VF8TurgK6nCW03qFUXF2KZS
JB2OjokRLkNdJj5l6Fs9VxjTphPo6kyTL++ele9JRGj3XXWJO1qkcDfPUnstCY3KMhXaGf+fVEHJ
j0ygD85BfnIoF/nBFakQbX41ZNArluDa0eBlzoI7OzEgFro/QfqKqW7npXVtR0mLQSqIPpiYIvEW
Z4uZ+El+HHfmTYtn/dYt7KScCCnK0QMEyhrTy3tED2vSrlXcGkguHE1qt1cg8WHTD6fjGpb7RF9v
jYdQA/Wk2wcrSezcko7NpiYWIRPD+qkrSXqfybFfiR3nFxDmYRQAgmP6l5qVLMG1ozP3pG3lXM3/
oWoOGv20DXb0jCV8hrW9Oq/XXllqVLMziN0ly8BJnVjQGG0Di7NTXuQlqpMXVwYNR094obZjaVhF
wXjJsRXWQOdHY78Rd5wulohuNzbIVikKNjRNBttWDHZrXL0DIltrRyD1e3SKSs6Ofw1nBnPhr6DI
IsOdcjGM8c2vDzUN58qjLvJyyuKfyJzdhmu74xRtKD1Xw4sXB7bckCppVQX8SS2VVPayUU3jagmT
bQrbZGBpeT+ePxOkgymGum0sK/jSeEbF7dTtwU6NQjiZktqdilHNHhYnZrYuFimQNxu98v08Z7NV
A5XiQFGNg+jKnrdaS+NX1e39Eb2+gvNnEjrw8ZckxgcuyY9W0pQY76ZXJ190jPi1FI8+MyUYcQGP
g36s2Iw+GOgCzGW1xDuAAsd4qHKxXYd2ZHmc/OELM5UxctYXGVzs6mGo8IwdJKfltBpVFaKSuzU5
tq2r5l84tkZ91Vx5Q5pXcpR63wMI2sVBZza9lobxnEkv+8yH06lYhv0uhjCAt4V0k1vljVngx4Gy
evgy1knNljnHVh0f+8ye2kE7nEPGuql3CySZRAWVbUyk71+e+otHMm1VGQTVEsgJN9M10Ufllu7N
hknz1BfnRk5sMbWjKu+GKem4HIJhikO/L37r91UyiV2reCARhPVs2/Q7tePvZMRvcN5sPD//iv7U
Sik36mzpho0TA5qh8aqmTZNNPCORNo1T6ovBoR8BxpBBghKcvEdvpiINfFwSuyZIBnQfXv7w07VU
rWSGagg/BXgW9/yVJkzilChcDbtVy3VhaOTwuGk81zCMbBS61B7+gl7fsgiID694k8x85B2kNISU
R2BE9IMdJF9/G0YKo9mXkyQbhubIS7iVS4y7serdm5gyCEIqUXU8VqFbTTO0avaedhkp0zFL1bCi
4qTF9Sy6J43UeNAoJMJ/Ot6pTUAVTEVEY5yatvpJfpTPIT//5eEmRSSmf/yDHsMT5PKBKT+/7Jf/
HJNvTNLS31bql2OGNBvMZePs1OrqQNGScsm5SzanOhw/Vv+EFZdVqggTWCGDvyZ8pJ+YS7ro1DDU
4RN6pH7Zqt4IQ6ZmqThU0S/CaFPTy4IX3krCAD7ZNWQ0LkI8a5kYeUuzzfxTE8aJ5CFW1FwU2M1J
quha6MqHg+4nfZfhkJLPo0jcBmG7GjgzgTWXIwf+zw+RzDFIPGMsbNy4EotmQzLZ8LHrH4maZlI/
ERCh3qT2MaILdiImqArjDTn7zsfAFweEVjv+ILPTOz/9jXk+o8agAn9WPemS4CwE4WjGx6ZJ9pTq
UHbfRjQh+4n4gvLMKun9YdLhJi5rbuESqmZIwXDhMNiepCkSQnDDjIKiLRobY3KdytIF3FR1RZZ/
mVhVmTLQPuRACTueVVnfA8/M7HdWMNKwW1V3FK3e/fiOdmrsGI4M7dJ50JUrEeTECd3c2v0y6I7U
OXtZ7Oy7hdXAnNacmYBFEPE/WHNgogbigOvEuCgC8wO6x2OAsjnTet0ToHTbd5Xtkl/cEAAgaVv0
85zh7OzBvB34Wg/3Wesknpn09XStdMVQVkBt34Lf1jhYouUfosKJNXvINICLxyzOqoJ08pmCyNqo
B87VJEboX5U4AfO2XWr2SjD9BOEoAz/6eIMVXXgQAZTf954QnrHBmZqhnf+YuCxhxz6QFdinjCNM
9rrqS+0G2fi97OCtuRY0+uSmj6+ul8xW6D0VwcGwf70LOzAJVaIeTDEXa1Ar4BXhi2jmxHdLXmUd
LBcsRHwJeG6Sr05DKbAZjqoqL+3aceeQ1JstKVXxq7Eke38zd2rOa291htQ/XJSkTajIkt7Lwz9p
KJWiC6trxe2ziIjRkFV3ikSNXkA8xBLK7GmXq9Eg1Bmnd9uKb7QrZJyRCm2/OdXZVVZwmf7XrDSG
usbOLnG9gGuKj5n8XgnlthOfowyBP+GUyXCFzgwfLIA8pjgIaEhegNRS5+pTLnPQrzeALY9JUZdp
aVWlG17J4e3kCoxDXvD14kRNLebGlWt0kKLbaZvaF75Bb5IlNvC6tHA5PT9bwqFDhoWXUcG0YA2v
uWZ1VD+uH3KZHGBnJCX2MDjoIgtqiuQt9r85MzoTNZV3S4S/7hI5ICy7cHcEbSUVdEogtFvYueA9
Bw47pF+HxgHt0ExbAy2byqkfGCDsjJUVFGUeVDiEf5RnNRt+ZbdAcFThfHBl7r1W1pMxI1W/2K6I
K92m6E7ULks5AvzVTtmIzqIqXOC4Fn+ntyyThqHSvV53no/2CphYpKBkrnUax9bnu2rASkc3hsFF
5ygdfuXNlJrPKj4X7gK2MH3kAZKal3/KEnnEPkgHaTgR6hFxI85B4VXc4ot0bVciuoDUrQeXQKZ9
tkhqq8WX39x1oe2DMvBQr2jwA2+QKcxX5dEXY76Z3TUssZjvk7jhJnTs8zBNqB+Sjk5dSFUeWezW
oGHfLuSwblKYH3G+FaWHGnKZ0jbegVZ7YAOfYsmuPpp7RqL7KNDNbDUpvQhk5kxFZSHZEAokpUlg
yC0bnIhw9eKEPi39Cl7WV7huXSezyW3p6ZWDdkasm3qdyUrld8l9/DUJVY7sfD1a30gQmNG9US1P
374bFWmnyIlvTC4Srh4U7z7SuPLx36W/2h2QqkKCfvL6Aict/QoD3v7ykdDLTZSrHbGAGHvbn9K7
qWwWzCOPcCBJlsaM7dKrJjsrJzEzATFthkpU3UKgqMb7HQBAcoe5dnqbfb+DRAkhPuV5W5JQhcrr
MA2fAAlm04jhUY1rE32qsI8e3HkaB56EcClXYGv+n1bKGBipoQhTQvZM3slt6M8ARp0jDD6yBJKf
ybBjE44bYeDoLAmlzE5dY9hk3gmkM6lEUXmj/+oiZjuNzWtZtNxYjMiG52EItkKH3x0Urd7UKBBQ
vWn8+CA3RJ0PbwdtVE7TWQww9YWGlJOyrYdcEn4qsUrkmPINZObVlHjbv4f3B4/aoh4T9JknReQp
XdqEd4ohvbvpM8CEwe6mYWo/qNObN/l5pKT9v0ojjajcQSqItReD9/WJizoSBp42jVTYP5qpA7g7
SItwSzSgAyAUxKcTKTaeFmGdp2o9XXzq40Ws3m2vXnReIs+KpXyOSBUzBESYso4kHxepYyYEWmf6
ZdP1TRO/Xe7TgV8/KuHSJKc5JJxJosokzzxx4ZX8cmw1o29/vKSgQ3pP/IBQB8127Fsom0KfTgKt
DNayZzcMeozeQLw6UWXSvLCJowSCquTO3RmgeB39SbZRugXZzkeKtgExLuCcSIB9wQXJxC25adj4
2bdZMORizvwbRj3IWgf0dKVx8WpgmkvguczuurMRdp0CA6EBZauFTPe5wsu8iijXusG9Z6QSc62n
mbt3Bq6JNVTY24BTd0mi8Mix55fEMluR+Hqy7BKdvoLYfju0VqKO34g4f2wxs2zF70pUSeDVg3GT
vxbNSqSdyBc1ehsWZl/VmxLRse/uETi0KJLlUc2+SjADRTPEUvwokMEX3XnSmigwFtMfK+hyxuwE
wRn/Vd3xTZ+PJFw3g1E25NckMza4WlyOAB39JHUrUpCbmFq9/NrBAkFCz3W6gNQaEDCtsPReJRAy
erloRDTizYy1TuuNvTngCzx6lAMXw8B/N3kel4jWSv+k/zMwCjljlthO2OeknFyTBZinifYI8M8H
QhcVdYTOBNSh51w5g0yFEtAF+azIecKAZTGKgyeyy8MJggwTTGTUR1liUuWKpdeSSadZijfd40Az
kIXTD91qo03AlRmkXIOb3xC8CvilV6toL5wZyrxoDtjh14gOdtmEPz930ZTVlTE2RaovBywZEiec
7p4KRGP/vzmLDgxKIgWflU0FAbetzZYncuurld2PPRkH79Nhlq2+EZ6k1VXvMxpgTnZZLLjznikK
AaUee3VCfx2JwV5aRsxYXjwVWP307KuJ0foJ+9bTCjICEpuNy6XxjqFw6VvkwfjbWs+Zn+b283Cl
hJjlOE2qx9Dyo46jEa79dT7oAKdXbvjVJVFKA5xl6ogMOWF2JevwfWt5hmCvyUuM0K2vQ0BrmW00
jcdah3i0GCZLB0jC+gQvHEBbk0ILZH+YB5jPCpyE0j0Z+YNzYcBjypGBNTh0f2Z/UMttkgP024R7
LtpbzQeF/rTP/j+c/RFDFkP5zRLJ9me7vba2uPPgDo5RNdUCVN2dsRd4jLzQIn9TTbL8OmkKXsxc
WY34NuNL9rz7cjdUJCw+OsKfCVJzovjRQZExQLTHcjgjibRzuJoEdpTPX84/4mz1F0SHbM0kdaoG
0G2euTGyrP0YTX/ISkfqJrkHxtVFY9W+8lLw5/pvSUlNP3rB6lZz5KyCKs0WPynsv3c0ERNin9uz
WudCZh8+X7D0Ax4XhELfyl1XZFxkeqwLph2GG6Tml4vbNdp0gnTcO0df5D8clEVRVW25UzUTG7p+
50G7T1cDxOsLi8H3Zy4KIIge8cJqIVsIwQ4gOKBvzA2NXM/ouGiWUaiw6sMTPFkdDNwV/YJqaA8v
mBe43Vr95auJu6QsSeZrh/olyToxwzmuUXc4TaXnxsehK35vgBpF58B523sLnqaAMt14ZLkvi7o1
juVMFR5a6AKBVcvJQAJmTLhixIqfOLq3Uj5eN2fI1ydxneDzj/LN2YNW6kmt4RcKzaURSMbrdSY0
YJ3s6Ja80BiO+H0Yz+ULpKBkNskZP1WmpQklYyc0tcTGgLlipFot80J9804+/mCLtdsJM9Cj5QZY
vx6K9EVAy3SoiMfBRGLqHd9qez1Xgow7FfTNmoKWrQ0MjpkM0WYH+IjhIRtD+2gZ9idfdklDPfOA
G3DKTuoqfwwVGlM2PNxposH0j5stWy9Om+EgX6JuhcwfOgnEaRxZlfZnYnoTro4Hed/qSN78hQIy
d5QV+PGOXYb2pYQNQ5npZeuuFP24EHgHgJ6JJQ0YWHrvpHhGR99ciiGSS2f23+TzWzcXVJ8KfvZn
QuEbcl0nZDdVeSbps669zTOpuRJMXAdFtegdFURfVOO8MDAKrODFJogbJ5+AzO6NQWwSn/QPhwBl
RrtjzWQY7V6/yYld2pRcamuWOz11flMBsiwjRSjiqq0xgNs5rhkV1fPxTfV+UpVuQLcgzvKDsXqk
PGkAF3c8wtK3yjZA9sFt8ZCkAhZfH1b3/jDQ+Idb109QfpOquSUW3gI323wt86FqhynBUjjMuje4
qb/qQq2uSSrcySHrZNqYNKorqUINVXotOhZBukiPbzo1QhsmKAqxfcP31W/fjV2bzhnUAT3IHniD
kdbI/pRaahiS0937FMYOI3DK342fBWXqi6ZJOnjw1QoX/Tq6nalqNzUPQFT0EsXy0NIVX/9jqzdq
A3wwGOZETMROLiZsi8qxDpWY1Gk6iToxUAYIQbyCaJ7Hs3vR9nXEz0woWYTiZMJT5vYK03R3ffPt
BQla0jhrQIlCTACquJaB0xpQ3HYb/l+ujMnlur0+KGWynGjtkRmoVXgR/KrrYktJxSBS38UsEsL5
yq700oBYmDkq6uWMGW0BAC2Jpx4ED68IlqR41REFpGbtd8NmQfuw2rmXYFvIlMHQQGaqZVgvBUA7
lM0kWQ162Rs0l1sjIlZRaK/Cek95R2m8OZit/w8hft3qBBfTNPC0AxZJB3iFirsY3NPKbK6MIsms
+/6IpXKRtcShs1NV8QwjtGNIJYCSXAneMuwEgoWTwny5hmTJSxNwnbVFqN8rS12I0bWVnxObNXNJ
mCvqecg4Oi8/DtYPZr3gIisFd4P9dbem8SQnNmNI64qUhMFkQyNw/CD6OvTw1TvbI9CU3f1U88pa
/JUDbELSjfFi5gtdhc4ZP37F/nNjF2hsTJjG3OMLPxacmzmvQ2DKEtAQDM8Do1oM30CGK9vdtYbe
8aeXS1EjUbOPmKq5siGcBExyVjckqNx1DHT4TiYbzHK0tyjCfEqThHv1lZCFEg53jkdMpCwtTc02
DRlBlFXedZBWcgLhDUhRjxdjs0ikpHfILDvijCAQH8zra/F8qp4DLVZp4h0ZYuoF2ptnW/2iFJeb
tbTNReHcx6r0O0IE+mGX8967Blud1mPPjv8yJqva4BG+9HvdliVeNl1v6EdcRuw6rH34bCAX7LbY
NnDy0SPFYknTdK2dIQO1Ask1+0cr5en94kAFsRcm6dbY8fq6QRnsBXK4kPfmH/CxR4CIaBtdd1hm
Sw6O+h/RW+BR5WtpvQBIJbcjcWcbfq9Ul4R+VmUzXrH99k+7L7XFu3uf5YIJnc8kq/FRsAcHd2gx
9ZmMa3Y1B2d8cHHMDu978fjSt9EP302nOfEwUbzmbZV4fxysef+wmUgP38xJhzwdyN4vb2tSVFDd
CX7O2OvudVPiFekSZtuMDG4yvO0/0+0xoRIKo0JB9pxN2/RCYmqNFFG2c3av4hfsGjB8pySpFqRZ
i6yfmO4+7kA1BJ743SrB/hsg4wZfWc3CDfwUZjO2KuokhHZ5NodOY51EkHnpVRiio28J+TYD60Ne
HxxFK+2HUhQ3uY2FKIkWjjDksOL3uvaiB/s9yG7Qo+pc4zCe0OgbTE6Z0ObE6UYiAgXNLFhznhKC
82/Cf0WHwroofl5bRjXRwktacbC26g/HVe/Nvslxuasn6PuGQn1/bmqukrmukf39syrU6/4Mqld4
sVnxFLk2pLk0pXpxg3Wp7thXPvDfc+LN0DtxCl7/5eASw75kfpxrn1y1un6cfpShNqRsDT4rD55f
TI2UsBW9YGIHhC/Jl3R8bnPa9XUCwwv1qRtg8kOUblxI909yQWKMw5nTn69+ie02yGXRLUdcOKDj
yz1RMQXIcbncjvHLZXkLRR5Aie7loCiAF0goOjmSavDkjJmATei98M67ZuM+rBMVrOHXLPFLcDt7
nb/COHNZSAFgtl+wJ4v8ublKON/3ILtyfN+lv4kb0So4dQ1dKlE5V1dfHTHnFgBPHnRKtTZzmVRn
YvxWQ522YxEuBHTDAUt5TuA6lTJ6yNUC1H+oFz0bhdeO0XKcbPFDJZIVXgb4O8vU1SAu0tNIGmcc
KjmXJ07Z65O7qL1o628eVvsLyy1Mom1o4TaZbsgQdX2J5/LTVKj3oYwE4eiMn65cJKlHup9xTOeV
2XhZcff4DkhmEjf5ZfT4+Y6ycgiSXTWviKJ9GKtl/0WtZIu8OpWusIHN/BjUjJbd9DTWMTfF+k7p
Y9gBoroy3Wel1YGdSdZKtAuqXvpH/kKUk6vg4ygJjhf9FOHEiJriIIn8Zhgv+bqhj0N9nJNfMIQi
4vHWyLY1ftrVf/4cikdDVCTcNKzHMWtOydUebuUjGV0Ths++Cj1VCie6P6pxC1F/aAqpvHCW2L2+
gXzKbZX5es0OfZoFj9H+WKpQfKCz/yCH+et7y1vSDVv95ANaZNHPMMKBt18yjlowvCGBNuc3xuyM
lY9ky8BSprmQD9i1CjbzfBPbid0yLjyki+PZgXdCVJyQfQX4qnp1N+HqY04vlOwrsy6uoWc3jZy2
3JmtImW0U2MfSB3eX8Ds5dfWAXwqHUMWTbBUg1FkmjFKt37dGFrEQLDZsZ+OehdLj0xBSjNrKNyH
FxWCW7JJzPQM31f/uo+q+SDOJJ7IYXw7DfTOBP1Pj5MX78J9NME85bjQrGharAJqY2RPLWiqy+3d
GhCx402sDN3SdmsPtvX3xCNCyJPhBLkOBj/96lf5YMvxG153n6PjHiyINImqqyNCl6bB9HD2pMFm
84ph/TzZ2dJBLHsAbVhCYAjLDLY+nVLsBskeX2A6m8Dwgvf9/SOh/+SICMHLS24PwOYG5yQNq12O
G/HiWW1cXwaFaMP17nvO9rynf+sK6Zbleaw7bMUipgWCYhB+IAPIOKfqJhONKNh7PkBpcoqYv7XR
mMLhcn6eM7XKMQXDq+SwHaDQDL3AjVuhQdI7q5hqrsWTwRQMqKel+bpSykwIXaLH/BCTxFsH9dYg
R5c3abtQ8aUW5Lbc1O8IRMgKiaZ5/5CZj5xwDcTBkMPq33FwCKHwxsJFya/6dkPD4+3qZ8z5Qhme
5kvsxGqkINzJn5NhdGYlXH2fwUqucRSNvZU8/H+PLlTOJ8FRYT+F99xRhuP9d/f4WpX9EutRzeC+
gtV0izZvCAoItfLjGIpGyUJVOnkeizrixvc3eVsLopPb5Lnb3R+jVmScTc78yKQo3FyJrDR/G8pT
EICkbHnUUrm9/uJZoqBSD9fYCitqbupaJ+BGAyz6bYwh5ojw5etCiCft4HYl3aDQyjKSssTGVydj
mYuJjy3jF0IZIIWoJjp4Zy7L/M6Fo20JP1fBuav1UXcKebp7eiF/By+4GtNAXtmarygzWPJ0JMDy
+YE05c6X9cKPblog36FvWmyPEWDbaaXhgf166cD5nMHFouIBUg+gE9/jqFVPwHP6MuU02jTKWq3K
rXF5nxLtOxDC721sNV0ir4++W87dsu+mJFbL0N0UrVLoXR0pHM26xoPhpDs0QDQ4xANX6MewzPOp
9DrxPZX893Lx4Z+TNhgHARRgyrFH7EZMLcpowJf9Jn0nr/pk0TfYLgSR+w547XkScSR1NxRGOraY
j5W/rjX3VKYo5bV2Lzbp/NVQ7qP/9k1Mx0YbUOAZiaqVaVQElejFwnEuv8N8tN91b+5SOY5GCEOs
+btwdviXgzOcRxAa8kqvFGX2ORHIopujKWRgda+NeXi2dmGlwjbiHVS4X1NlBNfFnLB/xOY+rzy6
tAWGDrqWWv+80WpIGg4zKm0Ayw7HIQsigmkUM628ZIHodz0Ldi2s9Tk0qy3Qu7MaxjYkvbZGwma9
BfxFZSHJG2q12C+QXXic482izghSFrmvhKom6iu9hZ3g6JXUvqk2zt9+KIHRNIo9KusHZahSKP4z
L4omh2Zqjvnxwno9DufwgwVpuT6Lllqz0wmlhNNRDhisyB/Fb107tXckGehH1wzlTxGtGy4Ct+E7
vOCL88unE0oyE6i6BDaSUn2/ZRz0RONE2APdjhzzOVU9tPaCs6HKgoPCmGKu5h68jdJX/wr3j1U5
Fua3Metxq1Slv7IvsCaDk2SXHxJPs+Gcb40lPaBYNfwMMrkwsM4Bvr8K+JmnPpGBQkU+wgf1Noob
t6wMLYjQ0rfbskuzaJfz39FIG9E4JcOO4cn+ENPUSgE1AbbLzjxgPIGalIDZB6g0MzvJ9VFW7N5E
h5IjuTpLpjYurKM6ZHjPv3TR21/glizb6FfiCcCfrkhkMP04Lwp7VoMmkwMMZyOd2b74TLyPYKGw
MVCPmULq7tYGVaYZtBfFcXv3VIfe8I5tc/wxnOocWTTNo1VHdAjKmBdvZfnO7dc34D7qfohjmqsD
VAxZjURSJAx3YpBbWBxgeF9KDEnTPAgaaRlJcyZYiKvFAG36k+p3ywbcngX2QQNz5rYmrWQhskua
SXVKZp7M6ZNr+5QkpzK43dF/aEtzaHYoymlMyJTPb+Vd2PItE93sDxlzYbt3uOdPr9riaLcevdm6
Iysh3JQUM227xEShFjsAdDMqtIZvm3WE+JYNpcDrnGdOHbAj8DxVqjmCZQmMvGyYPwCyGQzxjm0T
3MLiwprjWipGIeuuCL4zAoiIFl/7G8YebZu57+KXXQu0V7gIsUpnVdR1oN9jttSfxJgYYREayzLG
uJwxBrzMcaDpqpnWCT3OqVGOjT8XdftsyBxrG44fOmoAK4yqlU4qTJ53oDDcNE+rqSCOEauKaxSo
KF2IPXyyROvOjYk9jfLIRfwlyNCI5ANS67fvCd3EgnRbk+cw1xxl/UXn3DCL/d/u/pydEWBrZ/lq
n+WQQO2fOBjGYbJauYplensNnO+pxYN0mlBNWs49pI0mXcLrtBAjsZ+xvWgma4Hiam+ke3w7wAaM
XWM6vFHxpHmyjmgH1tAAu2sz4xSUyekEuL40nXrY1/h3WNA1EUpzES4KUryHH4rNiZxuQ40Zt774
ttezpbyCizK9ZSAVrmDUHQUGJFRud+OK2DQpqHKUR/OIlbyT6/mCEJ5oXtZJgm9KwvlJ4zjnRJ4J
aBYde13KFRpWr1llQzLC2cvVmExZzkAQaVxTOhyJPall6lq7LrFqJEm60n7gKMoznjTXkzi5gigU
fjtSIdZzLqCiPeIS1QrF2uwLUm7ZxEGN/B+V+0OB6Plx9oWTTwqLKzKW63z3eLQ8jK2odGQDvP2N
SYW7HTLIl2HJs7n5jjw9vhAGvDau2UhxvDpPsX6x4W//0famJHfQJfo5PJK33YD86IbHj9v2W4pO
w3gUwhgJuBIKCGwUYGSpXZPruz4ax4Nvqa36JGdc7FPMwsQzH4QboGXlIqiOanJmoYQRESVNxHyz
lK/WI0JNgWLu3HP7/V6ddYxmJK3r01HGuW0Ri7HQP1OODQqSZy362b4L3NH+OD/XVG0sCVmW872Z
H24P6sR5uNs2cqrXxHorJzCKS7xthApy9tqti939GO+tzHABKPHR4Xgvvk4JDEh4/qG97GlAAazG
N7GHldwFx6JNr1SFHL0+thG22DoyYqsyZI5cujPh8ry72yjB+pyCgYic7Myou7/rRzMtGz2ctvsi
Sv8zDoSBS/Uert0Fv1NwdqoVqZ27IzzWzfjGahXOJXaud3ea4AX8aIz+qH2LuZLOzNGS+Jk+AYau
SiukE9IYC4/o55XF0My6VNxy+ttYvXccYOqjM/iAcJTgdNiAPyvJ9PVSZNnqt5Uf1Ne43Lp3VBps
u5MWn+fbis0qOhbwivlez7vLlxrcHhQP47Q1QT/eqBVgGigOYLnkU0vXLYUaWNXzrGlZynxp4HAU
+7nLWN1qjC2NmfTdTHvSj1GQVck+xUEKWUP5rAKATG3Qc8ph0OFw7zl3c8Z/+41RDU34jYIcNeHz
Mkuwbq6jCgoAn51YxVO8cWA/NwtHn6aMB+BaDFlIOzWgWaTgbpBwB5kCE5eWWKUMOba3vuRNI/uk
LnqkVpSVXDfPdCG6R3MlZ84qfbgq+LHrIHOx7PI/ddMlJ9ltQTHSNTDuvEcc7/vLWT67kidsXw6U
y5680Iv8hkWkkW1SOMfk9tlW1pmZ20d4AgvmeC2kIqp5vhmSmoinEC77uc3EGU3wO6yd11sNmniq
+LC9OA3XHlKBNLgzV+zeN3dYwLWqH9tSk0PJjaq8elfDTjuKc9JQpNwN8QSAb31SHA3c3TldKqGO
WgGlcz7aI7RUyeb+3mxtgdKlfEFHfLlwVpDqrEVedVpLpjc53CDELCBdHgJnK8EXFEEzK8zQ2OUA
VsWtf/HePg8hEwhKHlbcXos29uzPi6qCrMxTWRGFtcdBgVztqMLhp/qzS6N3iBxnF5kWWzUIVWu3
yFoUbdgm1tQl6D/sjBYEjj+tKoOxXB9d+TZHW9dlNngrMfg4MFV5KqOZFSNBTDIbc3X40c3ZteuW
Cm+vHMrH1GoO1oNwQTvqOKYdsIAu4E4DT8nor/zfmop+v3cQyq2xrDtv0EY2qrOly+tF37P96Lnk
0/dywbkWVPfmKASvR+vvNqAaP86Ouq7ShrSKFruYG0pu4n3VcDijZZxgjSprO13Ashq3GGNAi26n
H5thF6XC+fyVvQf1Rmcg5yRtXuBL10e2ma3aD/LR90kFhMttkKGQZAQpHuvxKV/B7YzomRGAMM95
HnTtsbeniMqlaBjKUQK0PpzrXFV5YIjb4yjF9QzyYGg3iaEpFxvZ2NtJwbuvxeHkVMY8sSsjt5MA
72lMT8AOEIq3IGVOaXjmFGKE0X0sX3H8lwxxH+jXNXsAUnrgoKKS7IU6kSQop9bxAhgpDH92cf7c
HyhBJmvERIXMblsean5dLYEERE1o5WK2qtXx6IYHSP3qkWplLMSH6Adt8OS13priQVEIvOVHuZOA
blVYEp1E/18CFDz5CTKiB45Qk3q+DkbgFwvnbnL1qTgW4Rz07DDNvFIfDblUlUju9Yssfwor7ksM
fgR3RGKV6Ba7lnronzqFgQtlfL69lDmalAxxmEkcaqVbdOrzuowxzUnPtyl+HWI6OdtPH3JKXGK+
5xs/5Vjw1SyN34cMcb3hYJd7rkW6UMEVO5CLUPO/jXrCBesDHiKxrjRFnJxnuERvCjjZVCaRFn63
Nu3uCG9aa/kDyUCP1MctLtyeILaiLrHIicHJEEw9LUz35UhYS16WgxCoQFqroKFpeGlNXR+nH1Za
TFwrIJx2s0HHBQPlVAfaKo3Yu2zR2q6SQOuvIrxD2EdxhHbKYQwHob6zDBkNFYHGEpWnud1s9iX/
3KGTZaXLVgfvBxOS5HHDBw47LizmvMe47mvRLZaH23sIUpBy57exmBPz4YN8E5Xmi4Bp0eTwDhFW
vL0t2g6W/lWp58n0MTc0qbH2giuM/QfiE54pxTS5ZE85MmrkS0QJT/VgW197lD7WlOwDKNvU3SHf
hOUNOIU9evMB686zf9rM2EEtMTTfMsqE8AHSBugBbNXzZEdur2D/vgxtZAefxD9+URLsBfbiDwem
8A0K09e+CfhEaBb22Ms7Wfogz/pYB+i9H6VmNH6aW1DFKNlA2XpOUjY31lrUmV8/hL25kQ8qQ63k
JEGge2+wGQQzvrxNyQRIdD4l1LUkxehyEXdsiaFPMU0evJdc42SCPaS0+T2MxN/YurXt0Y+U0sP1
XHrhW8YMm7/eHH7bd8js1mC6Dl/z7XibYn1CX/JrCFmH7qR9XD+slnE6MOen9z0CXtr9OqJ2cdvk
KH2sk0Pk3EgpR0Q3MX2c8/FzzkJgsfAH81nZmFQT7hQ9CGIZUjOJxuu8XGSJbEvm928ih2o5WB3s
SlcFKQuQV6kjJNHsu1nS2QLmc+kx0HLG6G8tEldl0R6RCbOITVk/0dUyTex5cgwbncUXC8psdWUo
E50LIYSess8c8CfTvA9zWx5OPv5/25PFLktjt4Cx8Y16sn7eEwz/PeNuTyirIHZIwc2k/h980Wam
hppqsk9OAqNdS1eMfWKk0ToPqkoyUrW5HK8BRGDFIfNZhAEasWM+TlIzMuBRBPvQPNIpCXZIPdIN
1ehdhngOUOdPxggpmbFkPKy+NrZAw6cak8OLA+Z6bB9WNkwlYvDPADv41LbqsAKyupF8xG1XivIP
dckQmu6XIGBpYWuYheguxIz8sqF7py8o6rxEbjoxVFOgnPzU5jLmFsf/1D2qSZAqkmzlO2Y71NU5
XwA9PSv41KGTt4cfLOep71hb/ibPDYNHJnQDMieJalWhZZJhwZW06akHxPfPlV7rSUz4Iqk71hbA
Vz1UyaJQAfONSzxWKpQNl7zxguneTes6gCMURxbVvfIbKQha9KDrteAe6zZtVG5rfjnqukqkN7h5
y5ynTDTf625c9x6PXJfVaLKcCY7KRsOWDEUWQEKNcWKbtoT8ssEXKPDqlYjGfv3N2YWC9KDpq704
8FqG8F3YKMo9b60VqJ0tD56vkCSeE83pGnWk0TMuQ77Efv+p3LaZjhw8pHZ6PCDIQIVGTOSRYHpT
/IU6VogqzefQEInzKnikf1SDx1iqfzY1PSa2dHB/06WePu44jLg8TzDKDB+XYIR4iK23L4Z5wjss
V4NRVQEtAvBs0E08ph7w2m2VyyGugzB4BK1ablHXd3wG1WJvTWJAlbe3UnV8FcqTSwBwODAXoCGX
WP+4lbOA8SMzUt6EA7CeAJ5r09ixXZC8cnKr6loHcGQ25zUlhpCzFSmbt+5WHm6YFiQW8ugxhb5d
eNI2b3vTMIsgxsdqMgX5fScA90V2sjxVE43Zh8kwxzscRo6OYhnR1Rekz5N8x4ULD0m3Fr6Puf7q
mXGGP4eGlBsCgcsQ8LdqWtrIqpOY21jnDv0ARFxbKE3dFPl1ump13wiL3VxRJwnGSymzL2ekYGZu
eJkc4V76X6u8cLFMAne1447/KTRPijuiqSotot5e3BuTEB4rI/9A4m2G7K+SUIZs8CECmpoA8US1
45B2UXbVA2cy8rH9F16pu6jcl1+yIZNIyvf/WdCQdoWnd2giREhRPVi7gbI9HAtOsH+Aa5F1PqN0
P78QmlHh3HoaDeu9pvVEjjeC0Q/lJnz0A/H54lcN8fIiQXTwmKhcTr5YtQEU7bQ+0WXsruY3kdP7
jRf5AW4o+azA+xOB7oVvv6f3h0m7SZsIFp8KEaEyeZmUu0lCCkgzKJbJz5KLQdz3x7UhVhb0Zg2D
G840dNGDRVHAnqrO+c1QYSZPHVnWS69+LK7UZX7Ab97RglplYeSv8vgfDdFZtPpdYwaW6fkMZ6F4
H0qx74aH3/LwW0JYpNiBvDLkhpXNqA99aIEp0FfAekC7BLmvN8vvD7+TEW4st2aX4d1htslUVO0A
3NunECVQC6OjxNNIJgAFBYgSp4R9r79WMYuhwKiFGa6l565dzuHQW5C1saE1h3wrgmk6dyH6/i0p
M4QRyMQ5cqqqotvQ2+/APhf/lLqv5KyodQi7GNbwApZlP1z/Irey7pTX8O5RlAo53osF1641pUkr
Kaok01QTwjgGIpny+XQCcDiE2MKFRl3tmsUxb3NI4Y4IAjFPmAtmc+qjpqbAmKqeiZh1bflBugFC
X+NL7yCaoy9FD9buWH9Dt/akn82LoT6bsugcUHFMVehTHUGdIMOavXUTNfEhNdV3qipiRL6lQtcl
POArD7s9Kw4f8av/+Qk+UcccOoB48cyBRW7e9In9NAGbUK+F1oU74Qgi/o/KFh9UObdtrZS418S+
/0GRcvujHPhYfFB6a1/2Q0f8RNpQr5ycHt/qf/jd/n9jeB9ukM0/jPiHpyDHeFgfB9kw2nI5m8pJ
27B8SkK29G9Ae0xSPiJxuMRSKCO/FoHlDu51VyAg0Xb/uZkGl+alXbdHjMSjQBl7/3Ca7FgrdxpQ
I7IWPT3rgATqYfDcyWfxyCmS+Jv7Ir7jnIMvzC3UoVUjvGd0FxgU34L6P35GCDIqHpVGYNmOdKms
2SA4yz6ialzr0IUdGV6Z3wpWr6SY7srqODgCtBRQQXhDuSCoBhm0vXhEPHWCa88bZamicRdBNlCD
B/cfafxkfrf6bDqmqsm5qNNMyy7I2nF3W0QrZtfBbLoRiXYv7+Lg4XP13jA2lFLAtMb88er1Awj+
9XtnR21pJ0FnH3ttVwpIR8BDl5RsIBNCtwm54v6uLwDzI0ifxjYAPvT1Rdm8se3zG01M95zjnt5E
I4sbfEHLh6PrWzpFHosj/YFKpnToxY3w2woOCTPsneQHq4OU0WVNRcC64EshS7tVIh7OVG9164fA
xU4rGo2W+1HPNbfw3Z67GuitpB+C9J6f3sdXHP/oluH0blW9gNbT43CgX7/WRAaO12lJq6AgKglo
/j0r+icRtSxxYiEEFKPFwtwhBSS8ZWv+ia9EQf+EavrDDxYaPO5MEi2OJZl1O74gJ6hWNEbq7ZBO
gnjgnQxeWxvSFyZtEZgmSLGhLHaFZe32WhtRmLx51Rvfe2VMlvl5Rq5VEPOM1XFGA0HStGr3Rr+Z
25yordgknvTowlDq4zmtpK+ZFV6Qf93WiNHM9lc5GvBdC6ZHrj7//0Bczvk5GoI9hpJKV/3VQO4r
v5LAuplzdU3PW610z5NL2HHUk0VY7rdGJDxhQGsaW7+lpgklDRk816b1GSlgM2hWhBx7w0GedS5t
5+IJ0gCaLQgTvbge8B9IanjgOOGaugbFHR3WslXGRl9kiuiUbpk0Tw8cRr4NirasBu8rrCJcA1KG
/kB5A2iFvh7/A9aDAnUZgUSNLvnQnxGml2Gpw8VQHWt5YlFh8GSra958PM4006iGVBL9rkM+atVt
gOwyIwSEgJUD/9FZRelyCRefHqiCp7ZVQLykHk+6x36HJ2w913nOp2gXpn2nHxutUgMrFTjacITX
yWqr+uhtRYNIRO+orL8Vj70+iGyHJXvj4Quqroz5TpkRGB0czHuwSDlIhidzbJSg33V+9bytiziA
rxWDh6Xoi42EwtyQlRT1q/58Co3lvjvS5HBGC6Hzx3qs2/CgheT2lKhOaNUtx4oonghg3xmCD/Ow
MoBfzzkBxaqbCHkqJuJzaai/mnBlE3+zV6Vxu+FgtidCOpcwpYXHB67UohdcqMiWLd3aEz7a37mx
PdwFSg3npWC6O2eDMxVTWipXy8fw1VdetYxgEPBHi08K0I02yJ7TgOUBI6BuzHJ1a0MIWPUIlMCw
cDBfdYFEuyQxNjcxAJEgHZvTwEm5BlCI/v7yimqCEG52BlCkqi+y5GUzj6GAWRJaCzPqbRv+I3vG
ZPKTo0HasJYlDUe05H49Ha0Cdn6XYrVBzahe5ku21JyDPO3UfUIro6WanYTFWePIBLUeEnUnxu4O
LZbJCWg4raJvZRYVDfdyIqd6zKXucNviHo/0lSh6z15Qzr+/1VkJb3o+B2EpKoiRUubdEErKadTr
zQzyJBIyM58NneXaWMECUpB3e6QH/0BdX8XSgEZjDg5/Up58qDVHwK0EIZTHbSoAHEI8+rp7IUF7
OGPzWSy0dA7vfx60uqT2YL8ZTBPwmbbPRJJ897hfL9uSocth/eqat3EwSlB1Fo7eNYtFgcE0Y8Kc
QFFHZD4bHKkbutaGGvwXZp+HwaF5sUCCJp5sTGlsonYfdPojRfOUuMXl0qbbCR2o2A93dVKLepCR
IsmOL49NmHhbbfjnpECGEExy2Pe39KWHhOOPG0j4f/pbcMyb9AnfeTYgULaNQm1j3te8UhTWQO0E
kfyAsiG8ysbnFs3ClOsmRWtt1lzeZFODT32Yu4ybXIFgflvuFQXsChPMftrN2hAmxqnGjXHXG436
4Nm7T2pVr3Pnn8JjGfH5oJesNDccBUXSi8t3NZt8RQSoXX8mhtzuUcIzf79k+0tDbOdp4XoqWK4Y
+4YE5eNpxiwenzoKTwh0Do8ZtoovhdYTFzbjZoy/N0iu88V82nyYYF1K6+RawJsTvkQbusbdu3hW
78RpVV+GqaOOcY/12DV1nN6qM2+mdvlr3jzo/7i/+hmOE1JL33b6HIJLv7fjKsBn6tPDhBv9f+dK
hTJ7U4juTSsJcu1XD1y5wesezZjkN5pqnr/D8XR/4m+RhMaYcILl5QFniOBLTEilAmj367/Yz5Iz
rtqDFUzm6bIXRBnBZ606CZoc/M4sTaL8oHcdqo5nf9ISrr+ZXlTU/F92ZuT40WUIucwPWiG3b7wh
0xrEnJlQoL+zTuVcxPTQrfEaDcyESKDP3lcPxt1GreFJrz6fM8R1ssmaAH1jz+O7EfQvIVSpngQK
rIqWMONNd9iLz6WmaahRL4M4F0oZA8VbNviCZ+e9FH7NVqlA3gJzN9rllvtju1YHs6/+jSUGI/zM
OnK5Ebl4GQ9AvPA+KGaYAAgEU67g/wpSBXeWnC8RXW835zWe6OsOf0yCDIJW7zInU5Y1FYlXWXL+
UZZBU6ELwG+1rh9JlU5jLLNxOCCwqGEk7RuAet07WiUDeyoRiAxK3gJO35X97TUOlJNtO1DLFn0x
WaTOJGhMkWVOFeoKj5FSdGsUAvvT7CbexUZYHc/IRH+Ks2RMEY6p6y3+QFo4MTNqPznVhfUBEgmo
QH49uacSXOZtdm/ibHWRIRP2VpgCEGtTH6kaMKhBKE2o7KiQQcxOS72da/OYazR+urAsyv3qFAfH
+9czH/ow+OB8DQpUGel6V4YOWtR6GTD3Pxf5Bk6KCd2x4ROPidjFKgALN+j4eHqxQfaNI0gPLcmB
hnn1xq2O7A2R5bjzBqlcsl0ul4WTFeRxr2x2touCWkDY9AZtWgPsuKTm0zCb+UNSA3ELxsnSZmNi
8z2X0M0+w7PpxpRfAp0Fm3xptA6KD/f5jsOiX88ejhxLPWOS2z+JUYyjBnp/paStC/+wTJlglYee
2o+mhBWfIOdv8p9jUB69h/NaIi7ZXVJxhq2d2BYJ5IVgi6IuG2cgkFdwlD+TckbobWWyzQUPeZol
I3AW3V0QRzylvVyDYfQnEM28SJBwNvobBUw2jQ14qztRHQb8dLRwhi8sNQKFWwLU1TLHxZ3NUGoD
mKFHeLAJzt7gGlPbQ1bOAA9koMwZZ0O3uG/6hcL7L60lFXFeFvUwhGLBHX1a32QlcGiEuwPiaaPS
z8uhCX+TrdlcHvXUbjBWdafe8gVX+dUl25+Zk2HXtYv2URY/OWgvQizK2d3huvkK3vuKfsI+PDIi
4yGvQjiwXyQTimBmWS0TJ6Fy+Sa15PUgzx1tpff0sDnh6H2dJZp0H8IqjT6BH8eXOd6w2A36Gj5K
8/l29NgrO44EtXT9twOUWi2ME+By3aUU76qC47dc7L6caY8ZadHTBIoQgHIuLREH5X9+o0YyfW1p
bA3eX1ikLnSLeYQODgeBQ28QEw82/cgGn45w+zNTskzXlyOuRFxiX2RTThkxggkY3B6AifL7GPAL
b3/lfbPw6a/Pr+yNM6CKAvpZebQwn93nRfglDVyacPLOG5XQD7AU8wD8DZe//0cuN0rUVEGaZY+G
lMPDU5f+nj5E1Ag8XUt7WJ3smXj58Cu6ABIVRpMDO80VWRwnRgVao3xQME242L5s541jiDKxyhGl
L8nn38Xh3uqF6wWNH5kDP+41wi2H3w0jasZAcG4nB8Bmsw5bVUtpE3fnHXTwawtWF8sbLKVv0dRp
E7Qdvkgr8+JPpkwgh9B7RndLs6GpG06R6YDKXfarTz1PgxYqkVo4PkNt+KDiOS1NJK84idASsDPb
R5JVNETKt2LcJmMVGcOWgzZAY2D6lx+09xug/x/PDsdu79JL+0ndEC8LoaAzV5xqI7FaAalKboaN
pReh3Evc/cBniCgwcI+yT68+/obKGOYNXVPCVLJUMnxwr+6eSOEXz/Jx1kjeiPwHOMn9uhEOyeaH
oijSQojPeLZJsT3QwKB4BZ59rs3+Bfb3q5zHow2XojzcBu40Q7STZuZai25ELc/RYkpJEmIZCnVJ
s5ijl6jR8OKS01YzftdKXMgoiBxYSyZ5TGNOWDl7/sy6JerF6ZY4Pkwflh0JwOAwBA7y7y2p+bTV
LKrvYx9zwHif++scUOwQuV2P5XkcIw+wA/Q4SR/dzEHBg5Imk+mY7RcvW1dSlcjyRazPMgJMy6We
jk11gwiEIlhS30u8owmyxde2vCnW/qQi1u2xdql9E5pIQXxc7bG3+L7jlUjKcehn3pWMZojp1Gnw
kfNJRfg62x+dVIFvcCO5UGrFaGwv3wb31Z4Y8/IHO53d33/TlPHa7w9r+lW2P9c9pR0elz3YsxLw
jW4rFYPQiDpuFHqcgiEtbXYebkPEXfSDSoSYFoIk47Xa1e37v0aUuE9uJiJ54/qsnvLpucCc6qxy
mxVfQhENnrceRzJVRuqxXh8GUd+7Ilgz1Bui+xT7VP551B4K0QqnMskNc1Oo7jxNE5UwU+3ktma0
LZgjBcpT2ghzjhMDB8A0SlMPoff6ThT9retxF39Qlmt6XhmEJyNJ6MokZpITjaavsJF58sI/ds1Q
KneybkqQ3e0U6/xNB9Lab/rK/Z94ov+spYEY1ZMom03dxU3RfhG4aTR7wgfxtCZH2+zq74rk3Qrs
AuSZse9wYcD/QDVBc97uk39HssyMuX75sl7FVY/y1U2POA8NdLFSvu+nappN2KpNoOwl2FzRXn4Z
w/Ly0X11Sb5Ml3zih9h8aEE7WZJpu6Dny9NoH/adSEJMVlnbi6QhgGj7T3veFdqRyzWhPk4/3ECY
6+Cmt3tWJ4ElYn0wkZoFBp1FBK5/19Id4pHQD01JS8bmqjwYo4gG1CUXlJpTxYea8dJWR9w2io5B
MnV8VgEMe98k9bocyNeOXeSMEepCBKR4tzDjc4vCLVITyG5pwwYQW3IX60ScMPGVgYTtYp+Hz1k4
+KINYuyUsN7MOuVoOI6yfZTmOZ3nGaEBgXqyOqsBMzCy/NBiFO7jfChurBBN8xr1Uu8gqHhSVTTV
JrP7sNbVgjHgTLhmVKBA+bzQBzuK6O1ykuj2bGH7DAOMZL4ZVqIQDClE+hTr3bno/YKUxe6dt8Oh
bia4y9NXLoJYe9AeuvJFYArpnRb5L0KNa4UYjjRa3xSkWNvXJ1sDMNKL0bgvJ6tDUHQx6cEBQJSX
nZoW+7jC3UNtIM77Mcsy+eAeUAln6hvAXwa4lkAyDXNiLFjZbqgQ77+ZNYNs44RVCFCl6zAaQyPh
9JyJmumU6wU+KHNV6jvG1XBiWre/BjDWHViXA7gk/vrHekIwxWrC83MV2f/JwEWuCkX9YU/JXZ/O
deQ1ppryUImvQJ0H4msT7O5foQsy1huiSWTE3Y9KnhLNinuRoqspJWe0RvlRtM6zgbTf5C4+pAiH
s4TdN6aX0qGUAUuTwPVG5sxsMsiGpKtMuayhVMdIVDtH+0xLoqq2nMw+mVJzZjaSI5ms1w+RmuOZ
X6BTKvRzNwF88dhbCmjtln0IV4/lX/uGQGtN7glFLl0n/EGoq0R5nUcsMtjq0Py0/1b6xZmN2Q8r
zAsS5Jg/Fo2rMAFhRyTeoWxCq5OKb++Bg503SPSFjjtgMBqJg6Dusgw6/uSbidkWRJLC2R4YD0HJ
EIQaPk9YmrvxXoZ81NqXeeVoaCyZ5RpPKKQCpK63dHMMR/xdl57SBJkMOqQxXN1UMMj4+fqujJ8h
P0oQheBdzUXfz+G6HtMB48oNHncFYZhgNMbeHsECXKEJ9CZxWt+z3N0ctPQiBPTPlOX5/bDhmKhd
RTSA0rVFCnwaFZnExm/X8p+Zux854hCC0ag1OFf2eUQC5JfLDugv25/3+4pXrjstX/wvbUkTFo1H
yMgENoX470lh5A8Hsmih3W2eaDUxjDlL2JIITUbChatwugZQ5XnoQrWyOukP4AmxfiEY+eUVsPZO
H4ZMcoibMo1x0CzyUxx+Wq7CBg8ohlLkKXewswpKstmlvhv6lv2aGElaOz3aWnNrbpP0irM/zUeR
bQ9aYf7kG75EWGSLa4zxiFwbKhuhXs5rUyU4SGLvAe+DxEk8TqIix4ARpu4ploFAIYpXCTBUAg34
R/gAA59uajWgVU0q/5yPnE//tiDUCx8wmMBfNR+VNB3ccedmPicLNEGR7ZLqpE+/MKQqRgrpUtRV
JxTgrDOv+En8JaNbK5o56gatDTqZymWQ/EKUQQ0svFIISDNDzJ6bhsssWu06UJs5Gj+7wCEuTy+y
unARp3M1AT6rre5AVvWT3efSfrwxjQ6UgTPKyicBiEVGZkwOOmWnF1pQBLQ3v1W69UMdoGgj8GKI
7W9kTsfGxDVLgLqt7IgAk46g8KGrqC1sjSAPzJ5/O8eHIw/fSK+I8prnnXlwi6BK+eplUdumpbs5
BhNej6ZtJGevIrWhYxZ7oGPpb2Xpl62+sti6dBzDhLnkafZZE3ItXX6U5mObASndbHsGk1jfAEJD
jT15hdA+9fE02LZ8+GwIHRd3jQauu4w+fAqR1Px8VVwCMWM61t3sDvrmEMN/2UAuXkfibFG8Vp2O
1EPooCph9jnvqHa/Lh8ESX5R+vs32D4m3an5lGCr2R+VLmiKSOPTWFCPR6tZTsh+ZaiYH8jE7Pw7
bGN85nep6I6OZUc9Ud+QIm9HUV70h+kOSgyyErmwj5pRMAtw6ANO3sfz2NDhr1zQxpte4kqPeDGj
IwvPiO8ZJq23LgWtZ3MDMvvF0zPwvYQU9c/DT9zO48CDOoF3ESQEvkaISKSmevE9HWZTT04QHk7/
uB23p00kqUAa+aFvVG5XwDspQGZofXllAC4Xffe/IrEOK/yy3VtmArrxBIuuLmJF4FKUoxsSm1Ht
56NAdRMlH3iLhLcGfA62g8lP38DOZLihsHX9aRyPwl5El092gZkXDEA8N16tMnftNNuDo01ucFXv
itYoqrN6ot/pWMV0bcehlDaLG6bNOKkOGMP2W7b1+EGBuN6wboE8jlF+aGCrPxyZ3g3O04jx9kqu
P8xaiHfQv+izH96/TyH2mTwvyn+/N41BnSLfd8mSFvw8j8Y9i46fSLRSEbtileE2MyPFlWX/gG68
lz/wN7/NsgNy6b99NHNT1U5BK7jNZPPuC7RytiQa1O1az079zTu0nzJ5vRyvSlGsruteUwmBhVk3
0FCf6EBa972/Ea2V6zVcfi18qoG1bd6mw7udqx8FNmPgU7kc/zTo72Bm6tO7Ubd/hiw/AwmMf/7B
KaWNLiD409jxSRGrrFn1xbszpcttzKoE6C3950oDgYuUn9BkNC9r5pv+/ao5tDKaKzVQtuuC9/jF
nTVNKkBeoXMGoT3aMt4e/OK6woz9ZLe1Y2VwYmmphFD5n62BjJifq5V6MXPau7wkr0ajNTgVP29l
psSTMhbBBymumKkeoSVQcLla7rPbsVSmNUt5Un6C/6ph19yQtPv0NoclKUVkRxs+t7N9eVWcI3+e
04MHAGeIfCqusPbEo1wXhfKDjFzrxEgi2g3UWcDGreiEdiQKLmkkxqhBZNzLdSKXPOoKoy5WdOf6
UtKTe7nBbSz8ChJQR/4JzCWf2VM2h2KdYM5BRswTjuah1sc1D8kNI9884F2Zj6SsbVtivYgal77h
Z4ahR/rCVWN7jiW+Eq3jU2HonVTiAxQ1DvxXdyE5il8G6AUILHDWWj7hF20EPa+CsS1BPGuiw9r/
qWt/fQO4qA7uHvQCRXE0L34Qr0MqB4rQyMxorYSuxtd4WpfZRsgxjRYTFncMgF6nyKlSfYDeogaC
7cWHAKDLWsEPQrheSyP1VJHHdHfCpfOqsS+BalcF4XUjHjg4aGGy3njZ4+xtPScgobhK+ypeM49D
ra0Kxit5pPsxBrIADrhkaRhSs9M0YW5kl5RdsU5vT6FLU2vga3f8tshL2SGBT0u2vTCuTT4VnYVF
6B37pacVUKU7MyBpwb5dAXyYAA+E3SgKOOGizvPPxyosTbiUyvgY2NQBtfsQvlITontzt67xGfaK
ZLhMsPwL6JzGTH0Zl2mkKC8XUo6hVBWmOHC2QbXDKtbJZIXH53qO9LlS6K0YINoFhvD3SKTr2/pY
/gvGbgGX8Ru+4I+mimD92PI9OpeqRZSgVF0K3/G0UPhdHJ43Q5/gmJOLbXjCUmvT+TerHtqvrcut
D5scdVOPinhHvcysg5t0xSnQt5oQAJhJci9U2BK5v7HZlwVxFb8kgNzSA5jE2LXcrA93duCBqCRT
DvrrAmWtr4aBdXuwC/7STV8NHtpZtIez7U4DbDIUCdntjX/tjcH+Xi2Nc7IUbN13KQv+eb/Uj8Px
u7cDtg8rziasZRuMHuC3E1kKRv651v2xYsU8ajadU5tTZUTjLd93bLsAjSQxfc+1sMes2DjtZStu
AaOrYYzMsCR4NjaTT+mVuK8Ww9Ku6qs4bwBUG2SXLu/+bgBE1C1SYkxW66fJ+OFLE3KNDtztRTYh
OGBNXqmeJkMmgWN0qtMlVMPehUEc8N6Hn8g/w90w3BES120mJZPWGwHuPg58SdRNJmRlpJoT3IBh
kPNnxVJTCBe7rXPp28jADNcFvHQx5SuJlzgS9Dio1u817Be13V7UZVEp3jowxN9kbThMVL7M0obl
mr4n4RDQHk+VrTz2nD0sJ+EAG8peGXStyw+DdrqL2Q+S7DGjZimKvqiwmH9eJldvrM/Cg+3Ow32T
m/fkIKnkKzuaplNlQU/X0WBbmlCfqfj99btqQJi4DOrEehzaUnGHSWE3wO+T8azMikCSxrQPBF/Q
TB+FT7kxPgwhasPimANwlWzF2S/k4YwQZsQ4I8K27O6KPDJZs2GllxEYz4B3oIrR+jNuA5w4QXov
IFs9MYh90kHbk+rfvpzzozJk2rXPmpEPp3CWtyCidQiQFI85lqFy7UQbNFlfqDY9l8bGNIfxI42h
vNHjOLFfyRPK25KnRzMyqhwkTOgoUC4nNEPOtwiSdEvQYpveBYTUErzIBUyrFonb399sSIMe0fjd
Pqqt1tp0l2F7Sf9BbGhKjkMEughvs5aXyy+QF76cOPWiMllpqqOc6PUS+rKpG2F8wPuIzKCZdMLr
/F/XPLaCW06vqnaPt96EDhN8LQglaPqnSVRRFM4GAWkzpn0PI3M5/sDALqLMr5iFebOS/3i9dROu
8nwUMkJMU73mgOx3uK1+uJR0o9DDsH/McDvMS+t5Op6+gQe2nAnZNy7NKUaRY1K0llVgrQ+k4DiV
HEqfENL9L++Y5yw6+eDnbnt5jaDuBNdO2Vpd15UxEVsBMTeY5oQBHofRIQT9/vFrCcdvE/13bQhv
CK+OMGyrG/kwAsNZFY4SxrNG4I7C/xrnH1pjeR6Xo1JYKi9omTfaF07/I7+Fz1SdkNo0T/EBKsbe
gi7gU89KAexCeJ4+JPamZ7kwauzmUJmpjLZssDpW4vPTLQ326tRDmG5YkHS5QP+/vih+O4NqthHe
mnHZk8kF8zl8LP1wO2wlZrY+7KcAqACp1P51tW6ganwXU7vWp98guqyPRSwJJMN0H44hmC+6yrzY
sVg5Z8gVSeTDEkbtt7RA+WCVE89WsZaw/18V/KDEGKb0eqG/GwQPXsTWIZbCZLpFWUk37C9w0RCA
OSHHbCmZ9jXOavJWzYM9P+2y8RMFXHZXQ3mexO5pMKEx2KVTueSESn9CTL5nAX4JeUJ4g0weZAER
8EegSNyts51uLoBqm0EHmDkiOQc9gnxOFxyW38bxCvXZ7yKVItdXsuAbvOrPH0v4xcE4pG4qi7Lf
Ldof4rFo8EZ21oVc0tZCtU1nVY7nKDOc6RMyvGTxMoOuAIoszaDRowMVFKwch9TVIu4Mvwbt3iDU
MtkKN5E8e8A8FjTGYMRgSl7EhyM9A+oMFakb9viU0wsY/iPe2Xytxdj5XFR4y6xqxWHriyLLjPUD
yTeP0ohN+1p8pPU5PayR15yHJuM0D1Fnz9xPqenyRlDWBXfDaDjQslO9YJuJfdcdaGTvXUjnV+La
y9isv1/I2YsyfCuRytJ48KKyryNukU9e131DLhqLVLXxotDOeXmJqAv7yWIefjZoiZ/3bRBxuO3Q
143DWFzzccZlmQ/1gd/aAc0zHNdA8PPA/HdPORlSXDCYf7K7oC3AmiXaKrpLSG/M8WnK2CR8TiNz
BQq+tUvXElL2onRoWz6y4OZ7SM1nuqU/UbQHR3GqMCGqEY0ctdVzDebKcpucyTdfJFDAONxkf0OT
NJgyHYQ6E08HnUEspmUcJxqS2BY+LkbV7GpVuDYnUExGt/RXKBK+4IcVyBl/DsZjkvNY8q2MT6ac
GlVCVT74n5fmR8jPel+E0FqSxKxg79wZMzgoFWu9/Gphf04ysgBpLVAbT6dXer9JqnZw42Z2HzDx
56C7jL07mLCfHeqqo9GefphEduvgqx/x+fggLZaCNkbwnlg8aiPVw8QxjxAqKSo0thG5zNl0w1Hv
A8I5ydqxKzuYlCJXZ6v1LRFWK1QHI5Qf/oxPOrxtNQtC4/tnrD/dlAhjRli4EbGf/dnrZrp4WUb0
xIdySMPreI4W5pfZaO9we6lVp5hRuLKDMiykMQeKG3OoB8IVcM0F684+ckzJgGxNS2Eh/SudtvfI
r1F0O+NI4GjHZFySEtJYupK2/jytVFP4Js2Xv4tDt/ewz1sYxP8nHrhnXshCitln1yOpN7ED210C
H2r0UAExW689Uat8cfLjzytA6EuWTqfViqOiLx1v4g620WM49GV9/I6wb28siqfT4zNsfU7Fly8w
SfBN4yB4epUbh7DYeZC2A0z30d0Askibh17K5PloWnD/AlC+2ttJ6VC56+JG4nqUCZ7psHBCmP7Y
Te8KqNp9QZQDv8OJrVRLr++bBkW/haEZUpR1tvn2i8LQnrHmWGuJ7qAITI6tSYI5AaepjwkY2BD4
8TK+cQyFsLyqyBRkoeksmllSj15CoXdqCrUDL2C0rI+niZ6vHfsBc40XHjcHuk5s5tgXJlv/jSC5
yl4zwJJXutZ8Gt7PYbUkdPVrclF9AAsBkEL/WGqZrYGy0cY4D1BAF45ZrRDa8Dcbef5U9InYxa8O
RebBusS5loL19Q3JHADkeAeEPayOC9ZOQE+hiYT9OqjCQQ8Fd2OfekUDBelROWMsXpWtV3naAHej
s+2pBdhyCMy34lZhePSDJPhhsf3AkGzwNtoxBhXtQ4CNcr5lmaJHEyBdjkVBhKecd596mfiZhuji
DaMSX6LF52gYyAPz5dtYcimeyQ/+vJSmxIJSuBRtVgssCfX2d2LupCP3JCna0c9Tq9RHphGbW2jZ
GrwR2td0iaD/aaE/gRCMSq/67HqzMX+JvP5LoWR9v1W4sz7BJmLYcUM+cp/Vp1KWDbEcnZ3fexje
/NabuQCs/TlXs8Y/KCC+uuNJyznKV/z0xkEtx9O0BXSzQWAE3NgeXrZIeJP3xh6GBglmIK5KYUMi
zR6IB5FZ2EduWdG9mrQEcA2vDZM8BZc6NYeGzguomM4t+kAOXJa/b9iAilywKOMJSSgq/7j1PVZ3
bBwY86QfmPA4QWurIKOxQm6GTc54+mBGebJ2ev1H0kOaqWmW0IRQYNrQjchzDN1riFipMMBZQLx8
zOszNcRmetqjCsEvBTR4zbUpBop/Uc1bvHbaHBtYxazG0KSSs5SL+qbP8Cad4J4Ns0HwhIz4802R
aFf/1lMIxWokJTncqJTz/GeNFQXWWDVjEkcD3EUW5OeRcUSYh4bGlGdtdPqAbl7VBa43QiTYaqI5
WKYag9YnnFRXj+X7C+wPQvsFfH2vHNc0pJKgWlDpm8BuVem/lOktG1p35+/HKsRk3aAWVZ5MH0fm
JyALzGbAyLYkHr9Grc/JR+MheqetZ6jEBQGJMlkGuUxF84RVVbPPaAeLNrEqWbVZS6KBdyghck3U
NPOz8LU0cU3MRvAYQUQTVeoRaP6zu/w50NlLjMXxnuOUrgbNBy8pbc/tjz0i6cDh2ITLZz4wJCHt
6PBMIGmRsjVLDKUIkJXoSUG3YeB3cwQo3q7lucWFax6v5Svx4rlGqgwU0U1e7hHyRP9vR1YIthG8
J/CaadKzWcfI33a8tzLHN/BjBPYv8gT8Pzm4SWvf8BMbUD0pggfQoTaSTE/o0hVI+yqOpFBuIG1w
EOyG4jstFpf1JZBXPJpCJ40Ai5yM5ND7Z2LSHguQ0H8BewvM6UwUjJW/6iUYO86qAnNWXMA3EsZa
8A/e0+NtvT7vqIb6d5i+ZRkb7SqCvjwJV5tJDKdh59XW92ivCwulKuZWFvwxUD0QWOVepOJDeDMY
NZjMKx2+5q6294sBQsZrprL9YKg32cK5bx48gx3yT+m67gYEErdq1I4DYstDpeUc3PzuRqXrk8eQ
RG3oyN673ZggTcCNyPXXcdahb1jb3GBIOiziE1PJAsEeLJUjFoZATBr7gRmgoOvw75cBUcvjDVGx
T+snjK96Eeb8DtWbb7WKXe6kVpXV92wvVqqQIGqspXwq77BZ+ZQQKhc07LpCOEaYHKqqHsOaX+oq
r2g8MNcRqYKHus2B5o1GSm47EdQhsgF3Kx/2QEMRBB65n2yT564Er+9qLCB9UA2Ioz39AkuLPW7u
q1HgSAhGZOKXnPlYc5qwelmCB+JVXwIrTfi+a8fIimGpwMHbsc1y3k5lHMEgG4inZ4ecwYz3WBUo
7OIngutqXMunz9CkTfkVoj3UIeBxTN3iPxa/2Rdq0OAhktySNgis0Ehpn57y6GNf7PblYdUHzw5P
E42nnXw1hvp1WE29C7ZUXwCbnxY289l/fkKvYUWwVcpnX3Vh8GIHrRGnqGXGGCyhvTfTia3AyaPg
uJZvM66aVeEp7BPnQ5d40hZYm/IhoTf/+ZMJICfUAdzZemE8JYV5GH2TYHET60Sdf70NNItwGPA0
YSfA2meXwZDwGmyHQP4XkvzS40FfQKQ68QAFMcvXgaa0QDlZjKtAGEVE2RTbjMpLdJABpypcXO9q
PusBlvcXBPareVtmlb4CmKOfXGIljLLbtZpAWEebRAVqXYVUQwU9WrHU2GAxXZZ8wi+aNoV6dmyl
h8tdXnqyCVRKlkoIR62NPRDUHlms1fFyYow7hin+f098GO6ALwUHGsVEUrfdQP0WZ9+cme3T83WL
fG9vRGVAxPvgjKxyBuvePaR2ge5ZDfH8XfeKhLFfLkAy+3IwYvWuG8ranalifO7tNW8nzwn/OiI+
JdE5irOYZfbFZJyE4Y1CNaGedsK4nBCjimh3GrkxcXK2m0BXvW6/XGnI2Ff5XehsnHZGJ2WuqeCw
KDYSCuSDeb5inzYBjPgGaf4CdpQstfPpInOkIkzsud6TCcMaH8Mcq4Vt7tyJKPo41iOzUu9IzKYr
y0cXNoGg1ZbmViYTwcqYftoqtPI9Fr3j4hi8FVP43jKN5px16Q8uugWwrjG0OHFVM5FMwweiAX/b
sQsHwVOWGP3PnmpNUqQGGlbMKu53KcjpDIpzTS1584P9PNZT4uw5d3tvgPRJI9uyubJnFX7ufk1+
+4ms3ZJbTXnkjAOrwN+Csg3RuVU13Hx15J8Dkvg6jzKDhQ57pWCEyFWx2IwFkCQ9ZPzfXb9lbeY3
IYfqozH1uwcmalHDC89VRt4LdBeWRf3CCD4wucpDOwUmHrrpGAC2Pz2uFWdIIiF4OO6+e2OZQ6vV
+/l1SK8x+swIAUVYHnRJ4J6fv6bulTDtthbOddSawDCbXA+rqWuAfLU4YMP8NLRrcw+M75BWog+I
GjId/a+AUoXU2aNtODuDa/XBcGMjU6+kC6dWotzMBDnIxkB1MOKVVe6LFFBLtsSyjltUvZfohFzF
VG+oAr+G8hhYzr1VOxEen9z+7ifCnsb9y8VqTJdxGrmu0BHW+F4dJRt4bubzp8OLnPHsEt0LHVvG
sJZZtcu0i+++Kxil9Ptzt/t46dB7W5x8MHYYHY9Vf9bJwPlp2ykF9tBmRJLRsWhdb8eJpcfFxx62
dAZzju6BFoNARffZstuQvGfcmHo3dkWRSnColr1aSLQ0EctL07YGtnYXUOMjLABiUOfeLWhyJgYj
LvgGGRKwEMvEOLrZ1VO5QZUZgUywlBcDH2mfa+cZmc2jfQ6LjXIWghigZbaseUQlKKE8vxNzoSiP
GnXT6rTVncI5Wb8sPCrOMshuLMNSQ/ntm9NUR1XjpOFeN530Wtz7lvCKbk17caDCqeisxxrFDDYe
soY0nx2KFVmstcjepiXd5jkMeuRlRcHMmfGTEX50V+fFQmr/AtxeLZV/tH0IG6u9apQYXf5Xd+vM
M25RxKzQVIJ3mY+KqKcnRtBlqr+RYnIERO6Yixw8Rm3LO9qqmtOwS7F8nzX44TYVQDvwx37BBaya
bwr4+qrUEYhwvvl8yt0YOVcV/9hkhlmzBE9niu/wEL+E74biELvHSEmRP3fas/5BtNOgSZSzc14j
4VjiE9nvN1rvoWzEM+kb8THfUMTpoGKlXEdEcmxyVX/0P6uDkOKrWTinZDnt37dGqdfNB4t1Si1Z
4cnQMY+yHq+ZDLrashoF+qVU9bVm9mi9m3QvRQdQkZ/7kskdbo9xdVwFrUXlKCtuWVmJoPPbh4MT
JeMTZXxXcKRZGJtjvnprmYPVSc6IbHJz27CXGILaoPCAQKIbFHE5TG9N2sDJ4LaQGri58csGOiz7
7EDHcA4YOogIJSbiWip8mrsJ04by7jBMnbXiVDsDb7uo75/4V0AdaX3D0KcRczvJ2Bz7ObEPFhAB
sNa0ieoglOm600iO8foYwsaFdZKpYQMXphGSMh6lYsKoPRlLQs2woaYof+lF1x/tZudWuz3ZBOf7
pDD0nlXXzAshhYZdyrTYRx8gI4jXwKoJQpidvogIa7hkxw57GTfwnp3e4bXv5yFHZY7r5065vn03
45ln35HsM+IwxJZWLK63VXoXkeDZxP6B9p/MToHi9m+3rp1hiHuEzXb8ayO7nZXH3q20zAXVr3wl
5qTBI5snFX9SoHxWHMwniEmcSzqkGAsbgU5x2jOEIzcxE9AAvi4OG/r0LQw3U3NY4rMpu2CR5Nta
USR4o/QKvh4dgUSZEeoQV6R1lSH/EO87iGVnhuarYcwJlD2oIiSDtbvYMeLvnIweJuSlTKLl5Xg/
j40sjUU7/qq18saOMJXBPPiGTZ9Km7fHP9gItnuTvt5f/Mbfpd5AKLAsqgIKTSLx1COcg9dM/Nv1
ilAdSwFusHKnyjzHdgX9uZXSTUr4BigSOTVqRfYXDgHg4DwJsXFK+7SBCF06vzHs2881RnLGlJMI
RmE0XIHEiF7xPj9cpLxggXPqi6XIU7clJcalcCrFT/oNw0p3EQun0XiGPn5GuwfUJK2fXJZqww80
cVjglEiUgLb/Y//xJgIr/D0vbyHNYoyMNGXDd13x5ieHUL/nWjHSAp+BpKnbu20lTfN1XTSP6pCz
EvhdOn+n8C0utJrUG4g4O/+9DxLiJdoO9xiOu2sH9h6FL1OdQC6pPl1jH7lzkUzBCzRTmDv4LiR1
oPFs6VlHmZFPMOxIuv4e9F5zt1C+0p7orT22WL1FGM2PeQJmnUGS9uawY7HsO04RKQeQhy4wdggr
VI3ll95CN9iA5MH4K9uh0KI7sqEbYxgKzz8ZAV1ssNsmQA1+bfDoR6YVj+te52QZILEv99RkpsmC
sE18AHcMvqOAmLOXfyi7mWwpCEqTs5SDEE+nEsm57J6L0+T3fwGnD0B2xNO5Wnt2/uE21VEbCGiU
Uvr/2jqo++dDmigneGSC7x2Nb2d4fgiPd3vPVRHqSOwKQuzLMlKfc6vAvSATMtOO+/MpW3iXcBXs
rqyoVXkbEEhrXjIMR6jVEmWToNCrShxGr2cOwRdp3yZ4G+cR/rj3VwxR3UGKT4fQ1JEckUh1P2PB
hRQUvXqF6vT3/OXAqm3nA8AuYcD2PZ4f8r45/MoswrccGJEa7kl/7KocKhdd1K6d6abZ+U+VnmpM
XSgZ9xvnhk+yk/ANM46KIfRRZ2vRk/ZaP5+pM6wDDdWvLqLoCJm4Ctc2qgLHEVcY1w30WY4HKHOh
DmaVNXrnJ3oZKZZE6fdMJ8z2ekp4Mxc6U8uKsqWkoKJM2vvOvwbJYFDGDEsX0zHK6wshGdruWrLf
ckFLayeEtoGQlTnseOkRDmY4koeK7qakB5HMYWC5sptGdIsWRgInuEYAnSypDyMZXbkXqsLCMcau
37DGWfzCIyBLcoFqoSQncojytbCu2+6HhsqW/mQmV7dEoyHJ+Z3kX82lGwkuKQfFnowW+cPT+Jno
cJZle8MnBvcM6jmThjXR6MVzBMGtckCykJ7S8j7k/rKIa8AlMwE6Wn9oNvZ5LybUVhnl37zZtxHN
uKiOw5gfnS4zXW29E9ej8+PT95Pxa6yEsgmKhVlOdL7jJbZ3gEFbY1AkAuhuJT3TzMizy2pYZvhl
ZZilnL4CIBExyQhSu5GLq4vI12777xV/qx28uDhnVHgKtEsS36FSfaauTV8MR5dDTnMkGAqgNBoy
/WjubHBEsvfT0QqV3yDz6w3Tvn1aQgcz+Fw3NCesanVqq8CWjdajrJBzRLtHkQmQwKc9GFS33DXn
othCiTZpsDxGjMC6m9sLYBDK5DoyZt1WChuy+AB+5cUl80tuGmPYb07VzB3PK0z7oZJAM9PYn0MD
5c9YDGyLLQvq2ng9hKD4lczLLki0JKtM9A9ProxokL7IKS0z0MPfHM9vvUEeqv8PLSWMJfyh4x+R
Pjwh5TjaDAsHrzerTQ2MJejfRc5rphi4raaYMldBHcjoJ7P5YkNfpPnhkvbIOmIPmQ8x7Tb1UiPP
zCmAjxgYnPwSoeP7Qog6KIEn1gM2xtengui0jazyiwFGqyhH+Upnp1RaNRTXIW2h4C/YyorNdidw
kGPAi6r68hhLixXzp6wwwdkss/s3WyCzEVt7V8cAh9SmcXo7ddkxLl5+OQsEMwdyeBtSUFR30ReO
ONfcKe/FU61IPtMe8Bi17FJE514s41T7UXD3qfzvqAQbEudJg5kQntKgQjn5WQVKol91o4nGM+Yi
9k81vUoxV/p0eTiqIZExxHvIuWK6P0sS3MVbwEy4rJSH/8xT6AafFnCswTDhue/ZdPU83N4Kd3NT
WrLP809qBlfalG8oTaZ9QQuE3TkS0bpnt+8bzbA+K2XfUV38yM2T8dcbmUHGTS9guxZNTICmU1n+
/W/Uf2gelEIutYsOVCIlvVJSQ9+tBIoDLRbn2LdEybxNb2pY3uBYmmMeZbUFy/jD5SPTZw5I8OYM
wRspuE+chajq2oHcK+WR0VbMQFvOusqoR09X8AinFAA0LUN8WmblRtxue5nLLudd1XWC6Jn2yXYF
1i+o2JpvgFYC5glH12QLZHlKvaWhC4yRV8NpVLVrpzmrT+ZwXDapV176Xm5E0KZwMWqesIIROs/a
Wnr1E8uCC/FsI7BhPrenMerKRjSkT9G40IuxqDvse7qW7nV6Y8Q3U/MPQUKWKupbsgxnXqlB49JY
9Gwjx8Zoyz28lAke/z+lAF2NJuL0poXCHoo157sm/1Ya7iTL5nJn8gsdn2im4GcEApvaYAFrz9xg
x/Y4VOdyGuf46WA4bBgTaEIgW7oznPQd4AFHHdZw+Fz40MBCrGUuZ+H6frSo0npy4jbreMxpDY5w
XiP/y/8Pf0h7I+0tu3Q9MYFr3aZph1XG/SorY72Sa5Y3EHriob5twtVMU3lnx/3Il/tgW59l96x7
H4BERYyCHtDD6L38+ZqSLjFG2mrYXbbmv5ceKqAGyb+8pjw3llXF/sFP4p5/1TaZBjRuUt1qn8Kk
xJ7YC7GiBSxUVShWnbU/4P4nNYBreMkhh7xoCQMGwQ5m38UTm4XjpgedNEPyKvRw4QxI9Hj2EiMR
DClP0o3ytDx+XpI3lFFqz2PvcDvGefNm3pcSthzXMV4ltY8Gua/a3Q9NC6SUDcsTkwQZuh5q+KER
RQ0DsWnHIe205e5dfPltX1ph3AQoHWnsxn2TDmWhWTrv0yujP+LeC5uYl9OQ3O86cdVclAaCC1Ru
6lCY2JFWXsf3cqeLm1efPAUgyZdYC6f/qoyu6p1qHlxCo/JWj/aLT6fjXjnmc1RKZ+RC5AhIejH+
Om92e/7baxHWrpEf2NS1emmcdYpSxGJhmYGt67VnBhmOc9mxNV2+rqEf49ULShhkUIHW8imYclx5
sR/8oq76Nbp8toy76FnE931I+eGTm/kcP9IPMkQ8ia1rn/aS5vopM5cUB5n1uNngyHe8XrYKzZ3p
T5mHrpVUce3Gmr7rgDRmXtX+GXTijUVwopzioMH6RaolnEwj/DF3r5qUYy1BZ15wKqHSbLTYABcz
NCTRgNco9E8srKutmWNdmKhu+h6SPQdhG3Ysupl5c4UpHccDQSBKxxTld8NZt9pWx+p2Wb3nhjZ3
70TW1aY/d/uF5T9io3398DDqG+NPW7kz54gsT5tBldXxpNqjus1W18BBT+WWTBim8atwpj18/Wxn
mhICWjM3sk9MbRkveeIqf7m+m/4CgY7PPOTTE5Ynw7wpJo/31UtzE/B76TTFDNfV+mnQvxITfhOd
BvXHEpL/Jicabn+lxcLlYXBV4elnFM8Qs3B7CmvZ2DmSrCrl47Mm0IBemLk9fkgNg78HXb5EgIJj
avLMWAW5C2cC8PNzcqQ14GIK6nJL+2cQIBK+T+BSIZqI8iaZiplaeS7kVGeqG40O27DEvrWVqHK7
qPoWa8BSfAitabaeHYQkfuW0tpa4TEOT++ntJsu9G3YxSAxkiyzp4dEAo23GGefjacmUM60jkIWj
3LzKCgXZT8u57aTNtg29al7wO7n3uI6RlFLY0F8u6zmNbB/T74mfBwEcygWeO/Nh2rEbTw5L3nik
2xd2uqXNt7udDWp3fWbPE9iTwPM2B3aluo/SY5U5rGGptZagtSE5dN73JohAZcK5cAY5Xc80dxFO
mobxFoxJUzh1wSXWQY8cBtVPAXaSUZRHuAfRBJPltXskm7Kqkd+KTTSamlXpi+RvPd9u0p6eDNt1
I/LbrmLpBT5Za4oeMaNiItVYCMMo7yMGE/k2uznScmLHo2ej/YGx+En+G/ybegBYNykXK5P+9z21
eHd0aY64SQKWs1Oiojg4IUbSqS4z84d3y2GItXOAInj7B/guWaz9/7RiwtJusBCYEd4w/UjWfF2w
QxTExscoDJYRJwvMQjqUBGUK/58RY857cez798jaoaw7wGQtGy3q+wG19LU26W3oG7z6eVZxzhGt
2zyFpfS6YZsdmFMmvc02K65Di7gjwQ/7PAG7lMFUW9Mtr1mNxjJr2BKjY0d21qxm5bY8MAMBjb83
3kQqn6vQL/fiBRdzXJ/hqVH4CZf5Oi3xL/jKM5mzbFvHbEjMj8829SSdpx0uGaJ6pWgWjLL8nQc2
5ITQjmYt7HT46cKe3l7XJfP2nTshQ0aAh8S8wJw+/S3Fbwn8PIbjNt2CiWZSXkUhYbLqYYmZog+x
XNMujyNknXsDTT0NqHbOd78eoMk9EwY7jvH4F6C+frOwfmRSIVVH+9bNqNpEltrL4oSM6Wshi3nK
RHSkK2wnpvG3pj4aXyG/p+y0NRNJbU/VUj3lSTPYZ619xni+pRATxL3Jh8HslBSeAMQ9MtrrLq4o
KM/GMzIZ7UwZC9FyZv7Ch7Iw/9nfqBf4SsEg0dqYrs4L5kApy2UQJ8M79XduTdIx3j+hruxJiUms
4bDi39X+gzhwcveSHfNECJwHz9KwKe450ANsikGGJSYBroa+EFdf4iOERw0d2GzsqVyyDC48RDz0
bMyskdGNwfgXirVw5T0PX8P9C4Tdnmt5Yq13pvw3URcUYym5OM9g+MFFrooN0QbmR7+0mXOs45Wt
rGbcqAJNhbzH/XReq+OtWEKuM8esOmjqfHNuG/akt37quDSYF38JBAx1doN9nDeLRzR9MckW+H9t
fJzQsaHH1fnlW2AxGxdxTK8/s9lmmVzWP4jt4Ix3lwsOdVWz5zL/xwxglDPsypyrt4Ko0p/m/p7Q
I5H54e9juRbjR04z2s8Nd0nIsByHiXWA2Ed5u5lrbnLmckJf4ENpbBOsO1EkXlxoTT2ne79I3NPn
lIa7rt9jYFuDm0Ic6TybGQ1wOZ6iXe6V58zJYrfdzH4MNOXa2B7hAg+gbGlTFCo9z1OKbuWqFSVT
3nruXtzafprvWWEE2wYhWY+lT84bldf62nyJErwO4PDrlGb3F67P9qpQ1ph/1J2OZOwo1rx4ng+D
jPRG8SuXKsfuhGgmx2D5U1qsBIZuTS0gIlPtRLMVJ3VmriNI5oDkqwKkE4narWgmUHqRrb6sT4Rl
2Q0FofluI9rloxtl7SAHgiolb5fzn3qDlUvIw7Qzi1cuded0iRRS6u1MJ5PdE/mjNolYFNdHALDw
OtbR+qAuJmYl8qwL/7qgwZcdI87cQN3tetbYjYy1l1Re21J5GdGL06Mgz460CP056btJtbXqyhO2
RZ3OnJH1vBT9FiKPAicRr/3hgTxe9Cv1uWIPVpzPwLjMugv6kd5HQ+yZYJFGkrXsiiXqQ0vy2/E8
UZLMImtXoxhpmj+LddBqpQ48uE66IdrFGmnwQA/bokaDJ63Ql+6mJq7GZCaVB5maUnX00DWeUYUO
3hLJsH0SxZWiS63D1OmOk/D5qIASL+o0h/n1HFL/xsDxZTb4M9VtNwvb8wwC9PwunDQg+voUht//
O8cdrVbLPbgt8iB/CkM4ic9C1lEsyOOHJ+MhsfYCIodWbottE1GeZKZBFVRPojcje37BxE2QdWVD
awFVxfXmgXvZpCC12zIQtbYCYzHdd+3E7z7jHRWUureXf9SbDI+X+sO/r5qFLmU+rpbX4zK1T8BA
azc8OE7J0YgGDb/RVw834qAZWfGWXc6YnsJgeqXR+/58StS361iB5AyR+6Hq1mjAoeiL7Lkfv/1D
thkmr+DHebsqN0Io3omgNw7+QnIAoQqk42SUboec1e0oaFv7BCka5zNXfTaJpkd2HXunNYsYFVIp
sSDlnEJoZqruLn5Ch4kYng9mB8z9j9nqFUCp9CfTflJxyGpGgj/5WKsFxM50UgBemWPSdkunrL0j
DQaja2LlRVBPpxwDLBUW1cprQqS0Cakd/T1QiGPRorXBIimK1wZMhMeJvCj4imUnhz61aYJMZ3AL
W4YV3UrzPzAezchcaPlXZ8h38fEaelBkckuNpwRRX8GrLGUAOfIV4koZiqR8tuUqTILf221pKeu3
e3XKkMV91w/1v8A+Z1+rnDnjz4IkaHDby/kWZIr7d9z6vxMNhy/IyFEARL63hrWvgi+LmT7HkSiV
GwlSDBkr9p+uEy7dVkLZCTNGQE4Mfr1RJXX5bsaCh72ViCVXO/F0COhOk8mYCRJVwIWcRb78oqEB
wHSXQn3rGRo2OwTbOxCHmHYYzr4k7+bhc9Dlt+JHDnA9zTuzqGaA+u6sJIJ8e9Gg9KYV0XKGU/w4
BQfdQ7UEl1erJPHB9aOaH+6BUNAvZa0lhaQMfd/V0+LQ4p6NKC/seae8If3zYYPbU4xKAqQPLLw8
EjiMb+9Vbc44MVgzY+e+ofQhfpG+v88Z3PwOmSAVz4eQ60RucllSui546DaxLNrQZ8LUOURAkgYa
pd7C/bpTHQhF7I4eRhByoFIB2eFsodKQaZg5HMRa14P6BSZWXQ/6SAZIas8iFZw3ipfMorf8Uu44
adcnW+hUatxKZaokx/MKEqccLrv8qKcBDFZpbTlMXa23VcGA3s4RzeSZ7hhwa2FRCqe1ZGYeclsY
lm8QYRn3DKnDl8cUtmQZu/a7RAjkGtp6lVz+vEKTXHltj30J8E7yHMIgufDdQ7PdCOQMjPEvlVMA
sykfZKUmbZDmdfpV6Fajm5k2S0LXnIlucutGZH5ubTsHssRYtLASHD2m3LmRqLr3GkQDNgtAYWZx
/IuwR1pzWUBjsZxCJ6CECyNypShVas4wVtNBTLKo2DpomW0eHbBBfjQWFUZ3i86UaqtXHMsN5vym
2mpCPr0TWufnN45RWNITcCMzBcFWYy+rtSi2gGY67UcyZtL1grQmKhvfzYgUjs+KvkmMJPMcGaso
YvATdOtYNTES+3+Vui/zBCVME9SSxPDjl38QUcA6rfoHM6RTZRRCg1UgKuHL2BNS6MKTapWkg169
c+nKjakHXwTbgkbOxh+13JJ69U1mw3yHpmqfIEozwXeq/03/Pvk97M+WbgEhaUMnM8I69ZeAkNgp
4EllqFfNvEbP3ps+u9EAOBatjX/jxaIk/umaRsR7IY4FG9r+QZZbj+UQGKk0/pLjJrXP3jQ/K3km
fBMhHHFRir6gMl1zPsT+jyMvqjfw5VEvakNYZ3Uu3dJgSw7oQWt4ssmPVy1pA5o8fA0WNo3Ei0IZ
TSNgFr/v2SUyFhP5BEgOKs3P+/RqGPlTRavzq4yPFXrG7Rl1aFLuafC6EF22Q1/2vSzUjwVWL8pQ
laKH+myV0JsJtbhF/cyFp8V5yNU6/HmONoh3oaIME8EoMiSVncr6Tfhnk2z3BKBzgk6LNNaDnG1a
oY1RoZHMO4kFto1zIHpkzz4iHAOn9tKtNZbUDR5I1bImjmiV/gTh8N64UiPcVGZ0PXXPHzkO77nh
Xe181A6LQ6MxRi1iOVAWyae84fiCoWIpd/9hEtYGoBLm4D6NXmSj50wESejIJMtJ5zRVasUddFi1
ovc0euDq56bbK1GrGseykvxhktxpy/wPiZEm6MruYP8EfY1nHuuykXNwI4S8DioYzfeiQyMeIuoC
uoDuIXIsF+UPQtejaD0XCbHav23bDWeWciJ594C3/KyTp8KtccY4OweAX/+ILHeLI66sIEMNFyFO
QYxvi6jBAyZre0oHopQjrLJDU5mtqnJ3oBznBEkAY8gTJKawUZdLQWnEdN5jPTB8BkGz6aoCKVDR
8ehANadCZZEjBjC5PfwKRTUiYMg/DxIwtTPkvbzqpfFcgt7L7Enj13b8zUU2+EsaQsQXginV2nUQ
Z0C08ZFm0JXCTNBtf7xeVqHJ66lCW4AWxQBn46XwgWG1hb2srkzFQruUWGTt9GGok0RIUlljFzs2
woS5B4cJ6ciacyc6nplxHB60AKBEYkL2//rQ+h/L3ai5DwvMb8S597K75Me/YnFmcqfK/Sun6qGT
/yl4Eh/ovFVpeG3hbEndkN0xPMj2g9O4ZKMjcsX24elSmEN061lsxsY9IktusoaOH+0CG+kwSNzI
IWDkgxvd+tyv6X8Ji+xlMgQeyRjslNewgj7FzCyilP38w+BxgqZkq/uK+rWkAMr/ZQz6WjrD7dM4
C4efFtYaWUMCqd2tcFG8lP0F/TNqmrvXAZvMkhichpt/mzukRKb0/WD1dUn/0uyHNCrt+gjfNTc5
C6XrP24WskFudMiFGn/2NZvFVN+BFxRrU1lWGNGrwIX+92yiNFbkhO2XjU+DIsJZq4lhNWBD9y1A
npJ+HOguCu+dH0H5fvZPnSVetWB6EiGnONTtJ68sgc6l3i1QSuwT3ym+RbZz61gLhfsCbOTHkZpJ
afgKLC77IfQkCCMBWewVO9pYydS1/dPDNPNBmG3kh7rbOeFjiyDsBiiglpwNrHaUaE58fA5Q4Dd8
0CVkXS3J26iZf37j8/HzZCRkVp0kd7DRAt6VGeY19kdO7gC41H/cBarlVmDkWveHedbyqOaDbG9R
7nmrrjThDqTqCiQcWVevzkEH5lU7MzgeB9hlq7Vm24ob1OTzC54i5YyBVf0jQfvO+PBKG/tLYTCb
s40LRiT1JET7OlNhzfXgjMNZnGSH4pw14KzIQaVPEUTxVFeS/KV0rqDJg7zFFi24EzSl8ZF+km4I
RrTUKezkbTVLLdYJdWTRAKq0s4XNtUCV1pIa33vExEM1NrqSQLfm19VDhjHARC5X5+GQ1NXygLX1
9ap9kp0NhqhhVxY37fo/0jW1883w8sAK8JLosFPxHnu/0Pc5HwDmtKjEbEj8VdkH/acFV+3XMW2v
A/1arZYEOT0CMJCA1tm3ELcDkU0o9lpMJCRMO4VC+yyJlhZ5OD/PMUAqfWjgOg99ObfzmgVsGNDj
FdM15ii3YnbLDvnwlcDqlZZle8b+HE+fXX+YkzVPRo2tlLedr47hs66Gs3ffbyiRFyk+gO9HoBYJ
2y2K9ghemUABaG29E3QKQDiD3AKnWAXwh0s86YSrz/c8eXh1hnf2G7Ul8b7rppmFgeS9/7eU78VP
MDSD7uSigqfxEe0E9rs2WqzXSUf1jYiptWmlw44d4bMu+JsE5dEdO51aheIttllBO3Nyg5mpNke4
zGM4ix+ceUn3Igpsde8/srfO5P/JmqTbFaIlJV2OEJM4FsJBWy4FtB7DNAaP2IEi9jQmEpkb6vlh
Fl0QCyE1U2pG5I4MGV2f/vq83+TSWSaTuzycySFOQkZJa1H6x+VCd9YU//is3IJtKCYyjdhiiclp
a0mWrbFfMYPxac+E0WY9uRjVIGMfTH6rWvZ4nBUZxp+mLYaxU9xukyj8P3LEFg/rFB29DrX2WGfg
d/M7O6JMmVGqFNZaXwE/vgbj72uDoTd6vgPSpcYtV7aBiMNHcDYTF7hBDN/5sJfypnFGD6l6zy9z
NqtMw4u6N72RQz0YLZOgPBZ9MiaMm/nGOobiJT+gRCbaRykJS/+f20qlppHilKbpLB0TlqVi3GKr
j8pufOESj51yt4lT+niYRyeug2pqWd0nkx3QLrX5Saa0nXme2fm/8XZDyIidksxmctHKwzmJ8Ee8
DiuWcooNtvq1CIBV6uLHPzfEN7S1z6JWVi+z0S534Y1WP/DWQUjqpFxZElQddXHhmEJS/rhOnafR
4pnu4MXyJ7zJvKdc4t29IQvFqacUl5FJTEhGuAW/HvPkRGKgEdLEHE17kfaIOsQAp1pD2X+OvAvi
EA7/7xNgXx/NZ/TRQOnrk7pjoFS32df0wMkDdCsi/Ze0BYecV3ypI0L6C+Lh/J2tP5rWDJ02MKOk
XdLaZA2nJkWVxt+PLRRhvoUpvzSJjoFzrhUhjhyo/bjmGJFYriZwllYzFls39KnI/dganT3fqww8
pMAddCdIrDC+ceVARFA29zwqC2fjU8OECt6lygEiTe9SAhD3ncW6Sz/QW/HciycVJp/T9USvu1q+
VcTzbbqkoOrZUo1fQeedw4Rhi+mSVtkKML+GSJ+FX8B+eEsfJ5voP/L6/Zk5WRbDMcKm0G7Z9IkP
4yvwJY4+BWxlrd83LuY4EgNqEMhD2S5PaCYWWv05zh5FEpjiLjMuzTckirdds+FVxSNBKHBzY+YL
xz+xa+WUYBLfgToHsqXxAjNbTnlF38vU2OzObSoE8xVBusxdtjHtdOJ+Bgpp4IeJo9qupfcfnfE5
zMlXFmnAarsS37TxEYbixFingzEou2FFJSrmLzEtd9VWV3+UHg2GFVJa7g9RF+au6ipZMyiHgCcr
wJcnKOAkjxrxiPsxftIJ+nGrNhJPRUDkJJXTtSGWsIRBcP3IedZ8UFM/EDGHTksr4Ot0cjdg+q2v
s/ZouRbVMdAFUG2OFEv208NjIix2y+cAHhAnVNKFkL4Dy0L3C1pYcyLHYuxueZrnGHy6PgHLtkbD
bayy/+DWvieb7+t0VZslwApYkIZgK1+hUWd4ciGcvtnuqGWvRU4ClfirIc2FmGQ7wbCA+k16KCy0
h2MXmxaOSZwRzZNiIbMVWoEOAP080LX8L46kaM0t4GiXTK+qr4IKVMva/A3h1KaDXUxLjhlbuvuk
xm0k+/6ldOtHA+9r8/serV9VJiGpEXwdpjySgnKI53GW8+AYdOaCnzNgEPExzXsXrt+lthP4Stp2
tQGyp3CwyMfxiRgkpWX/gs7MiAtw1btN8MgtGHHmZdDZj8zyX6e49qUK0lQeNUQzErhoFFrlscU7
68iB1SGTNAx+qXbC4ObdBzjP2OSJb9XdakW2W6oZIPJRm/BRuzqVpg+oJcAAz5KiBYl2NHAPOMH4
yrmW2dCae0jlksaVZL8LNayKml5+8HkMMBqkE2rQZJvv0OPKq0bXQ834MY2aHn/gCLoTr4IaICXS
O2X/Qs4gGEqg2XBfqN5JMBznvRY5HB+9qTt5Km9tnjpoRg4kQoegCadCqOntA/RYPgf2mGAouUwO
XSkB9EUZgClEeY1PuriVmOouEY8ONmLXfh8ZptXpYxX+fS/Ln1W3nBCYoZ/Yl8Vgqyze1iL8gr49
Em9okBr5NMyVMYJwzMd6eSWb9le+AgVwZ8D6ZAP8vi9uM/SV7rkwPoSbGwrNVbhkqhEeu/k4+u2w
sZIEPprQU9IcLGeFCkj01WeBv+Ezyin2XKN7SHvmvzEqCejEDmbYE4uOAad7l184/OtjDk4dD5/4
hjzxygp5MMleB2YFnWo8GvKXb+D8mSc81HZpEiwzsF3CqsTkKAvXKwpkKC4NX7980QFKNRZanIxx
+BLnslSUIovX3k4ssOG8eEvzFjbHdTxZYf3SOn/pRN+yczh+V1HP+jUzNibLUOLGTSyk1l0QaBop
hKH7fQbljOdxhwOKrFgRKJlzaQYgCI7F/Qx53P+hZEPLNb1Wvn8rKdy3xvdOt6wfRvugWXkGyZfy
dz5+QXOKiXTTERDyoRfRuhUT4vvOv/tRUBPyeTS9uhrPp+QqA/54FFN17zKjtVfg9To13M3yQr3V
7XFQg3AReQEge08meW35I6tM+pBA3dPa++3o4qIB/Sb7Ka5G0sMX7OX9h1XUwvrVuhadkC8TZYg9
gLij/T5VjVYCeiVtl3uaqWOyRCkTby10wMZW52p0MXNAyB6PQ0Shd9GYv/aUm44WasuBp7/Tf5U9
Ba/R5ViPrjHDk86f35J3NAki9OaFkZr6u8KiIoIaWsRiVg46zBdM04g/pjzDYZSV6hUS7EKrieUC
S9pAWSNrFp+oOShgXhq/u1M4r0ipWrhTop1bzWsBUzINzDl1VaJW7nFy404g7WYWgbPyvH+tev7l
Ru9thz+K1OGkFCHX4KbXfMzbc3HJ4LYCHiGzRDo5lYCtnGdYDsQpgeulCNAzTywnhED5veUssZKx
N8ntxKaOtqpMIXq0cLrgDp8o3xfUCBsRaDDvvt6KOfyxRhpxJdKMhBfE7ZqlcMVI14ipD/NH9Vq+
qxpwGBFQHQXtIt+rhnZdxj+gIP78/Rfsg9q3F0CRL0ZW9Ra+z1Ieer4duiKZEXa8Biv5hlDaxi5j
SHDhI5btLEUgflgyJocMfJNVUmeyGQmJewtzV4VvhbzB2sYHYu4Ts6alCYz8FBBNjoHO2SIPDooN
B9ayyDg7hQ5Ob3GvAgN6sTJ+7SiuCnM4VgJg7ra8w98vdSHAMk5SMV/aIxANLJSaafHxlhgrTAVg
ts5mabPEykwou2Zt7ZD1gN6u1LHJuzwf8yb+TshjLXh7q8lvIaiOnGxmz++d9DltErTNvzI+pfso
m2bggD8GL+jx9xuVVnueXLflHZIVGVHOeVeI0xF3I3SH7E14DZlIH5tAYDh5eDmmbeTQqDIhSuQT
C5ouAgEWBgHJgU7mNsk5QKk3bkjWuhYn0gz1AdjKcqa/5q9igKdn0P+YNWoTck6cK8zJHLjyeApn
6IbqACm4gL7wqmDK2EXpQVPodZk1kRRlvs8Ta7ABNdWsO3xZL488wdWfKB15Qv38sSGOrSvjkiwi
ql7U5ptRS9nKl182V927Q0eTqBzULhoAmQ0TK0q253WEccXYdrrdrbT118kpy8BCLhMwMico3x9w
L4UIn9A0XwDxJCvihdnCMriJzBO0F6Gx5WA00tOYXZX/r0UyyRsllcTxhwpVhAUXh96ErQx2ZiIy
jpp75lmMDFCmD9d0a4TyndRZ8QlOYfD44PLkDbor2OO5KqqokjdKLjxLDb6T+80i5RR4+1ZW/CDu
OIY6WUURzKmtyiwUC0hB8xi5JPnn9aqP1jRI2GmOItsSIW+c2zCDytb5XYTIqe3pbIwIA/o8xzCG
Ws/xvPC/THPhnKdHCmSMTdKKuEutLBQEOEC61weWDza+UlD730hqyierCt5cu7unMH9JN6l+RAm+
OuhyjrxEUlTbWTxLpD/mfHKBn/yaaPRG3T8FBHA36E2dcKpJBKMhCU5SCPXx3ZGZKwL1If0sLUjC
SJCFYM/1Zj7TbklvfaPc/lIRFY6sy4UmizhmS4HDwtobM+XfMj+BNKUwG1AUSXyqyqrH4+ZZDDnJ
fhffFAvA9+AT59pfZ9dbnHtJoPYMwZAuc1nM+gDfYamwmabdo1C/qt+nth91gbEcLMFZCwBHgsIA
y5tDsT2DhR2XdoKBaVlxFd6fsljC1zzXlYfnWbhIcwwfrC3UQz9mXv92JGgBpAKuEAb40RwBrJXD
rmNH9wklsZVgEMNItW+YEcs9YTsK/1fOKYySnlQ4qEhHDOgPy2xwvnK/8gAwWoOapOolHR7qj+7E
uH05ovxY4qQRtLOxfNWBw40ULrPE4gqV9SsiypCBBBuYwXvT1Obwifne2dawVUtGOI1x0b7kehrb
HeT7h08HHx1WPVeP03k311jPwMzWwfRh9XCT14C7s+VVAlXSBhQo9UfNryCIyCOLSM5WEPxAlgAe
U8BmzDDDomy/DaljIpCDywRtHWQcZz4y6wVqUkecB11/co8lBJG2ZueGFYSaPlTCQQCQ/yfgXLdD
NMCvVP6wMfNSvjZL4H+aunAECV0JZvAf7WWw1aU5KKMcp0FTh3ha4KnAxE3rDynCEWtNqZJhoM+G
SW5ta5i1gw4aCA76dbYGsgojJIabW1wBxF1tUCT3shsoAjp7A6WrG3PPZLjl0zPIOaf43lsrKJpm
Uf0vhqLddbkndTMypmEDdOn2nMUp2haa4df8GG4FwTkTdbgCFI7lURO8zssfPPppvPv5ujYup+IW
JIYG/IffZFMJ2R9tWybrjSGFGLiiPFew6B70MK6qxzZjN6KM6+a2XwMeknwTIY7czCcnjOCAZDXw
C8vw/Ie1Wf7qyHMVt5tOrkdEkoPuMWR/8qoaeQZv4E1Y20PUoO5JryL82eV+/Qolho9znKeqX7qv
k9wlGHr1hGYAFR33Dw5nOmzJYiJgqjP95yMPKzbHPdcWuU1Bf7KHOfCQ0pOZjDXj5qM1+5S4IuHJ
Z+14nC5CNYCNFVIxccGD3nXQ89zUOHN3lZpkgMprjZXhNAt9ZMPAQdxEwi/fRfpW78yQpUPzNhUm
W8eaei5cnh5NObJbINub1DWRz9ZetOCx7KOgHwll/+wkuHRlzU/HBgRwDsRha5fnOlOHQUR5pxLK
Pcr7t5MLeBccaHv5WESaPokFlQ8yhE2ARp473502TNBtvR0qsPFwBJ0vjKUAiJD4kOJQwNaNeBi1
+Y3GYZnLI0d9WMFB4kbWEWKLNuhV9mvssW0Ta8/GJcdnYL7kxDIq7ET6V83KdQewFG4DTNPKHJHd
0dxVoZF/ucbVBonj/qL+zUlco8nI7n0nR4Rg4/Ft43eq7XC6KHt91IIrWSVLYF+qCou+KjKpFWjB
WJ4fPivtNqqfSinuWXK2n3ok+hEzuzb2gOGhcfLRlv3Uo8xDw9fVA9c61KJ/08ew8Kq8C2iD1Jvb
vJz9yoCJVNLXeHVfL3eHraEZD1VsHvRUTCbJvzceCqmUaP/yCBRMpJ+z3xEsM6hEUdFz1dRzvlpM
lcnizeTAVjNOr2Zct01USHh3EFBdMKmVo4smWIdzxokRsPOvNT6lX8yinr3ArxOVx9LcZ/S1rKlz
9JXTRm/7pXyy7L42hq96w2ZrSGUmdtmuFGZpSCS4ql4yVbTw1I2b0CaSz/Gi4XVBWfmww5LDFYcy
luFGHiKa4+EjlVe5TR39Nj0qGfvsqnW14QoevonX6t2S9/TluZ5CWDDQvU7UM2vPqYcSvFLqiMwH
/C0q0Iy56fZL8zn0pFgsiee2yJ+VOyWiu+c1t7KxVvB20NE9h7eKVVnm4xTggH4OSZuobfMnzTcP
95w4xi+TKHoev2ok5PpwXwNk1Qk7KAKOZHIjrb5Jzn8921y6G8/PNe6BMUmf3KghUhtvnx/D5jXT
b+kEe2C9GOugj7EytLzSNIipepe2iGr/fXYALkXTtmFgFHwMmCsYDwwHv8yo8OvAMuYpIA15ntGd
CCQx4Hdbpq9NNPaAx8CSum46LABXiPAshDJBWcot6lEQiSVEmow93qQHzqOi1VFbxgRdQNBcgNpZ
gp/HYFlWNv2azoiEENdb1E23YjI//CuIkKHh5LgOc4v2V5RbDNo9awfQFn92Y7Gty+/jXekcd7hx
EfKgPBuoocDxdqjN4dccrehs8M7BObe8rkSeuRM7ZwX+c1qpmDsMONsrfiEh86ZSvp3n3mjEKP+1
OunBZ8VrQ0+A2gv8RPPt9ztgA1Scr6KNNhkd9d+JZuw1mQV/1pVdIkSwnWWO7M900tCTJbGQ044/
YnWJ/30ngLTFZ2b+NX4T+OmHzV63PZuAXHwsE5p6n3VVrJCvrmvypO3rx12ruOYBPHdzRuMfSOgk
vnYCBn3oM9rR3tIBEy7PkHq+LfR7whRAMPLaUZ7Mxh9cLlaTn+QFZ/DyLeEjbxLpWR3tCjrfeAn/
A1B3qWqsUfEvZtwu1FJ4xz0eQAjtbXBAaDUbbR53rfR/IwklFyZ8LASbrpkkCtT/TXKlQW1i+BrF
8ecjSQeYal4cxofih7QMQfv8EF+hYBPXkxlJKZoDRw3SWNCvKw5ULyBu4X05o9Fb4fcT9ajY+aq/
/qzm3mPXCzZ9KPGFXy0mCOZUcTvi4/OGiujjUVI9uo4/akpGUwiYD4Z/LztN+aCqZZwIkZVCI8wD
pdZXhrstNUKAk3eKbmhf2wob1sZVSLb4WQ+MDRZKJNpt1cHOz0mMtjaCmCfn+JA0y21fW+otSX7J
9O3rB4DW1HYwHfITpkAN3OHE0nC3UpcY0jwI3HQgegEV5HseBzerEk2ojGWEignuPWy+G2ZGn1/R
68ln+rMeUJOzPgkhfOkklFULqjUoHOD+w+VErlkYzLeG0QwNyJBnMB1kN4CaNLwCWZXMR9Cjil2c
QwFGdr+TaffdjasmZET6A6GHe8Sx19ln9wMB+Xxv1bRgABeIX+vbY3wDgZy9GJwu/3UkQdYTEZZ7
9zyNf2i+gWJ2+WLuRnyhEMCpGk66d7Ph5cQXkpe3CUR5z7VYL6ujvK24MlBW26QzwNrRw8gBc4HA
EOg3bnfc/vx0Tg4XB10yOBCR8VwdB1lgtCkmlH/vy0Qyzhfahlm1xIIvjwFCvLHkzDTOO6A/aZQk
PyvDwG8Mak8BS3iZKj/hBfeHXPfsuyhBqpxozlJUsm/IQkWN4EIp6rK2e0SfEFTXXI4L6znt83Xe
1kx9QBHB2VASX4fSnbBUjhvLkN2MOdDJyQbFbq3BvYlfRFuZsqNDWXgDzH81LeQUg4g0UPhT9Uua
YX9xz4WlFf/63kfDcXg1wbTJ8AiJAxKRbG9bqQkrz+LXn9dvO8C5Jtkyg2+XX3MsCJgCJvRm95Vg
gBjkrLBh6We3cW1HT8DSABw4/HtyZCyRNdGzn5rKvvV4y5t6QmzPLzLXxoiKy0yzejYghwRn75dS
8/E6Md0+IYaIr6HoL7HHqPyvPDW1QM55EHcehnGtt5vkJTRXvQ6qoEVAyKclL9ZKe6EN+4YUd8zS
qwi3YbbUVHapkEimpG3pSkJgr798nnje4RoTHvuB7UQaoqkn3U1nzZ8OBpA5VWf/SkSmi7+wtzpJ
o3h+Qmgmu8zMQ71wDT2imTEy781Xdx+XXiDjC7BCUEn6iqoLE3t2+QN3YVtmwRqbIR4hBoeiRcMV
gIKT5du2+6zXwMGyx/i4Vrvv/vYtnCgXyfhaXf37U+a0W2s/Js58mP0jeiF580OOyF/cEoZbyyZ0
3EtYdYsaNKEc6OkZ0eeDmxrRWswXMw+cxjK3UpIIgCajCp2FrxD7b1jRJIAZ1Vc7CPPSKWOKQSFw
vfTD36pwYMyjIC8NJxdfC3jd4cAZjbQ9Epm/usEDu/PayhPgv9nLTvbRjHiZ5MO40G6snYsP8gr0
+GKy3h++Cfs4mnQ+CjUdnXPjl3/8I+8+QCrLELcnJRXG615qH2Z2nk2S/tVqDT+xyh2G3Gv5jP2o
ebDClNA7dKCC/DPdSQUin7OiLtYgYAReA+oXX6bauWQtS3l2UmWtsjtLd2BPsQe4Tg6BmK0mWC49
Lcj08G8+HbBL3nJSl/pk1hpfg+tSacZ0gnGAHHtPQuigHgZ2De35AE8MlJ0sHFLWkN+S+sGbkZY7
HI0JOxxnEc4YPE0apoOMSbkoXisMKKgy150Fkkf5cXbKpF6adcpqBMJHea9PYi18xTnTBnEcdGg9
Gt+bO+ZuyqQ+KK7573eXHxOJp29MzEtYwRH33TTmVxIbeKiy9Jkpbvo7KQUqzybEnVpYoslemTA5
1NFb4Z4zM3CZkb7N3Mxd9Rt3/wdWV5wE+f8r2wDAemeT+5VtxH8NoOigFw+F+/DlAD/jZlLYYEf9
n6tri+X9UdDvEd67W1kKxr8s0QjsODl5kicACU5OWPFah/H+Hrrs2Pa7qmOjGWK8IVi+IwcfS+js
qNGOTnRriW93MQyUoJvVF3QMBPIuKn5imV5tNhNR6n/zOecWZJwacIrPs4AtBhUbo9y7f925FPNq
tXKvptPekJsCtzWxqir4l1MzfnuGdRueFFi6K8gAPmjmnIHzNE09CG4UKlekXmVv+TWczLLibjdf
rwL5WC2fYcA+sOdxVbm6+HcKrbQPmoFNBditjtOo+bZhgI1pXovxNLNWjF2tAIK94m08ipOYcNhU
XtsMFOxTV5HmkX/LuC0nAF38s5zxMra6kbhBex8REs3J1uFunG3tKlTJK4yfaZfEYYVDestE/NiB
IUhbsu21LqgDITg7YPLvvydrIpgoljQMMnNjVQxk4wAZbV85k2yyFBKtu0v0HRp1DyIS5sCVEkFg
NLZvXe8ZYeJ/4BqYi6KfudkbTXEHR7Eehc+mvotrRkiSUUE31GCjC7sAw2NN+fwEGNHaT8f05MaT
32yweBLsE9drFK3hdVUoxulzPcJXCkpFXr8LVc6cf0tzHaJa6Y0zYyUjeErq6WkSxfG7ubQiy/Sv
pG1SSMObFgEubTmaTqHp1XjNSJD1sxz+Pj/M793aPJTMCFTm4utWX6Rz7zMP/yDR+RkxUVD6aybL
IAaHVVdnnTlnrxhL5J2J8gE63TgKaQ7IWCJH6Owa5upQqh2lwUxDKMYjoh3yPM1L04CkZj4mfTV7
QLSUJzteMSxw8/dI+oPFFQ0MZZq7xN9MCJhVOCkuDtNCbYG2xDADbj9eyx5DH8eD2/Rl6aQW7Kmx
BzYl7F9Ross5CXf5vw/0pcLiHFOl/quHX8cw/10YrZb+s6JK2S+1l86I3tuEaSY/u+vNypV++0pq
Xzfo+4OEB9HTrChhro6xQ6rlaeBGNZXQaimjJnux7twtKfzPCvwb9fcebrp8Jymf+RR39HBlIz9h
oRxGtYAkxiApZH/utEy5fIV5GNtCD7OhGWjNnMesMsTbXNPGPoYhhMbqXkLJMS5Uu7hT2UoVm2Sc
g/l4hnM7NfmSMKyVIuzHBnJSttlVZDHt8/G7/xdVpCV1yNd64HyLJyRXbzE7wn5GOoNLuuMrMpMl
CAbSHVzhWgxKjA0dWNRiOPoOwhX9qft2yycdqk5yb/jd/sV/Gxl6f0NfIz/jOQg2RngY27Bk/SCz
9ot+Zn8q9uYBgcHE4GA3SWju/6kQ0Xzd/8tx8QL5flFjXAxI/NA0WEr87LBM/KYHIYbG3rQ5xEa3
+7Ew83DL3NJjxTsciyf1utcRWR7VCqIQauTS3J+1npf79S6mCSqPNP6429OhGC5e8tPImuCqES3Q
tY8FKqbKYvLo6+vx4LGl24mrQ2w9HnEGCX6zC3r50HSXBWI7EEbdfuVQ3H8U5bJa7yVvwLeOCxQj
+iu94faX7tVtJTnqlY/urKRWHnZLHr//jLygTRV7vmYu+rxNlaEmFdt0961HJkNdfn1pxY89d8Q/
tVOSAyiLyy4oAAubMmTidaa+HyVEedKwvcG0MrhakcNBDaAxloYPykdMbu7qD69fUujGZdtOJGt8
LrPbHg5XkM/UM7IgE8kxbzPepLafXwnt3e3yzDAWRbQkKvIcFLbhLJzUb2Kaa5Pk+aDwEghjcY90
XFSG57CMNaN2zqgKZE5QVCMeNsJ6ymi/ApWB6bAErRiIufac9qHWptmbzPb8ajfmf6uPPKUUTP7h
V4WkCvKD6mMEL0wjreVecLlskcStKXi8o1o4kobUkbGITMT0PPqQjUtmhHF07PM4Uk0Bl5My7rau
cNHaWiz9DfN9ofqsRcYYBXdm1COndVRiM3PZwauTovNk9mYZnb8bQWZUKwtaG2PxND9xbl7UqRqN
4SO0lva7WZAlFIkLe1QCCGkt2WswXYe1RrRFoGixbqWid9VNotYeUpku/LNx6GVHyv1WsRREpLcS
UOjuvL+uCYEPfYFPxWjLAqPRD28OW9gs9kzMdntlZpBuTJf0Y+tJi6EOIy2TzvG5d0gFODo1ZD7O
mWE7eF9RoYQqka7eEITy4EOmj7TrKV+Sqq9pPv/KD+X5W02GKSPJx8ylAm1bKi3fJWwRANY4sMiY
UkzZjgsOx5usj0dYPPOqH+ZD2JTmNel3PFc445VUZJNTnofSkfqOiWOP/vYOtPCpk2us2xG6POsb
xSERgDZ/QxZvj2C/g3Uj6V/QIxcV+3ayP6M05Z436PaD5Dp2c2pLJ3sRiwERrc0EdZQmMjpcQ/iK
p+RqEFCNNMxU9PZoTkgCB6Epsg9iV3C+bLW3QIQBcBVEB0e8E41AAxx8tMQ2QBEmcyAD4qdV2YYR
Su0Y8D9T4AYqgnYBZ4YwgXtnsVBgYRBHDM5hqD8bOG9Wk90ZMNxZg3J1ojBUjf2dlXyJ8lttr93c
QfNWWhQMQkik5uWe9sbcSgwLuCcgbpje/79m/E/RDopCvhaZoPxQ/rlbprh4QQmTOjsuQYldhAug
CFJzvVeIxv+6hB6csaSgnuZrEYTJfFNi37g92xAgWducB67fdqp42vxNipdnnq3r18b+VaQ/XcVe
oJY26mluZMNdyxLr1eP2UsIJ6y9ucXxItk2YxnhHqacEcsbOB8W/X+m7vzGoBF+cWMbwjBwDoGAy
ZiF8y4Qcgvg2am4dTLryXhI6kH0LKgwuFiYs8dU1smxXWqC/ahChmZiWLuq/M6tjF3Qn7iK7UF9C
/BQcJlzJZhctdFPjjQSK7/qOtu56thUGjVrtIxIfoR37tjipnVrXwSy846I8Ys/YtU0XiFJGhIi/
WqM/ddYldv9tVd6lXVwps26SE+zhA94FhKsuiUEDo92Tikyg22MawMTF7l7WdBqT/LaCkmvLF9C/
at8hWjamkus6Pn6SNb9Mx86AHZdq0P2Ha3wDVBU15RtYrzjGvjXQMZnQnaDvUUddvVzWNhh4ic5q
oEr3U59byQZRLrB7EbffnkbddbYBnqi2kMy/DjrBcWr/cKA95YT75acN4OpGoyGz+1jNrEF2QNug
TpgcZYW0DfM4g1BScupF9ZVDaf2nNt06m1yXfPpA5l535uWT5tukX3izaVUcrZ5NDwEjvgUzqMbs
AjprhmmcdOwpMRr2KHSpRNGj+OB5MqRXS3SPRTEGC5Qul/xV8u1tigmTLuSZaCEGYM3/W3baSf5f
fZeIbdY+ArfxXiX9hi5RqF4YWLJi3WYMqD5d/yP9diIwSBPta3xfZ4qbJCttCIoJDPH3seHUuK9P
tiGDQ+cO+ajClLGslAYf7iGTTukLHs3xQj/50ijmPuaINSg12Etvf/YoWrxQ5u3XxIRVsQ2UBEm2
9a1IftEvoAbG/bBoqw0EkTbeyq7JRLxWh88LNdeNjOt+9SQQ+TthDGuT9jj/tJ1i3bUM6yExzfS9
8a1fFp2+jkC3eNul9hbx13IICcsO7jFTQC/OO0ovplAClVpHtFsyF3BNT/qXyZm0j0nZwmYjnvon
XklPon8Ny4CJWvGJRcQrbVBjB+T0L1NPInm+XvDgoibDhjg9OoodJ7VvvaWVSPtQRdnxIe3wYGfU
WhP1PuRIl6TRDEVdMMDXFzWqpEMvhCTDPglRKjee5WohZB8bStaGGZpXUsHTNa2+NLLQafKQe6oK
4OvJQIbVICiQDx8KQSb3MJc+thFVeSLUYy5TGXNcTKNC95uTJCy9Qh39yioj74O/l6PhI6SBw+Y5
Dq2F7ERuW78+k9n2qOis5rChAxP42cOLpgDHM05Kakh0tHBG9W+Z/NaYi2QLvyNztHH3qPiJAqjW
A7ohADkDP71w0+E/z+F628zshrKnfhWb0ALgru9taeYaCuRKyJeo+ePslAo5inNvpidqWCrC39Vi
j+HzRPIsSDV+FoAClq1RAJmrWN+J4FXwlEJ7lO6oVUvlTsLv4ZJ4bgk5zzGpBuClJRbouZ8vPBgP
Gt+7G9LNIHHFUYT96WGXnSXO1lcaOsBlr6UVFu573iCPGr186Jq/KqYrfmWvS1O/zrrcd7N+AGiN
xhLwuogCgi440Zxwqa3qTcaTwtQfeh7+SQecd8VQ0/hAb4bNEGEWKX2PqPIyvQp7hkTvsNQDv9r7
64SFOojPHeuVazcwTe7RmVc+4FLaSbJgUd/RmIaXfaJiF9T6K3RcSioZgfcq+y6T+BbW7ZW9ISkB
vRxCPBvaJL9/q1t4gML0EfC4OxbCr5dRW1dJvpqTxI0oKENzCJ9N3RAflLKXPqOKPIeuLpmwWgUf
IaJb9nAahkzFEro/39NkTRl2fI4EPpCfXGQzMl5NIgqklwwX7IgTj4y/BK2tGz41A2kBzP5xHUgM
hlTGscGMd2Ea0FtONAroW4Vu+B7qWou/AfTC2CJ9UDanAnct6q0St2sTqQf7995kEHMorzAddLCd
A0P7IKTONeW0KHDeooRY+E5C7Rzbn+suurz/AnMavUG/XDf5RPHO0wSf6lHJALmCiQrgg8BWLgfE
EYaXS1ZsmzXsVdCW51TPX+KSt0Yqm8QpH8Xq1J9lWvFMh83h+pQbSmWOqx5U5+eGJ9pgyU8RLO1b
aeZVJk9eSxsHbDNy+MNorYO/lLn74YfA5+rBxdX2GO2329aY42d685Z1iKhX/0d/ZpI7Mx0oSa20
n/1zFzgxMiPHJD3VG7qGDBW5AIS88zeWqoIHh1w7iGpkbdM1sA8A/B32O8HcDwZMPbR6iGWf73pP
b2IQRpFiD2OEry8kLoNvdJMKlf8+NBH1QW0BkggFUkC93uKLz3xvX0eGtrx1PG8r5TBilw711FyI
X9drdimmkrHAMxLnFgnWPZnqCtB0pv03ePK3H47WZDRETXnO7+GVFX31KmHLGKpf+HG/9jvSHObH
nW+ajC2hIaZx6IzzN//hdz0NzH/L1KYJm9FNfkhCT2m2gjpYfDWGh7GpdH+CproFn+92Hd3qiNAF
89jY/jJt1HTI5eFXMjDwMAPPXT4M/ed2bVjyVQMDk54bQMlZJset2DbzwWlxHYqdizhak7OLnw6q
5R9MJWeeQoqYz5Dg0wCmdZw/4ZU7hsMJsxlBWnSTj9IUClRvBYc0ac7rNQUDzP1D//J+++5h1tsl
32inx+0JyFqg7Q4NSUVD0VoUULoSK5f2GWO6rzSqMcbUFNqJVc9tljiIOsCQSWG8PCZoWZ/aEdeX
RTyCVr5Xk2fX7UhmnSnnBpPxMvcQgFrLJw+ctdrAT7b1ycYmfmOYTrd4gJvZfxkkaOSroZ9okMFV
uPXy9hGIduTDTdhQymsiSkU61+rzVg4gQU6qnjZEOdJW9zRW4dsYTZmhfG70G6ER3MFsRyZLw03S
HFkhoTxNQyRgpwl3I9F/vvmxTXJNdiF6f7091S1XnomcFWUUymR6nQFj6p057R07t3p0Fni2fg8i
AIY+kT/+7eXrOZC6yWq282w21aJFjChEJdncPdimX80HlPw46TAuP7po0ERCV3Ggby4be5JYAmXP
myJs9b78wcfv2jbzJxISLYkOz893s7MmXKKe6fKdcsFgeMU/M8GhQ+1hZ35pnzEy+yNtMTFttXAZ
aXbl0Ri0gr0EpyRGPfUa88VMuwBRhR1yKkXhEMNUfHSW5KoaJoBMK2p55EBH1cO/NYF9WVUIZkVp
SoyjOapgWlG75rvQTXhPp3g7gIjo6NIXQo5+vaWHhq/mgNKJVuoL1teBdvD8yXvtXBwS1id9CPEB
zd6s6Updc0CpPAHUNa5caX7Fh7dgtbqQTABY+MiPGROk1uD5e6d0NgF2mDhfzcPP2pvXZRMCKTxq
9IZymUMUjFmz0oQG8/yu4B3/sI5cvs3nAXo8vF+lDEms5En24C1T7SedBA8fJIfWvi7HxJWDq/FC
LpdOOxahOsl84b3p/Bp+5pl4uNcgCdsYIOOqoqHXm3JhKG+k8t8Z/KiyhUcFNlCIh1B8+IjHMEUA
RyWAvGVD239l4pv801yAAaGsRLDFAu/UwmY3k0c4z94ivGgB3ec16lVmPbT0+0xStCLVF4XixTU/
YnnBSIxDM7Vzyz7LOHwXLuk29+5IG/lOSj7jyG8VW6EB2xrm+1iU3gbrzcoda+98X2x/XWGWvWNy
ted77dbwT6W8g7rvIO5c2UMSNHIspHoTaF29XUueLIvCj+Xe5oNbJLIN7/l78rnejsJSwhxmgXkG
Igvyd+Ep26LzvrgiR3R6seJhBXCAPhqvDzuNNgaXhKz1q1BEAKPGjFIX4b7jjPgSYarjz3uZuMCW
QHh3e9ppDYi25az+/ku5OJfHksdNMidk1xEAZDbL3BuHPxeF+rykUKH8nNw05Whzh6H2d1o4ytPu
6YNHkg4MHIKH0qEnbRHrwPfpvEB5rAxwWvlwgO97YlNjyBkBo0V7Pih7v8I1vIyz1rqxLb1NBpKS
y6sS22jy39eFnNYbQFedUXncpRKq2mecGru0pHIhRZH23sjGEcWxnr2HQ+GZg3EQ4nfATpcsLik3
epzhFN1l4kJvnRQYDiN4OzIULZEz+1fVnUa9E70H6ZrlDdMazoOBDG6KncxJ1VYDGtEibCe4lPv9
zvXFG8tlpKQ2Sei+Fg9mwg/bruRoUjrx/pfrpiPL1JKgwixtBM5zFoc3wD/WX8+Garf/UM3E0/yU
ISu+Z86UqRHxZq/MFBy9B2M9AdUgFixfuUVpYaz78LAucxkyHQG/FkDOV89kcB0eCZF+q6zslZfq
Vap89QXRFLCQzFcY+pRfltYuzgvUY29Q9QMNb5lHXatUTCd+la9wG6s18RPk7Pz2ThuQacd8vLsE
DlZXPK+ySSMnPaWxdyJ40pawjJUaroj4a23Gj6Deq2W6/tn9f4/LTYAYVIlNgP2nNbHYspUSrgud
R24OPRsMGy8iHWhdlrRRgyXPzQEZflnjh76DMPHGK/LW3rk/lb8mh6P5fmW9x3MD0v66HjsRq4nd
h2ruDKx+NyRGOFPgszvZV1xJwczrj9XTl7fj2uVUX6kFDwpijYvDnnGgfwK6LZEDOd0L0LX6TSn3
E24m1O1cB7wzydSn5LYJ8WbxuR81qSfBdanJr/EOGseVPVHdfeGpUmpsnZR1Sw3vLSX9HpDSqQp1
49Bhnei/zkRni/zzGbRlNpHtzRobpPkgxEcebnCO8VL305hDsXpOinYvvscOu3gr0pz3hR1UqkaD
uULgyJ63scdhCx9QTv+dbBaNCroSOXpf2rXfxsvbOB7lQ3OHbQMg1qN+KJjA1hHm2wQ+CGXf2e5e
DUklHt61iYTIbCSUlwfdC4lEGpKIBcu3l9Co0NbExxphHC7z0IL7iXfprmb7021Ie8JQudgxtUfx
qbLuMys++oBV2yPEBzwnqcotlA1b5fQSRxtFbKGgMPfNdK/J/WPce7tI0RO1LuGYOARjLkV/sJ0x
piaTSHWULCT2a/46rLbmSz17x+bO82eTX/3JIIc7QlKKrYMPyoLZXFx8xct/M7vyLJBe2mxUY5DA
+asjVERTg79aQIRLLRH8pDGWFgsSoDY+cLDl3iD0KbsgaoHI90YZ5xxr44JbCdM+mCb/cjeof4aZ
wKzcEza2wE3//buk3i+uPnNxHbQ2Sf/WSDdxDFujNjsBIDNgdgYEq/ypBBfjfB6Yv9l0EdpYMBzS
etom4nNhswCrfYxKW3XFs31yd+IPfhI+hDF20Bf7Kc5wGxv4U/KCei9aVmMawgR6jHSj5xdmKgnT
Q8kvK8w8dpVM2wDKVPzRU2dJbXr+mDblIMJsTOLF17PAFUgX73AZEP2U8VV5F5aW9WzZ4gSype7/
q75KvBuAI2Rp1mfFizYSjWHgSJfdDUZ8BIX819pToZ2aSZim6NunOqwwFMt28CMutk4VWgvWfAlq
reM7Uw8m8+yTg3hFH9+6J8mfvaabw2FMNKzwJAI8tckgvFNRl0RxixwCY0IxUw379ylU+6tMn/k7
WhtiasVfo/6d5YyIuq5mZoMMfiHaNiKTrpQBCevrrex3tSnw+oEgfM1pw1CuEMaUR+RXJEi8u4sw
aADu4XoCKmNk4QsTOGzqeiI0/0TPtdkNFcwyJKN8GIUZn+UizeSY2IZ8IfhuogfVkiGLZCLfrKEV
g5tELDo6JT1R7+5JeHBy9RvpRvbWQT5Pu9eOIC7xIxpCkeDIyOIcq6ysdwyHS4AglOIf9tz7/dQ8
V0AFmtz0D3b//HHvclEQDRR2b7OgxQjwEbWSJckaaS+isOCmiW05QSLYo+XhbY+2OlSZs9ITliig
7Q0F+bAZdN2fY8NwLzDEQqlJowkF+KHhDC2zCfgMR6HUNHgLbLs5rxGB+DzXVxrQ7qcewFgnRN9J
jffVTVAzYYvHKHwjyyiCoyPNnc+wg4jk/EyAz3J6wWShTbTDGYrBrMboq/zXa/97rsB0S4VokkDv
EEMK6GRyJ0gam4OTsOsZAGX3n06DHPwK0Xuwb71abwDdzCVm90Oz03DwgKPu0EbKswl5g65JChKJ
ICawRLKirjQ2cmq5fMkfEwkqdoq3MhXxDp+U8wWLiSpWRdm/BgihMh/3jvgSJ7XYCDeWfJc6mN3m
/EwUYy0MGbajODWZyOXYfxKw+UBOo85AMjWuWbal5TMFU4cabSH+68tON/Ikt4EXJuoAsxk7p5QY
oViLWDa4HCf/HuY9oFGRIX9Zt91ZgaVDRPL6wrZwmstmNOsAGLXot2ktG6AV9oCZuZIRziluROXP
GncUxlwuWqJPE9xxiuZBifZXxpEcS3q8Rqt9Yq6WzNGiSL0+UEuKgAqlinWLKnbjGio4vhQSxQE8
J8whcC0MQbMYnRF2VB0hLSnrvwu0q/pfIAqOA7HGgw0R2iBZokeuedlUGip4Zpli9KHfUk4GJtvF
OJb6DhgVdwiUU070sFjImbFTCNQyjgEVKky1BckG9QDOFKJEdTSlW9jq1p9we0sXFkZGBeR69ibo
8fJLG/FL4BZmEH1EBiEp+Szw/ONapSNMb69cEUnTyEQ1w5idDMfdoBUxQeUvWyqVLxf0Du1C7LQv
QCLbOdtXLsMMKx1rbFjiJ+D/qJqAL6DTwEKzyx78ad6OUTMLjYg6NSRIqDrGumcBJe8gfBsEBylr
6LObj2oTDHviKFE1/YoxWmd3pOPbQss9u1+ApEOaU57WOODG4C0BCECFCKm2Fo0ty1m0f1uhW3Td
KXnoK9FLF9KQhkQPuiOfcL4eJ0l9ctKFg3v7r5PibWOVX4arco1yIvskNtFzX5VMxUl4UX6edDtN
VJ64E6VT+NCNzhUSXONiqEnhmT04EDzA4af0yeeIiv5xnHf+Pzax48tfQJwdSzTg7QXqqfF5oZo+
wd1GRmUQpCAdQphygN4fGZM85rXLTP4eMLN7a1B1grt8xsZDySSu1tgUTjvknNA3HhbpnOQc4Gdd
kQuqQlEtTbtpUu8SYZCz2edTjxEPI18qB6j4GJN84c9PNcSiqPaGiH5PgFeh0CP/+NeqlQEaxPoT
z4duqgs6uSauRdFYsy22xWWJbvtYFffbuq3yK0IUGYS3uqhG7ZV/g0Olayyz0pr1Av6qd8tuK0qR
UC9jkYlVGU85q3OQHsqUWx9jgUJ7AF1EGK4qzICozN4kPiuxNzUpRN1Gy2D6oMUQcKc7UT+MBZo1
0BVivvDNxVgyvGnrVPgFCQ3Is1+GInhWDGDNDUTP5pIzLedJ9TouuFNE4ZND4BDvxOL+68nwOe97
Mctn8yNBYIwvqX7XBFfUmjBdDNVLr8zuBQ/78MAbZnbjYCMYmOU9v6scpYsk7WgcEnSVkgj11EJN
0xwdUM0d2s4d87AIj92hODotSNMb9gU2FAdm9qmlCUZ3Bx5E7e+ooof3C3YOCXpHiYsxGJTRgZ8m
S0i+wyP3GjVLWTsmmYneMCq1HZfT+rY8uATFMX0UMaG52vKwDnpf3toUJPQFo/eZ/YsxXl1gr48B
TYcEmUl4NLBaTMEl6CXLMw8Igw4pf5KYcCu+jo/xJDMP9Bu3nMpQV5VpYu0wKmbgC+iobInTkBjp
Tx+1Zo2aBLqFS+jtSO95O+SsaelUtCUsAkQinhiJtWgWdxc5wFKs8/QGweCiDfRJVHcMYgkCRwhC
LhwWOX6PyDXk2d91eQB5x34lMky82fyeRQ9OEUCMtYUD8VREh2l6fOdGx01NuKG3HK6YYmRMzfaM
JVfiYAaPFDcXiojHgbFQVEvGOrxc9GtiSfREDy85yseUxN8UejOm1nVmcoR5BtQ+0E/bJnB5Yop4
1mKNFHPCM7FPqIsitFQjeFGTBMYcisIA0TqToCxkvs7pmYFCKXZK7Lnhvf5KRngi/qNIJqADDZF4
+d53MOjjZ+eMlmfoLSKU7ZO1WBctR3g5HtiDh9f9k6Ea/5QtC78plvMUErV1NPUpIXTTnAK/0ka6
jX0/JvcFlAKdgX23krpnS9TEk0q95Xr9SskocxSkdG+qDdk/wJ3+/DeqbiIHd4pZJSC1ZREbLaTn
ultV6069OvKxPf8cHKrK2wqf8xXH5hHYTKZ16oO/O9ZddZ135cKzetC92FYDQIeNUDwipxMJ9scW
bJ/BH4ISSSGk/mf9Hid6wS+xMoVjfvD21XSLUsjaFp+qvy0/H2uZ4VkKw/iO4kbAuiTUIZ5dU6Xm
zSsK480zNqF7NTJKOB6KrQX6AO3/WLDQTSduu8qpn6nTatcaQxVZyATM8FVrKGbma1vHcvwSRSCm
MYP9f3aY/KyK9urGHKOqRSYoI651ffETMSvBCzufIBfrzMpGRNyON2+iVUC8MJ2jbD5CsGE+CzfL
yVI5aZbqxMZk9/liKMPkzOYj0RObjDrRYICuvrp0w/n1b34CYCCa4QQPCf2x+vpqYb0yIZgiO1nH
4uXxJ0rqwUq5qneLWZhdrbRkWcxcILKuM8/ydwmryqJNmJU558JGF/eiEYYMejPBMX3swz1KIMxU
gkCbRgWpe1VIQ7SielmWT9NUOJNjY72WES7/as7OC8Id4kcQFLqd/873FHajU9E4hjQ8DRw06VkH
96ZRW1Oxr+4T3SeeQv6n5X7OhHzxiAE/uHDcFFMLok1vMotwpQ+KXMdozFCX9QJRhJuOloJHvHTe
ZazBlXSbgwJkLW1MWUFzhh53xscG0IEj1FF/OhDAjBPZdLUv4XJwW2e0Ko+ShIFzhDkYO/CgAcyl
X69VKSczt80leCmYd4YfUBkODJTajEBbKJexWBSewXToUuoumFpqVUUO0UJbwnNcdGOnvHTiW/bx
3MiXlRwUz5cnBRAptyYVVo62n+DLKkQBkZTngZQFjGDB6IMAsJFuEE/INSnapCefPgaqNv0SoeU1
F+ju0cI42MVyWokiZolxdJoVRHsvu+xrpPTkb08+yAFEazJKDD/THNcB0ZA1bZ8uHZ+gWKZ0gDzA
5mWWZ5X4HBm/5xDCH7ifTl0nuY5TkJteWI00f5PS5ECEDNtOW4KmyHjOj5SqufQAPEwhECdMZBRy
5ueUercKXqL8BHla/owR4BbA1C7GsxRq24GbuqWkhXr1PLRdEumAsArZfo5XJEUvylxgU8RhDyMe
E06mcNFe5snEs8tW0G8kP2bJ1FR0ljwVETAh0r6wJyjNMvwN33umlHHj1h8/xSBaIe4cjphUJ/u8
asVk+XxoDZ6Ue04HXUarccGmW3+QK/RA8KsDflSq4XavqM+4iAvos9C++luYZ+1TkRrVURMKWFkZ
+NQpiL/VQgZ7SOcnFtarlX7KjgpwAj9loX8Yk8M6XWnoZ1EB/NtldFg5G9fHTHbX2GvCX2sxGlFM
hn0O4xIb2qw9DdQe6CuroQYzUcwCIuvJrkKTcxTiYWSaGFITqeHnd6ECx5UO8Jx+kSrHYJup0Ugm
vghJvSnOcjyxYZB8FFcgESPt+OJUxBUjLu8HPJb8nJ58CO9QYhFiPk8gkHsG34bLk2mrL0sxSTxP
MviDMn537Bt4PEJo6X8smOBVoe0eJqiDrpg+4s53soHyzJYcQqYIwdnTtOgPxIZnQd/MNhS/F2TY
cx8WpbK0eGGKWi68srsCVkcpJecLIUiBsGlHzKbd2brkwhY/9SNYMZltZ0o1v70aHDmDi4aCic+B
DGxVDFuDKIpaw2LAbnshVN8NAOhp7oD2vMn7OH4f05qaUmBrqRBmwpV5r+E9W9RFRljBq5ipFOXz
DzY/D8e9wzf8sHvHdMLPxfyqKGzVb3+12Ni2YzqUqNYOoYQtGWp//5q7Eds1IbyhKbdWX0ADH+lr
uwoksBYoEx6qqGrEC1EYWjK3Dpr+J7nTp6wkvVUs2YRRRrRlFXrEkaFVPyhcyXIuDGcsq0kn12tg
NMFExEb1nKnsUBjc51H/BtFwfj7lKvwx45OE7b8Uk8gQzdOLtkOFITLt5lvH4CSY5bOYSlnYMq+x
6cDibFv6amStA2nJJxRxuckug8giKgU+ipX1lsGMfh26EZ6z0qUF3rfxp3OyHouP0waGXjBe1aX8
yjQVcu19T29WMqcB3hY3AixbZ3o+Nd4/LaQWoTdtJOvpo/jGZ6rb4xW7bJ84uEGzhjhoQkDG4aQP
j4wMwpp63wjeSJNIJ19aXQXiPNz696FswVuEW4kKE4T9y9K+aXtMLFrxrfVCbNb2K2xZH2Wqwb2G
3+a7xuubAsGycWLN218awDJOCJc0miC8gv1zSVTVdKgSPX5AJjByxba8xFiPzxMUrBBqSFQANmwc
WD9KmpcyZHNshl5ZlE+QuQBQXGG6DTqB05XyZiLIGjT45JnzfaR1nNDQFhzcMJcQ/mThsixuwtDD
bvlUfs0PLCd3poA+TMG4c0Jb/gVvsUZHf+1S0Ju8s8L2msZf3yGqKouBDNxNz5s1c1zv9na+g+BG
hvgEtSGCpbq2J4+x70e+DJbSce9pAevNkBcYHNutzJeXxfrH0pBpA/oqUnWMzIXZGwLMis2xJUwD
K5PCd0XllxBY+lCg0MhTycAGQM4ByMmWk9XAtI8Oi14gOx4w9763AZ5yoV9YtODkUHNVSAdEtrQw
zK79Jg4YzIIAAxLNPcQu+bOzIfECm3vzOrdzW9sGJ79oMi40aaIrYHxO5jPq/32MWHgQM3JPJJz9
ThBCUswI8GCI/Q5SmcnyE94tvWzx2TM8hZaAZ3/dtkpYLePuCrxRDm8ew+p7/islK/bsU8lSwrSJ
CyKihhGWQtrvuWRkgcEAoK8MDvQ+aq+NHxlIqHfgu+oFrqTz5A+s9buFQWyKiBwVO9oyxvHaSshN
y/D4pWdEp+/Ac3H7ZjDQmU4vuxYQJJL14s8ZRkotsPyS+5Sg9OnHY9hOGQ4zeeVUAyIUHZgJFW5F
4MkfC+Ms3uxc32QV23kC0P1KM2Wfak0QU+GYNH7ZtnThJ747gBzfgIlx/9jXKtWjgF5AFLgYolNk
Os1eeTVnCbqqF5t9ZNqBq1C4LMy3ENAacpJeYMjDQRtu68Cqga0SXLUHUpER5NW8h2EjwnLFvtpg
CSmdQKzFWzuOtaFq4kO7aRkz++pKB9TAb3wI59mQkQbLKdltppnMTBIFSxDpZTeDCbMc4DqN7eL0
jKcpqabreK+n3Rv9nZk9jJ9DPm4cVaSrUyiHT6RvAXfcCQ38JQlpAvwW3Zn1YUqzdaa1PI35f190
YAxOugQhUfIfPZfJAKmWhOhP+bOms6vF43fjAK3T6aD1rlpof8rdhy1BYfZvzWUHeU1dFvW5j2st
l1aCLus6YlAUo8t3MjSY1baN5EYtOMrCcApwOnH5GxC4/wBqQvkC7odIvB4iy0HMlzmd7RxkVnLu
EjQOe7nLr9Mzye8vfB8H9y1uJhuj1kwW1oSNc9LXKs/fBtiMkD9PXE56Y7/6YiNTZbfW3EkZFsdS
zle/ybsnG1eKUhLl/se0yuq/IC0CEWmk6Yso/aqjk9O3LdCBZ17+DWVERSYm0aSZp7lGAv/K+eqQ
2XzAOSi5h8h0MCX8Tc7XfptUfo5O/8LUHT437bRrRet3sQStvvNPDSaMHVTFK8yQFKnb1VmlWM+7
M/5mWALrZ2G56NsGxKpPnpC5VD5Cq7kPr7kewN4dZ+Z1QsqESYuQgAVFjMCNwuInmy0mk0TJOo73
PEKVPUYX3E3Ai8rOkwFz4L+m8u05MwTwKlDoY6SqlNc0cNTv2HsZawC4G3a5ZxtelRFEHCRPxpYP
MuTIv6OcSk9mZQKbAkw7TMsyHIK2CVILCVh7vRhJoCbbMHAvsKBctmegzywZAT3eN6LnxW2yZgD7
+N/tvLaSujfH45PfhQN0wb239dnuLYjOhLTLIek82L31qyssGS9D8PO9VqTZJ6WiCVVfs0Kwh9RO
XPbm8ckxryBokJ2gRYQDk0v46P4RMia3ET9U7G7G9ygckbVcYOtmeemhYqQYpV4BsR5WImiuvLJM
MzzR6+hh0UI1ltbfC7znZZv3OfpC3BnISNp+VjvC5oFrFHU8gxwmg7RDR+zoPGjfCC1ERa+0IPfc
uo25zioF1pIjGkKGWZqYiJDJ6RGCKIGqCNVNN+PdLJtrLSl6hJ+KW3gwgc/w1NV0X6SguKCFUrZ1
9l716TmYJEnO/KO+ahe5P+Tb3mKdZ6/KVwR2koacPQCGm1actFita/tpzerQLQGHXqs4yKAQu4FO
25N/aA4IgU3R/1juupeiYqAvJ7o6NSyuEeePhM7E5EvEZXkrdIiKSP2DVXZfVHX4j7eS6CppIO1M
rgnBFqzpHsldiCZVVtRwKTxir/lS5xbdu3qdpIXWLur0Qu+bPPadATSecZCjba1vJyCGOxGRY4US
VBo3WLujaF95h1EfWr+DIN2PXsLvMFqhI9OySuATeu290CHicO45tV/BuaqEncTMMT9fM5vOVQ88
jhw0gf6dZIpilzWGscQasJUENc8tt2cuXD+NZkeXL3sspVdNcrVVHMk7wXRFPUvDXvuSIGXkkbPu
g/Ct9B23OmzuQHu4CNTx1AU2VhbhNN+mJywXkLhv3TIsWGT7h3NhkAHR3HMdzgV4xxhG4oQHsPuk
TBWxBMGpXF839RdqC8adhLbbWVqAIhHA3CX+qZjkYSeGfses679MuvfJWSjW8MBfwwJpWIdH/o3b
j2BuzeNm+Lq+KeOnYIl4W5OJOoB4JJa/AlyxzAcFte5zXVxRZSAbgRRLItdwPK1/Aurxf5pUVzhU
70y0A7eTT1MBnyUuTMwUgQwhi/4mAQcrE0rFizJ1SR0Mr+emLakm0bKmqagpW9FDXsmHLjrcOB8+
w3WmLpx75IB4WMra5TMuI9xZ/wHgfPtscnHdk8Ll+g4QZ/SPUYzlGOCF+1Qu4+X2r/ki84m2R6sV
D9tkq+nkPEQi4g7Q6Ph0I+d746caI596pjt35cYmvGGtL5Nv5hb1TxxHjctRcwUXr/Y6lv4oUXLY
Nl0mbM8wvhQQl+Neq0MhUvnRCUMXkQVQwtgNtp5tMsGLlL1ZybV+svKXE61t+D+uqOZ7wOQOArZ9
3mHCFo9V8cCXBI7brId2DbQMeaR+NZiD5iwkAfykc59C3IHUOELWRuDv6YdYmXsl4DUYQi94j4Q1
BGW0CdVXAYtXK8dugeqH4bR/XQlrSmk/bDbhrJ+2Op3DKSC5StCeEGTHMqqhpsd67k1GP5MDti7w
H29qvqvbK4rjQg8PIj7nEsPQGFKpLiVMUcrAL8WTArK0k5i4B9FAbeQwgYDHEJ4aEYcWgm0/Lsks
6450y0GI6Pcql6dd5oi9Qkw/uflO+Xupyb4tBiXjXrhpgCLFU9K7VoYC/sdu1PC2B2npWZv2I0c1
1WK2PlTL4zC+HLZwh1q37c0iy4+O+o9V75tTbx4iPc/xrFjmiP2w7JiJnnrOYNiv5kvA4zMrFEvW
Ea+OsOEBZ11jLJChNlsonW4iWy2d/6VvSUI45dMwEpDw7AAlXpff+Fibq64LccYOAvhEcfwEueYw
OK78jL035tvbTyyFvWxlii1m21JDVYn++ZFz2rPSqLyd6OjXdEmDnfcrgPrg27bSXg69P9ONCHoL
KgLuyW1GoRlw3pvwdkKrzEkf//MFxqJm79SpjhOZpiBv4UEhlnmbCrvt+d51S3YWBxDg5YoexjOa
BSUvs6eP8BmeHrnwOEB9V2jYtXPggpJ8iQzmanqqilW5hTzGr0Yvg3jVBSp4F13yOE2DH6QgZP4Q
flNJ72n0u4/m8IcjcAP6lJ1IJWjKh21nyDZnKkor7FMFwmud101qc1c6gPvEnhEKaEMPI5Za9fy/
67UtUGtBL1BvoFqL5tS7SSsMc21uxncWuhB2Qf/G9UkBKW759yEfT5DYQM2fYRKuDszLc0fCVLwa
oZwlCwEYHnKsqzFUGh5bI+frRDBdZp0L3tZKwQgmEdexDoZDwo3tpV9YVZhi/TIitg9Ny2zNsJAT
e1K64JrK1UYRaEwa/59gPcw2g0ZmhdsAkgiIFHB+T58bJn25uLQ945+GgCzOfmXx18WpYlkLJedV
eT7S6BhFe2N4XKjaTWyEBrcHUOWOmRTTS6W1Tm9ctQ5dQt9SXx8BkfY86SyQzhL/u/NozNJWTc9c
e+7SmTJQUs2FY5BxskYPHv7oPkmmuQMUzttItYqxtLzh/2nVVM00t+b+jN2O/PjRoVq/PtnpZahr
E88mkDWVoNcHLAAwS2EXAwo/L5ftH3joaen/ke+6DpFhhFLeM0RxyqVTFqLu1B52Vs1BrQLx8OZM
03/tyivGUqL92tpyXeUXd8Ap03xc+HB7XraKqBWfpyc+pnZ3Eelb2OI2N4FLW9Vgv/thf7N2Yz3C
0efw57tfEoxf5uwsVD/5v7qbCl9fA/7d8P4mNd+Oi/4pL0UWV1EVTxBWWdajEQnHyOq35IiqjV3D
yYuIH9D6g2XtN1HBTmYGTyCvVwJuJknJJI7T4zE77EnhCaPDrjeEx3j3g0MYJy8iRHdAd89AWDnJ
SDQbt38D4r0JJ3T0YQibuAvGz0DaHaZcmkAbkMN6ArR9yFWYp/UVY3c/TkIMCQJe3yz51kkjLzHb
y8o6VuLpt1z7lzmu12SpMhFJ1jLNMLLCHsakg6kh1DRKH62dK7UBDwc2zD/NlU0GcBIDgQJFI4dx
OMIUqWPL6EYem5YYTYWVCTWV/mthprdiwC/0u0T92KDBnEkoUWnqorru7UkFWhBaqk4CGO1fz0r0
txXouamLWSmRv3pcpBi/r1F9cLOkR7jVCSt6H1BMjFNcZ0wUiL9N/pFCFGESMT8G0llObdblIoiF
4VlrM9KYyfQVsnSNKPo20IVEq8KItOGWorLjSOP+KY/hobV4XhoXqrp6vErs34pq0VI4c8/f0oI2
xcFxa7KmIUUGR+53cFgwCHxSJCrl4OStYIuMhfaxdvQD1+KHA6ty2FOAhe9cMcBdGf9Tj5ALQKpI
yQhF2dss8v7fDBGLXrhDInZKXFecLIWFQo9YKyJ8NCkZIvX1pRkMA6xk/I+bYe6nbjrx3Ew2nvoB
fjRekN1PJnp+VzjyEP961TeM+Qx174NPxfZ0gXwpy7hwfDg37jAJ6Mg2WqnKjyL3jRNCkoCYJIg/
1aYcCfJp0uz2O2U5NsCA6/wNnLXpVtO4uRrHxBDlgnwXwT4Z6gtVH9y02rebt9E32n8M1RJv2q44
c2E91mxJxErUS4CEWcsrX2VJwMGhwvG6KQX5p0+iFENrfOmHl3uQJFC643qQ488qUjShDF9VYD30
g3Nj5Q7v5v3rk9gpcHX/8rbSC79jUFhf7Xx/7MdKXpfV4QuDfbKRFlQrXCPaXVP3V3FOg5da5Piu
7837KqdUI6+nwamwQ8dtD4SNqDtrs4Nw1L1xs48O7wh33wzS6mf5bXCvGoWQVF9ukmVyhalBd6wn
F3+ojkTBE4WgONE1C/0roDpw3xEO3wGagUiwLN615sdM83ZxGD4fGf38y9NAI/82cT2F8IYGGwFN
vmy2YAbDXeXGSmso3gyVzTsD450mApLspKZQ7mKuZQlcDnXgS+1IUlwXOjFnNGTUnNElzI4GBdp1
ByvNPreCsQm5O7YDKgtmvqV3P4cLp4Ia5AWE/4hEZEhxK7NxXMCnnq7TKwDIGbjHLPe+26n1+duS
Sb4ziKYSXagIX513DZmjaP0w/RGArpHM/MvzsDfAnu8r4Bj9kBWOYowdr7rd3HjElUgoDHRYrbg+
bH4xtd11xdGEOO2z4cw7y0w17oXXgH3Dh+4rkadPOq0QC8M+oEIsJ7xK2hTPm6UVgsqjptzbimqG
ranyPycs7mE4p9rvKneH4s2yHWj0N0pjp5ilkMXXGQHzxWomfUj5stJISw6Rbo6t4rzwGpoC5lOm
+lVE5EWwIsimeB7r3uuF7UIr3++CN95oPCTQ4GZn449aZknIFEDWzNz7HVXIMaLcYv9rzD2EOhpE
83PbF0/hdC+m/omjsExsLTtzZmsonkgdir2+xAYXWgVfs3G9NOMR1geZosYumV9+iz97HoxqYz58
gPr+TlNbf8AqCGSGfXkZsnZT+Wp8t4O488fW1fZ7guChAqCInG9P8fqvcrYmA5MDXxTVpZossL2K
Y6QTXt6mZMJi7X7LLNrffWvPGPBZTKbdIOk6U8emyzR/tiw59l0SXDODGPac9ztVaXhzEtFoRBPH
ERVZo9nNx82U+Hozld65iq/gZQzu5NkIGWFDXXYvMY7VHwMfvA1nTt9Pw7X9f9DTtAfglZpUT4Me
L7i5/J6V8VuqG64PZvmRH1qXIQNP6WSp18Lvpl0QRtRQT2aok8DOuoqtCHxCksQmeRJSlKxQSWEz
o7ZpIF+EDvJscTyiaUbVhRk5hNhoZlTEhChhHVjfTNYLX6Z5Gj8yzrujFDxU4V7iXWvLSLgVvRYX
j+zGNidZ/ZDoqCHzK3OdM6By+DciMeVRFt9daayLTh+SLKJRP9WLrvIVSJKIITLobLnpnOA4Et7m
lbUW1aN1cc3I1rza0bpDHyozzBGju2lf7AhDinS4qqNCTlfPb5FclN7rsCMhHKJUYBHrrTvARJsF
WDEnr0/GmpNoFTGFEl4pEmrK/vDB2ZTmZr+dLq3n9tkZ8yHHC2crzi3RdFPgpgXcnuyAU07h5oc4
eRtqp3pGOdqbtwA+Vmh5qDPSX4SSa85S4KkTZQtDj3XvkL54rjluDi5PWxOrapfWguSC+848yflc
FYCrbVOjK2torJECFN0ng70eNBnkq9vVRExjEgURxIO/NzKMrj9xFsKghN+tsycJufTSPtbgMgLs
mFERhzNvgcdApYHAhG3zLvJ0lEU5IGQotgzpAMpCjKTPck/PTl06cw+ln6fBAxq6XEkL8y9rZN1N
KKr2NTxXZMCO2LI9cRVB/gibu3s3iAv7iC/fRexxQ2PawV5dgGZSwtUx9ePKuVdGzq2CP9k2yseb
s313tcY4kl6TrUjjNbKRscWZpZDi9RS5x+wLt76yQeKQsoAWWLKOSIB/wO/R8kWtvm5bbIa/0/GE
lA7Qd3OrwK/55hIcCV9vmgtZlqRBIOuctQ8eKq5rhYsjmVIfMQXb38y1hHnBEl+LJaH40rds82ev
f9kJutA8rtG3V4blEJpeqZ3PNKF76YKZSSM+fN3THK+S/pI78i8Wy55b4wUWY5QDlTRMAEkqtlMK
91Vqwwfac/WAu2zD0vVLwn8fz0OOflO8yg8RmqnyBfofMCUyF+KttGX3U3U1h+ccD07xIPHft335
UDuIjVK6sObjNw5J+ZwVK24L2aFfkzeICda/i344t0/F0e5WzOwn4HpMWGUXeJT0JjsYXRqPcaox
hb+Y3L4z566vomFfR0pi5J1F083jaDZohrQFM3xjGm/6BXyqVqsGA7G1Bw+wt3Ih0G//G3QUqCH7
lokQZNjwXxyAZXSA0vPOQRJaHzsqYtqhJKMr9kPyUDnttRB6iVvgFJ5byV7LsJ6SYsOZipgpA3oa
FRthjAodvIFRu1UhhsHO3BwYhI0ygVZZAsM0kl+DWQYl+zFQYQIr3nYim6XDOyD8M0SOV0KZoOYB
3w+oBGTuAv5qwby8ZUs/x+Z7+FHGByejTHeEvWPxY5fRstc/2FULUv3qy2ZRSqz7rwiXKfwd/qtM
x7giXsOCJFl41yLNplqX6q+WQL0iKV8ucVNbRJ7EFIn/908kq8O3yIcTnSNAyVspRDsZtSgvPFLR
oeKeeI9TAdyfR0f5TV3VccGaNkjEfCPlt2nnfnQjxvjO/SJUF+vOWXuCHz30FMCzB0L4rcWp45wO
1wHsmXFOLRwSsXeP4OJdgsXZ7MAZPr5v1AoimhaM4s3PXGsBtOMJyN3ccipU8J+BGDvSTz1JIIjq
GjTStRM2u/KJ/tcBHPiZz4UnsmHcHbiXSmS8invY+17JdK2QiFtcF4kQZtA1KxuvTUIcYjCT9fEB
IhYr53DhKWAf6eXf99Rvy2vgHyXCBty/kcOW/WeqYHxsHN1KFvhj+4BX0UfSn5QDzZ++FcwvJfsr
A3Nqb3Nbava14HkOUKjcN2tJ0AjNZEbpBdNGOLk0q/lLS7thY9n7rDkVI0SpqBG+6+ePEDuiRKkP
Jd9cEVVmaqEn0GQtxweiBITwipIlhgaFE/S4r+xsjSQs0PNZj85Uk9m8WC4K57npgyH+Lmm3zL83
cNB3HSrK8C9fIw09TzU5RSrVUZuuEGe1Bo370N01uECQr4KUD5vPP2qYOnfEZLxo0KeqLh5PD/D7
qzP4P8Sr3QDZ5hAwa/7Tgu3XWPcjL2RY4798mT9wOHs+dtThvDuwLctUO/fS0BIZxlQcWr/OLavL
EVseAItFz32Ym5AsGBthcnMsu9w9yqwD/92qL91uk6K+wQyay3PC3XTKOmosxtRv5Ec5yfZUFI2b
goh5QCTwj2LvP5BEnLdA+IVPagJoPs1QtSlv6vMsssM/TN4kToHyuCMg7DVZcI4aF1VWggkYrmBN
zzqGR0ZycwYwjJavOWqXqh7kv/vRaq0ci4a1hlUU4R4Fnvtoy+lUYuEIwDzQb0X8E6wGL/uRUm6I
FsmpmRJ6vw5CckJIjeWZjDET5jEvxBU8ymHCW+TYI+jAXiYc6WIHc1bM0SoXPneRam7m0d4rGf5H
ke9JBs3S0zqb6SXUWZ6K3yEkEUZIOljmgjROYcN+ySqRRNxkavUObj8CO9D6TTJMWnqPgVNyhdyV
ttrLa7DVKG/e54MnwRWUVsWnv9FefZeCzahdxrBoCg8mEpUTHo4bKKHY/KS3RmNFBG6hJUF7edCP
Hw1is5VoPqG1XtOiRd198cKwWUNM7+siV+Y6mc1tlXp11VUb9u1PwIbCweNarLBhFFJ2rAwu5z+C
l3BRqefEVz1/dCuwIu2N2adBLjU7YfuwGrwYIzeHb51v5SfeQH30OI9GX6MpkSKNC5QgSSogEAf6
7ahRkOMNwtvmHQBvI+0wThF40i3KG9fcymHVIfYi7lH3QXEYrFPxPNgsQKNGlYGuG6LLvU2QqdTN
3FFprZ86RzVopT5z9ZVX4nodvGlJ8HRkPr2UIDN9RCX2JUzIPcAGMEJ9nG04+HThvm0e0l5t3UF8
PKOevPSlp4GDrnLSg3EI428qTLx0eNwLAI2oYVMhybyHtT6eNJ0A9ku2pOnlYiJ2rg6hYQZIxrct
LoHv/F3Xi5tFoDc0MiM6UVVzBxPPM2TLK24dskeWoKzjxT4QSDIipLUbvzJPJjOSavwRMSYVMVYC
mnVYcKAZX3oLyc7CqzDbPBu4rhEy8yXnrOX8DegzkF2GdCc2h68SVKszPxE7u1eh4MGOh+NzVzEE
Oc6odKBreD38e3dfZGQhRWgsl+Ti5iQM5Fo4ZoURHf0LeMP45R96q40khcU2Qh+xfoKnWmmpgNVN
Gq0rQ4pV5EguKez02K5sMPCioYyujDfeqN2foI7GAJCtZQKOYIWFaW5JKhTd7sV8sazjwS8haVfR
BM4sUxeBKuj27Awf0OvFiD4gbi1n1TZUjjEqk/inwjL5+Y0MEx4MMfW5QCLd5x+HjHzfRX5GALWa
T+7DMA+4lO+EKLbq8E9vw8j55+qpuN7MKw9WjyOF7spZ48vbLHc8AfQfuwrgsqTX0CD0ZGS37H3e
aAN7EMv2MEfuUvsXtxRM7jCin5kGpjKNGpLxbXnOJmqq8CPujn/RH6FwszwOD6kmvWwOdWiWI7RJ
XYjox/kU4rzBafg8OjFYSNBOreKzbzQXETUIu34IxogNiZEMoQf4zPefHIAR5HA3ffKOimI0P8yq
Nl80bpnbHnMNUjiPEFGJ+xVXlVmeAZh2KF0JYQ3rbAEXO2HVO00CHHc+Yis6Ikmh3CxkCK2ozjyv
4njh2/N978oN0SghxJWFlXlcKHLzSkzty82tM/B7jo1p2ZPrhFBZb9/Oh7UTK+hA62u6cUeFq2hD
1cESaSshiXQkg6MyYXbkpHrX8ynf9RWzIErudBnO2LqFSK2N+pdGB3Zq378Zn+Rd4K5Z+99Uwcqk
KHOguV+uVid7djq+oEL52Rzac6AOEyuTwVymaaLWyjKsb5zI/0JfOe3adhBlgiZJObOQkoaBNHT1
eRTBtoMrqI+IwdX8QZQvxMtLuq2Pj1WgNZx6tAspc866s4wvwKz6oVXb10alPJ047SL2xGc6nT2g
YBUnCrar+9RjORSkpfqCd7W5aO9Y0odPM/U/Au9pkclWsNQRxX2HswgKAYxFxWqZcz6IrzNH1LRC
ZlS+XHQA1HmwcklUmzL6wdWD3Tp8FA2YBxOdcnJ+pEnwgpUhaRVnSnP+ZMwHoiVRwz3f6bsAC1JO
ZE6kfmLmbL9HsYEHkxnhbp08epo1Hq2hyZSPwkOQ9IqKJ02S4oeOBGVCae2mtA6uyXnsgD3shv+f
W8myxzBW1AOCLOWW4AXhZ5U6fUb0bCFxJwzA8dfOZOZLih5ja5PDwxoKNoMkqEEp7a1gh3RmqzPe
knynNC4pwKYBj6LOGziojtZXFgCowCtafi58BdUe79iYqnCRFxTL8JKNVPu9yO4nWIoU3VUZK/1B
AdMvz9F/LRsOCkCU9xoJ52gQutWiSwjCF3ew9OdlcfsNqx+fCNtC4Wzv9GEdbiWk85Lkzp7NEb+O
W6pEeKd04rsMZnweyLSogWykYEDfc0b+0KTD8mR0DQYwI15jo7LO2uJKvuTaCwp193AJAzPySVYs
IrW8jezyq7JjCX2yTLtMtW+99gInr79ODJhh8c8OAhz00/WgVWMObFN4kgk9mIsFv76XliJ92ppR
AMinLxXZdpezy9izCrK9+plIGnIYSntJmPS+9/jYUJ1k4p3Dktu7DHFI6jWREmueSYV58Xo8H4cR
1fANZCePA9+rbQhQqsjdjVHbwXSSknh5IiYkDqlF6qtA4fSGx97Fq/FJMajgYRpSj4Eq4vkvMPGw
BjeXUyWByhrps/TUathYwDmI4utH8JHoC9qkpQsafw7GBFlge9wJKmOR1YWEpbVIYTNEyWRdD48J
MW3Yi+Qp2/EyTqpW5PFmaero+/Ymf+YSNV080G8M851gBjFfIGeZ+t0VnAI4+Yu2MQcI7E+Tb69V
vQ6Uhiyaitx5A8A7soTJMi5KoMjARmsH8gYlSFTaRfOjiTIOCRnHrkfg2aU9nmcfQpWXHP8Tc/R/
axldVJpZP6syg4c8hiYliiXu0I0rtqw97J6pxSRUnJEdpZsPKDy9m5BOoZQ0OIZLNKc139rNvhfR
JDT3jSkOYmKWHlW9zFlBnSaa/sDAddGDQ5OAfDvvSkZ3RJ5ct3GolBzsi4BPqP3MFF0L+aXhv7lR
Sawx5F/UuDHLUBRnSXE68GRu5REl31pZwyx6A7HZ7+F/XrlJiAyRxI79UPiHc700byCMRRvyKGdv
Oo48Vn2F7qmwOztW1iN0WGOAObvTawpzaH6SyHVg4ccwXIlV7SqCtCzSb7M1Tda3MZMzAoDTVLvY
Xv2JDnZjgBjsyIp8j2PDp5Fb2DZqZpUstKw7WB7hElxZcSsGzLmJAWfl8DY2oH4XrhgxblLg0IP1
BOj3vKpkJSX+kNNs7cTlXErH4KzLBxlXNSbiG7a9MMH6KND7re15mhomUi15eFaHnxPZQF5sJ1Mj
TRHQ8M75PMZ3en41jl8sRVEDbw7whpNJejr7UKDLTN6zvmDd4F+JNAyxrN/TkYNdEzF60Cel0p5/
ktPC6TqUUxHd7jpkq8Mbx87NdbHsZKiA/9vm31wRVQg1Gihx38ssyStPlh8zuxuNuzVwJP6knhfv
jrtkM+iBivnrzahize9v6kZYVNxC0+BnuT5dF8Njdh5EIVX1/R572QiQyBpxbvRGGTWkWFQT9CXh
q5ZN9f2Vjg/9Glb6NqHWehNHEvXVidZNVvhtF3y77ZrgHAoJP+q28XARPMu13PuWNc0pioftLC9d
X4V86UQtADd8p4+1oughKLBNLHUJDWe8V8mecqdacoBIuIn4sWGpMsabEfa7TJYDu7otoH+occ4m
H7u+TPAp9aIlbAqvjLzOM9WRRh6mVS98b3Avzmhic342ei5HTUfl9iAi/eF10yshEdezqDILqqgX
QCTm3yQDg4fWdk5LIgHD+px8QCIr0draIIsZ6Bb1gPEHpx7ILX+GiBqQLYbS3pGk0oO/c9jLHNN4
u//N9QQ5BPrWHVOhekekQJC8nzuniqnWUmmMQl03NST1QP+wynWK6LCFtwEPVpvGN6CzTNraFutq
wyCx4HrIH5XZ29Fzd+M385FVf5dEps/e+14XQebHoiIn1ZVKi6QDwEs/6Eb80WquRmRANRGN8sxc
q3bnHfh03Lszv8psdXRycAgBiro3mGkvAFGX7+3oarK4Nl8Cl7oaeIxUoQKbiI+5r8XZ3a+Gs7mh
WHEGzvF9cFbtiSgW+wMoQP/Pe6WbDHwcfWWx2VljoIo2zQIVN78CcdsxSo/acz9Yzw6lTW/1aNgW
PXiKD5UDVFdL5joXSn75MrtU9gCYThUn8m5c88opOOLrHkol0Y4LeSYLO/mOds+lo2oyonGt19y5
IVyoK3CuM5v3sYapzTqymRAKvezh4Jl/dh8UbVvsSF9poddjS2pUhY1bBzlslZFhwyt7oTipqIpb
vjFdMYIW03z2NUAWaNc6OdtIf+0tLxmbyQ9HCf24dYYR9myI95HZIIQFj8w17KXEE0HYjVAYkYOy
4/z82dafy7KQwjWc6cume62+IyIkkMFlC3Mw6YN8TNjEmlT5TocOSm3IrbisCXNE3/TgOGHPezFx
PRQUthQctg1Ihro4szdt/ajXYV0Pp0Sha5mtZAwe9Bc+SXf/F9KbMgHaefqGqgcxyTT/tIHldslT
J58RDQDcTpsTi7JATeT3ZLeAkX2WSes4DYCqszMdKECw987TZRqSBpwRkvR0e8ogRuPxFZJ5JNSe
qi9LcKXcRd7SKlTklbR8ruwx+anoi/AD0QksnCzyTzgz96bN3+1P3i1+UfyviiP0JGRYKloiUCTJ
qxy5NIZvhq+NrRqwXgNAb1LVT2cLNg7GCDrQy5wzMaPs3JHFhb+cxNv38+JciJET4zLLDepqsGr5
ejxA1NqK9C7Lz7+J+HJOpcyYRbYW/I8lUdxmDDzBzr0BGoDAOo5T9fXwqO+GQm42RYaqR+GcCZM/
+4zGUgGWDf0Mc2O2cU9TikrkLpHR3oZ1FRGeDzwZn58kGa0+3wauQyR3hq8HVXsYizFnOb8Su8R7
4QSNmnGgpt77jGGHbV7ZuvsALKE+xWlnZZ1iYhQkzuHcr4vPxxa5720E5GFn3Fc0RtWN8tgEH+VI
+ICJXkdzwt+LbylB6Hv6BC/2CTCf0OKhei4cSuUlOvzLvlmTgVzxFCO3RRxT+ZJMyvXp7/CYW3r8
GWFrxpFI7TDGBKYZk19JMkV2TLxOiS3xxjp76BiYS7rq2I9QHPuA52o7X7tPSabNOKvW1UT7dBya
g0bkfp3A7aMsnUxs8uLGZz/zwPFfidDT1JAtWqF8y0bKN8aKyevZloNuj+AY8NgbgD0YO5jmSdpz
zAgAUsfObJvFfEuLhTGWmm1PFu12/Egp6DrtksqApCC6dn85F7u7C3nlJAjLLpXkWpbMcNbpirUY
Y4QtiO+sD50QVFgGGv6/yIfrJMVUtZazdGK7QCQtFsAnNK97h7miJ9mL6L5+03BB53YjmZeJy67R
sU52Zt7PSFHEI1LUuNEYsnIzkpysw9g4jZb1yEqLsNCDycCDmkYURRk1PjcBWUmDzLU1dOCO/Yni
LYiQCj+a0CRJLqMkW9VXzcW4L3H64funp8jphrhqNTqndntw92t3F5LuEL7cRUclR5ZdclVxMync
5tyQA2ipxoeBzuqChu4gN2+Pt2OuCZvIgxaw0i/Oj8+rfolWSCX0anLeVZrO+Xnl8WKv5dBU+fVM
iD6i3RWNFeXpd7rhqlGveokZ8Gu6DjDOal+X6fK8ZyIvs8zoIKmbN08A0NPROjIXLuj7f6/eOT+P
yo2E/z9i4gLRDUylQGY31sMGwU3sL1BwU2h5N9EPQsYsLjG+Yx9AVjiPaGa8QENONKtHKOsWFI9s
2wdMX4saVVgUotf7cat+jNMYgpqTur4CdcKhg6rQcbnCoDfFhhsjML/MdUWkxuc7e+8IbXO4BZzW
z4zP/KB8Vugb40JLIul9JhE39cIMSuPKP9AqApV9Xlr0n1aVviALuaeXDKj7FdwKGxs10iFrdFAM
DoNjzHIpIA1xOiVCLwVuiC+9GJh5y7IrarNFSn71setxvMIRubjPVv5gReB/bp3hPF11KZF4I/ts
Q0jdE/jI+Svfa9kqm72OqOLzraKNQfLY32ngmbvWTkJZVGulMg+Q99MRxsYIW6Y50hiX7uIB2Zki
/1YM/Ulm6fOMQT8jdexGfcX/wjHmKvWw3tsaaVhNWBFJe3oOllgPECgI0lXLMa6L2Z2Q0RO4UTgE
ZvNm1lsCzfmBbZSrK7JO4r/v/AufnwY5kV2vjGureEM87riU71DvctUk4pIPV1wOFQBFOy23r+nA
YUDyEDGUQCT9xrZitG5iEneBeLelXgQ7METMf//epRiM3ggVwhx9ar2ajcXXew2tq4LlGUn2/CCy
8C8B6o7hh57NwQ2anDNG4KjL43MZSom2lmOWknDNw0NaBRfAcp5QILRlZv8MChYIcw8UaOrRhvdo
hf0XKPgA8Nr+7jdOfq/06JFqRavP4JvEXwBuRKjfs2aBL4zAcsHSKtwRMkFV0b6MtzGKLwRQKlGa
fWyOsR809MzoagdMxdd+dWb6YQ+4lef6691m78ESBhOi4dGzJ95IzpszKnG6307SfADwOvsk8uZE
5BqZGGqyiWlC8/utwRs7R/5lp/wP8CtMbGu3tOF+v+avYFf0OhmeCeZRikLirmdc2Z3cgIIFQXeI
GmWdl9DCV429hZUGTB8RwV8j8Fasp3yWtod6qdT/LRUeTI9vM1TFTnRhy4l6uhcNhBOSBrMND+GK
TTiyMUItu1645icO/8imLZV471YFEDy4PrEYpmW8nLj0v+05ViDxLRLHnBInyoYUxhd42v9gDzP+
OGD5QENb1y3cWQe0856ykcaGETPF3XznNBCJEfNjaVIFa8Hs2AGIeSfA0Gz01FQNh00tRLzUEPGT
AyxfrB7eOcgIuVRruNBeAwGjS+ApehHjfMxOvhIbmji5e4+SKmnWxi6T2tVoggHoOsE6YFe3100M
X/eUz5GvSOpFrpQDXxKDlg8t8+DKqaCzisQYvPb34nSAitKWduZk5/Jyc92emWxgt5MerpXneSGa
pBMZ+KOGwusaD3tj52fYwVQuY87e9hbBVLNzf4bfapD28PvPMNDeiyRK0gFF6jMUGKUfOZ81WstB
BjrwsKfckYXqLFeJVgrqKr4ZY7MVYhS6XTPvV4QN2ycU7osnvschJL9tG1wrfjebr9sdXITvBvEK
iKOgpPcXshmqBJIgy3n08qkjQEzpIhtDSxei9FPXEAQsxvcVO8C2qzXN1188gvE8kXypDDlvbYBI
ck+bflzsdQsrUhT7PltfLc6uIzI6aZk2rY0BsUi/hnopLFt2VGWDtPOrS17kUfv6XyB0cJ21XSy4
A/p9V/v9wKXDCyw9xdpFYsuu1MQSUvZ52SvKFAfvifZVCVkZ9BiR6Aoc3pikqDlfvmERcrNoSa7R
IjE5nvLy5RgDGO6IMcAlzgSDL6AZzqZ1aUE5UxfVhiDUKIgSA3/qAzl0VfxUv5xvRoNeogjmDXSg
baUwR5/dKHroczNsi1tBVGJjac2OFpADK3UFdtoRffYAyrnXphvSm9dj0nbiJMwB57vhjENRXSQU
J/jPx3Id/NloJeqh5reI/HSK6z4nuIO3Wj3ny3NJZGz/UBBJDivQHI9H4PZ0MqCugLdae9Rfjfav
rvKh6NaNfRi77GECwZzW3g+9gdG2Ai0Bn3dYIKFTIDMgTo343z2BaMfpmwN8UlJnlIXP4saSqAht
MU3Qvh5ETwrnlqjhk/ovAv+FU2N5gyygQTGnQXOEOgZUkyY104NLuXJThkzFB3v1MaA67kk6nJEj
8V2M92LkHaO+bS2x7TtcQVddtQL7vE6fLkzNcXgyI0WNdbmbJT/+kCBidiK8apFuiTVqH2QgjytX
3JQCyU8QslT6++2JPScvCNFubxiPpKoadE3m4Rw/VJbE51Buhda78gDi2/EJY+esHOHZHOgIqUxI
UPXyO/8Erub3s0KcUk/eGvRiCRjtUugnclF/Icges77VPz29bxr+MLYK9JaXYYhkndwXPNTkOETw
yiFYwW1dQy2KOxGYnSmS/x8CX+Z/0MUiWG14DOyMJ0o8QiYFcA32eGfcgFhu0xIlyRCCRF7d2Y3a
in8lrRaRM5is55Vt6+NF63DJk0D/g2LtuyH1SAh9FUr5gORHpX7oHD17pbloKPiGByoQ+hABDBau
4oYmhDtcSHO+PTUyVeMmYeg0vvD6byOLxcAld4ikBe9bQDed256r/UePuuaAHzcLbbt2qM2O896W
v50Fso8RGafq+1hM0TMrhYbX8prUC9wCyjihF0wVIi+nMI+ubmFQGPeAq+kLOHDjGZ9kAftdcFie
3k9QPxlBcyVUa/NKNNmWZWfPIT/AjIHXB9fLbuNt5u45fYrlMkD71ITVTkXAT+RjMgbeQKdEgCWe
yUCYmBRpdTplUDM3FEJswZfNw+7SeUq99yAnJwYqksTJgj8nOsi64NINCc4J9ese0sUFhlQYbU2N
6uWxcdAvTINldUiDUYYOBJkmtd++fRcfGn/Jc1J0G/bQ1GCXbUFzwTnenTPhvXLkSfixfg8sl0XP
QGFllkg4M5CM7ojBemRT/+yO1uJoZTdy6jlNzZJg733WbMBxGl/xT+PNzeroL3Lfwz/yKz97xfx7
Ix49l0Kr3Si34ywC67eZa7Y321M2bFg0aqlhrv5yIslglTB7wSmWi+D5zHpdjVEQ7iy9ar989P4o
u8z/OpDFVzAF3UXlwSCfDiIaSdNxpYx0JeIQ6SdZKxujvZBGzHq7vt/u0t+QHLYfOLJFiE5Brvxy
SmWv6yWICtIblHbl9ZxJsMK6spa/CurCbmBaUNf2jd8KK25BvINwKAS9H8BYR/dzAq/w4W2yqc1T
5r/6SNCb9LrbRjZe81zoxVzekNxPwDxT0MeD/TUsaxPcD1J9U/MAboElMRoUEkOdqoH+WYswLT2o
5tcKozI0t2xnPLf7o00fevInu+x5QbE9UF2MVPpIZZJKOITw3e3ATnTxnvmsg09SoRfj6x0TiLDt
sXzFZFzynZqDgfSb8BdIoTe7V8nolF7tL2Kzwibwifmi9duxUp+tKlzECsOM4Pm9PrsX13cAvYX8
yM75kFj7wYrMW/iFGsKt7blUM7T3UZjoffbwQ8aR/9sQmRqQ53p3iabOXgzFA2FlKxupEHv6LV5V
/m9yhzxVToWTUz4j/3zROLyga8dijulxSrBcc9hsWUWTiGlz3hsOoKbdJubDcvP17VcWAqqfnMTd
ybyR/NINoOFzaKu4AncMVjhXT8ujcBl+CVWPmHkBTJZGl5JYV4QNhBQmrSInGschERA3FCVFCYCy
mNg0jqynJ9mGQ6vj0X6L+AmJ03CUh95vxsE6kcTY9K9S/N512t+k1Q4aqmh6q5L9fHufOAFd4yob
1fXA4jlt20LvgW/cDG7esOAZmRSZ+nwIsimu02ZxddIbSKj6dW7thwJu7GBczzSQ2y9GVgt0jgq6
l8H50ZfcTJl+wvhXmnCuq9CbUCEa5N+U7+UHk3YOQFjswdvXTNZR2S+721zxb1ITKSf5LC9mJGby
bXxgPQPxil8CNJfHERn9b+zl80wNUAOauGLYnCxgwktWHmcV6tI4rhghwvbW0FCetsTBibHoaL5I
SYLAJ0YJDmcedM0VsC9rRgvGdTqc+/Ssx97ktAD94wPXdRTQMe9stSTkpO/395su40/iu473a2m9
hBh/r8WDOQjMOIHpGz+5TsIkPApcyHqbmjnj0FeDSyEhUbhoCVP4SGy5H+lXZLGMJMvuExYzx9zP
ABi7mOtGnZ2WhL0buggeukMCmXVgZOWzFgSujs+UMKQ1OKxLrRlLA9ilaxs6dqo1qkbHNjf8/fJw
AOmw+jE7OBI9yxwFaZIAgS5nzv1V5t/G565ex5l9GeCfBZ957bM7bDOKI6ebN8bMpRBDPCBHOBRc
W76sJ+1qlp3Y5ojR58no/HF7JthmKOIlEClXKRbR234UFU0B6QN8/qdfQ9tmvCQq6lyuH3hOiDxX
W1ysNEJalrcs8sKdhdKawnaTW53YXLf9DoL/VxkN2TdWKUxluYySmK3QVZ3P5CiflfDNZmg7MGsU
9mMAkBpzmep6AF5wQ6/l3T8MM686zz4PMl8ZluhwvEb8gPMigukyZ0gXslkzYz+KypIJFvJ6A6db
GYuNmMU1vzFvDfmb7ReSL772VH5/GoA+FNtol4PAiVaWN/u8dLO9ih5jdDCh2sg3uZXIPB1c9WYW
gA5L+cWNX5pq93wX8+fnyqD3CENO0PIX6sxSz9o0th9ARZIdztqarevP4B9yumd6jhDBvl/pAgPY
cPGxC/4UDLFWwolha+5M8Uta9XusjZ6JTDbSKaFxXLjqTzk9H+/NZXJ0WcYiXuDURgZ9AjdLwHdU
oB9QvwWfeiX1ACKGDoKYMuvDUvOV+2Q/gDCIsQ4obpjDgI34tZtBrdFRRdScDK/mlU8UvrY3aGVt
qoIxt/XtoBW27byzGKp+y2IDmEhmO8QoRLnmOHOZXyYFFaYW3zQs1RomCgXYfWDNFUIyGAILDQyc
svwYibQe8GXKXk2IxiuOeycxgEriTop9nh2z7qUMRYR9YGWMhhO6jvukRVvERUJm4SBslBfZdj1j
199JonYK+cYvj3WvumKb5pNWYW90FbfV7YUsSOZ3g410IRsba7SWxRGvLy1NBJC+8H1jtKYMyZhK
hfwNI6O9othypO4AHNvDI7vRya2kW8jzAj5RKXHKHhDDOm9p/1cPiuLX4lmUfucMk98UiM1FOlfE
+eiN2xfLjEiQ1uk9UfII5sNgJBfP1VjsDo7ZH5RIR4tc0FJ6zO0pRCmKQc3b/5bW4vc4mHzopSLi
jhawkuLgdJhcgZD9h7+JZFMZKnknp5vmx9sNZ9fgSAJi6oZz8Z6iwdBCsNsrWu3FkrzZdERqFumv
KmjwITvugqbFQqnCVHwJ1GKufDoMmkDZ/fKGfsOYHSh2hQ6Ewwvn0gcSA72CREn54hQsCTSWUhZJ
dX1j6JZMdIqm+PAYacdRYTM7MBitQMUSQgHTJPKNNfRN/Py/A11vgBmaOvkRuJKBPqbWSQvHB+8q
T/IfaeZk01HHxynVcT9P7LZn3E0pesfPnHMeIjxL/ykhv3mwv6KJJOtYZRknCo/KadkoxaXvB/EV
bJz+aHZgtp1D/cx4VFhJ3RE0YwbCw331DrMXXhqYt7569DyVk8hYtp5VAZ3dKh0OoUuMIqoIGHGa
uqwXIJcg+EyLJQN0tZqnj5mEQSu7iuzBcE9cQFtiXtE2x4Vd3N/o7dvJPbrJHU5XUWp4Wa2nF829
3vXSDhyh/LPZ++ZzJH/CvsHvxZOOW/mjMYPT/hG7QZrqB+UjcF2yxdp0O4XOWswvSknEqGYzriMR
xKqrXiOiUnW0OWVlK/Y2x2CcHCdmPTS/LKJX2hM9oXBQ6R+sm8fsQ2mbfBeM043D/ztqj+spH43/
1lhDzoOfw5H81zdkU6jWWAf10NxiKm9E3kqqXZssPDqHGTa6KaKP5Ws46edZiC5R0EokKmiWejWD
bjzsbR6aDPdbj/OHGgjR5HLRIxYWBavS5QkENuaUwdp68660O6Oh8+HRMKas7t85V9Cqt0S4gDaT
ph5cm/LkI2/0bgjQhVVG8jQBDlzDPsPHMe604q8agCA0QzHmfNwvvSJuzqvex2ZD2nvsB3gVcKTN
I9k7XczltuBSaej/AXGE6LOJjoX8ALCiMt5o/99vX1c1Jvnl76u/u15cz1/X93NoLM5TGZ33mdxk
4WCK+uRbNJxrU+V40l7Z9zagcsZYZmEHeBCPN1+rOLbWHZdqiPYZYSDFGYrCxSPAAm7ckibKSFMj
FSq7X3aZS8mDkAA6KXdN4ln0xVRghLM8IShRMgqp7zENlWTghe/VXi3au4P6DoKjLjNmkhLFR5p6
UpzLSu3J9GJt5F4n5F9z2ikRKaGHWY/4kmTS+LvPXep5NQdjJPuyEo8+c01UFAv3EXMEw3uWO9yj
nK5oGPv+Uym3yOLvdatbUdEGw8iJPIGWWD4m9Vn0Ka9q9YIElMBq1+8tIfoF0/jAbUYMDvGhuHy5
pp3FYe4ZPPSSMxnYXVkmJ2LoQepXxjBC/OP8J4+NZx4dPYoByV+ELNI5nSZZdVWxuFaKSe2cWC5s
2dXJeIVRu6l2Dib4nQ9PltxxnW5yj3DfRBZli/Elk3WtOYvIlkxsOVhd2GNJLfL26I/8CUy5at83
59zM8b5ZAla91TuOyLft+JyCvNZeOoM2Kg6X1MKKR1BKphzpGYljp1HM9Ck7JvQW0A0yB+YCkHo+
/5n/hQ8vB9W8q4HiSOmoHthpjOYvoazYnN/PiLZ3HM1ovaMA3V8VIOXSWe6uWWtOxRImGZRYIhT4
zQMxOPN4HPnEnFT6sDAb4EXXMkA7QpFTh2kmbwBVIyHpy7CT8HmDMWt2qtUDVKuRGgRWJbcXYh7V
tefAgGO3BiJaM00aIb/e66hFb0v/EEZn9ZHKQC3udlsob29BFE7qHYwR1hHyXm2BepMdpoAykWoW
jOtOWQHBedH0x85EudCdIFjpz9Zcx7yW0PUdd/YBUljappRwLJWHOjpkfjGcFeNNmPYr+LucUHbM
eWaATmemSh+KXT/0IoWdqKDuu/jjlvNf2gtXeVCR3K8qNs+eS5+PER8gtAN3f3JqD9Qw9zHi9llt
vsjrjNmQQQnZ/S07DOhtaZ/KaXnS2CgClv1WevEJcTofIJlJM1V7kodJZyFLzD97NpkMH30Uw272
2IbrOHvej5tKAgQl7vxK2eVy/AKbJB+7Z7ZkYLjCpnk/efqHQexID8XHAusqX/Nc8/H8tNLmyRPT
xvw4s5J7oyk5mqPims3HGrjmuEOl5xT5b2rGhGXoTxvTkF9BWoYJfxMYQKlmDQl+vxjWe7CQSP2X
lW0C0vCiaEo6mG9g+zCpPQu13peKamZCLiwB7ICkHbZm9a9cyVFgBMmlgCoKJHPbkpB+7Z9n1znN
8LxNTKqKN8UpZzXeCJdm0cWcoqXQRayphWBP7/KHmcWgAYXjZfxyvyKnakAFAJaW+/VWs35oyo8l
KO+zDCCOKa7AUYpcy2KM4rVJ4oRAC1pYRdUG1eHppevadJeCutpQ2dvFJtAGGFeZ70vK3gUThHgw
V2sXioiLFloOeqQvMGRnLLiNWJtbBJ15hyeHikaoCn9qIJI1mhVB4AGsmxyuYjmFWmegJFMTrMTx
9sd8kKk2s0sYfLb2l7Ju7r+Q0twhEYxou98t7AGhPqFWiMlvzHw8bFYYztyK+SxyGMTBVVm8dKMZ
cit06uyWOXg0YPmm1W7CaPn3XJzYlaWQIG+P+RAG550QyVssUSoCrKh+ze+CXlfeoaEu5r1AQCQi
T8P3ih9Ku52fURJgI2XeX7G2reaTpeXSZGxBGExEz2nkidO/WfQRJf5UpYXZNmzsfkg8Ww+gX+cG
61Cp/YJGAmxQbq4E/68L2p1vhR241RATQspoGEX8b2zNN8CxY8EbCadHlGwkyLBfZpUuHndhkug7
wMqTA3NC4LqOZul1MkrNYwhj6MsBQf/EzBfvLmjKajcUksW5KuikyfhBdztGcKj41WlK1zq5cg5G
0/4tsM4+GdAoanDNA1HXRPMGWtrrlK5UzMvTFaC2R7oBvfUB4D8Mt/avWdKCfhT90Xu+sNC6J2vm
rzqQSE9k+5Xs9NR0PtmUKtb7bJ0wHAXirXlnb+R6LxO3aJhb7tRpVRh6BsA4Nfmwy+dbZnb8/ehl
nYcFqCSRBZWgppkN6x+5xJGLebZhtspkaWbdAg5QTXOjyDU7JQJFyg2/2JUVZfqFcXdKckL4WUcc
JULRuipZmcYv11vKthMjyg2OyBj4hUHiVC69vmOZE3D8rFozlPJ2iu8m+8ry8kd4tNTXLKhIUX0H
PPSLGLCUth2CiPCLVDHXAg9IhO9PdHsoRIhUOeWAKCry6dTQAAK5krvaFzYClXrOvlF2QVj7RIsQ
pflr8H4fVSvWSbZ04fYuI24UgZBvcJHXnIkVSGe2x1QDJgkvUejM0qbrrPasu1hXDd6o0ONpZjmT
9qSTMjn6ANAjmPF3z8dHG6PfwAhlglyrxET0hWdBO81WnxtXPfUSGnB+sBBTmVUXAmvMCoCVwByN
LJP7yDTDVo5pIhxVLt45EckLMsyT6jvf5ec5sGK6i8tLmNHCKvZ19XJZ1KlL2Fy/VS/UfZCX/c6Q
zC7pdii6RD8tDmbD8eHBPvWObcQpFghZbnuD2dywiliXBqAecTiBvE3ZbuvxXA5KcvqcBA56He1c
wMnicwZQ9BhLGL3UDRmFEQmksQSgKSjKkG7Xa3HHWCMP7cbfAQ38KKs50kVFp70j/IJ20UmS3Mam
aRa+T3N8wmhZu9T/XTarrNRgEFvhgMsM5sDvq4BSaezUMgNSRE1vb4n1q8V/nLfidgQQtGnrEIP1
KSKOwcWkQgTTB9xGs+mlBHBzgnxkG/luyyVImNOC3dYTJ/DVB9JnFBs9MGfuIauOEbmwiHiRMv0Y
ll+4Otzc+DOiR7OdeuEVh0t7BiH53sHO7sWze286LcXgdZxJtPuthFAxJIuQ8Y6cgj+xEwdSzVFM
qRWtMfvr87R4QIQl27Z0q1F1FPzT6NwkB4reczgNoyUjdTcbn4l6qzU5t/QLGrqaMUoxnFmqLpZn
EvfjXM4yuD5se7zbfhueWCDs4NzlQ7O7wsbRXeuLsWUfiNuWkJCNf9k0+aN8Mpy6XdkYzl8OuJZI
evvsgWLpp4raBo2CZtWCJMvpNLJQ8zqvwSVy/0AT99qNrczpbUVwjb7zI5PD2xO/0SgFSW8jb5lA
/3rQy7g+CQI/1Y3tAo12x2fr/7amwQKPTWPmM9pCsmHrmys2dPHm3kuVhJS+2b5MPwABgYv9OQNZ
3e98HfiaCJGhex2WyAckt1COuNq5vLE5mKLLZb0zS50ui+2WWrkYzOoCBuFUOEZRqTeog2E8MDsB
loKv4X1rwMOHariSsEcGRXo5NVKxnpfOtpgMi6u902jaeAv9Gy2kx4T9hWPFC5V1z6rwdA/Dgti0
zhJiZt76uGKlNjSvnjgQIhD3GakdXSt1l1PJFdoxKnvrTEZmIr3cQmZV/a6IOj4j1uJGEJRABt3c
BDIHbaTiOWPeFKaKE6I6PL+r7d82g9PmtqqGGjb4mdnUDrHeGazrvDeiZnKsbn6lRZgPA8WS0g9h
tyksylGvtQb4KckksFzibhwiY27h7CsRlaWUY4dm4LLzyUQUc3Rebe6L7g9s2OkBzwpAuU6z2RHw
6PPU4WiTpXH21nBzORqyoTuYhQ1NUYn8qCXqvwuxyY/n6dYbSn4jJKgpBy/CKrkN7WhNRxPqSHZY
bpXjC+VOvC4nN6rwx7w7sGcURPNMG975BieBqOPROkUmBI6YsbUpyGjEurZcPZJTCHi/JhcoSFxz
d9/p/dzPw4nP+DoF7tumkG3RqjJtsya8a0WL13fyqogsfdvxdmd/lC5DMpVCnM5TcUZBKTOWamAv
419LnAF8IOnYbZ0W0NS+WpN/OKhVgK5RPjNX6iZRQ1BFL/PdHmrzsaXVgOW7uZqguoaJW5pDjhcW
THWbRjN8sGltEgroBOoMu9mjDHFJoro45kVNUkKkTyypVRfQSNi3+liVPiaKelfZokoy3q8+mQuS
isDAHvmdYZawMpRk15lV94Ob6g1eXVUDzQtmotg12LXtIS4hbH1SdzGdlmxqlE8/cn/GiAO6Czsz
TAsq18OwCGMRcgU3x6Bip15npUBYNu/wu3gospMFRAJBYyArUSpRplpofWJ6x+7GRsMTfpz5F6vw
3D1J63OHQz/EE0Om+C4SlI2nLnQx/jparQb10L/IG231K8HYqCL/UguSMfAmhPIpFOMqZ1/xg7RB
LcNJs8EKy6blNgFxzuMGEOe2zUwrIAS3NYnv9Xbgzig1SH/uSHmLtsw2HsNaB3kEw+5V1sDuWKRS
4M/qqCUFnypKEWCF8Xblrpb8rDIIKaPHatQv8O+nU+rG2gJ8N0nu6u/Wf/TXCukrldKEdulskyBO
ZyVnPHiOfNcNEC7qTTxItUdV+zD7j4IWehNfYFHN9cVf0ucQpmMM/bX2/9FK6BRJCX8+R+VE7dZN
burfnKR6lafYV7qLLyg9/UwGaKUY+tYEdNwzMIB8JpWugkR9tzYD0PpudhI++Hqdd8UlqaisT7Wf
cDB1nANjLxXfDTArsvqjYk3Vzp9eaG5WCOhmNY9FvdAUQH2fmS7ypDkQLYXQb/kujVgiVhZrorPf
ZXIN8677+E5Q8lWHRPjr8fucOx03wgtbaE00vD6Q89+QKKIpBWRW/eoxOWBOj47zbR+fImNv3gbi
WQdgCvTQjvxrefjd048WeMOCcq6vIqgazQo6PaNM8j7D+Ki6t9euK7Rge70kc425oe8xDnRZb4Tq
Lbxb+pVRrUr9HsDD/AKu+YyNrYr8ZhRWpQnDVMA0hUh1eL0ooudGr5gbKs77Pho8xEfdh2JOlbR+
qH3a6UBrtt8/ePhzTWuI2pJGYG+6TlIexoMvmIMrcmF/9PrfnSAGWgC1FASIIOAui6ar1KVCr5Lj
TzEMLpYHiePUc8sjd1Tky6iDxv3au6utCvBTVwuJ9T0xQnlRI48N+0WN3YOCcJkVZSpSzcmoiPEb
x1b1rsVbv2IJQb959x5XFanSQcowGTqmzHHCvKGza/RhEQW2hS9/IYGK2wSft8Bxs1pqADfHjuHZ
JgfxOrBtaN+jIs1ZUU4kgpFOs2z/n624E2r01YAh0skoPeAvBC3FMO+7DGsXPzaa1wH3YmuqeqAk
lAAyC87j7G37ljiZYZshGrFXS+jhnVMueWzY2sCU8AGfmx0rtAjzVKC0i0b3NWJGGuK3nIOF0t1v
mjKbiET5udQ06sW8Pj9D+piIvexPDBmstFCKw4DIguVEjLGCVU3ZdaIslh9w5yf9VVy4AY5B3hIR
p1c8Xfy+at1G7tXPVuYKTwIUh5oWb7ot1rSP+q5joe2Sl4rC6ZUxZaNC+Dc7nY4JYlmTWUkGTT2Z
PxYamAOQvP0LfvkLn7Ub4uNYtXid9+1JTvOtMUePy3CBi2WUonHIW/AiZRSjGpbE5Ok5xnXk/hXi
fFnnC6RHQ9S/frs0JnuEvp9Js0wQDe6miOy83Fpcg+Ff6cWMlcm9QHb3TmhlEVQPcTUHFxS0aAMB
y1PO28BlyegUOs907NMrZv8zMSXre23QwNAhsXuWfoudalbh4OgWmQWOvnI5ouqrGhasj0ldpRHK
ttQGcvBnK1LnNjX11te9nzt+IMWKPRoQTm/694PYknssTBFm/QAhvPYReIM+4nFfcwj68NcgurAA
eJa4zWmpaOgKe0WLkbi0RaS5uM3QNGvj5IswdslY50pyfZs643qIrnqaP4L3JtpISFTuWQg2V4fR
tPiYdnMNgfC7SBAfnNUS6kkKXCfZe0djxYZzVglc8NHKehjiJUqKkOrdZ6FBhY5lwCso9M/Or/wE
KejL7TwkQUgGbkxAtZ7+USYyyFns2F4VbPhxVxP6YVPi/phg0dKs/nx6R9pfswLsc/XdEvka/Nz9
1JXtX5vwskgs3DfVYWh3u1jmq6+ESv1BtV1OhSe2jlnsnmvEDvQYR7BNury/LIxdS4n1Y7nYLei+
mMaXO6rRYRt9j+xOHaGQ/I5+D/FYu17zAeDkYatZBghMH5daH//8wCWO7Po0XW0XlLVJ/RI1xhSe
C4+JvOEb/6beePDI79AvyHfh6gKbB4t6DHfY/LXSzmapanVvlSAgvhVdXt5AOfJfE6xNSVKOCKeS
a1qghfYhrBsX5+4YLP3q4gY3aoG7UdV5ApU5tdG46gznRNfzbOsIER98ef7KqlndfNR9Hw0a5VbF
n5OluvtEnJwVZQx+48DiDXwKL1rWOxQDHjOmlGg7c6YnCHI5F9Mhl8AJG+QNPfw217QWAg3Kl7BJ
eArSkMGcDnR61G/o5ZootNM204IChii4sXJvjFNyIznxkaSaPyRdfDfkAliWfK21rh2Fw0pwPk0O
VLDej7w+9L5pZXVNbL3FXOpQTWoaLa+8su0tv0o6m9jbbs3ZLVgZSFS8IONrve2h1/iKugsru3SG
IGcjPdpWoQk9+U5UxJVl+U4upBGmDIv08sal0T4gDs6AZXgMxJDrsY+wB5JyV7WYvnzkKCt1Gy4/
YvM0gSuI76XV7Y1h+hwXym9cVH+Etrvr9oLWmPTjvaXnfCL9ZRTxOpANv4p3IrM+FtlcMv8P8MWj
kOimoJQ85QH6822thi4ExvJc4Ye30R9F7GeDc6alJ0oS8MzFULRTMOU/bisVyJDd0XymIC7UxtbZ
1mPRf+7rDofqbRwgZc6RPt+LQdSju/5oz4B7Cj7gV7R0U2mu/iMQ7NEFTmYQLlsDnC2/u0hJ3YZB
hFwNahzyCPR1qqx7+CtNDU9EyNYSt1r8G+5x2THkKn5efkNQ/h+vQ3zptRpSGAHHlQaZNVxQ/PHO
z4Vwzq9BETiS/K19Vt92tTmf33rWaJZnwHoAJcpydShBUAUMp4HffxeXow90phU472WZVPEoced3
au9v+fNrOMsABGPGmnVW5apHAzx/Np8P/zaxFNZJ9099JZFjpMBIxQXCyPB1F2Kdoc8hNyzIfPok
nXWTt8tJ6zFMz5N9p8o89zwOhk0MJNvjjIxcMd3G7YsLoL7VL4fHY+eMmScuzSximdrglhWDYb2O
OJkkXL9HIczowA+TYVDTpjsSYKcVF8V949C/vDZwODP9loDAwAny3jAw4FX3YG2CyvuSnlkvRVJI
oEeWQp+SjEcBYjNjWJvtTul3Dwqu43Y5c5gP1BgSAz7WZClAnuSF7hN4PciEGsCtafEczTWWRjw2
4rnmTppWUuLqxXtLhvvXDHoObJrjqZRMON6xfJVHpi+qXCPcIX2zyCcX49J+Yhlh2zyaP2WW/Wt0
9x8SRYKjXkL4J05wcmE7/GkOXe9NZg19xxSxrWHY4WZ0TbdAbVSRO0gKYa3N+MtKzQq3pv7I4SvY
xlylEz+UxX2hTV/BMMuWozPoCpXIQIf5uMkLBxY5p7tqJBGgB35w/T4OeKqCW6QsHCHgo8OeDaDz
DMEl7RYpLJV2i8+qtBxRQmgOHc+hfd5/fqsfFNyfrm8rAmpZ8YhfCfow4Y6Kpo/J65Kr3uDFrcFF
tSviXl14aYsnaFOmkDtIIzGdsd1S5MxriMxQYg82y07MoLF/I+NrCL//STloR15j+pWSruq14VQH
5WvcaOcZ7KpzDReGjdEFnf0qcmiqClF/r3A7NHPPpo0/ty/uT8jTA5bh4O/v9RYdJD8wLfMnSzls
RY6TWkI9ppYrQjSmcFbLuNykv+mvSoqQ98VuQwWqBn2amJJHOB7rhJJKSO7mgpQnyxUAdQIpNUF4
yhNGBoKZ3cIjFtEwZ70Ry7V/ziPUyxWTz1qIBJYHWTBSTUMvS8I/BerDaMTcwALulafyZxIJSK6N
uYB/EmzwywwC3YUSyNbCT1VOE3g0JYPNP98n/s1jBR0AnB3s9J0dozCG4YITWsbLdpM4iY7WFYDV
0iVYrxMSNQj0rt8miEoo3fjRQoBZTiFNT2SytrQs2FjhENXy/Vzt5X3to+disuvVFgrl8MUcEQKk
DDci1V77bIyo2oxuArzkK0/mjoao/3NXh6JKXiAVWgz+pfcIfyVOmz+4FTmXFDgWcWblYS4mc/Yf
SgmVXjpSRZbsJE71igzK0/IZBYayGPfg6Q+OBdqOP0H/qb1kEQGvUcQRMtptJlNLH3SAym80TmIY
ips8SikXTPPeOourNce/LxZDXpQxUKi4w60XE0eVQMXTs/2iM1QGJClAI2p6pcnvpTCwIrviOc6y
HB28aPbLcQxro/3TIuYHyk2SBfxIvaM2qfd34o9yM//ijunr8r0V5X0wheSHHqWp63SMqJwLkATE
frmJ6Vs2RJZXC7JBiy5rh/T/i1dRXMSD5EAZZHa28dMQrvfxY+wZdAOhZDC9Rlh4DPbKOi41QI3d
K21arACTI1hCV2iCEtilKR6xnQBCgH2mUuB3o61NHjr2H7rys6L110uyVHzNUWxJuQnDZp5+c5XM
/qYHMzd+l32N3HS+7qohttIulLzbYFVLmtON7L5Ww4ixbj/1Cuu4iLqbTVKuwDqBhKOfvCmgYBNK
vIcJUTA+QR8Bk1a2sFQC6TYO9rN95e3PYmN4zt8BY5J8P88G7VB5CPhgf2Motr+N0ImHhS9YZMO1
+qATy2+pdXiXfsHgR3py6TMG9PGui/q9UzabBxI2az4rAnfu19xO4fFh6dZmMiKNWD6OEuaVkvrA
Xe+FFd4o9o2R1qDhht6dt9IDQlHmhHsdkPF7aaWDT+dRZFN+1h79R4uqHqR8uQC4ZG0h/Pilte3E
Y8OEyGBbBniEcQGhKoyngkUK27k3gtypgTwR7eEwD//vh6aefnRzrs4hKAZ0NTtTsyzrAGe9ifRA
t8n5/k169zM2rHK6mfgj6t9oz7jFMW/x4k9oBatC/neIhfEVrSwTs2tcgJFyiQ5/abow6rhBHjRM
Epb6TyIZLDT5Netf3fmGn7bUZj1YUUbK/4c7a1rIDra0o2HsOediwC/Hekn1FyNr4ChKK0DM7KJI
Cn1Du00Qy9CEAsLSbexaK9Ac6v8c7MDUNbIQgcrWzPgb97BB09nRvpbA5mcaUKUOu+iq07NRUScA
osnzo3h4d1svGLztAqWKKAgTmIu1fWTXhgga5r0zUDf6Cl/Kxk72ubiUrKiRm6/vbkUDKl81jeAJ
vhsPFPpHnKgz9phOTb/ptQNO56H22yZb0zqdpjMOvP3GqP8F37zJIAHN1cZq1RhE1hIZKpX8DZDN
y6+foyFuFBdfQJ8oGyLjZzqPQ9PXGujOTqFPMmFRA8mF7tU39pRNaFGRJPh9ZXEUSpBrBgZgyBQH
jf26/Sx/LW0Cd4FSbOZrPj4rYvNebIvRsjd4BhJ52sGFRdbyeQfNWfkNfMEQIZr2ApCv+VX0PYPx
KHTLXlyEhh+kCxtMr8F/MQftST9CtPvRfb8x8H+O881cgOHdufxV48bmx/ilhJrCsZ+bZndykfXD
2ElM+300YXnsfgadZ0AuXvk8RRGuIoWqShfNtFUk8SrbVoklPWA7o0mMQ1rHfXPxsJQ/7TjHAGSo
gshcFT6deetK/sOGpFKAomAM9cSpSuKZdEWufC5zPG9szRzjAmSKwnvv6clJPtZJfzHP2uOxcZsD
qX2wt5mVwL+hgFDH7WeXWCm4SRmJmvK3Noqs4npm93tvDeY2if8GLLJZLk03x3BWl3WgSUmW4qfq
YLDBmoCzS/MqC5Uy7lRhSkUkwo/xK9OswUUpL8yNj7U6tyJVLG9rWzZ2zyJYn/Phcrf40K/ik0Jn
0ABIoMjTvZWsYx246Jbm/bGEbuHaD1vETattQPUzJQSsIYpUtL5VlDL97tOavkcxKqaXihmPyF0a
QfZb0+A2/lTSJJS/Wlm7EaVF4ktGl2fWKtgJPnQw+6KjfWXNv0DJ193ZqjKbVKOBXtq3NfrjkxEL
su9dszTVR0Cud45T26UnHMUpRhLVmq6XK8FxNS+Q4ahUd4uW2Su2IcgaK0+WwqT36Mi6cd2Cs+Oy
urcaSBrhSM2WmmN2bhh2+7igfKyOUosiwwvbbS8LCqh7iYZjwbleQz6j5eXAahMZGOiNtES/GDv8
QsNppwCSbTW4lYQFqI2OFbOkELUIUJCeAwrCoSgr9+LOntd+lEOYoQE+CiDlr+LUo2knv3SI8c4T
t2pHH+3yH+Q5yF/skeuob+Rs3ElyA9VnApHXTG7aBEnYs0vRP7cQ19ZX/2ml4yO5U4xmEt905VMJ
57Ph5K7Iqqsh6NVh66HfqEDUblO35MBnZiSMW0eaGxcZtbBlsEdGbEml9+vl+ZGF9YOF5Ob4w4Ug
FqEYM7mbWhZw7KrUgoCDglHCXszXcQA1uO9fsDybuVROvhIhbtHaqpkaNjj6gqUXLjS3s2IeiW+a
cR4eOfzmSt4ag6bBvXSe6f/R/3/Pun4HD0Xo5Bv0+KKHRtL72o9ZOy1pc9rABJz3zO0dRWH4++bw
EICauRKkedRzlwS8hGdzcnvqcOwCSciUHI9xqP980y8DUDxpI9aufVH9D1EfoXExfteUqqFSBHQO
GbZmyM7W0azEmnzcsN5ul0jpGYOKAf6z2HbH+SLgcykL6+jN8Lzx/CAXR71OACssEAwjYZqyguYq
fkdWD4RiVvjVPnbENchsWaXeQ2G0Qa8gpv6Q+3ojsGZMWi5rnO29Ej/UHTpgcKTc5T6xcSsl9Fcr
5Vjr4ztkcf1BFRzKCtiHz4Q/gYPHW8x+VGaVOvCLUCvBY7+BAJNiq1RSwLvlhkEwj7FieVMow8i6
VhydRIsG2mMZjD3Egmp8Tkmr2TvyEqirETV766ZGxjyz+qzkYvL+un4Y9CAPM5TXj7BBrT8olmHY
a298fSUtGXVjLEau5rE3oE+0DMZEaudAfvVw2EtKB4/x7dyd7uYdgSl9XftCwi6nDVP2sdlkMyE+
KB+ySMTgDSk9zqyo4QGPyh1Y6EN+MkVWGkBRUIh3GPJESqAi/b1hnQb0oxwMbf+q/X+Oq+40YLAR
vwq2tg+gmyfASnUHs595/oUh9C3lDmDfzswlwA3AOpeAz7Q8eREs7UIBdJaXHLfBscuAC5Udj8b7
MBfpCpB7nOOLJxUmnagWj+sjBqq8zTcVvPTBSod69YMVSOWBBMxPNLAMV+rMVRY4Johkpg69Vv2Q
j18OIo65ZBzqeToxDwb8KoieHlwaiVqT0vxpVXDMObLmhiQNUpW5aazccsVwzcd5eDLaRAWpc/SS
h38Kvo1Ook2TGlhOins9dEP6s1ynGuDYPsw/+UzoDmSJebZ61OygKn3tzvO5AUECIIPFQ9zBjHkx
B8iZEkpgDdbTZC78droN3GRKtDSZZ+PEvw/rnMIy5d/0scTHw6ofr9l5BGz0VioqMBp48sbkJ8uU
3hiOkwO6sJoLq5I9BTs9F0SSFVhYfMrQLFPzw5DuNVzIMdjdnjJKPH9ddzevj4Etyy02vfRPT6ca
R1wVNi6AaIoPxW2lFhAtXL4t9Q6O5ayLMsPxtZC8BZlFvh89LpLf9ZC7sOr3+4cvKUJTPmE3EWER
Nvhq8qE3SuasWS/Bg0sEC12F/fT6TMPQytqTkUJJGFR9U0bErpDANA3k7yhsQjSfBOOwoFWiAeA3
JS2mIffyHhK4y1tSfHmCR42c1XgE1LHwPtI9hRWsuSr1c0WsXUYckZJjquEYL7ZiopL31tcM9HU2
onhFWjctvZD3Qb+K2uL0gMvcgYlIkTUVdnvidMTy5elG8DaSMhO8dOMkLHvBLW3uBMn/R1uVl/Qo
St500oP+DEStlWQhp0pPEXYUgI3TJgpIWjarZNDY5TqHkqKehSTGvZbeGp+AD4Hlk3m0fpjYWfOQ
HHpopVV619v0Bkr8ZGOYXg6hgR6M5bS5f8d3UtG3Z3tJws1RUEkImP7k7xy3/SI6WJhrAp2upFT7
PKZHNDAhtKbPo9/3dMnWP0ThGjkcfcMeQqo1zmBKSJIrYeCq32KArNdTE+FVJQnw30t7vKGrpda8
ATol1mdM0ricU4IlKZzM+Ppz1EtgJdV+vipVwgPA5TZou+o04LYyYBH4pLGHA7+T6W2PfGRGjTPQ
Ri/LNYGNNv5VHGld95n5IlOxM0WP2p2gyWRnOBoLmVfOmfvj2bDheBxBZv9pJlwmmuzS8g1M4A21
YAgrTLJA0050azdf3jsQ2aJ0Vz3Ukjqjgkx0pWOTGitldqqoPLE7cwiI6GxT6vo9lwaGcAQKetrG
jqdJXYM5ZKWK5E+A+FfDlHXX2uMHtgaDtEC3MVfo2s351CEASTgiGxa5TvU+5D7hQmf3sGIqXoKu
4uOnAhuG8h/ig/X7VN/r2QYQH3zPriUh6wF5rZPpKP2oSOIzdVUURVmbcgAJ8kstW5P+nM4fBHf7
bgEuUvBRGTkBkp7GtI4TJ1GkP1Shssl8du0N5Baf+8jz6Nq2kTXpqS0t65vNsdMOazLyOVVNneNa
D1MyD0rl1nhq6lbJWvEsXwkFW9jSANJayF5Qlcei259qEsune4VVfjoUHTyPNMFx4ecSuLmO9r1Q
XN0a9Ayz4Nl9VlxPQLXJStuhL/bBj+abaYg7Lc1OAcUw+b85CdcWlqp0wBSpSDLuRIwiVDp9gknq
JBaSdAa77EnROlWaUZ8yaT2t5PHgIvyLYSP/o/peBkU4oUgEDKgBtsbvDuHdTUvCggj7UwwvtKmG
e9GyPkPaoVC4uCe9GBe6bo5c1wYUiemxdBKbjsxL/tM/eLTFJOIsiVLXLDq2SPedDy7Gb0XrfFK2
GEhOGHv+d/QlXuy5nbJpJH3mWW/H9OREJGehCJ5/CZ7/TpmEEpx/WBxvQ5shdPNkrBCYQ+YKNJMR
b7YMj/5eyP8oGoCulFIgKtCcCWF9wnCn+zJ7Uc5JKdKIj6zlMxRZvC2Q6mIHPXfWHeBroXH4zD4/
0OefikOLVEdzo2WjSH2rf0Fu5XdHXCCChqrFm5hfEf8RAWsz2CESa1fpgSz8CAmMdCTyXoImkISz
F4t22/KSJ+msp9zTZEWiqMxL3+S8hg+VUQTgm3mu0x/Yc7PaiWsqIMs+eH0s3URO6aIxZKJijs2N
ZQm4d9DLOHTt1OKhEc/lkKrUNFAYeoE3CimeZ+A4VmPDPPzsrqhgsjoVSX+89aHUyV3X7XEMhmRe
vsl5NN70xw9i90sltnxz7ZauhXNwjXSbbYLyVmGpLy1yO6tTR/VajpOh1MYIBfc+sdVkjsh9g2T3
REYXHDinYH3nAKWv6dCMf5XrXzLu/k/fCHBMfgJAn19CPbjouPg5azVdLz24yMchBJRlFEiXopNF
PUq1iQ3C0iQHfmLl0NcbVwG3Ht2CQUZIMC8cCh+hzJ9Xj08A+9l5NZcdrnKcHjQrSUMJk6HEcwxS
N4dCX1muUeNc5Am+i0kxQJ3UOvq4XanEs6etQUMHTR2UzvRyGgAJIfS/j1TVxYZRvW465J0oWBzV
w7DdqkxGcn0lyKVR7njJcj4s86WpEmW68qffEj+rkIE0bcYqE0yte7EelRm4cS4N2F4YCNdQ8sAg
Bl1/slpV0d+mV1f2nqEfD+LuaC8iXNw+q9AjXHkTvG2i9nHt6jjVmZ/239S9kvtNB5Mz6jSAH5Qn
5DYVJpGWRJwdkoJZk3l2C537tbCrMo5dzSzqCRu4Qukb6O2OEIn+8IcDlgJ/VR75DE3gQF45XEfd
dNSa/y6aGNlSmvMSno1YsZI2Jv0IHwhmRZEvOIoNRZ7UTlmxMid5qXZC6ZVgqkGjKThxQtS0ZhQ0
wquPz60QPN5CAWlRhOvq1mFK/IOt+zdGaiWX1eeyW/rh2XkBiR9A9H65ImhStC5lQUqtVHYPvE8Z
X8pRUUS7uL3aja+VEZhCoiJFheHfmI5A9Ppdy/2wdN6LZra+UCvth+1G6h5EBOhBDIiL/dYQXth5
FKQ/N1IDG8AyDMp2Mh70bl22sfj9lZJqHJHmU1oEf46WU8zExXCqpv7H9y5Iwi1Z0/FFwDJj/reT
cFMkwEd5rH1kaCCfxgS/EYAEXAfgDLwb/9Edh4VAY7sYCmv4mntAPO+kUnajvqgBEiHgZtvlpMYH
JZfwb80ZqcZrbrH/nbMM6JPiJC5T2komVO2UDmOp+KZ0uM2H9eh+kb91o2HPklez3+pRqZ3pFBvv
ImlvKJVQzIkj1FMatJPiv3ddEJl7H6xTH8vpp5Un7iaqqIFDDM3As8ImdtXcB5lwRuCrp4cqFD+o
QPjBxPbP09/o3q/LHR7hHx02J9CfyCMXZN53/S+O4JRwh3UGxMfnCj5TTxnaOHC2zb+DVmgmLIhp
0N4yJV2UYaqp13UxmNNBMyL/3I+HTwMckZQAlnzH0sOVI+Rmu7AbojnXIWAlMjDB4p+1rvy+iA8n
x447F5a3s/QYN0kzjmw+qrFTruHyRQ+ZUrjkHQx3GuuDnfb+S2hwxRGLwJTpvTFaojB2zFojUsRs
9wG+7AEDgFLlX5zNrbrItJNZF8/5U5OKYa3d70SFetkTsNcrd1n7fUlC85KPsJn3cSpFqQ4185pI
GZejrrPBBz59Qnt24oreiCxVl5ItQXxtgK9ULO+EqA7nXQohgHhwbqY4FAzdRKcuNphOCxb5F0SW
DJ/4I5HV30z0AqBnxjaIvBVD13wEytTrubXAxpAVQL3d3FHldHmpT/r/lVA9Rof22IpuEv5Iw9/s
8abmNhWPaO3af2GLEWQHg+IU2jGVG+irTpMPTMP1GOT3NOMf8tlfGYgZrTdTorbjEb561lFDNdzq
M4I1sJMGc885lB6KhnjKx5YlRb+oXWEC2u3HsZkgKNlBotn5usyS9l2GgNV5CkohiqSOayyqRnw7
FH3M3HwqDFW1YqmxFd27JGi3txEvRTizzzE5ztt5GezPI7Zwdu2BKv7QtWDJoCbjpLB6gymeS8Wi
8tg9wpmRORW564J4I3nW4U+RoaCnMTHxQudIiZz+KKj/iKV642RrjNgEoduPYBLDoJq7eeh0gpYc
oiXXoF0/c3QNptQYcqj/RgwiJmqp0q4JooU6uBPUqboACB+77zPQVfI1nQl5D3nBylTUBTlERPhR
K6sEMnJze9swI5T/StgXOE3j6s6apVSu/XzdmArOGPU2Jt3+ZuRLe9vGODRAuYRTy1OmqBM/RznK
tWG/NkolfDLRzKdFFyzj243SfEM73FW65oDdBhARFxupALIRc4q/+Y2CHhMvArUurHKbbR8nx6wn
MOsI16JMWssjRppvnx1H7I+2qNi2sEfwVbzTWgQsOWeP01W3LNjlNGGpTUK4T1mq7yRirmvKgcwg
2r+m2wTNKyclHZ3S9NCLBsH2gFwxO8qc5Sjb4w2hGuExLHCLK7mmAS2bPBgom/nhwz6s9aKVz46h
GKI23DTMn2dE2djgG7WtxFn3oGF/lTULfmaoHlTAKFQI1SkY7YISYvLfMnSZlzgPs3V+wFx/X45X
GieiqroXvivsZWSpNbyIRlkhfV6TcQzEsUXoxEDIZEDao17D0lgpc0ursUuBYAFVT7YvLF+zdeEU
WX6hNXQLp+lmirwIoclDdi3yg+Wo9kxP7TVnxHQLVugZXEWT+7Z3zWMOObL10+ZxnJHpdXrIrxg+
UMN400Di+w1YMkiYy7355gjV1DT2Yl+rb7E78A15A8Z7zdO9PHOR9Q0UvF+x+kUvIxYz3sbWZXXT
R9I23kLXCok4GRcCG2p8ffNWAypY43M4y3hCPW2vM0fyLlLkZIH6fvR0Q1PiL2TVqGLHXE+h/nGL
/XZ36K0H5F2kTzjNlmw7gFFRksXbnhjL6AKhTo+5vIsDxCKk4VhqbPA4uxYg7WHYhgJW+p3cmSN2
2mS5TXpBsGjhkgxEFbxYrDUBbKn1om2mNapBQOingEVYlb4YS/oCG5qrDKESINTgVN+SCDPXDBsM
CdVDxXvbWq2CWJcwY+A+ROkah1IPhrDF8I6Lhv1kjbJpqINgz3gqWt/RZjmRzpsJKQyu8WcrwbVV
0M1wgQpUzLrzP/hOY/Zl2aH3oGZgoLtQF5B4Iyeb0/ZlnZ1eOI7jjiXFHKxcau35qvTJlHFVynxW
z8wQtJd13lHFbDU9rI1vAaBXNIF4xQaaAJBtcnGE/vk7u/OKzbhTx4yVNfoVCf9BQTYkfGR6mlyX
lXNahWBLmrLLaQfhtQDWvFDYUaKUSFmDp8Q2P7GLecBvBQCLKxtlw2tBWWAZ4HwtUSZgG0Fev7T1
w3GmGp57LcGbEptsSQ9+Z+L0s9dLUbsp6uJT3ZffyujIdcezgbsk4YwLWoohsaAe2g8tr3+bzaCe
vFWacEY+7jFd/5OOIueX0V3Lp9ZdeSUNVxHxYYtK68yNVEHxLCpd9qNxSBTSAdyd/I7AD0VtrTt+
Xov7gKnTZXO+7eLSxXdxn+O1GVvq8zxSPTK0fup+Y9aaLvvF8P7N8nYtSvr6KhBkNJQAECgwwl1k
EDYr8iNZGKsxZd4FvjmYZipFmSa9xmNfkp3vLEaIPh8XjhB2fivI+UJ+DvEhOXzqWooTX1Ytzsuw
o6SOMG07AT60tGQ2fNbH0erabZKfodCnx80R3ak77XEiy7wfeb5krDHp6O77cpl6w/iNPNiS14ho
2CuzqZcwoQ23LL+w+R9PJghJbFTVYWZzTwpYRnwTg/sNs8C8I8GM5KYCx5z1MBfepAiKP66K5Q8O
kkxckPIqiRjgcQ1ozulJ1U5rq2L3tGqv4rlJSkDszbAhcLifZ+BtTKaQlVQfkLQbOd5BwVvGly7z
/00qURyj3nvwMa9N40V2p4LBw/UkjUBM6JPx250PtehKJu2FkqZ9+HJdNl1ZB/EELqMX/bfZNO2f
6bu4Zm073MlBTBNwosGk3RvGyyFrdC/TntibUAVEvV741SVUyRncKewa0zyZ2dpVKilzqJuFT4Q4
U0V9sgBi/rID8DgdBSG3XlXAOEmRLCd3V44n6hE2Kwh44vmw+vbok/E75MPa32NIQ4iPjVA3Elxx
o2nTkAV2g0PMNEaOZbwUdTvdGbDymKgtuTC6nH7v7tWR8KX45P+FXf9B7p6+BYGCdh/XchM78+kU
pyeai5KAWnYCKLT4llbqNhiRqnmaNE0cNXgWT4hFV6+hWzcl5gAxLszyt/CD4xHuOVWrsUYI21Vl
4eHcfTWJO1Vj1c+Zi6nPzvMDpZ4fjCoJ8Ox/AT/XzTuGy9MzVfR5GXlReo6/w2wN1v3SYXZn2Akb
9BitYCYc3yThpelXZPigMTy7dM2dyFsILV1Oa9yS43tAFi1ydGxqTqXyrU809yWpRmEJQKo9lOWJ
h9tREhEvT0ctNFjvGr6/TCAHibJIxBXNS/o+fKL9ZmImyMvMxR9oIR5KHv9bCBphN1a2tbVHicO4
SuiL1LDTkLkzSX5JnYTYVnJ32KXAi1TPRMRfh9qkVnfg3+G0VhD2eo2s2CEj9fszeOnBDslpMqCE
YUGVplsbos4pcJw/vf3aunHYpvpOVJz94sH500McB8cVNXQGB1EvWMZIVWQVyNioedj/wLhH9JW+
Sa43QCbPoe57cjpboiZIhfIHLhLGbge624VcP33l1H1o1pOaPItPtVQm2ANN475ZE4W/YvSQsMZ9
RpFaeRFxhLGZePoZVi1J86uxfDYnm+Re4Jc4RQZBzlFD+19QkEqfrkWWAhp5HpF5EDuuPCLa174A
8zrj1qisyF1DZIbJgF334zvGRyYbDKcsafjg2qKrJ32CUMpQbVsQedep/fRB/nLlG9tE3uRQMcNo
CyWJdND0X6uijnRMeVdX8fVZqHYjaYKLMN2a0GTftgP6LOwJUehE9lG90S+LTEied7bZ62q4Rlen
y2bM7Ck5s06ddFRp8kGOPWAFM+q/KFYpU5gXOdgywLXxLWo4cKzXY8dSOMq5P5vDVyhiXiot0EfI
Billd7QEa7q8SH0Qs4q9Sgx8+aWjxcd6BQEBBPhnrzZHaxuC6I3dgMeck0f64L5ewWPIQsz9Qlgm
g2uWZlyEU/lyLt6/+hpWJtGpYr76A01mnwYmPa6W95eFRy9LLj8d5R7e3GHdUPzzOQmx0J9tiDEn
SDSqVcxdUazGTLcNW8iY5kMWFBB4j3WLwOapt7N0QBCt9WUet56IpGE+Yg3TcZj3Z3GoswDbzCXY
F9W4k+48DKDDuIAmCrjn6o7LD18X7gDh8cSEiJHFi+DJi01T5AWJExnfVomtXFDbvzhKj2k/aWIw
rgb3e/k9uCSnYJHCB+D5LcS0kpg6Pw0KGsdsTgmphgJOQsOQMC3MtLie9E5T+NoPj6oZ8nrSS9r7
sMJKogrTfKU7KDGHPGG/dvoHI/NvJIbfIpvz65xC+fh/hQxRbAFhr6rS1svnuT3f5RVHWXMUsGDA
/yRO/iYQkkpq7FymdGJAkJWaUjpOGYJKnzYdBrNE47mJy9Xx3jXXJ8zQuJaaDsa/ErJ30V+TiOn6
+OFfWAvrzotuykx6n6cIGc4ut3KLS4u3lQbuOF9hpH3obPS8guJDAvSb49Ds9IypVVAdRKnhqcz/
7HzzWl9wRddW2hctmihUTBfF5hqRrbuQWTutGP0DJEdcFMwSV/MjlZiuMxr3QNMV2casfpOBuTTC
tcVb6iyRfamcKqf4bijUWNPL8fMTGYI+erTEE5qUJqZFjM3UbHyjY9ZxGPkc8URQScZt63dbC7M1
2kRfyNrApa6S0GxJ9V1qDqiQA4TENTP1IvkU1PLetjaR+tADgbwtyieh88Wz7cD+3l9LJ6yhMLdX
8V6mfp6uwyOTunChwDBU63AvT3RGqlop3RBVrCgl9RBDW7ENnxTqXxXq7lI76vuvQXAIg7xuY8ue
XaPDNmo8iZtHp+bZ6Dv1sicYM4UBbGgnlEVa5GX0YFiKNW6e2b8/3rUQd7jiWrug4miRKE9Lz89+
DHXmWzp+YnPD9KqSr0eXxTZVcr2ZsRFjRStzuqx7M8l0wKKzcL/ICCZ+ISaOXUZg2kFeC/TSjglp
Zqe/dV7KwRASYYcrWu1PCAjwUDj9HI6Vm66FwQlyNdp7I6ui8ai+pB7EO8QJpzzpcwdRIYRHYCi0
WJdQfRgNdEi++q0s+6MweeW+wmWkZITueJA3DgPNPhY0NwdaknxJmjFdn/fmUHYnWTsqMKtj7IsD
tGWpxtLTdOiekh4XWToa4di1OSH0ZAk68viQS8ywDgDbnckSlh8QydrhuLRnjXrGyUEvsG0XdyJR
zoMo/Ruup5msSlv9TMxpkRSoCKreZKeKRHcXt+F+P9sOVsMgjkmZ5HA3dJ5EaF9AlYIsoElWLmb3
9ftn4A/2eLCZYxKRq6HQ1vJ0+xmZ1vCK/7wrdNOg5Brkaz8APSdvoThUtgfFWKowHppI8SJfCkbF
ALzPVZ8OH0otPPl0TsIQDWZbE02RHDAWyWH0OMzBHHxV/Jwxx4+KPCHUXK1UiBSg81gkpObHvmsD
v4ftZZ0WY3rPw9gV31HOmPjBqsk15TS6YbasJM49+n5+/xfGEWhTKhJbR8zATIxXl52VhjflgDbK
OU05mPk3n/rNw0zKwoJOFBV57WqSPOH6kIhm5h8pCBD8GxjF+52PvNgHFmWm0tKiYknixtJhHBE9
lEXrBB8jXHaZreS4qqPp9piDgMYtFhEnzD7gYFdT3mjkdzhU1wGOdixlqC0F+0+3yu0sAkUY4Xa4
MojpEYGMlvwY8V9qVqVMvDv2hu27BNYKZOyZxwLqjodJVuEyf8VjsAc9po+GOpK2PeehEt2OAxTa
fsVJqx3TdkdCxgT/KigCeI4IByUmPAJAyFymdEdb/kcViE3ujmZ60/GRDAU3oh1qIQosHfd0Xx3y
nXhh3Evi2ZLPi81Ha8N5hZ/ztN8jCnV4aBna8W7iQf8zs7KoVsJnTAqPuM9CzM01WN0YAg2diour
j38fqWSFmzpbv3gRFTsjLfoqLuDMowP6kw6vASdBGBAWt8U30ovizHYM7dFE18HP79G74UCQnnDb
TZidD/w+wsf0dKo8ukFlriXav3vlVz2JNi0EP4X0QF1dyr7c9EItT+0qnU2cQ1TvdzS+NDbq/t6y
GfKooHRD8U5WSrVoI6UcXtl4mVuRdQlGjFI7LBtdmb4Gu4gRcTjMgIsSktYNxXqKH8dh8veI2dUJ
uTft2EtIZnCWUTvviFm0za7T6irVrPNQwVlMuhXE/p2BTExTvZuBZDq9O7WTUDsjpZPvuKS3qhzd
Mzx2AKYwRHH6FWgLigxbNp404eSCjvXF9E7YqXJju+NkEn/Omm1sISs3u3GU/aa6twwBLF0lfkiW
FPmrJgRNZG5XniAkc/9KfEdg/SFkQjZO4zoUGszWhh/MJ+Emam5lulbtw8hfDMZ2DaesVWeqZ/3L
AOppoTCx+VFynkkGemjYrVjKP/ch6ucYslVq8oISsYD3y5pxQ6vg48cO4h9h4hggC86yXfGCRR+F
n3GlP94kAT+8+zWOnUa/Thqq6LwWrA00zR07KYThdn3AzVsNOTC6IUz8pJxf3t8aQMgecJS8MpcQ
PWT6DO0rNvFuQtfv3ONvceeJgGCDTI9xb107Sg4EXoKf3TqwiLKvcgjSqWZ/I88JMnmR7EcqdGD4
dnS9PEr3gwXKjYCNS4sft+tpvVs8Mnzmn5EsZ44llUAo6uoiuUmh28xdN2QkwbBt81QFyK9XfkVr
AmBi8mk6OS7cVFgkUoL+e0NQslhQb7zrocAx4QwZfiGujNWTE9an8QmVScJCpK1u9sIt+D39tPbu
83MFnqf5ujvcOkF/XOKYJpvVq6+Dxp1XQP8tpLyG3fFfY+mu7CAkPNwrzSBUEQR4akD4p3v2VtZ4
cG8jV4J6m210EtNVk4kRK/DRZPP4px8GAmmWfF4zdYWhXpmm73+VIAtEoUiPejRAhkAFWLrAfuKl
SV9Wx/iVAEEGGT+5ciaDxXCBVfuybP2XXTpeczZG9t5GyPBuR/KZADg4tBxTPyS30LZ6pMQOq2ak
/0BHyeAX73sMNSJw1Zc8hBnLBH4sJlnk92DYesOQU5xq2peAtl5u5gukGwzkb4eYsKiBaZoH/qhS
HHEdXpNGciAVgiics4GDcrS0UG6/QGM4Nfk/PPSD/BDMOnDwknkaFtY+FhEWRVjjcT5g6A94+bvy
1T9LV2mEkeQNXDCSs+GnDB7oaItm61dZ+veM6nds2HSOWyLXf3wA4e10tansob950G5mtXbAV57v
mw2ueHa395TTXg/sxzLsZ1wsb48XCQAX0vcdSlVmhM26I6ZTcPZ282URxith8uoFz8v88k9Ozgve
GichaNDjZV1HZMu54DmaPa2RDEgx5b9DrqsXH6qH2LYTfLIK8RgE/twHv1Jej3Ol0OeIyYYgBChA
a5AjDYoVZbsPowTI5LEU16pC1KNALNplqv9TYbblhO05M3RfxLOcNREbBLbo9q1FuxfLXjKiWIbr
RXe7z8q6oP7NW2GnXRCf41Krg2JZJpnePRtJBbAVJv3pnaxM8zpzWc2iR5/v0L/zTMf1/4SNh8Ah
eTieXCia1pT2K6WcBp9eu/orhXJq5U1UZREEL4PrkxjSk9PkaTK7cjatSfrzK2sV8SpI+N26qQ0g
PARu5SJ10uL9Y9oc7EN9inIR7pa5i2rMQ6z+vkTuMyvLMxItejJhtIB4mATC2bZaL507Jow1cuQN
qXZ8G04tiGiPmwysmPYnjTaJ4qvWg1tIEjqc2hl42AMfl0KPxvkNPebvIUHpXg92lXPijT/SzC9P
S7Ce/6UAQKOVDNZHuDNNaH3NdL+aPaBOhptwNpPoKn3OthQjjaTnew5Kzuj2y/h2ai3e4QaVmSfF
NOfB1FsCcYClusKGUdS17kY408OAXGBc59X53N3RW0CpsfJmM93EZnaZ+JrcPVbVZGqmt2zIbXxI
37NwugoGyPs9zpkAbnI8/rMxNVk1pEbTtBQw3E8FuFkUHSeGpT8GVjC8+p946ovPdcqMFoS4KNnj
fHGNgjNRJZmAL/NkTiIWkvRh+zbRLgJdOfyTCILKgLzHwoIoTq2Iz1niQ2W8DJek9VMoTiZhWXLn
zMsr4DhxI/puGQ7wwF3aJCYkY7+pH5WalU1e8x0M/XxTaM+iYjFxCk9L05dB6fWKUo4XK0g0e2Xn
gh2IHG92zYrDw8fUk7eRo1fX6K6UbzU+BcsvSDuEoXjfb8mVVl7eakU6M0azewDgtDlVb2ST7Ci8
W6WivRh3MpGAAnEIfiXbO36qfBLVI2fZHet4pEhRZYzjuUvpvjT6qjqh8COSVCq4FB3DAGhJUec7
934/hukink0sNzLeUWDZu9mtuc1/OxE3dJ1XtOT39ylpaP/Q4OytA6mj9us++FBaaBV8yZTBobJv
sWT8P9x2WMUkWznXGHI9Mi7md41FhsF2Gvstne1puR/DAWhle8H7dNePeCmznBpcMOOqx3Pn+WtL
CYv01LkSHxaNyet6lIv+GrTwXR7FepQ/6I+12P727lOOyYwYAnX4fiXiwV3S9lRKhGvPbY+i4wv4
dlk9SIEmfH+kUrcFkBkphSYqdu4o4PfaD8qA80mgY7yNvBixwNAHOMiUVfXiHlCsMHfvgiQxftTR
1UPQ4c20ndyLwMvMzYERaFuycmwDjDRf/8igPRjDKNwjtD4S45vQy7xL0dkgK9tUJkGf/SrGGIx7
L0k+nASMIKvswe6o5rKqABOKSkmiGjG0a304X3LMNS+0tTeGY2NS0kiu8EaF5SDO1iyGmgnX7waT
419y+pqN16/kQr06D7reuFT3IwPV0xHVGTwiRvfC+fy0Y6VFkYtEWpnRJ0CoSghe0wk+q4t51ErM
l8Tv81yelpFmyCMnwY2v7ucSUQeNpNWPfFPwSfPwBCa0crzlno7Ivl8psNjJduJ1e4d1UkpD3rZi
DLPOXMp2A7TWb1dUvnj2tZGbjoJYQWruecGqFFDUiEDdQzIfEo8JtGVkYadeAjJHsSRnci4nG/v4
00LMWJkIL8V0IqTCx8UY8CSu9fFS61Js6XLs6J51Hq805dwXkAYzQ5SjV9NvI21iS8qHjGGCQtI/
CYN9xLBdgAtAir4Tkd1r7qg5z1grYRTQ24aFWxo8W7rthekECgu9RN2gnwxsoUYqnH6x4cb8Jcie
H0MJa9LdWfdYW7CPj6+Vkoj5jE+WCkT0EK5vcBoHvkS2a44hwEpYXuBzyCWT0QdCXU8tFbQPKLA5
/ZSVB0UWSSp9t2K1bVZCZH8e5II2FI3WFSow22aR0GTxAaOGHDBX/tQGlqWMFJ0B+KviL14oYhul
eKTrICrESP3ku15QcNkQWkes/Xv0L1BmDsd98QaFJ7Rh69fKP4BaLr4nOzWBzGdL/0wm8tGCsBQu
gTyr4zCW7fYHkSmHdHWGUemcftO1e9HAvp2tkaZ0VpQmhID0YnAMWWlYchXFkUKgIUBKuZ52iZY/
IKjEqGHUn1IArpsn3XmUWhBioTCzWUcnCkC6IGO+2DZaHWmc8wjKwO2r8wbamWfi747Xp+h1Q1N9
Csh7D5M5TfTdks6ydN42p0XKd1DRvdT6dvcqbdCN9SPMxrJN7nf4M6Wkis5l0BiSApF0VPfFS9GR
gDWD6NRmI8HE5TK7WBVX6JM4siKNiKF6uUk0HAu6yc4UJp8sZpdt+j+P7JU+H/sAucW9ZdTI60Vk
68RSZ8d7lcDXKvnzYy/nr96adSUbemlcHq9HrGO7XzLDArXq1kkXxEjiO3I+2o0fYC0K5ytaLfMU
zpnOu9jRCatidCgSwqczZ7/51xGEZYvPqRSuOeimkCAnx67g4zxboiL3wc7XQ3XVw5U+PokJwcM7
jaF3bV55n88xfPoHXRERoGDmYFZlYNsLlwpy0xUB4vJOYL/hjXSsvGyHPdHseDgSVkRLhc5tzyaa
oVspMoq2tI0mkkB5SAaxjisp6AHlr7N0K5CCUcKUuoCetI4tVQpjFxU5NsokJbXjeRQ7qzyq+QMZ
XYSo0FCFfqxFuNUl1vx81VWKoECA5syDjHPiRaEpDraHDeqXHXEng0mucgPxyWeSDXu0IvsLQuhp
TBQ2O9bZvNEsetzrdDeb+zRjwHsqiuc76vlduNl3bcfvxiKeapO69BEikZqGjORAmeqecTMhMbd3
EYNW23f7f/2784q48TaMamfvLHw6s1MmTu8kTIP0yR69ccEHvMlBdIdGsUEZWsYgF9ZPu02FTSPO
wKO2/ybjME1WdVDAG3ZMNwY9WvDP4TYzmdoUy7ycolnn8ZEIL147jYXS2rDLoXEsiRgzoaVK4m2k
agSu4Gv3nYOSuldo1ricZH2zbHfEaqcjIt0d9fP0tJL6DKchFlxDenFkTEZejRIHS0kvlVPRShyI
kAGBSizBcDLnnZxkGyLXTz/O6VLgLq89dxLXi/+PDxXIUYA5l3iIdTi2xdL8NG2fJ7xtoGoYx8oL
B/bKbklEYMeUurR04J9ZdwoAF1LYkVn+qrUoCqfMD3RultXToC0ul2J2T84VkJj9SP/smRQW1PBi
o4ipPNV7GsRLA3aIHfK4FkNHbcK4z8K3XrJ1FLM/Si2ijCcg4204/mRBP2rmkcsjO8SyrF+YOKFN
S69m0gVL7qLwhDmSNE00R4nVCgDn9W31LIhr42ID3daEGraEApx9WK2S8J4sP6AVXfy7Gc1ZBR9Z
M17iHOok2+8ZUhNMnLgrASvykzI2MqNNjXvmUmGKdclO+2hD9Y5frmTB2ECvd/n61e5LXZofvJxN
7m2/PccVa5O85E4/JKnyoHOdinybJjZsBXrJtjoSpKBjSxEkiykubtpquvz5+fB3HpdZuA48hYXn
l3C8yMo0JGIYUGpdQZKxPEAc0kqVfetIwJR91E5WqqIIuULuLBOB1/P8ahqjeWzLkwyUyjMoCg2y
12PNv4RqhqWRErCGjdvzKb15oms3HltRrOq2f0dSzOAyf7by6zbkZqV2Iijs2o9O+SVu14d0fDWP
0M50jHCbSAsRS6P9hsSxCsumXN0PCEkaMp6NY2pafPUfxfqoJl5keMvoanfwVeeJWLoGmZEiDh3g
G1lEvvpFgL4DkKbfkcJqNtqeyuFPcrha31FsAol2/Hm461A7t483tXLUsC6BbgPDlMSr+bLXHPsq
LsFIdGBrp5UReJbRVn1QztVqRoH0twHouR6oV9GgdHMhcXcFMhczv49XzlZfz6M7dsDoTQMTDyep
yXKgSKFdY7xRH0OTQm/+SNmzFjh+uUpScBM1xNUJdcvNLRoXu2xcBbnWo/IEaruRLSUxyRUqflVH
xW55RzBG+wzX1sPPMlK5I43fvnop0fDCV6NTDvMjDhqa6gOVRZS27yraxP0FJVLtMf7fF3nU1RMY
dHeQSVWftW8pZvOlDajQSBRYA18stJeyvbJzOstb2bMXAXL92yVlSLg5/382RIIGCFZ/UiVW0PmI
xnLM7X7wKBVlQBiPvRWxjIzAkkrQVi6lAMCeJPLMYsYcPV1Ptx3O7YNaDaua/DwCtv6C6wu78loH
Se4PnDs+5KjoG5iyOTGhGCs0dyeIPG8qMBggi9CQdHgH3d5Yqqb7jj+qfkJLRdQi0gsw4IF01jVr
j3KjPpmyS4l2L7IZ6N9tkAW9cdIopragGkKWnr5uwV22EqA6OP4DWA3wwAOkYbt4RNLpA3RM6qFH
AJgIIzk9cEEG4wYOTb8xzRMJvVqSZ/bw+f0woH0sGxlLMgbqo7k4l4rZFuR+oyBfOEmH+k9IQpSB
QZ5UojNYteXxk5tx9IM3NzB5Tf/Gi5dV7lKkthkHAOFkQiQ//9Hn1rQSH/qK1t4aviuheRujs/Cd
1Z9Keast/gzRbVj/eWyhD9y4AyIbPwxhY9GW6HVa6SUbN2ESEMlRezbMBOs6LFgD9UxuBZMUVAGA
J5u5FJm8L3hqwE0ENY4L0GLn7aM3YAVxMKzFizTCDFfmrzD9oglZ3bSdWK4wTdi3SbnHiVT7x4ww
gHEGSdf6lkiWBiRjnL7Knx6UH6BwztbfyAfmtE/AkySh1lbk0vtWeIeLQqRPTBP25M5TA9PqYzMC
mjRVzPqOz9UDeXq3WYiGiqkuscHzfk0yCYdSQDn0aIG3EwMS9LK1ddRzNw5WSY6oazQQVdjHftnX
NzBgfBA5sIL/q8nFmkVEL2m41TiVH6FqzwNZXj9nOsED1+q062W3jT0t+V58k/6O18/xx7CzQ+z0
5xxRNRjftF6UqASPOF/HJWqBCCYt/hSdjcxk5CANKseEurRKX7aWkCL/dFPX5cTp65+xBh7FbZi2
seiBqg/MDc8Sz/InaxqrBp0aNUQXMbREY3+SIEbbCXDiCPO3Ra2fEXkSfWl5vIxiiqsoaMC0N47/
hT1jy2GXj4CrCYjWlDCszpViknE0d5RsPxkuRV1TVK4wPYy9ewydcmqnHzt1hMmIYdMndkN3/5AM
DVhDf/VHN67pbrjnywplVNPECSyD1FMm1+wQYmaEkyK8DNlsRn0l5D2UrFFWbh2KBwrqpaGIp48C
VWj+nEuCe0Iv8WsFkm/nttKNPldKwkDgrnD5xQAwO2I+Eg+BUhB6BoH1NjiNi0l1kKlGlwmB0ldL
g1ELK4hJG0+Sxj5Kk3AZrSRwrZeTGOdUBUUiymW/4jFzI7G5EN4o1GtpHTRuq+4bcqcDgblpf/Yc
wl097qsz4OOMikghuuUVggPap2rj0g+g6HLlqfTHslKgQFjXAEFlKMXvDknPveDSP5/qDVOuS2WY
QOBvgIHHX7tfYVCDxsoiFU3dpQhd7TG1N80116qRlFzV/Tes97yKmlCFO2yScNK3DueaemtCTe1V
Er+vMTnWCJFlqDy8V6GRqazC0T2ghAoE3xR3tIlskBSggoM37ZKiN9bAFWOTNHuES0DpMwruMbfN
G//fEe44l3cKpyoX+TD+POyJ+Fx0tyzuS64fNvspSCZ24iQSx64+fvCfpLQGTuD1mmolAtCxGFRu
mrPIqZRNa1GdsycqpHOABtskJUd6u6zwe9xBiuERqTNMoFDeubm+1uKrTahQMu0vDOJeZi0cheAQ
evSXGgLXyMAP4J4JCPa0ORKKip+muDnBdVi/d+ncdZZk0YgbP8QI8n5oqnDIf5xzVvQsd1OuGFAm
tRib/nY5Ju7Czzu/xUErewYhQf8und/xl4O87c64BMugu/xBwYkAAOBpJTc3j26iBaZke/9GoDgt
vGQQM+q19QdLaTDwzDXTwGT2g4/meoCMHfDbriBgaOPalZDiLPMiNlxKcBBiYFozqeuaQl4sesee
2Hsj4ZBQHFsIFrEdUK0CwFrmCrwA5en+J14HMY+UbPaz/6eh0G5Q4ZgeoJyNljIxebS9He5cAuX6
NpTS/2GVee5NpnjS9QlOPMmr5FA0OlHG85xBJVbEskaC7YF7kLe8jKlCd4l/dBRAMPVmDSceMRi2
8s137362ndcV/Fa0ymbtLBCf550kWSJ8yREaqNhf6CEBeh/eA3IIu+wtpbLnszM7TIHyhpbLIKIw
Y+yz0/igcEdfu5g4RckD7AZmAcm5y1mB9jSVR1G2IUTBuq4iOAs4w5tvIEhD8cWtvQBNUy3N0yLF
//HFYmt3jfB6P3Wehr5FoYp+UWjspNMxevK1B+7l8d2iKiwPdIM7DF7WSNibKWRHo415s4ScqQqZ
clXiQl1ghjaXq+hfbHAjQinCSdavlP7gX/zPWV0Ny4Kd8+x1MLQqWXeTedPSg2dD+2Xvmd9yQBbn
4l9qu/FxuqrYBkqQeQEFvqxmfABwbcf45HyaT2ji1niEPu4ehIgd3UhkCekPC1wMbZ7po7kwS437
jinZWt8sq/hhCvLVqt+/sOThfmbVyo6i8rGqIlkso5MkOshksNvGOEjHMpdCUV5/GxHU/oLJskeI
550jcgKyx4p89qMAGTBly9NnX8bHCpK7AqZBYQhMLm+JH0OcXk1l0blhxo8as1BWKP2Ky6Ty/+Tr
RgBipFzvLnGd3mLs2g4q6tjmYsVVpRWe4XK9YVm3WSE7U7qNTbLlsFcvYJVh7H4tramiWXhvbplX
7wlc/CxKEniC1k8GfHSAVcMbaG970pW/H+KSXLhxHZ7mh0H4ejzE7OFArd9QqRJc9e0qB/h44cNj
pJ74Uy6c1CmFl9y3oVXIEFEG2dxfvhgfJlIOale5THGyJ3zcitQMBEeS8g/M2Rqlep7x/G9SryJM
WWr3UMvNnmsLl4okiK34p6nA59vKSxF4wb84nTndwzSSMFTn49LmB43XCcgZi52eLRyRvnwvOdgW
6X6R3p+JJkEDm5SZiM58TbZhMJPbBE7Q4y2LpoQDzMno2GAe1Z7V48EkuwZlJhIaRZaDpOOu1NEq
2e+xwFOW71M67Xe1pVaXJwWCnt6iMx9JEU4TCqyV3so49c1gGyBgpzU1zLadxqM1KYsVsVhmMBdb
j3wC5zuBtZlu20cII2GuAGCZIkl8PxidTsBxk+54RonHcQg8tOUebnd8GsYMG1BpPsyfczXKvtWE
Eq4YL1uIayPSyJkL15umhZhCPBJTO5wiKiEzhobFk4euHag3n+toOTsWmha6/yA/iA9ROi5l623r
PBPQW/wdDNWiWspDDUlvfU9wY/FZE1T+q3FHGig+Zst9s+eh9lNj7yOv7baL8Rbyq8oeg+UCfLpI
cCfNcl87Tlg3kswlC8B6liuwoeRcv+3ha9cII1411yCqDlBtgjsl9EUPMdsEK4ybkXo7PQAUsF5j
pfw+kahPQsz7Yuspdu8xUmbHPZjjB5DlBwyg+AI12VRQygtp8x3MblPDRV4Dd9Uf28wMf9wARLdU
yToUvyqUd0rOi2KWbXbk5XaTjFRndPytI5LvIaj/A/6xQxujXhK1w0rjh6S4nq+DtaxelY1I9pZQ
XcvXPIpycq2rJQf+tZSArOcy1d7mfFBbqZ1dB8xPmP4SfRjp5sTsdyvwcexXT7nuvmOLiAXmCQ32
YvuLQon4fka1BDG96zVKKc8c7cjQZG1RyiGElLk4E2gB3299bzmd0DtsfJPJPP83KbVwpW8Ujw8T
2Cfgx+K0t1y88s37gScTgwEr8NYLcDE7u8e7K/fy9OeNLI0yWYfCX9NukdJYtIcCsh9ioBxF8Bu+
PSkPvbcTTRaP3pIZwC/I64m3sFJ1O3B7luJZkFxm4HuX5yWz4E1bNyTnvgPtvDxfl68pb/hvBNji
FCM7E1uX71xd/4iJqYse1LlJRV7/IO+TWLDRQekho19KCNO6qhr2MkCyzFK8+APCByJv3RO7ILgc
cr8Efy7dWHjO+S3UknR6dVJ96vhV9/5p/LfwujcETAvzSIhKDcDNKDyphbtITG4cNReQFltS5lH1
FBxtx7e8FK6+nVygGhJxp1R2FUQUTA6gEsY8JcmHpw3ADFLdx6H4In96QGHCfRo8LiWIX5V2KdVq
hYwdbnVNnwTGpisNkY7Dd8585uD/IXnv5SWtcSmz5t7+Unz90rZZmCr22PIIvMwktLJ/fOzRMAZs
OHQANsNNQpWwexBYUybrlUBNRevPMdA2DA1HTNccDODRHAU4/y+gEMTNLAS6V5hnMFMsCfYHFVMh
eeoq1phdkWsYLKSExCy+xC/TVuSKbd7iAj5v6WeVDZCgsPyKOsWhkpDYFzPaSL2IOMqzZx55Z4SG
5fAPWP6uISt2M1k0du2aS6e16cfib5H91ZxMEw4yb7b6+LVfyC0eJsIfR8/9vkKcEjsiw1xMksD+
Fx0hNjIHfBab+3FltABs/vtxWBSlH0zJyr2ljEbU0Ob1TsDvm+ER18GFnbGPKpIci0yBh8g4R8Hh
dMm+eRF4aGMjJjEu/Yre/f5SVJNJN+rlM0KPAANgOWJxgvNrA2c9cl2OqShvWWaLfbNYuDsyCNUu
GBjzkSIUx8E4uzzToWABhVhXGDUGFWYEqIacFXdbchPS/TmKCm1C9uLLm1kjbKiMVwq2hcd5A5Bu
MBF265Yl1vRVT8eyXhvZHBMOWM/6Li3XPFGn0/vqCiH3ONlOWG2wG0sfqwxrrwEyYOXIKgbfP5BD
BG62dNyBhBbm9FFV/hNynCfkbrKi6Qh/rT4A77Y6fP5rvmQGaNDF51NMq/lWTFmUqgveHHELwnfb
7ojXMBF/npAVxse/uVmgct5RwTBULBvFcCmVtf5wfMdAkWim4RJnkUn+JLGkZf7G7HhnMWhz7r8a
XV3RsfIK/4veEQiQFF3Ms7asCDdhRarCJHWeMilcrt85CH669f7uk5v11vS9bGmQb7bxVI09TSs2
Sz/SIWSQK/KB2R7m5Vg2Ui92XV6GgnLue9uNX0PtiZKnn/Xx1dAtZkZAbhZo7qzrnfawnVissW8q
SG/8rbK6DM4wdKUMm8Ys3YfYKBGcLPBJnXVWxeXm9MBlE6Uh+Rp1fNPIeqBhJWra8ItiF5JVaLKU
tkwH7s8olzu5R+uCRlsFntnVueeN3eF3wt0ObI5ufaDkjrBwLQg30niwqgeQH/ORny9nDwlmfYfI
TE9kphyGRIoGs94ClJf9ENxWgrFSBl2Z/jizcR31OjtyFsvxs1TIJ4hA8ufiisYWmfR5wgbWJUwb
4git4jvqPa2rP9Nv84M6WbS/zv8lfn8HIYNO7g5KstOhvaddGnq/HWpS7w+iqO320hSy4LTwBBDd
gOMiebJvnHMtY37wPtSKSAvBD38s1LMqYxZI4NhK6DRWM6P4G6lJ+BPRNlR+9ZHebaYUYCaVFX5X
3ep2/ldesCLCPh91v19w7PomJ5eYDSl4wdIYtL9UkBAfmz8ulXhZQ8UVfe315VM6fEG2S00HdTLm
KdOXarnMyqBYwDd20+eF7LtHh+zS6lGTVcxqz5ww7ZR9u9EmHEuZemXisgvAYG5blVOc+MnlJa1h
k+7p4xV9JHl2Ym2CvxRbiUtaOLgb2bZtnAL2s9YiA2/ruK4LxKOGnRouP25RWWGmI3mgqXoMQY9Z
EImqdUmodJxjB+bAj+btSy+cmE5j5qaE/UycvtqVnmqlAUGl8ywMqudRyYiu9ZuF9JPG31WejiVj
nSuBizqga4tLgMb5kTUFrfbmCzafcvF4We5pnL91qc7oGfs30c/+mbN5/JyUL4l7o0Pxs7vGEX3s
Au5WpteHoxU1G5aYCs7QFXMT2nU7KiPhumP9us8QG0BwTYUPKO3aiQJDNtYtufuO+1m27nSBF+Mo
9U5nDW5Un04jtNGhynKYSUlAkumhkOp2C09AvgGAV2w+sNF99EyeaosBQONFMdPB8HIQHDw64EkX
2oLo3VuciXYXCPOT0DlruAaIYko1g2mOwoKcEnNplMLl9gS7YMyAXmqBKskRE7tBX3/VROd8pxcI
SRHXrKqmE1o1SElULThTrgnuY7uR/nQUxRcP1YS49SoHUWFL/8MYka2MMGHn00SUK6OVDaFK95J9
9syGLLCtD+R+35bfxXwTfd/eZWMjHMa4UlhwFIJ1NI++u1FcHQvc2FZE9oWeWvEsR7zgDj9KTXss
vxAhvgOrtgKXfHGE04YAiFuCK1C+gPngbg7u7nWIPuWYDlQh01VfkMF1zmw+bEQ6R9PWzwzNcqUt
TqxJ7UPFmH7yTIM7scTpBKO6mJkRcTRE/ujRmFyrjUneT7VGzn/lIXW9TUPIrntCEMIVtdgle3Vi
D5j5vxyDaetu/GC5ZBglMYF8UVnIIr8HdnGuayxR2kpeMEoJmsA9inmXFCPLdMheEL08/Xr1UwBr
FuBMXbJOTN5zfCtb+qQ05ll1lUH2W99u34Y2SILOnx5xdntjrNb1XE7ff63YIWVat/eW1L53sw3O
Ttfs2AsFqQvnAywshC75BT2RPA5N3W8PFvN+ImrTXYCGag7BI2xO+NBsU1hVFnvsZ455LHp6+9eK
C7J7XRGwOLqNT8t8eJJF+czRHZr+S3EiNHBsmNudvTVwbIBtcoVaDHjDbENGT9Ynd8gx2JjJ3VSF
W1pu0hLTA6kovQiHhjxLZb4/K0X4eSj5FcyuoheH6sYsF0yKim3Ed6DhlwAxOzozqom+xPJJhJ+y
suHMSKZt3nwOikK6yqC9ChdfKAe4c7m0cumeYXkChCxlKcQtV09un2b74km5VcdYKADySaS7eEHF
PlIoeozHhoRWFMnadXw8qXoZU/RBHEy7CbbV3G0Ltu4ZpHbdZBHghAQMFM9XqODFPyLMmaB5WAdu
M1iTWvXVbIKStWd/fe3pVYOvVf2lSSsvRSlDbAuTnPEL+7g2Y9a5kFFoMZOo80cpNOZ5CT0DFTCK
dMeHO7k9XFIw59LSHt+Lor/q+Kjyoyky2edjs9FLDvBlZ8G7WoXgTnb/AmlwshvsfnpXpF/D8kSv
cU29JMu6imWE6zJpaEHTqoU6+++8zFYuXEU5ymSHcf+cGGN0sGpnQptr2XZD9XsZhcElDbdDZ8UU
YGHDVSK/FF+/AGTWokzONHTTxE1qIkrlX+Q4CqEjcqhIEn33l7uOgUTBCkJfu/o7gHnJYiYq4+lI
djoRFT5gwJBgdS0xWM9n+NMY8yChIPD5fxDNB50s/HaZFfTWnvybw8UGmv/sVXHJKHAhTrwFKc8B
cRryq6SnXjXJn/2yN90G4htHG3xbtpwkIOwreoB+kQjjT6eUDUveqrPtpmazERlGI3Ug1U97wBIa
F9QRz6NEv26uIP9cpQJQ0KOqshWc9Ibz7cg6bCxa0Q970r/rG0RSRsLebfO87fcgQx8pGTw+JhgF
s9PLSpkxuOlzTYWQzZRXvAYp4axT6evgB3tSFClYp8cXyA8Aqsi7pwu83tuPs1UFIcYmJ99zTAAY
l3CMSyzNjFNxnfPQ5du4jtud1pbc7rXVMzoCwRW+ZuHrOdgpem9L07dJjl7UtYFHtreFrHKVdLqZ
YTyvN5gLabaX625RPU8maE7VjYtCwD60B0kGGgsA4bfNF/NQ6cEt5GqSiaBkVGuOCKVwG9/Fta5n
EL2k8NqFyyCVNf5LuHjMA4IsH0GQQeS0e5IIYejczAZYfhhX++aiSbiSyIqeMWxaBC1gXSeSv9WZ
FXD3sTbYVbBtql2sAhC5JqyT3MAGofmX/SpixePatUyv1qonF8sLM+8GUUU/iH81j5NsGQcIe4ne
R5K4lENhepgddP+xg9vhy2iw5vixLaSKUqAHyvgP+A83EzdianszdHRSch9mjMUNvDvWeSQ8Vs7U
XC+zqUrIibMDhg4KeGDVINgrJ+n+95kQc5Vb9I9nsAxMzLaia5sziakUNCPC04mX5eRBmV268zS7
DtIa62kaQ18QjTlmBb90TjAY6DpZsF1JE+x9rVNlk3maZV8Rx2aohFXGLdJ5WBck0kUSQyjW61ig
ijxOMbEyQR5JvSyTF0Z7SQxWx6jGV5hzN2Dwq9g0EnIndtSllCDjIFqL/qcOyU+jLEnGHj/E0PWY
wLFQg98zzfMcqrizIoQKGJy8+z7xhfiA725+cTP6yejHaH1sxIomzWDoT8vEdAV+l7/vB+7iJtmF
bDRJtM8yN9fsgFp3C4F2BWdVP0ewt4nBCp9rJM9e+4UHzzoAPz3yNnntTwKcrvAtcddsLRc7qQYH
jTHcLtDKGcC22TBciENdj307FsG3iMQwB9oPHzZisupxPP8k0s8jIQkXo9p5lLTjefoBS6a99JpM
uBpXlUTtt/FpISuj2dm0h47AuikKGEn5dgWKoN9AGkduxoHFYuO7G+4MErqwOhdquUt2DZyw7aNL
7chqsKhsIBv3FdByNWElb3/bYA4mgZWHO9C0njP/UpEnhR8BM3Wm7D4KbcxVoOeGK6HL5YUIqcWo
I0+QYEZjjcJVvuwTvE2oNg7Sz2hKa+1j/WvBeXsnBuymtwZpBjPUaXMkpqSE5vzIKQX6TXI9Qr0D
3sLo3qlUk9sshsUY+EdLzYJyiiZeJuMzfi0p44O7Q3pvGhMMkFfK4eIsSA8SwdH5CpzzX6vYxUjR
7Bk5uQsbD4L2TTuQk1y3ujexyTrrlHHyrqU31I5vxOu/K/C3Zgnzk484Pl6B97qIS2VyGfuhkURp
OU3BB+3T4IyKPuUTuNPDZkGHBjzGWyTrcaK2DGV2rn2f/kYvCbBwa2JH77m+ndIGyPZfGmkcn1Mg
QYtlxvvWjnb03sLVCswgjBuCpNZwkSJugBVnxjEgzPhhBaGAF/KQPi4gdEv5jf/szH9AOfNKAfdm
GFKQUs9qs/xvpK7zSTBiKI+yPrCx9OBEu9I4ns1Gn2pop+yn2a1xK6Lh3g6pfFoaZoNoVTGRm/sI
WprGCZHAkhVuQErQE0ZwilCP7bkIRMVutG22Rp1CliZWwbjJXT7LcxYB9vWrZcwFLY7Pf/XctwVA
13yNxb57n+a8ORMvHVjLS9Ho17EFp4XiYpr3IB8PwXCzTMf5XBsbx3U03yROm209BWSubNdstbka
6J37CYlKeB3xfqDLAd1DqDauLIW5AMUXM6Tzw1XTrY96vmhMJaKoBBnU4gGrpy4b9lnzjMjHLSm3
dA+4xbUKyFDQzSH/PDFdzZFfBodvqDHR7aiQVPZEFpK/ids2pfcNC2CHFoabzFzO72ChDkWzT1aU
HMvwkDaepMBIP/2w+0cY+lmqdh5wsElE/ReA1Ytg4f6m4xnWYRc4nmh+kh8qXubuZ5/vY/YdPlBj
Ff2CnDv11p/P0whEqIZ5r7Z7IGS0Tm1eTZNgLzZWrcXlOWsrPzdklpVqb22gylqmVdUBbRDBnfvp
XLZneZKTJkadpLikRtzJhQZ/EVHqSxnLwVkakuBxXDGhohsOcDYo71r0egOgPI5AaRZLIhkG0Y4X
ZOgm8p4KJRrpQeGipnw4Cji3PrzFck7SuQpCzuwrP8Vw3UKf141CbCT4q1TyAJ08MjDT1Q1mYB9l
OS1R1lmQxpdqDF2JpTHJDhPKQe0keMRJL9GJgLt+cgJ+/K4SZsY6EUtL2m8ZwN8upnlBm3E8KYYF
1J8kKa9zOe7u7Vu6FCRQYgmB205aNQ8k0vthV2JQSApshyJEJcjNoqYHACqoGr1ppoV2Sm0i+Qrw
6ohReZigzgE58Hbt82XSxNMlzLTS46aAoYHPvRlpDF0ZMLltdfGrMUgqpC7OHZXOlVSlKP6vYNOr
XUR3ThhbbUdDrPqSuGI1Pc3caRQEAnimfE0bzSESiBFuGKYESN6YI77OSxoWZlFj0PDkoiLvjtb2
9ESbMWhEjandoVSt6I7LHqUemHIu7I8p7kilwtrY53GUNnJlj9Wtet/Y6hnj9vpbxa+T7d1G1Mfu
V1VMW85dz6wea5u0ySyYDompqZY910m7iDUmE6u4spCCGiW2VqdE/3HqaK6pa0JaP9WLDm9aV1tc
gGBw5K/gfuuCuikLXiEvGPCstUIVk6iubBZNWrfI6luY2jISjBO9kxpf29YGcHH6KJqj69IQ0yU+
RHAwThnr3h8B9BL9eH1sdfAKYbJHcxIAN1glWwvsF+4sHsbJxPSI1RPVHXX8Z6/7z0CNvxVQ0mV8
/YxIMS79t9Z2mL5w/sV9rlcCYtA+jMBA08mt+X4BZu8ELNqjgpvNk1SkaIYFCArG83asz7Lebtxf
8S+h/29wJQfMM6SqpHGSAytA0/dtfKr0xz0NA+kPK66pvCO3CgkKgfuA8rgpA+2Xbh4d6KbmrVjH
fABskbo5XxF8cnrGK/tHPlR85Kd71HJafFNNKhyEtstmcRneCuU0TwDQv0OOFibybioL0eyO2CEn
/CEngcOOS5s0ZIl3oCKkkJHu0H2ajH9rILkDDFfm2+hnz5Bo47aTlRRUnpJnPrChcHBUSDp0cVgB
6FaFn8T0iQKSlYkYr2Y8y/SN0tMpNueLiFZdy5DZFaDak4yUT/wkJme7gsP8r5ma0LHwmd1Z6fu1
ZsnMxRq/gOrCwsOCPdXA0iOLqOmsYYoCJDEZMRq5jw6Oac0IroFA9SbQWGDyPTmTFqw6AmfpXAfz
hM2cTgHTCNepKQaUrz6VktO15ggoCAvgymt8R10cjsI5FpSQpDF4u4mDL9sLOOR7IlwhKzYXEVlT
u8myXcfvU2KsgcRzDY2DQLlG9nj1h54annmFvSGwGVXvsIGCN62qWtxWcrzZTXGtO4n85mUrJZNY
Biaz5nUuhpRD79YlwEy5EaV7Ubj5Wks1Qb2SQLsrD22NQjx/GZm8vgXdCZdWM5/zHdjX6Ih/lZGx
5tngyk1vP73Ujyj8cVuoBrMSjntusWrhoEzddztHAtzi+Z7vGWQppIoEl0v2mq4NcAbPw6VEEzIn
pqQD+4qeoex1CQdFf/I38iv28fVMTd8B0ojqFWQdNWginV3jVMQPLeTvl/jhFuTKOxYGFIrGGJXx
i+oaVlyPSE5tUOuUUKZfkACTFiKrqdCgLNgjmEaqQwfhNLY66fCWFqAgFtyCI3/RERT6jRT5totz
a0FEOYkK7pu2xyDalUYJdzS2fjRUhfugH0I/4Y5MgP+kOkTShPbcFlyCetORqs3tOx4jHr/pVEwk
SybweRYLJ+7S8FAWPDPuSo1s/IYj3aGaBeVh6PPqouAeV6OGQvthh1kpefuR/wPCaNtl95GreAhO
p68JrzT55K5gow4HvwpqHFwwKu/6toAFPUWdOikJE/cBjDeXu/xM06lemfJ08yoPEptqs7o2VzPz
FBK7A/xv5DBx7fN2unT02IM5HFCBTgKmd64xbKhz/oPqP01zCqlg2C6kLoBKNRUX/MzqgnpbZdR0
wuINjIIxGYdluJOUuL+/acUWOp+UOBhJR7QTh/DX9lEU+5l3GYHrzbZ1sKp9glOB5r6Gdwk6q9+t
ahlUFMRYwlKMmO6wRM1VAtmecQKQknHECeIAE35uSpwVukuWK/zjwNDN+3NFFFs9zlm36982VYC0
knf1mtbWPRI+P9G/08psaNJVJ1frPwDHg5n38YzCly30yXW9qiQ0He7aF7NEPEQA9gbeHaVLShZu
eEz4pTBp2c8HLZ/Zxr6t5Cg3ZPyMrliem5k26hAvUosprLBH0WNCmCmFUgvbemi9Yt3LPfUl6dGs
Hs6xSgxHlRdCRDdmhHRF3jHLZoaq9al7GCZqtyQBPutW7vbNTLTUwbzrFKJhTl0vTsXssLH5FbQB
rotxrrZ++Dmxv4oqP1G2htgBDv7+xPU2F+XKwcYrFrIa+qAwO8BTgjX4z84Y22x624OHu6HylA9m
BE33buCBOlwgA4gaOV3BbkFi+PzBLy9TCTRV/UGNYJltBNqY/qyFxWFPeBBFjBc+5FVjs/uYwprT
r3qIjnkUx/GE1YyHXZ4Fw5lVZe5qoyohDfwKUeIIlriL2ZUWKY6vbI/kgEeGikzwHj1oHTj/mpJ0
ANUGiw1lxcf2Z53Pm+nbnyeaBm9AaYDXDZwNO7s7UbmwXRNEb+ktybBnBsHzsvbKtMKNzS/tUSP/
xP4CQfraHFPaZ7vC0l1TfC2zNIba/VoxZdf90b+tzApJwJ3JvrNh6FgYlTsBHwS7LxCI4jEBAlxg
0iB8OUsE8u0flQbASLIT/f5IQ2pxDDoUFS4E2FBmO+8IryV4wDJzK3jn1JpDxEn0H+9Y2iB21pBb
HyFT1jVxWsCZvrr0XXw/8tQLhYfRag9MC+fY4XOaFJT+Zm2/oA6jtoI+oLbGvsmbUp+UEMR0Og1n
pVaz6+TqAwarQti4IEUD+9dImqdGeEZz+vcfDtQS6LkSTRwgNBmNeoHIDuNvJNKH6Dsgalwm8pUv
nrNXBsxq9txnHtjHuhAA+gqRphFGpQLVMCUxKvE9OGyAZ2YsvGxe2VWN6v1V6CnfKQXSgNjoHFJL
XZGnb3bWrrNk+XTSaGn4QF6GSmBB9BRzkwtdtwlxC5M7wIEn7LNCV6aytgEIEhcaNtevZ2PpBrEB
jVQtmr3Doznr4jDRIxL6I3ExSBKYDuhCEWttL25+jIioyms3Yp1Yr8k5uNqKcK3kyTnBgaprIlXV
qulltvcFSyOGluYKd8UaF1iHZ6v4q71SM4o3pkNN28V3Qt1GaM/uBtmkaDvcoEKyu3UBYt4oJx5I
uYPmm3YhB8HpPQgQuzA394wrSGv8nvZM3J31ofByCAn2qbVQ2Y1SAsY1WPqQ6yxBtXlGzNuXtV+a
mpldSJnKku1xujLPFEEJiOQ7atGY9MoMtiZZyQVQhj1O8kTfZBvCUyVU4RzyPs+kRiU3kUzh5Vfq
pC+xokbaDGwK3KrEsitTWisc4B6YWCEJ4zNBaTrBoLNT9G2Tvn2r4v0hLU5QZResYhR4S7ss8WdP
o7+Q65XHAXK9ZdI4HFUQzS2WcFoBIqrr6LgzXTQaEvasurn3291cCWKq6+pAZpbgiGaqK1xjV8VW
VIwWr8nGh4PUGUJRA32gQ/wqLjw/oYW4dNlsyaPFHaFv8Er3huEcJe609y7R2v45fuK73Vjv6Vn9
5Ukh/J3+bxq/BsqBfSbYbXAPnJQ/jUrpwoDgFsdziOmMrIBj47lGW+Y2sfNlbhlWmSYD/QhWRe+Q
1qeGWNgeNNPmv6WzamKam2IblASm4wihSCLHMCAzNAKcOjgbhstCPuKhBoB8pXCS0w9mzpkV3tJi
xkXDIbVPqu5MK2yzXeE1wXKdP1p6ycGxL+7CE63mPwaibjQUIUprcHQxGbBl69TO/S4+lqpSYEAE
jQrhOUpfao5QHV4zWIeAHpmO3bVeX+XTqdOYZnx9kv2NRnfhqeyCV5alvZ5PeF4aviqc8Q+0rzfi
fmDYr6HQhW9h3fE+9MLuOvYPIRMOWFdh3cKJKELTFxuDhuT85zer3QP9LappcgLpcpyYcy17fn/Y
97ibLt0uVwFtP88ERpu4xFpdnNCZ0ntzFZQJI+EVjtCGbuTCcgGH8sGYz12LvlCZE+FaxEzVgUnX
c8h9xVARCt22UnEq4YfSOabauJWJ1mN2+q8l0bMA1E0iE6SuvX/6mcUD4jxp1uSFWayaEcxOFXDv
OqroXf+cvnx1D4ZOfNVPAj+GsMY4iroW5HZaj/C+jSEjzwVUJoFmUaOJnp9DgRItWfh09COHnWpQ
8RHdsEi2pvFfOcEMvliTibTDZwUWKuO6WuANA5nwV0Orem6+w34YiJokIsg0Wjo3zeHmc5ng4yZ1
NtvTYecU3Um/Budm77kfZUJ+jk8+kw7/9R3WfEetM+7klnMqTBVVdc5iyzz7TmE7UOhN5XqpXfMr
6zDKUuVMMbb1+BEsQx8Uzi+iqrqKe2VZ7mflHYLKbpffzzSPhyd+Y8hprTZyn2UzgwSWpIBWJL7X
9alTcdRFR4OxDuvBu8AOs6cFnS5YygqCT5JFa2bYGM7J/I29ZRXTkcmU2NmQTPwAIp1hJ86KReyi
+traGAosbIQ5JGvPVMfk1IZO6rZUgwE/MSiiSYsbCLIAWeMk+eLJDR1+KTijzGfM6YwvWzzUERkj
3crQWkA0JPabUtYfwEVbhIz7TEMvEkKeXSL5we9cHb4RpkT4diIZlbzHWPz5UhL42Sv+SfXvFv0d
Y47+GdzxH87LqaRF4zWwK6CVxaEI+4m49L2kCKzX582ZTKS6rheNZsdxQQR+2lhlbykksKeHqkIh
Q1aai5KsqSMAYjHp/Rkvk8l6vvC+5TyeLuwabQ6OXQhweZngXo96TAixbfz6DAd/XeyGFItYKoXy
AiWwQ3xTvYP5NqZI1/ntiO1ebcL60OOA2co/79ALGVa0pjB0hbYkHF/8mcXSD1DSyHGDAwxKnFYF
evJgR7jn+swfN1j1oa1nlSK0GH2QPyTrjd+Ku0ySB342WpQNWQrhjn9U4mWF05sr04xgzA2agY+S
u0fGHlTGYeqvFW/cWeqnfXzVJ6Afh1xUy2QqqrJCJtWPXIhEoYm0dkbZjFWIcW+2rmPLDO6TN8WU
5EXlLrjUEM6wWvtG+nYM+YyrSIa1/iDrvWpBCF+ouZsn3hXV7HOu+BH0+dgvh3hwHSemyQ0O3eoE
GRChIXW7Zo9+7RCNFQyZDRkMtHz+f2xU/ypLOZiDrp61Qbl2XFvUBZlvjDt6QiNc+hZIMjt/e1Ak
9ZNioMaBZgIXcRiEm5UPVqGS2xW0cY2a1yKjPbzwsUMqB0Tm26y1U5Us9HNmGLnAZFvRxUz+HuqC
lFpiPriekB6uVEgj2AbNu5bZgZdZ+rTc4JneKOGN1YsqaBscAYYXprInT4pUuKZRzDdG2RgPeJbT
kcTNehG5IxgYr7lIqIBqGXLpgWG2FWFtViyF9BIwIJnZCMUAywqBj6fNcqKur1AASzkeevj9MJ+Y
DwNRq/GUQ9655To2B0MB2H8YW/hxqHcpThqkVg8PxA+kb2EaLUpAJdZSsqEIexkgbda8gbW+C8I7
vil3269M/zFDgcHclOy3Ma7dcGdRdm40oJvDjn8t6Y+rEGHCLup751ysOmx61O+rC2a9iSfEqiMN
uxtqqoAuRk0B7ieWYUcAFtnc2yY+zIHq60vTfUaqgbEplnnVE/2Zi996TyG0lF4IuLLZNRU0jsCo
/4HnNGbvgxrHJd7ftwT68vnL1HwaGii308YYSLdLm/WhPQwyyUUa+Yjjy5gJHfPLVSgYdi4QhxbP
1bDJJcCD9Ut3hDMVJbMjKtom4bN4Xfd789jPi+EMjxq/UjiYoo7Cu32NhrjxHrLGF45A3nXGoSd8
Mx9NVFSfY9rxPxCgZZd+w/vp+gt2Z135Vhs6S8kTj6vXLDFH1e36Lgb3ghdVpCd0IXjhgP2S82Mx
JRM0WP+q9aBVz2qnPSL1vtSq9pbGuD2+liedCzOtyl1pGjARFcuHNhvSleuYUhDap5pS9PNzgxyX
C1HOH5O2koXMMe1LBk0kzTbjr1R1iSxvgcJj3xBQLQamVkazULSw0wEO2o3dMYbxOvKlmaKMX64m
fYvTrnOIGJEsFLye8P9+t+bTgxSdV0hFXGAtluYSsz3XlKKFX9eA39M3V3OKPvOZSJL/RkIguCL7
//MBbfTwPeLzsgZCBj68JrcFU9V3gk7nMRPKiIPryJxcGeKvy33Bi+62xzsBewqvTLR2CE/yv8q9
hFhOSvcdwhDmld/kA9dTaAE5b5p6go0NEBusnT//2nGCYgY+Kmt+75chwKxi4VZ4s6sqVPS3ri23
sP3k2JV+YrplOLLZ9Ou28V4b77wApWRKjGcLgQQ46XzvtpsJHC7TOGcYj3IF4tYPU645jL15Is3O
4QtX39bFVv1YZky1RsBNvV4JP53DgtQsfwA+6LG/aQPjesyrOjlff+Vq/r/f7+34kK6lX1d8QINK
RjCI4YJD4SDU9yFGN2bI0b4pKNSSBxvsdF6uQ9TYdyqs3X+bCtC1sCtw731FZFpqxygU0SXQ/T2i
93NFL7PVQJtgHBid/IsTIyApWKfGCUvekm+w1EJO+ueNc+nUAbF6k3wtxZtuWZW6HFiTsOTiellU
2Zp6ZRkdC9qJvH0pj3qp7gYUB/9RKI5SwfOT4mWQ7q+sxpAitYxlcH1u5YIoxAyUjp0LsYchg0N5
DCdnEKIW7J1Oxx2t/8VUHKHRcOrXGKCGz9No25Edglqat6ZYIyvxqT/Ig+PSuUXYrQXcHXCOTg7L
4+005OkDuwAzEEQeAKdVF+VIdB6i5uNXpgd72fP7NNn4iIV11MvimLAVh8k4bimqNUmbggwGNowH
m+vz1bBH4j9Zh5R4E/bkV/chKl157KTd/146dqVzl9auaz0QlfRB6WZMDVxJGwhOGmNV49ee5579
DgGoWiyenTcmIpAvSsXvz9JnuhU5UNJzXG3jYN9DzTLcvlTMCMyvzY+mClNO7CDOmBX9P8hICXGv
MvTeGm+KSNOieIvR5aBGtxYJ5n9Nc6kLRYHBM4bMXwbGTK1MPWsl3L0l3Yb/1SwlG13VUnGefHgf
FClR0s8qjPvfsb5AWFQQKWqZ0QGuHrgb0W8smrrhA43RIrvk+dZOjqxcRs/lxLH6rNd/O5yGlCa1
1sQIkMMNHVQzutON2dpjfBDlhmktGqizuZ/O2eJLL/xh6vYHDfDsK+JV0EYNp57nzCzJHKyIfFAf
VCNsOeixX1dVl65P6r2PxPFTSjvO0JojUmB8lP4S4oRp0ExLAveVQMpPv4cY1FffEgXUdtlDNNWH
jjEGDdD+KpImP12MeIg9CgB0SSJGrYc/NWXUjtAf9UJqCDNcZzUg4V0wAFuWU8U7D7q/nZ9K4clO
rEt1JV/v7jb/vRxkJbbOB5K7qMorB0gr9Nd8EZg5zpNNhaeiZpI8QdDx875jwFUeSx+AyerTdMTk
cKefpPiyijziuh/8jzOw1YJSU1o989Kp97EXRh9uykN83ANmJHcmAoNqIAjq1Blp4skojSgQrCWE
Vdv9EIbG1g9zxhSNf8hRWzSWJVOQa1C4yXCkTE2UbJ3St3Y6fqeKN6iaRISTqFhxJ34a3pV1U2I2
oQvSWKQwhN88KhvLMUbT7Tbj91gCphQtlce47KvmSEE0J5WMSqmMlE/+G0TVqclr1zmf9f9003xU
yjkFs8skrkaRAPfVfzLSEbRv2FktMfIVnkeTYh5qBTkk1+T6THMNdIXyDHyl2uIrLLx2eQ+b8QSM
W03jXwpoUYHhU7yDlqhE5kv2sTXCWwYfD2tNzvyL+jg5aipLhHFcq8YE4inKTgCdy8EeO9/YXL4/
jlURGGb5Lj+P7g8Bh9do4NUucGjrZx7gD+AREWU0HaijgW7t8hM2N84Ob9GCFcWkJTf6G9++Emtt
SrPHLbsl2Tf6aTm4qRqVsfuZi+x4txYFHyvWG6N5oBu/j6rtGR5R8d6ISt8CrEckrOeWKY9uBsDS
AwwktWgPxtXK3bbYZ4BI8t+Ug9Gq9+6gXem98ytbdPfDqaczgeuJhRB4jm7G5Jf5hrmSQaznM7OG
bJDGwWPTG9N5mCMqYwEXO+KdDQAv1F+b6l+7+4GZCSUeYDRb4M+YygNM2RAS2GncCnclH9fbLLAg
1eNL4a0bdueKkQjSR9BjZO6IiIoKM5BJ/YUNu9R3cp3BYp7cqJ+qiDpvNnHnchuv4pkxALizscgG
MuhlH0bSwzew+pmmxkrgYtQvv/Cn+u6hqLv9Kc8C/F2ohci5pI8DysTLgGt1v2tyRr9hjIAeNxzN
rCtDrw4GYKaEqgM5nLJs7jDoOYSfWcm2xI9Qyn2uM5x013/3XzlU+5++oBSI8YcjmSZNqxxoYlL/
2AhKhDLNITup61TKRdkXVwZMeEbie7nawSscQJU33yh8uCOsxxGpyE+l52/ynbEPJ6n12CNh73LN
/DzIbVwkA6a+7YE0JtSxdIItTK4SmYlympqF8vBgxDoJWAlPDFRY8XF13jPpo9E5PSdc2fAixiyx
j5E9b8bpH7vd4R5Sb+gBhbvUACg3a3LbHsupWCj9KhsJuyRbUGjHtvRhKL1vAWQWHao5Ul7mhiPO
I6vS41CBw8NW0d/zp14MWYo2udUIXajYRvZpWVRJHXujqu68NiTBl49iN1v2rINzoqvq2JeDfLfO
u89QZD7jcEvXP8iZiWaO3/q3q9j7zYYzdj4nryFX99eeZJRuXThxI2eXkQXYPNleBQncxbyBtWgR
3f/JJmr1h4ArfUHDrw9mDJkyojbYR1KyR5CW/lVTtZnbvWwlq6mxjsgQUMBqVHFAlOpHee2kVVBE
QQMt54PJnEvqIvuR1XglHJHcn7lJhLjtkJPSWc2k16dsyaIaDPlE+PQvs33jwAKJZvzLZZSYt0o1
lS74DC19/+UDwXxCMvOaTLUNxxK6o3ZCW/6HYO+PTeuqj3Z0SJNaHecQ2EDoQzuqUpN0dsZ5xjM8
NdCqMBH4veG9UzZhm2jgTY2reGs0j8p1HJLDAmRCaC8gZ2q2SEN6uGMx/AElotoXsX7CuWz5BUO7
Vn+c18f/E3HesHqOByXEockKJFI0+LpegA/iIsIwFmOxoWx54QKvBE1E9aPg+AFR6eEnOAC4GfL9
Rxr+0lB/KIousHvMd6CsF71eKkOdYJyDhtYx2cEAOYnX9M6Uu+vWQRaswSIdkhpheecrIOwMqXNf
Svj7u+xlneZSQNs5H3g1YXHjZzLK/4EoQtgokrovTaDvLeKSEa85g60uOLJ7tsWIqpYixJQx43rb
IHJBu33WJM61OXcqgtx2kdAsXsVb6NmgX3olx7CNJZLasPLSVB/nbsRomY9gVpQYUfDTnBMyoJ6b
g6Y/ALyevIZTsSUnKWDytxQyuKTV15BydgTHaj5E9nez3F6UudE7T6OsQDX4/FzIBkwbUkamOi/W
x0GjMErFV5VQgXuGwtCs6QQ4+6aKRYzB9wfWEDp+E+cHTomGSeHXjrP2oa8FeGz3sypMhikLZp7x
gHAkUyTvScjd/7L5TH9wOV6hwaTfpgBiGdR5SeOaIET2JWjetap6v+g+NNZBR7CgJSb0O2Ji1Eml
31Bfe7hqwZ/SXai3Gr+WYFkD9puZi/iqK0DqB1H6bMCnB8KhjEgzw++eKk63QbiKYNhULgd9rJ0J
is7a3N2LpfJerdVZsGDZ2puP4ZqWQayzXbz0S6XFTqbL6JVzgd8HJ+0wRvLXD0N53crbzPr51y0K
kRFReoKQcya+x0+ntULxYKQVVuyoinxEbeYZR9s2qZkgO3VlX0yw4oXR2EJKVci705+oxkd2TUlO
wXYLC2AQrkAWWBKdGdCAGgPQeEYNPp2+KvjVAyIFKPYsc0r2KhiCjOMF+YPhKvtkQQjzbewZtj9n
E8ElIIlI+p1f243JiU9h490c4pgP7DdyILd9W1BfVjYdM0sYYH+FGhca9OPkPFRVgPg/hP2fGAXy
QQW7Vh2rELYPVwEm9y/mJ8lIEWmexCcsCklWZMAjRDKKDbQCqs1iuG1nPtlO6NHWQnd9i5By37vv
Y/HXxwCWAUxduvQVIXiMiRu1ZidFG9TeGbejWpFn6MRD7NLbcbxBHlSPIVxu22QvPRVnOjAz0ZIz
FtWCD6S2mg9Mf3KFOLbSKucn7AicT7MiEhDt5uKs3gpmmBSo4DNhQ04L0SwfWQZsodIqfiB4PLQO
K6yYxrpfr3bxnGuAjc4pCwsDBYlzOi2O9V5MWl8o4A70h1Eon2QNDPiFk13xHuTO8sxm2LI+JLNy
keopaJE+qd37yeL4FvYvLE9SrF/+Aq012PIRfodSJYnPxiIU5wDEpfwvXHSlmvKfRA0Kb57P6Whl
fi4YSJ8IXTapqU6Jm9pQV5RH4MdjL06O8IW7Ll57fauFt8vSLpXsBKDUme+Eip7a6cta29BPUNv9
YtWti0mbPN3TlZ7ECdLl7CmHEjMY18tT1xixP2jrBY4DNo8nY6B5RyKrWXSeHPkDpwqqgk5pHGTr
46Xi9mwEC0CY4I6cBlEjNLc2BquPgvPAJ203yatJXnip7W6WZSuQD7E9X0pUHvwgVqojBF+arKbY
AxoqWrhokXjoNPJr0JdD8aGIp1bAjefMUhg94mPK/WElOMAf/vxMM0CGtaqv+dP0FlXSEurXJvGS
FYsjNT9wl4l6AE7wnpBvvsFcjkIQte5hM89ErpVCtDRYEeKZ3IOtK7aucaQDjyrPttX04GR9F0J+
fNu2kxelQAsL0bGAs/PnM27tlexUOAs+7HrwYJRWlEjU4oxp7FBzgDdSn7N6zwHjWq88SBY/elug
3TfmWHMce3nUt73bXj8uV+VVb25+ib9Cmz3IN0HyZrR1s13wYPCk5Sg7dlyGzVOuY6xaiFR+RBJc
STB0CXF/antFB1/OcRJk+ivK4pVhcyz3VwbqjebviQIpUbG6Pu/l9ueYXl3Rsaet0i7rH+zGvSFY
yNQozzTLHqnFFJVhRgcwP8DGURn/tM90uGvGeGUSZ2UjN0cKJ0tN0ebyXNeEY82oNAjnQVVfkQN3
hFl6CbU4saZdiyMr6C6MKI/0MDil6od2H4Wag9tnIMghZ1zEaTeYjxtvvpbckghr4hjujl1+pM+k
kY+g0f1LB13t2lRYJHj+rqGOGyaouGl3qpdJJj27YWTvsw6IeaNdJawUNtkPcaQ09kySle3UaiiE
CTgrXUY5oyw+XhAyOOmy5K60HbchexKDAszDFxnw35LnU6w8fNg8PstQPrKAY2SxL2mWQ/gMhHVh
vV2A7gRmD6ejh05vAHtPjmJWY+uyBJUGEkL7b+niPJsOPqCwmpCxrPvMgFe22SdJ3mDHm3g8hiuk
P8wk8tksX2p9EjAKZUManOIwHLwZobx19b5/iyMK+jXAhbsGme4A0K2NNoBhIcmP5K9dgMftUZnu
/E6gRVh8AgAVI32idb25kM2xponATf6WUUIQ1FHTAwzZTtOnX+zUblUcnoG2//0ft0h3Twv9t1Dd
sHGyb+63ZEUj/ptz2O9f7KIAUkFkAOdBdhLDQsvHV33mu8UEDosbk/af92O8QlhKVjFLd404z710
3jkKhW9SwgZwEUuBumA3h2RWqLZoZvxlgaslMI/PpgWpmtTuteDt3TuwQDSyqT1SXtEUs3b6WLI/
uXCUEfeIcanql2EqOmYUXdi1tyNvqVvTP2vVnSLvpcpW0bX4h7KblGm348V+EsG3H/UZDKhvBnBD
FvuMjNwj/DIeH45A1X/YMUk1VE4ui8DltzlgwEQRigtRU1ISzaW0YUaMWkaVEEcZhS7xNPvmjkVO
WPKn0YhWxXOtpq5VO4JMiNelwiD9FXJfz7RRcOvnBYZnebtpO7B5xC6hNAHFT0N0NH+q1y1KRkOv
3YOlnYtdpN7Gh5vq1Bt6Lz851bNhUHl3pE8bvrXPc7Tw57ip5GAeLYzWhAu6ARdesAEVWfRG9sXS
zWY+epWg2wS9sXm/qkK3ymWCdaBUt0crqdai3TWdPbevN2XSiU73njAcAhSSE4HdXWOlChyNbu3k
2ZNWRIPRbB3uCF5W/6exP72ZQorR+0ukNUGOml6cFQwwMdYA1xvj19DmkynOQ1DFObuwSpezi6qt
HQWZbQl1UbFWKJWB1XcG9lm1uRBPFYxIOLbjmMHC3d6a4CwEIQxBiM3PeB6LVT64fYEwugfcZgwS
gXUnu05fV6bW7RIsnBWEsgLQOa6F1I6ojlo/43c3IraVesfInsjcg6NSKUcl+2pJE0x9ghM8opE3
skJXCnqnDzDuFHIqS3bd52VHkURY8gAPkL7hZB1AJ7KsNTKlDWc1Q+JzY4LetytnPboT8GJyD+ev
rFjJa51ICnbtDQ+03cJS6RRhruNA+SwfePwEQsaKj3hkwNUcGhU4KVKTwt7gz2/5GgvJc9vlb9Dj
pKMqMr1bI/LjuTI6LPKcwLVtjLAOQZ3F9VQ//k04xl5uTjhFvIDQ98NxgInJhEeL7dxyi+Fzf/xx
B+8N8WbsFks8k/iEtRy/8gG6YvSTjxunhTsxvPVPbP6gLw9CmpagTSVwaL8ZCYBu9IojzFApi7MA
/sqC1TLiN8qSzDPmei7+5YBXSm4kTxGXeNbuOrJjjJgzhJYr52ekyJ4jAD3hayd7YQ1eWmr9fmHt
z+DY7HWRu0uoEun6WQE/vcCNKlkTW1S7NVElJPlbWbmUcWHVDjMUcxjc88bN5eyTRfoL16mcIP/M
9qnFo5PGq4rzNnydJJMWPV9IP0j+2190dRpRGpvuEzZ9PqEmKl1jFfEP2OyiAXpdiD66zEBmPu3O
p1ydJMv7EKxBEDTx0auXDroWhbsDIESpaaVXjRNEblzoVHiwLEIkVSFZv5FkevvgvieVgadPKJSK
pKFP5wM4DBSkSysyiV3I60hBdDNx4qdQM3a48xTZDLWEdX+aufDGSF4vLf5Yzpx1LsC4OsUXYaxQ
xal4I+IN3phgzGtk1oW2e060eHpNmM2LB1G24R1ZWGozdG4zZVicnxFFOXRNxlgQDrTrSv1K4L0Q
2Q2eqrDF9CkwY0cXodD6GwnEGOXSjDVkCcjVSc4d1VYd28ywV0rvJS5PLvULCuEjDCvUAoui01G3
MlIQhF79uAulyXBVseMQLc6N4L0WeRkLXaxZsU/XYbKcnKsaO7wtjc/Vx7xEaXK6uM7NAcNOXU1h
49PUMfI9jETmK6JKvBBs4kvOCd3yXz7TSwiPxDFw5x5gfJWpN1IuZiFOJq8ZSv6uAFkLSWIcNkMk
ZZ1BfomK7qnmNEvGyKxEGhwM+U7hX5YRfRbctZaEWwZu+uoxkWZsnGKz5IX4B8jgDiVQYTgAHOnN
DOwjuy1rIF6SxqWws/66zcig8A1hPaovegm2SQiQ4dsTtYzxCYkEZzpsLOV4MryZndDtrrsrEz3I
pFdalIZj5+iGAz6tLqpOtnzURoGtr5dMlF5qpF0SWUCrBfkagwdmGNaUMFwkmxICSoMaCFzvCwFC
to8dcnaqh6ijk+VhfByJiDF2nBMmhgKT18Q4YcJW9hWuXOymyO2AmRsWQfOxjKpfNerXhGF+kQ8E
xC9mxseswlFrua1QGFg5YIaTHPBeOpqjmsp+W8kS+2ea3J8hmA4qehOBH3nQB0ASc/BWZhlUnVaa
CJ5dpZoB2jTm6kkQPsPvrRTSNvUvv56urz76sNbauqj5QnQBUbTZAyp3/UbCywWGoPd8CHO39yrQ
WRhvCYDO92RMz49h66ntZ+iNdoqw23U0HY1h67ksJY8UPjj8vGKs+6/XNG4255YHp6UpZAjknih9
uom0bIjQpz79pTlYAXjTWH6TAdWm4qtZJzVLhllWdRO96vB1+CzWTBtb9x2lEyqmaQr6V44C/PSl
oEjy58gdlLBYitYAZlR4x33d7zzKYw4dLomMVQGStBdlV6/O0lPwNbC5n54pwGlSBaoxpVviYAuK
HHqX0/Ntwnk2a6h3RwaZ6ia8J1zJW4ojfXNrLrdDY2vsUvwvIew34LExqB9mpOMh8wYlIkT+uTYE
IzD4eGJcnnXGaDLT2q2/opEryjoiKn73WkPwDGHHTDt2nJQfoPnFVenwGh3Ab3myG+onam002rEH
6CU2Wni+uyplFr4GDfmg1Y55yUU1wCzP6XKcqjInuIjTN6Wjf9V4jbpUL+6itnv34eYtHZRPbmHX
QiDuazBblkDKEaUuLaif490SilJah9HTUHD4IfVPCDTHyDRKiBXAh/uOVPmgpUNNtumuYbew4a1L
boouDd729BiGAnfncidZ4G8pKa+Yl2Gz72xC+dQTPPlMY9l6UILTtAG1R3ESZ1FCC4xv6s6kftbU
G+6eLlzc3ysrwuzOUnOZxU3yMQx7l8TGUQx3MslNFDnQGrmDT0w4/iN8/6i8MJnIi4pnmN4bOkMd
iIWKuWEHUAFFozOqbmf2c4ulw3tiHdhaQS4N//VPCV31oO4XyTezpD7V6ClyFULf9+XshUwDhHo4
YQ7vxb43OQ9QGA6mCNumIvCM7uHq3EHpO+F3TdXBKMX9yGqasGlKYi7shBVfYjYLGImel8jvtQyH
wCNl94x3fS/GqDjV8KPkN5oMGu1w3Vbvd6C4j7gAgTYGgkMEbdeijDhukvImpFFtqaaAmT/otjYw
KHPB6kC3tuqAUr9psCb+vm/MDQBV9W2Kwd/2DBTIN73JYS2wajHBw5NEd45QTOazrHxXC7c6glWp
+2oQyqvdyeMjoqTa9bS+kKU0lxEHi/fKui1jCEHAN/8RrVyidha8XbQLLPyW9Oi5V5G9/i7KFbIp
2Efjkf8SAwxrnEh4crhar/E5Ls1TIXC3paAuLdwfCIeAky/Fvnvkk+NrW6O+30H1UVn90eCocpNa
isSNMpKoVuYX/nME9bzHjzpcRx0u3C2jC38gB5MgDCFCH+rVtg54xBU0/m/lIqEuKQHhHhGsV+kM
KS+us2t3fAfj7WESiqY/eI0eR4tW7trY9E2dmfsAtKtfflROQuIeEWEdn19x32fhdBLYaEZPDNe1
V0YJRWW62i4yw1DwcIN6Wjlu+djzlDMMxLPyx3ryNPfh0KKGLoGpnuWPuMY3kVZFOvx8bk2dHvUC
npvcZ9db/3nH+iSetVJzt1f90cH9/TuqSDKIU+fH7AbAl7Ym37JQqK5rVns5KUT4uGxazmcIag6W
gsk6eVT5ByaZkx8hdO24+R69JVCH0islm7xQbwkeEbEfy6UMCor8UBx4io4K/BzsexxP4exKiz45
Rkr1Hj7257/v4spwQTagtmnIJELkttPj3qytu5gtyAsiAyUdSIoObFFoueZMnMNmSTlFCVBSqATb
pZFADNWgdBAtrpdS9U2NxN0W63C/NmiyPclRUMTsjP20eCoXHlig/FnoTXiZM1azbKk8XnWmW0A/
aUEwQ6oZ4vKnp3tjuQJ1EWjVKImA/Mmx3pn1DswiiJxXDSaZsOJ7BnHOWXnIUoxWORfmPWP5vmD/
Mwx6oHAAXIZ1HZRG0vh5ylCz3JkS7IFXC7XkjVjR2f+bp//Bu48Vn4x6GcwBqb91krkmsp4IxcpI
DcVJf5Sb4dTSUXuz51+o4Uxtfh4lVFcpwoFS+l48uUQzTE7fDs/w3fDklazszZvI4XogW5/7qDk0
h5qrGdPll07FyWa1qaBiwXVks7B7u4HxfIpIYsF0tSpgzM/2g21Fk5VckFUl6r4FCzZgRuHBfr72
Fk8bkJ48ymOIA7sQHhozDxApjCec+VUxCIQ7vEZmG8nEE7U3J8WkaQT5nJ1upuFdqV+zKJdGY1gU
3Mw7HYMXTsbNJ+HDCVKjBkIHLYvIrBG4zZ/8VgOcrFh8cBMfqZzuljFE+yVoqHtXMKRZfRkEJGXR
8eD6XQjkb3CcHZ4eWLH4BLp9VpA/6ZxtCgIE3BrpWU9l72GKmRaI91TANMQoBVOufk72w+ZV8DHj
COtjz1UBvkZmhQDaHO0T9BRWIGJE00IEy/Avsc0G3OASjV0lF8f4bxmeA4a2lX1yBIVTOW2dwm/2
3Hkq5L5bY1E1tL+2g61371qT7yukFrpV8/GNVRmEqc2TxZNEjZd42S0WsFFN7+rW1DIEDO/p7gZX
aCJ8JQ8lTzSzfBp+PjeH/Mp0KTxnqiC6ywaRew13sTb7WKovwYFwNQ5JBcDTS8M82C/uNnrdJEx1
IVhVP+V3Qf/jGgjQ654HREAg+b4fAC0zzVrpKz0sUNapvexA3eusziOnGhlJ64dLhqYVhvTfV6vZ
bcr4jvCq+eCMTlrd+N8Gt5/+iNEuAN66HLN+PpBsAai4sjg8vdgCdf6hkZNxdVrfGjRs+l0CPucr
UubFlcULowFcH1lPA2OXpn+GGcLyiN/SGpF0ayVLTZxaBskscKL7KkuJh+Q5ZCW1+y0UuyLdT7SE
9loafL8y7eB+V4QT3GXZNhN+8y7fELB1FESu3TCl5F6is2arZv4gRO0WAegXlMidXHda0Sy9b/nw
pFjOKDxi1HEBmMtovnY07qZtqPjkut56tDR9jW7eRNMOu5IAD3ue8YB3VQC0RLPKS7lQQcZC5crM
OZI1gt8cUz+B5CVC2k5OKqJnevk6gmOkCI8n9+Xkpv/TgcRk281M+DxryMS9ZPFwBlxYwKwOXJIp
hMz3Lv+M2r5YYjlrzEKNZzOi0BDolxIRf4rK24fp1Vji41bMUI5TXWP4GfM0W4+Qbv560SKFA9Yx
+O5rT8m4h5iU+SacDEqf2xTOsKEuXrptPA0mlK9XzqEfkykR0xX3QMXmsVvgmR812calRhhXzR9p
Fm47f2gRQaWVx2tXwxWczi6Qk64KF8FzLgZY7PdkA0dmRWbcV7f7FPfEoU2GA0jxv3fHeZlIuBiL
fyHPErWlLby8OSw2WTIKtj3SPSyvfLC9FPMvqWqUSOoMXQ0unxn/9CKhbd9u3h3SEz4glZc4hTN0
yY7aT+1rxTOi18E3z1cEXy/UQrn17IOu4+fFZvlaVbueXb9/ziswiC17jKhMoZcEP637G4MrQ0JF
BpvOc4BKAKx0ClS5/O09gTeMTJ+qjZtFJPCwkaeTv/UpwTYT8SboI4kL0ICvCSaZTG3LqAU8ahyY
W2rkVPVAEd8rvuuR8FfPyoW7T1nXjQIfv5Lk3OPWjrrWt3EVN/AuoUuaFMNsuU+FPSRWg/mfP+KY
9IG1g3OEzVzpJBFd5xcZk5Sd/r69Z6oTH3hcUkwZ9+qvWAqv5zK+Cvd7SBA0+5Jhlg3ROlON9UPv
Ci2FLut+MZuN/hdcYAS/vAKqQjazjCmJaOg5DzmE4rcKlI+IVjxN77IEOvRn2/Pg6ntjGilrFS1Z
/OupOObYuto8AKjYMpfCkqmyAjQNJr5cieeArvj7SmFjsXEC8ZZcxF3k8LebGir1/Gl33fMvRdJ6
+nksqB5HzNQ0sslNCjSxiGEpEhMPlssTYVxKsRp//XvdzUhxmVudYSqSnx5zEM49PVh9x3caSuM7
NWmfS0kZ/pI7qHtHJuf/zwY3UkpxSCbJbIRfK5gbyZrfZ9Q4flmj9v0C84xrrHXE9ajYnWDcIOQX
qbaPzaQJgH3vLnL7P4nzLmvN9Y8fe8y8xKhYrCwDcSmu/7kDyzwNrZ5MOCJc3HL4UKkbPTyR3UA4
vgTaE1JUENLYiNw4b3gRoZlGuhDmLyvokCFstM3uAqAu4hN/4TC6HUXKCtzMiPOI7EeNboB+Xe1Z
KJ9XyQ3LQyvVhhLlO8L3/vqjNgiCiCaVYJs2SlOqEzBtC+DY+aXTJiRnn8+m6jJPK8flSkFLOj2D
Pad/hu6m47O3lB2QjKK6jAh0L2oAxw/UN/EbsHaGXiIX/DJJR7M7C22Wm1TT2EmEPyUvx0nuXzuL
sHyA3OicHXa/J39RxBfEWSpE+f8L5PoojMOnLM0THdO8stvSaH61FeGnZN3Ko9wHjDXS8JkL2d2y
uLzrK+ZOUp2m2jbWJNwMDU5+YQNlwSvqtd1JCwi/2SMZvo7yUyr62HgfSx8/ciXOad1jTAow5ghe
hsWAYvaTNoY0SWUPLES1uvjnd272RpshZcGW25buaXXtWluFCfQ5XQ2R6BTUbacc0pbtdBlaj4wM
MNQzX3CTaA+vtLRGWm0pRsbu3on8HXN1XerB2H8o4RiX34JwCIeSkpD+fAkEpEComvVRa2Fi+mZK
OO+O7OOgw19vRFaQrTb52XEofThWzizxP0kjh6cSDG6HdTMoLP0kI2p2FLQtURHxBLyhG+IwBRsU
TE73RrTPQYhxuThE2jkzJpPZWw8ikbMKgIypvU9531HgYo564Co6ypYGWwPe8HCiFGDVItV7dz4m
vZgwH6YnLD3SMx4pmiWSVVimqeRhI+vOVde/c/pJDJdtUgfXB4mbac+xR0KYj13X8wrUGgEgi+pq
Gq0UQ6EB4UlXkE2GxgNaKde74Oa8rkf6vU0Ri9tR2bJlHI9CgHI3eiEUG4JNpqgbaJyAF/vO02Jo
20R8IvWYyVc+KE4aAlCHTK9lWkYkeoxhbntl1FnaFDRy7Xh/YChEmPYoYGMhM4Vn/blYsrtL4yyZ
MSonW2ZH0gaPhpKM+lkU3FEip5LR+o0hlIAtWkDXrJi1sAB6eIft9WA4Igz9fMTtM9k4QwtZshy7
j1XlOJ+fPYc+QdqCNMyWW4no00JaHnoc7HQobPZ35TiR3a7FR/OUnAONAbxkZKI/5W//z6mz94va
K6D6TGjEs2xm4OGP2g4rTUh0XVi9k6GMEGtYxC42bkguNHJ6F+FdkfBhFD18YRYHJocJmv7IRZ6a
gj/7TAW+AzONLj1SkdDEPK1ktT0dKbI5cxyfWdkr1ORtbpIp1q5AEG8WmLuFhLvQRIsi9WtAv3R4
t3NvPnRS2a7Hk35izlVo9sGStvlrl+S/It05BJECPM5ZyEqLpkqaFeyjvVbVxhMJOtpWVxkGspAX
J/eZ84936JVY0QQXze8zKVwbdMTHcusVx49YSzu3MxCfvashGp1oaC80XD8aAuaFgMqJayV7CEL3
9QUnEVhpNBifRQK84HCRKhOVP9WiabZySiWvnm6hZ2PlK7XoshqKf0LufvcCRxw90b13m2kCTirg
cIppwr6aPQaHcoIcMmu1gJdYCZvBCcuhNXc7ZkocBx+kENih1WMPXs31J1xxGtMHZmVG9G8RE48F
m9xykOvTtzNXBJTG/qKzCpIuLzx48iLmx7WuG/Y0EIW+La8qjuS248qxjj4gq39gfX4awU+p2EFp
BZdF+f9wzmyWfpN7FgQ5/maMt5fQhRDrD3TGx7Jc+Fi8qCzM7S+mE2aLPhi/IVSQ0o9+QfnBC4Ec
dnkZ0+mrlfk/ElqGJYibmezH3A63tmB8PMD7VnG9uj5hP4OitMrNKIFlZpyTvQMlDEvWValBs8yc
12ejnXV73psak692tkSnHNoP37pRnDsEfohHlRikYowW0BThNn5I5MqFRZhVoj6L3AuBW3cxyw0L
0S1pAbvrtLerItS0EW2yLoBtXF2q/icDzF0+dg56L1tqxYRGEUwB/Q65xnhFl9ee+KpaUM2VcJ8k
xYDl1e/VVBbXJZziVrDRfNmpQAH5rPdp1aDEb2hz82/4Ii8mz1NgLxDKKujEUHaiZ/MjMyOT2eJm
34ekzfWWTubSw4/pm7NQoS5yO4jpguBss9T+vHob6EgTZQqrOjhtiWVnV7EzxdvFwpYXwlJYWvlX
pO5RCAZtiYv0zH/4wLsdQch8VKzIcoAqrplY5N+HOeB0+fUYaYxdhqatBlcwNIFo1xyEvcByRgWH
dueTJmQziky5/UlxFCDHYtbdTAD9olkWu3J06CpebKK1vMh6jQ4EqULjw8ETPC0REZRDB/xdCG/g
0q2D9pb/nx6kAGwB+jqNy94WRWFI56bq7vUyDc0nKUf8eGtiH7aWy1gR/cTNA7Vjm7/hOeL2QA3c
dWhP2Vvx19zMHRBgClktyjp4ep3Mi8XSIffUTyd8cTeWbL6wfctQEvEioO0O5JSGkgUZZwub0xEz
xEk5kU7yjvFw4+nGA+byWpEyhiYkPkXx2PYwBvKCZ667UWppA/AVnpdDeTU7GYqpyTHBxNdG+1uh
NpqXgMsCTXZoP2n4fBvuU5B2Td7ypv/sY2gcRsPGYHim8oOomQIJ1C+9VANcDbdNvZviD3syc6ak
AqQ9Qor4ZVR1s546vNKf27s1AgHb+J8R/cH1PELxmF9ZSCIzgeP5C+RuI0mlPnJX+36kGzld7YDn
W5DlblOcyTV8AnRtshhdIYnB/yZkJLJwyh+fM3xz7c3ECAphyfJrJjWiNMkVfXCZIjaPWpJJVhn/
YC64tpFELc4xI2Vtv9ABJDn/SWrI6vOCjaaYxJ2eF1ahf9knP1NYb/DDeqxcHG7O8hPa2Q/fZudx
vawvj5PoGxfv4LQo/RdhHC4jSbkhByxBXuYNFj7VxnhEO2A9YuUWx8O6EZ1dfFZoDbptPHsdh8Pn
h6CCXXtREWfunbtuxvJbL46WrEpBMswohIDm2ji3C0oHwAhg4F3h1EckFxd8XndgNPju0RTLXcNN
a/DQdvqxYoQPKD6/bcFXEC9WhxYhUvk+oBMh0EEVycCJWAQdubcUvCnSQDIkoTQF1KgxYUn6WjU7
ApeaI4P/hfkffNGuh/GSdq49TkNO9DT5IFowVB8OPkH+33TrdA9hxYSR7x0y+XAzxPkM4gmYN82Y
GWgvemTerDrz+EsHsxU6ZxZULh6G70pWrIgCOtMPhBjwZcoOCgqd41e8zPxukJHLRd+2HwqXrY/h
9jflg6Zo4ErvzL5ZPHo/bmeWl5xIllqPEYbVlLIHg24vP08IZSVSIB1io6gjAx2VCemMaN8j6Lwh
4HfzfGLxICsBx2BOH7dyx8aM3k3UJpArnruv/chm9v3BiNeJgyFm4gqjSzy2wGxom7qX6ooHwWFi
9EnAE97iL92X5WejE9KLHuudq9uBOvIz8g7ri97fzo28nrulrJLlU9bvUiGLpOminNfySVo6t2bJ
tDGRC+xKNSXT5U3rH2IX0hMivhgdXxgWZGSTkI0C7a5TA7GPVNS7EKIfI7sXGbxW8PvA9htNmyei
zZirVxWrMBjT7t8pjb88MGh20TsZrHDdH2+WesUrF0wnD7+EmIJlcaohVyUD5+AG9nid5xmobKJK
xsQ8J0kWsZBoZXymPU3p/jiRbvp+jk2B6DuaLQswNsxBK5qUHfqEmodF6BZeXioUtPPAUAzu2T29
g1YNgVW5ICs5OgN32EI9/6mLfkJ3h1OtCwRdbavOUK5BCPRZOGMWBWid8DnWW6SNe5+IlcIyrUDl
HEIcUpR1+API94DGtSiAuQ6eZYgwKT3io0yGX2YcXuRtEb4lYnNpgWLs48M+MrfySrdhWlUkKMJp
wU/4MjP0jVAOauhFfvJ7wv/csihcZliKsylWVRaIpd+ol+CaZf/pHYnMVye9JC52S6aqOhwWsxIi
9rpipbKguQm05soBVhLQx9j5orGjwLhmsuO0nU0D1LaMnx+ZOBA1zK+2gCOvFyUNmRhkmBrXfqhu
H1Qi+ecUXZEuaISnBIPhGS69R3zlwegxFYdyh1m6G3+mMcz0FLy24IRLIo2WcEo/BV4j1UWw+wvD
YHjN1hBnj9ThXv5wO3OWD7GgesVqmkNcWHC90Wc79OvLf20mpogvCCtoEaJK3p7cMteWKeQiTnGu
EpOE2MilNyXCuA1PvL50TDkGVrrFy0fJ5/QXRVm1XvNJK4ZRd0bLWEzuvBmdZcCal0uQyk6sKN4Q
nsIeDkjhblfXFXIlCodoQrfWjbhGJXIoXjfCy3qqqlQDnMEHzXisj/TUIb81cOfA7y8oGRVVm1rP
2Bt9mU0CEY+5p+w5y6C370t9HxXx4aObuspYxHQGzHqb1T7abHzb2zpWVy9ZWSga+jiZk3ncA1wO
r2p7gH4o2umllSVWV44uv9wwEZSLuoqJbvHPL9DlqKIXiK9fmjGqDl7pAhig5mAFfRNaQ8vJ+j+P
EYV/yro6z0qGr0nuHrijKR8QuCU41NMEdpe8zwX81WxYf4DNWLqe7UWneLgSbRE0023AOwHVGvk3
xNeFV7cGudPR68yuK+Pz47eI7UwvMEjMt/PUaGywoScBV5a/Jqnsb0cn07fFGGKzoFvFIjmR6hAz
C0oGcHm8b7e/CjJKGCKhACCMB4MdazMYaK6AAhoFg4O79DixHq5XX2wC6E5vUPJ2I9Snd2Qeax4I
JdhRhJthdRos1wHnLO/6VaBSfIxaJJtd1NjrgrTKZu48C3EkLFN4j+q7gsSF62hXAWVEdfEbmmC0
Nsv7ibD9hJgUOshdja1qa8wOg92co1Mq5xaRzPwmBqSeXAbnu8OOOoagACVvD/wFg7HJL7v3Z/Pu
HRg6Ptlb0IRuACSZ67B/MaYbSI1Zjc2j5KO1Nw3By5JWOs+VB+HEXF4pCbd3v+/+l+WFRv2EfM56
8YeObKKEy2VY196pXwPywcD9ARiFvVyCuDyp2+4TGl03xVr69ss83QtXdHXxR05kCZGqamRBs//t
PojM8dxAlZx3fjCec4yZeSU1kv1UVk6y6lNgjuV1XwLSEjolr7j4gmqeBAjZu/3xfkah+wTXitRO
kn5T3Fb4Z92uNnw8A999HoEDZ8uuOg4wHDdiWlhXHu1znPDuLU6hTrzykm+gSyiEHiA1edDTVdT9
xSpPiI/qEWvr3qWFVq0YnaWN/v0uoh+LTMuan5A7Zm7uYzYlLCk/bl/moMULa0BdWTOQEsODvmVP
/J6Hj0Kg/1BQdoA9Bm9lkXPU+DQoL5YUmWqtBbM66TTSk/tpc4X0Mi6hy+PXxSDzfkjVmNM+sW/R
CWOh/juhZYke9TpDem8GTZ7go+52s1BKeDs8OsuVjFiudf7P58VdBtld1MfCzBJ35xFRyyTeeap1
xBY4El4wHRRUQHTLVFOxgJ3Zs2A+CVF9Om/CcmIh2qQKXGXhEaoaunxtGaCk4ec7DeHRHp+izXZf
LaX6+YPqcvDHTFqy+u3pzeY4nIU7kIYCmfanAKNJKdJM1qItiYonzYSUM9Z7iLDDgt8UVLZ7GePk
OrxG41KrOzwVnhC+vyzKua+v8ToFdcw2DlcYsw16TKhUVIElXKBw3Ic64BnFWxVI8J7detbnJTh8
iz0k6/QnMjkdTesrs9NdfcHvyueYbKcOzo7T2xQF1YMuLVXbUuzUEo+P6BeuEi1UCMUb66DQKD7f
EAvfTWLP8AFTc9A2DmbemUpjYAj54sWxn0hMno3txRFbIlx/hBapL01+4WmoVrh5qNhwGVjN8Qh7
6gv+48aTwlYv3cTBUKTbIM8ANIfm9SwK+HFcz3kniWNXUcCzryGwZw+h13gtQXzWMRUJU13ApvSm
/48n22TGJJdahOehfo/X8rOwgLK3RsDFXqSGQ+UMOPF8X8KP+1TlkwZ3rCb7m+cSn7lrJ1IyYgkf
ZkrfjZoisPWyN/5O6lNQjZyivwNZ9jHBiv1sjEyBFVEA8IVLfU2Ffkebjn6N4LN8BdbvKh3vuAiX
eB3i0NcqtczkRrEdP7Zrt1VUaNzvRtIvv++KdkX/ZyALqkdRpzPny2YM9YEHbCM5QfSwgaLlhumT
BFkh/opag4H0riQh5N8xy5nxKshTtTI/JUjRqtiJDETzRny4+9yY1HkFmvtuHwoaj2dS9wG7aTsv
lE5h3Kc6whrvPi4M8R9VUPLpkySREuW2a+IPo/CB6sSFRNGpaV1g6yJPe/ScsbbvjnHDjQmelI4K
9X8e8uoeTfFoUipYqyB/n17qulCJ00LHP6mUPGQqrmnblz6UccMWaXu5xDQJVPvDFG3/gqvPVxK3
aXWWX6Sn3V61oPM+Ve/Zzf3xv4vHn6TzMyFepWrEJ+gA5ERia8kOtKuh+GxFYHTRpiSUl5V+xOQl
4HD9tnEcXpl7nlHpBpw67zXTsnQFjlICkkUuDux5SVKaMqyd/gS+ZNn4RqPiis+tT5dUdxSI57c0
BcIp7LlDrXxG/b68gofuAtk70zvdWgRoLsm6O2aIdbb2KSbSrrNelula5c7tV4/IOncJBylrjiq6
hEPW6WDlD/zWTwolwkVu39UxYF2GZf6TmkDLWGVK2qMaKn6oijNzU2SabkeRdLHRCqOhw+F4pLaS
giUfW1SQ2HA6C6qF0HG4XEXGDnVMq2RwCVZlZ52bO5uKdh5Avz2+hn127H/laI8w2lilWxTKANnU
hDqF7rrAR95txbufn88u5y5CyDs/YeyQlk+H2YIobjjVeLoPcK64CXcJgSGVJoGt9srX6PxF2EKZ
+KtJ3W/jubLUUz9jsqVw8xqxlf/wE6xKyMv+mxyzq4D/pnStOVLNSLjd8A31AMii+eQMaz6JZ6z3
+2xiunfE/ntlUIxn6GWdY4+dj4RZgj1tRXbLGQq+3dCuDq9jfrqIdXm3RhcL3eidtKf24DVYM47l
/C0uxygC25ujnwG3iR4V6TMCf2w5wAnqrrFIeKtVXqILLuWuliQbImkyQBPeNRk+YiuIp7ih2O0J
gFPXy9f2G5fCjuveAVwy49Xrse5fwTCkVkB0+JlHmm6RvzSBYQM5I56P3tbelZloNOWUpNKfOyyc
mjCo2gO9RHX+WKanYtykJ5fz7FhbQgMk4VxozeN2leikZAVHPJOKK9D4VzmU6kgqmym7Z5G43kOL
Fof49LRQb01b+H3oLHI705veoj/j1WKvD5K69mlhBXLH2D3GPgNyeBQU0TKsl1Lh7Khfg4ZDpvgQ
JxpmUAH6Jd8UdbuE7fmKdGGvHR9PImx7XEKv2gtuiIef5oE5/G1vBqUZC02aY9ivr+iGkWITDPBX
+7oAkht93SgIvqYglQppo7ozFI/iOwvdCc1dmkcdn3F1pDNz4QOY4Wq5q207OwzJlD1Mn+UJmcyZ
z7iZNn51GebyOk8KfKQ8Cnb+3/J2AA/UMq9CAvw2JsOWiZ0W0vcvJKL/MWhNUxjWVmkcNt3uFt2V
OpmrEVedf+34bln2WhTGmP7ODyUdOB1kwnjpav3+DPFc43DOllsqwm3BxYICYDPzlZ2TAgq/IifP
SypUMmWDtn15zmc5JFXKx3ZhIxgRtejYlzqbj8fKnaKQM2+E9TwEjm+akOgoUXPnwgCk+J+rk7uE
BIWwkvgadYm02QI8N1zHPTi5jsvsUFvLSKDPucpK2hzrcPv5g8bI8exxxvL4vGDfIie97S3PiwhF
LCVDp10nGcKygrOnZ0YJCeLtYppblOkEoV822JZwY+t6ve+Zx+2rR1h08ZKBr8f9SZ0ehKcobW6T
HplKgcHpijhivm6W+OPeh0KQl/PLKcwOp1p9FHJqQ1boOHpf8J+mWOi/LCOnSIltKUaMqs9o8mR6
yN2UWQ/EjNP6qsx5zDRnhmLl9NoKdM39W9/P2pcAaqjOa0pS998u8fZpdPMhu4DxQuCejLpNYVGa
y/r3Tlu9ecrpyRED5uqezrCLKamVVaAl4MVH1E3dE6DDdxm7/HxfFei7dvuh1WzF7YsuoaanBBWG
NtzN6ETZtYHFmF0HCrGpku8XByHK2imGHkdqmjgznJsjoEhfnR+5u2H9chT+b1AC9X7kWZXcH/jt
gRkMpruAynOIWgpkYd+gVIJ1tml2FDftAcIx0uH3mId4wP3HZYHnWbRVxP3xNll3PfkC1hxkdLGu
VF/43KY5hT9meB2tkoeI1besY8R6Abn3+Kih+7xPGt8epGYlEXaGyd9i04t3KgmdyrfV1idVfQj0
06rECJjR/mmiaHXRD/BOGuj4Wd25u//A5WY3JmS/mT/mwf+WKEOW0tUcauXI2ULQtO3ej7kmZU27
H0eIQtsMgd3zkaZrAHEQeU6XaFsOVsjqQbAWaDguuLVWQAmChGIGkBTQLwIfH9AFqyCEFDWWBpPK
rrcLMauPtE7JH1nuurwVHpgHlvd9M2ozSY07yRZp0lLA7UZa5nfRxAlcMxDTW4L5ar6TkQY7Mh47
cqXwZlPLKGFtnTFV5Bo1v1W6Ji8wn4OgOi3locKe3kvkD6hmuteE4/UXmvQKgQBlyRaiFf4rkaGy
62Af+jU6KdksurlOY939oauJGYCx8VJf+NVCd4obNpDlB3+PizQoBb9ujfkWKcj1c+1jBhtyJdAR
dJRJkE4kWbcXL1VGJj6jsD/0pz6IhjfXKclcOvzk7Pvyx6DDKnoLJhsApZ8pVgNKNi1MPQYKyxlG
wBwJJ5mCYzOqu3XrJIY8qxL/mxBRc2l9PqGm9JaYEu9oxLSX4onWkeecBf5D1AUyruuT/H6ov00G
c012vUO68+PMSYNgFVszA6Kdz457KdGxh1ZvyMmZJZA6xQk6ORNrwcThTHaCzr1nlIQO0whoRwgi
al9odeqvW6sjqBRIO+9/73QjKFLOn5iDOj4qazbKw5dXmPfxKmbHig16bAzVjKT6xC4VBRE1xNBq
3qxA6EuVSXpW8Q2d8pr62kQR3CcNHvg+Ew9jZc5vOZpMoYXD3gYNCeSFhhRO3/PFx3S+NE9Zq3Kv
jHLXntEwTPYMCPOIprB9nbfGvhGLdV1iHJ5eQUkkZ+BBDiteAFSXwNf2Lzt7sP/6/De3JIN40/ci
rYrAQR77WfiU3/4yL6pA3Zwm957zACLN0e1o6qZzJn0OvNtllJvVFQZRh5sJScBLDf6bzRpZ4FE2
tiu30X/x2r0HzNrymhWpAImy2KLlCXeXeN/mNV1vPiGUfVPBS4h0rczotKr8DqqGVM7+5bYxUvQ0
XtkLtAGDFe65/qMvJ91H8vPpWZqdmHzx6uPkCiQZ7Ya2+Z0p8Ao8eiiNJ6+Yf/F44FfCiAuRmQXr
RVl91pCmcXomRmA0sBpAE+kfvfeiDC99/FiZ6SwKptla93SzLO42LGeVSi4WArdXgx2lqMENcSjk
iKPpOKbXUyU0ShOmM9MwnJbRbdJ36WswFnUfmGB7gUtjcbObKZ5aSLlfwXgA0HJD5qGDJHlAYcIz
jXIcmbf08Tj37mrecDrZ2sfsgJsDhPBAP5f5QvqHVHh5R47eGrPmt79lsRABnd3ryg5yIwqKORQC
G00KEKbUY2i6TseBPcgw8ElpyyfQF/fdUFiTaR8p33IryFgZ7rD6wrU+gwQHrjhR+U2LNHZUFZzg
yyzHM3lzZIJKSEVvawJgggtYEVDsa+W0/OkiuHd0WlDkSY8H4GeJPec277LITjqY6xTMyeKFWm+O
9RGf7/xiFG2H9UejNfb2gv8t9XJaXWm/jSt9Y3xbqil9IybglG45FzQJXb4b8i/KOmJghoBYJX5S
vFpdR+7IY7mALmw7p6Nfz2RX4HBK502MjnnRDnqdODLk67HL3JvzOU5XWDQObNhAtmGhjRsVfIT4
4aFQZko19zzBvIGDYcdEx0refgm/bxYM3IPaXfs9pWsgipR2bJ3d2RfzK8dUGOvOiKZ+Lxqux7Tq
mgJqJLSww3Jwj/SGdMcmZuW2+JzTi2+O0jt9mpeewHYV+1vOIXfc+xs0J0JOcVpynI3V3cp0UPoU
xG3rUKWE3rLNAnjbCIoROp7sOaiQ4ISdtSB4QEpsqvQxnox6lTeVb3yrPeU3+R+jNe1+c8Gu2M6U
Fl0oAC0vp7P+ncPhX2TUdERu1TLI69lDpBXavYA74/SXZ1jnCp8o8LogVl7APsm2cYjJjLiQ8Ms0
jM8Vt9l0Mx1KXL4Hk4zFPs7WryNYGqoOPJbFv01yYm0z+RVosM4PryBZult6omasmdm68yuNUOK8
/kmnVpCsMmG8E7Szpm7YWG1ji0i82DrWcUNCvBJpOhtE3OMcsGoN8KtIQJPHPPDlOZPUFJTJBoB9
P124O+WxXAYwgtQPyQJdNVPLefI48vKxLcLVRyOkZR9m64OjSPoowigvOJYbZa1WmhtiYVPoaiBh
PXGMTwS7XU0AV+2gaEc8s+KG30w985gIKBSQhou94cf/a8FdYxBwAlKi5MvZAlYgxvriQB6Uf5D6
FsquLD1Ae6eCkGVDuE0TBgTMvnxRQ1JOnwJ17lYZihzEWIHBWNxIwDqaVYrQE49mXIL/m6eCO8Am
ndBhV0S5LSw0QL4W+Ll8fnFc6SA1cDDCAQGk/xkmm1RIonnlXDWjoBtft2y2onIwMU4pSaJx8H+N
noQ6n04V1ngb6kLlcf7Jqd+p2ujwHr/0d5/YPslv21b+d60Uo/dJ8M984MPcdyj8Fav+qidc1CxL
TfPl1grY3TFfKA0d6JFax5ifYC2K07+vzt57iY03e/TrG/YQ/xN5cXEI+pDa33Y6b85G5er3fL6k
OG8jnkQa2WWTPDqa4N18sPnud6b0c2Vfi6PGouQM2V3CmNLWdu/rSWvCWNL9RSwPf+Gm1O2872yJ
9m4Dtx4JECSOJyziMmSXNDm8THMFJQqpyZ30FpuI99RKG6n1lx5qnwGYlhSU9XtOUQUpEn7rf/uJ
cD+wXNZQv0xj+afA5hk33sO5rx4F8d3GgVvleLNbvMlSBN/hfN88fBginV+4rI8XJ6ZFAKlr8q/K
pQNMb16wmckepikwDFnSwOJeo+7vUz3yvNFAEPrpWUEYZ+GVqVFReqmLvm1RQdaLyDJ60qU8A+5h
+5nOEzOncxV0E2JYHX+8P25tSWHzzMqbdlz395P7XJeXFZfQf5pAFQcZZ9poNpC8CEHo+Jr1pPg6
oOfOrYpCE/UJrvDgCBnRq6c4BN2rTn+yxkKe8yGx9854mkdxSfXzkxUDqgIcMm9w+b5/AbVeFBmm
LiIf9f7LdM23tD8SMNwqMtbMzA65kIq6ne6GlP/0lYxr7fSEeb0km0Zig5vsY0VWPbgJfg4obyfY
z7fRDrPQduug0w+aAoRiu7TR/CUcEBlH2F8XqcpWOL6KIgpqEo73UBg6AObDRfTKeyhmuLUw6Skc
9nYZvJonUDsVs7BON94HyGkjWXMC3UkA7O1hREcRIXE62W30BnxORLn1zxxUN4BRIXqwVaN/LHvX
A5J13YCHDiZtyUUtITYLknmPSqlv257agTntBf6MjoWX7HxGMNCfOroqkMzmhWnOCgX8VIEer/xK
oL+7ZAwK/jJYF37lS9U8ywjtcYmreVdqVAq8V57OoRzd6Zo03w0FqRhx3/VZT4DqAjRYtquXTi9t
smYZRBad/Cr5c7Fa8HnUhX0zkfHyB8tX5Th8bU6q/SUN+3/8TDMbibWtBBFZEAOEZOJVN5W0RLQn
Zg/ioYu8JnU87utHhzxfNbP+Ac4knJD8kOU45XZdyzEVaSocSc6J9N1IP8Hw+YtCyoUFfCZxxngF
tlLMerbRAYFgBrifjXu16+3BmuFDjf1LgORetxCh9P01jHL3DbJE77e/G4X7AShiLaUhxTMsg91C
DaHvxl3FUo2HfX8UvS2CzeGoGJTP99L3epN2LsMTdQ0uoEyBY/f87iFlF58E9ixMUtFtPsvboCN7
p3DXL4b9QtqJLFQjgzJmdPInuaZFbB/Wkg7T1cBisvoRoEyx0IUPwebBrheqRb8Ty5GC12l7Nler
+k4dGTclrCRdDojJCj2HX/XaI/DuCDPJLsG0vg+Ghp56S2cO3MuACD5cP+kDW50mHTm/RCLwkRnt
rXP2L279kHCkKf0IuqWDhR0q4tpOENYPOf3p4DvltJb0knFvoMPrC8tqZlgkKSx0KcbVd67geezG
PmbmJKHzPhe1Vm1rsZr0p8NkULfImA8gJfhiU2ZOL0fBhCx25mNyl37QFTbwloSOyowIyqTcXRZe
n78NR0wDqPSA/3hc5y1VRLBL1vodYw7hV/naEeta2MdkjmDN2jmVlCITYAmNpr2uehymGpf9yRkZ
LdkCVLwMnuhB3NCGJWOCm+ehikem840qOlKBT1san0oQqQlcuCC34shBHOatE/sqRgDnlvgayPi8
5BgG1BRw2xxWGcTCZSvW4PyOd8WrOARu65a3Y+DyzBY3iM0Ax0d8X6wrqq75UEOD7FR7fAcfpdie
Bq4pkuEkf3dpKrvlSHDPT475t0Hp++cYClcs7RHAgzNvtHNRl4+wtt2L/VmVPzmOdmXBlGnGFWnO
IPWrja8VmCCXBMKS54B8WMHxxMgyGVk8kAnYudCZya6+LhR3Ht5YTN8FvKP25/REZ5agNVu5e0f9
1Io/fUV7UKOmCw1OXRsBtybQH56bHkhY4VrzNoB0WgcDdj6AMkINOpuyb1M920mdTr0jTqoL+QYh
v8mtu/4JGlLuC5SRh+GMA7dodAptxWPi33g27W9qD6P+eLuEFC1DFLC3ktXmRfxGH2hKmg4tbJpY
b9z6pfnvEdWULFzDfxxTW6kg7UnxzFD4zLJLWl4WDOafa2yyFV7Om52EJjPtunP2iwfV250LawP4
Z26MfyXe7VuhWj5yyYC0eOYbQk9G9UTTguu1s+y6aa4nNnSXHejviIWbjE159/o0hdjxxNTUf1+n
jPFB0QR0/sAtZYrE/9A0WGVBa0/Te/xmBWKfHdr4gx4qfSXm80Wlh42TVDv1t6+T5WYPt+oN1qhI
bQ9uDgZsGtixy1Q+AHU5ZOKVxoKEpBtsd6I0s5ywXGqwpjev+U49+FIw27AYqXi0reNyNCRiEQ3x
GagcWtZaFJ7GBDoW/xfYypP27IzbluAPPeuQ7nCSqwvI1OcXcTK/6jHRACtbLSCCYqSWa0u2Ak01
YgBTLCTlYSpH3bQ/lV7opfwelXwxKljrMTIlGHCJQnilg5o5ZDlyPhq8ls7OY/FnHUB2e9/U+8tx
hW2GX579Ecrq9kNSQSEWjBt4PtV3ej5968k6yAFxQeuSKmhzueq94nk7tCKXw51bvqaDVUUzP2sC
OihN9iQH4CtSo2Vo+aOTy15uzpVw+MJhD/CL1GXiUfKfGxEIVnWR0NBQxyVRfQPpmVagp/yqGUaQ
eG0/tLq8nKypUdnfDT/paiPI1ymiptq9bI42sfA15ceosJm+By95gpSmM5NkE0Eokj6t6T3tBp+d
mq6IURL6CnNcwGrD1QPNLUT8mCuVgbp2cy8z1LlaBIcmV4MXmBnFB6bYsKTfMgCW8L1LYDKJalin
JpXHWMBL6BnKEBrQrkhV0uqfsD9DqsLkck9/HY/m180Zz8phV+plubM5vSuVxmfZzqXiw7UkANU7
vtaebEp/uNAP1Wtyu/eTJYzUb3BYe5XA+EaA++xgxGHKp4SmbE1IM80O2y8/i4obnvdTr5H6dPxR
La9deGtVmpJV5ov8lF2a/cN/VDzjwQ7prz7hFpRulh3NAELvbGyyyuZg9MrnX0wlIL/58htFDZr7
523aZciFqMoCR4tmfyqDC0XB1AbkCddV/2I7zFhVVCFC24dFevDYN6exIV60VYrIMBI9bHUibIYZ
pMzMKXYZo0XxEk6wgPHgWwJsA1bHg55dC6UjX6wb7AgKDrh9TxqaNNmbSJoUMIkbO7I2HxpPAbh4
sjfEFOAtL6oicuBessHkC+ns7tN5+Wiz3nlzZlRi3zc4wqTfm0wO4zJWJG4LDPEwQAaL1iPGJoUH
Slw+IoV6T3ImCF+Tpx/vkMff9dnd8Sd1vdQjzcAoWHSQUsAg0uI7wYFzPLdpUxf1sejXvR+cJoxh
jayBH3+tZF1JZVBCzCyE8REgcA1Fb6qXABVjmZwrsip7V1S9/zmNtyJni+wruod0gh7OEUdIkDf3
tBOOHmu72RC053wbZEPGHMWOrfaR9XEFBKxWfiyi/IuG7Bt73M1seu1xx+eDWuSr9MJWcMuQPYkj
kO0ICVvHEXEPruPiCYKiA56Y9yGWI1PqNXITuQT7fNfz/E5avSsrdp3SDz3mAp1vfANH8+aIyE/m
KCqvM8reWMJOx9kdcBa8N4VS7/ykY4Tv0YNtdyq1Jl9SxzPh4uKeNar4qD2UwubtP4cN3hwZRAN2
M3p0xYRRps2gM+cJtvhXNZcbWHNcSq2hkha3kV3fTWPLb4dj97TVgTeq/hVzMRcl6hHg0fe6ug41
/Q2+SFkV7D4TipJcYI4pxfUvdOCQpqt/AttVaHLwnWHqOI+DHJVLbdVru090FURJTWJTRDM+IPFs
+RKG9g3rRp3L8DVNq0r2b89G0/QlNE8q2a/nyUD4cZVSMgOxIV1a+Ww8wQEMYUo0TIaADrRMDySw
dpGTj9zCEWgeo+Gd5jHQqR6fjrnu7w8DLtAv6WK2rn9O4SXeEXrev3Q4RblMMMwpw5W1Ogt/6NTr
MlewCD7X9dbkqSUjnX0AyvStgcrccXnGXzxPA3UgCpG6Vd0obEAkYDXSPxsUVCqVYM4hW6A6SrJR
cvuilF0BHXEjJSi7yckX+Udlgb43ooyRCMMFYcT8IirlBRzK46iugy97r3FC0IOPBo8KyQVjI/MN
oPlLErP5PlT/lW3nHeyO2ed3pGtgzAjX1YOjQyfk/eEsI39PUt5HJyGGHnQQYp1I5tHMIpsXGur2
qVTlSq+2Q7SPKKERwKSQ0FnaQFD07vsrQWYs6ykswte0iRo8sV6brub007zMOnsj74uLcwr3jK3t
recv2SzHpxhOQjF/cNinXv/7XZMJiq5IUhzO8Dl9OMZgCaWDSjd8r6qs/2ojs1PQvNbEZEapfgZo
M3KykXbAkH/+On3Js6+zUn3tPlBOgOd6rUKSooyZa/JQLBWnl6DvpA2RHGcCTKOD7ejvJN2pJFkg
hvfTBwaxYAQCAneGQ/pMuXTBgvp9BioXM9BFQoJoOZV2zNbT/pbK92xZ+pIBnYRe/sx5wVynI40k
OZZrsw18n3GlAt6jhPHEiUs0EgeVX0BmAwLm5vKFWJyywQRb9uCwLlGU1FVODI0hzCMHFvlFhCe+
HQTY2EKEAiQxBZDnZ4SzFQMZnk/i8bEcxMKUyHqIXxjJLRn8UoMu+9CRJuAEBAdyXDqGFsnu0wOh
smnTYEwxYfl2GISWw6yqOfQF71y9mZam13G/baN/iv73Q/cVE2/yx2EYalF0a3Jd1MP60ApYFubY
TJQBt1VWg33yWX4Bjdd3xI9a3FvfolzMJ9zzdYMUlGMRy6Z6FWjw2LqCaqubgKGpNZbWZayItOI9
/EzHKXXMXOO+sD0knSm7uJjzDJe69PD02h206eIsCAKEKe92iuZvVxZEqCd32mgudVRRRNplZNYt
ahKltN/U4CAK+algu9GMD73+OuR0VuarncpNnBgLYKhWGrz+7XYbMfOthNi0UNk647ZKwfO0SW7R
UU2mXQBEy3UFuTYBoUlZPyP36vlZw02xdoWpopltDaIIb3oIkuaMEeP+ESTLVm/aY8ZqXwATKHuz
0S22td428fMWSUlx72J3Pzcjv/4TAVh8lG+Jwua030Qd1j7ce7t9rGeeKzt1xzr6jlSQNyoUfWxO
0aTnN8VghHTSAuw59Zgo7Pl6DGcgazm7c3N7yiMDP1njLojzEkj9cF8iM+WiuoWjfqaDhbiSv/Og
8iEntpDMI6tHOiuP78ebNz/PMadyLVdmJgnsX96cS2hJ24LFXYMOhIz0/rrc1DX1tJLPiE4qD3Ri
kpz5/nOCq5QyKUOEX/Pj1I5nI0bKZLWP+PI9v+PwiRLmT9YAjAG3fmSdyvrRsqbrJorE8UfdPUOz
thpbply/UcfSgwht3ZZ0THeYBIdFKOs6875LQRzlXXINC6slgY3QrXx53x92dUN+2PysgPjvurIn
FZ2ehtk1/SzUP/dyFoxgdmnmEnSg/UczBxSSIlRGRM0J1tW4qSWl9zgQXgt83s+VfBn10Q2ot086
c2HdyZcvP0BfFqt94kK+9EzocvKKLnsWyLsWvVyrD/Wbuei2EzTWs/Mr9BSp1bIXhY2RJYCEZNkf
F5CxbAbSRFl3zFUH6pvLzZ1JgVaHjJl/z2ReX6kElYs5fQTBZO8V6HZ/sp4OoE3UfbP1x/uLQvWd
Qf2neQMgsR5b8xF36U7RwaX0Rd5OzWaLEcQ28xxavJxGihWKtkJPsKJ4fwfG6DYWnKNuNIrZEEpP
ye3t8kc49bsTSHbraKVwepXuFqWjuiqyNKIMyOYa8ZtIp+vc/Fzcth8fEslaJcFakFMzU0PANLkr
ACj1cMQac+TYi8kTh2xtHtO5T8+MZNj09XwwHaU0tIKPvGsBv1T+6Tnxphrc5TvFfJ0Ote6h0phG
ywlC0ngL9ypLb5zy7f68VscyGLmwEX/ZVDW8vth2wESUtSXcj3r1/d5NliJgBO7yVkCDz+/1ws6j
YUvpxf5olpkSZWgNsRERsEpkZCdDAJIDYkTkwgW3Kh+Iu7QpzFlaMcOLeH64WFVdfNNQLwoyGd2z
idyA5gS2boJdqo+5FcpFZdU30SdTSXvUdK9RHcm6RKFrPBIWjAAhML2j58EBLS1SY7diPIyg97GU
thix5BvIiJ1gZWBmYEce440cdegW4wMdUZcJk8U5yoHKoU6BjbHgNNRnFrrbEDhZ/AkH+oDqJ/z2
VLUa1J6c/+snIurmG2F5FsdKITyOtbqlbm6hQWreBF8sZXNOXbQ9EB/Cjf26tJlxsLc0OYFvm6rK
q4dwofi1IyXP9lMvQSiYCPdFmTKRpw1lxhxigoy5Jz+Z4qb6AU5RcBSqH0p4YZeMbHo21DYnXqEQ
cDK2h8PGmjPuLyrYcU5XuNLt1CPuQfkFjg9Wkh7XUMLcf12cHFBD9JhgTg6wliiAKA2J280fJ7Zj
mBYq9WMz2dPPzUxA9mD56uL3tH8J053WlZXwuIwvwToUkFMh/7Dvt2PCeld2ue7LWAkTqUCf0qeR
VXNtbFFrFmjPXoSn9shCzBvGM9Fquwwz6PQb+/jbLccq2GAah855YFRLCTK2iXTU1+/skzLwlsXD
cQsLzS8odd6CRufDtA3haJgG6+baaCipcVLDDwD6jIkwDfoj489Y2jDVv9DkBJs+UlfroAopem81
KKfgpicbytI30rMFubUqN37hp/CAwFeTdMyrkwCQZ6UdWbBQ3USoqAuZMCy6SmNehRU6EB3eVi+u
jKD7eVdli+44T09mx0PB65ZFp5jV8l7IsVeZbM7Epsj7Wv8IDbpl12Kju9v1wwlnlRMXNH547gA7
eG/L6oNENP1Hokr+bLpTR8lqlEFoTwsFPAw2j5LQ3gyUeBAUFVqlNFmayXkFUT8CIP/w+kTDma+L
JBL0PqxJADOXg3r2+O8ZYDFPnFozXPESgU1wB7Uy6Ek3aXfWG+YSi0qqDK0Cglot7h6XNgpqJBxO
tsJzbLfAJbfGcdOLM5eiBoBT3UKkkFNm0EmuWd0lBnxKQm59CdBqyI/bk+F76iZKeiPrWxSlsti2
rQaydsiklAqyCzciIumgWwUpapsQtv4z8bYIGXt4jqSJ9NfRMkS/m7m4EgkF2CUgx0dGMbItcga1
RuU9ta6fUQkoR7JQb+w6TdGre+rAdEhIlLCSrjqG15ovkS/wXdtP5O1JVQhGLqDl55XrdM03XbQV
WN8k2IB+RFiBgrMiNia3mj4ifRjsqNbz8+FOVnnHlRdJh6RcpjqNkVpsvqi320L/Ti8lnK+ZANun
VZECOUxOGOhjEzKQ73fCby/m3vrwIEUfxgpB+WYQiwK+xNwut5mKcFCYHeHS205CN60xe12mqH8y
ghcRXqCWmHueXJeK/iE6O20SHMBII/JJZJCZkdYU9yRu7lZqwxmSxHdGB9HiH1axPwfffP+W+XhT
bzYctZqmnBMDlmox5wW1UW4/LE1eyKDpfokr6qrbFBQe5nbw3wh2+NJlU4ScZZ+7jDa2KncmLrx6
+/El7z/ObYc5tzZGPhiRy81ovEyVPhdciGD7zLzZcAbfCFsKhb5Hx+QKwB0aH9YhCJGCRvY/FzGu
uj0puKRcCpZbKphg4FtaqiXMytkK4kT6rcpboWgMSMb1Ltu74izdX/dwoaIPYwFuNxenCcwk8zPE
+mmbnc9yJRkxLvg+5Rq/OvRkNR8jjpC+IUANIuNRCOtajHgO48eMPryO3PfE8uF3eSN4Unnu8kwj
G+9J1oMq1gkRJTIyUCkLqOcdZ7rd8MhpUAj3wSHfL+H0Nkivannb8WOwYwvytbmPfWucsAH2c8bF
dd+RwFwgsOedkqz8sRDFBnXWzyGoaKlyVmvWhgSEBO8aVavdVanc5JoE2ehr6od9Xh6TilKfba6l
ElGlDR9J9CiBrNtkifKvxuvx5L8wsLi5SQg7INjGb69kWU8WghbjWcaE3Cz2+h+gguMgZp7qypP4
VfoUpEFHGvDW+cTgD7/ylDaFsbQFCgDHYrKWc4bLkvbaN+rc3xThk5hEuvwwUMiQyJhRb2CCXH8P
7UNWdJptuFyOZ5vnDdD3UmyJ8F/L6/HfFIjs2UHRQGSn/EJJuq1MWzFEAEFmzponzh5+pAjIT+Na
HOwRAkYMLj+TS255XrTT/bTMn2NLgTazFsZbqm2tP3sbbZOrs6iPVFfezmWMuu6C28np0KLaDJkQ
f0PecUrE7m9S+NhcYa8lsA2tdei43MlP4qyNQikCDEGTEKMQ2UU79mrUU/xaBTY77vFrxK5skOKp
s/7mcLuHngCimq+WFIYBbg9LKqm2W14l6wfcsaAEwfLV3Re8mggpB0C+2PPs+aujUYXWAvPxXUyx
JlYRSmmtZYsKJkm0m9+ckv2iWqyjLK5G/h7BgIHaVruSJUSXgLvQAsXICovcF/SUtTV+8IWGVyX3
CCIcDfpgl6Ac99ALzP3wqfomPL4WBsKOzQX8d9PZNjMV2nExGEK6Jns76Bfol1ANxqTDd17FGjR9
SODlCuJUNrSS8Ia7Qw4RDfR9Nab2JzgZy3+tYvLWJ7FLbA62ot89X9v0dm9Bscvyfw9/jBM0tmRg
8E4Od2aGg6GQ/XwafIt7NDQ/ZSM4GeW35O2V1M1cqrnong8XquJwbY40hO93t6MBszm1FAoDR8BV
DDjPNZ1fEoDImnLM6IYja3wyBrkRTo/ipgscw2d5M2riJoHYSf3N7cEooIOuXObjfTCKoMS3ovEI
lW5DiKqlN0tbcH4gZmQ1mjKhPIdKiC8n7kHczKFB8Oeirg9f0Z6FKzdasHq7CKfIcV79KDyLWrjp
r//CrmpUfo2szikCsYteT+1wJ57nYnIjMqnOsp2E4b5PTRgFyXqIzV3jPX1ZQ0Fq7FNy6aNw1Zxj
UitVF0PZVKPwD/D6KYZ0yQ38hIIwQbq8IX7+SIWTmSYbBOPlHtykS5JmyUzyfRcjJUDjG0SzqAOz
OnWNdqSkYxkXmHQ0YQFwMedornd2W1DH/KACbtEAfDTyLWU/tOSylU0U/XVIOwNUoLwHzBYJeP5a
YKqC4G2tU2CeQ7u4yf4+CbCIq4IgS2FrIok8nBfKnj5NKsP/NQcgEamnFDTuCTlKoKJYRxzEvarD
dCP9m9Vy4O1Hccjj8Ue6s8RrAPxiVdqfx9nmkreBOt/DhWoUAw+rAGZ2JUV1HyeeDGeZql2EZOTX
dY/rVQPBbCkaxueEX9buk5DSorP9Tr8thwXSspMO0zhKMgI6TIAwwWHgLL0/Q6lcryM+zaHgFIS4
iImOppv3QW+tgSizB1AVRwkthnRmesr1myZDxyr78BAGWwZsuLRxBDd+/vUaqnukSqLDwwpDoI6g
RqoY/1qqVp+Tcdl07AhOj177jGCGuocl/NVJdA7c6/XyELCB2FQO2l9DtlrNHyCWeuiBzsmflZlu
g0gtj/f6plaJgc/dwTsjRDYoG4Z22OOTph1sOoA2BL55PaGSUisqcJbIkwnOEm3Rno0A4kn0wrF9
jnpDnj5816zaKo146BLKEI1qtP2n4qaTFxXH0rlpm17lZrIKsGGyk8GV8qB5nJe2rnvsLmz/F7Qm
+npIjxuq+sS7FWkg/R0gfq3vJzbkp5SHi3a5AbbTokgh01rISzdL54UYIDGIBuN1i1ScTNEqGQ1a
eyUw7YOmEQ6+1iqgVUVuDJ89KBSgzQamCsJG2b7MW8nFzAd8hoTg6YGBYMirr1PFtnV1IxA798nH
YffI8QCum0mw0kxoZrmATW0sl8nDr6D1wcY4ZgmsNd6FvommGEp33UoeN9tMzhCgoAuLpuZUroEX
CnRG72+fYFh1i9xkUwyQeNTnyk69DJKyXsGYs7+9xIHHxsuTm7Uh1+/y5f9hfitJQyjIklDUYVQ3
FvHJCNFJr+heIeQf4VaK/ZvsGkFpzjRUo5fmcR5g+GRGfYQri1iGmybffkFswyfLkrvK7CkzSWfn
QyJ4qP35mEXf6/n5ScCpKZk0ioflMHV+zUzKSoqTMDYhanCl2HDJpvexpJbMCNgqqcu0+lb1D62F
rQiCkagzKveXR9jPbIhWz1yTzOa1fMsWjX9A8jZb7Ee4+wMigCXEebHjbH9Isp8p92PF6bW5saAq
EWehO1Hama5/eAUd+eVSy+Zz9N61rl9ziQc2ATvWp0RzEAM5isxbJz1k+o3rA6kTWgVjS8saNzy4
NFLfeliv+YYXSFwKjU4gB+QWkYziwWfrtuIT1Ss9zhVQ2/x0ngOZPYPkmyXHXJTPqWvBh45ZP13W
BnTe6JrO7Biu9ZksX2evAldIn3jWt448dmjSz+C3QfIj7T4L6tntN4JeV74lfBZNZJgiw4wZy79B
fTehNG1GJLrr6nMIgdjfVxKqBgU2LcZdOTdo7sFNL9LFAYkzzLQa7pN4vCpOnBEnoqYolxLC3my2
sPbYcUxLhxOzg+qTls+eh18jMgsVGuI7iqJzPbZlV34DLXIA82sYYEbDABFCFJCsv8AeQpnum7T2
KuC+sVzP/I0vMJ3LrHeflM6PAUa12PooUb6mK+Kmr1RT+z8huUXomC1GBmS1W2OLDauFsn8LsbX7
qomkSR2zimWgKcOYD6+EeBWtZ4POIuVwk6BToq6YYn/Tna2c5OH/S+xdVkQGyB0ETyt81n+U1gsG
GiApv5mPgKGpmJ6BYCX4fvxWHhTsUhbc3QdEeyC/0RrlPVy4duRMLECS0I/qa1XdDDkBWWmiqKZS
bn1UD0r+ea/gQeu99oRpdHp4eWQYD8wq/8PD2CoYuk1voxy5mFzItfNUE+mFfJHwAsXO00XOk7fH
dl5+ZouD9Lt2ZhnRvTFYvoaIRNa8Nj5NSnqqubstQ58/EJQjsTJnDIEO111S3PUL/BcwCv1fHqgl
eNzpmRiygomHyjH4vOzLl+i09OPVV68g17qfE8sQmadGZkaS6ZRRWhbxX+4AevFTF6cfFbHm723L
0xMEYLliCUrnMmhlyhKz7bL+Cd3uEWfTBmP1d2QZiORtOPGxCBHUnv4GCUW9tzOkCh24zv7dfKcY
9ceaJCyCOtuCVhPlDcl1zafZkuL2Da7JeKKNrgAhcKl7EmQUBwH0rdmxX2fJ765wjDXUNPFrL8HY
EIdStBWzNmC3kMjVIpX05t1Mv+ieUjkr+rDhhGjULSVbP4n1vdHQD3JSsp0jmOMlEwVxaQ7V437Q
mzdP+8Rwwr+Z6iXVT8jmeBzzKFVon8Z7alGUe0Qvg6UiIhaRFf4QoklTEYEoKrp8OhJFAEjmaeMX
9Cltw+wNd2GVfflKZUgSUb6vTPL1K4CWbPjsiTHvT2aw6RAaXuA6qakJCnrNW1CG1ttf5miPdzEB
FECRz5upaBtvOP4wpsPckSMPHyavLsmPqeKzpVqFhQ0uVwwbY7n3YeuSw3QVNfU8iGmwdDBkLDqU
NDb9yYDN6Yho7vkWxEyqpF+1YXj7tb1P6rui0jB11uK+Uy3qgZCWH/qwbIFjk+Qp4ILqI5fhYJkJ
PvqIRTbXc0cD+HmQRToLsclJlPMACOPB3/IvmeGmDtHjmF021IABxmZN25NCRm6RDUWgfmH25B1D
H/N1YzF47NMuqx2E5rfp5cqADsRY8GSsh30qpp5SJ7PAfRFca2wie7kPE3SLD6c7aQXl4lelE2sD
Lx+KVndUeoW3hbBPT6eulih2ueodCzwS16JWTOlfrMrCuz5uaE2MKxRLhxeJo7gk9Tq6jm2U7PUn
4TDUZZFlJxp4Wl9v/qWVuHsmciKsvkNpJXgxJw/fpfUyFutn6kLkdmKL55lizDa84GP5GsnTO/pE
mw8yIE3u9Tau1KxTgMkXNlGSXYHfEfubqMfcjY0GskUXW1fCoFCkgT+01RhtdtG1FQseVqLKEQv/
li3dMGk9vlifPZLMNqf72pGI/oML+0BOCqy78pWeTzeXnDkEzOXmU0C1pWOrKbHmRM9dkl++4ETS
0dlOnVI621RO+8ym4KeToVeJAZZBsCmGbTQkQflIiFgk0eAwoGSvDc0n/W/WBnBwngLJS3qY8UNI
icWWdRNajnAdwqgdtcnQdfMQ64vSw9N6vUFQHnNS0MJQZgLM8T2jsn8DgYHusU0IWVZN8vrRq2y8
Qh3O4pjnUM74JKHB3gjZLKwt704pCSwmbaBgXi9LmTEZ1VjBAv7ZJvKkBRjqNNp3OVPAl+RSjT9H
/VNv4MMfvt8rYEmkVG8V/p2MomNaxQ4WxYJma3ayXZR4IoUXnDgx4LSMXELbMsgsOU1IxY0vBnqU
eb7SsiWrYZ01O23ubQn5WoBIj2WnSVyWnaIfuJzxQLahHV5S2m5TF1/86xVO6b+CbJRHyRV7iHS3
q2/E1iMZj7dhXh4udu9yZaEuWGRbJQAYWwU2/x2aDc7x2q/4Nzbrkgjp52Vg1wxJWbnVTCPHXAGo
fLSbrF4TPRaRdw+WW9ThfU4sv5RiTtrLtk6LEhUrVT55+ocK1OJiaZ+3hVXPtjZepcbt+agLO+rn
lQjfi0Mg3oOa1EGRDLIvnOMromTTZpSh6FgHeBIchoOsASImficTtaM6FAcZBs/3CLkIzBrmx5NE
8+WF45/LTOxuR72IFUhEzuqWU/XEwIGoANGhUq3+bw/MqApLR+BcUlGjh4HgC2k7Hd1khpcCY3al
2vwZ3VnUbUCTfrh/QthFnQcFjkR7Dkp3puURavoRbKO1GvQfysvzaIJ39V0ZMzvb+iCEEAfpIh2Q
Kdw0NAPZisS/2ovfLc0yYemy+Tdxpk9V5mAL1lvVmj38axlbVqizBHiSPcmE7nHH4eYFKGBcMnfk
X5JFKchNvkEPRgbAi05SqbfPIJ5Ns2hP2rJ7B+PJbPyVBhcxpiP4q7j3enDJcoiP7OnhEp4uTIMB
gt3iD70VwUid5C3gR2jUA+MbboIA3j9HjiN2cJekY4PnoWP1cCtawh/j6Sn2PujSn/CFrLTUNK4v
yCnJOMMYXXt9NtmPLDprOkmCZnPyguRHmqvlCRqlUPAk4A4u1fsZQmYz0k0yt+VHz3qs4K9+CtKm
hY3d3vDPVH54/aG927mZXsQMMtKmQ8vpa5lp5g0qmOzmIX1j1g+aCMrRcmFakO0bwFM5/wGxXY4T
/nxQ3FzJ0SMvKsXVF2u155pV/yLgCZr3oyvrcxb5XJkQO8D7dqvtVwALGqfIMaTd5/CTrWHQ1qiz
NWqCw6ZAJANU4hvgkGKgQnTGq/xRd8Oe/6f+T1VzlZEFcrnofGCdbdI9fatqDHEh2E4/UWII4odW
eJ3xUvYNulHXDn6K+ViRVqjW4X+6xE1ulwM9EIk//Dgm9luO6BQQry5vNix/PtKVlO7JRUp5UfBF
oaOPRxjn2V6aUhETZIkm8TXxV2DSNznOhAcMquEK0s3Gj9NdRbGqUSIIZ0YS1AADgVVB3YMK3GJJ
M5+SL2wpU56rLHpcxcz+JFpkUCkWQGch+NTEJeNJV/ObbbHvKdQUtA1bUNAyMZ+EuKbYBiWcvt49
PCEdZwmKdPVdV6vEbHdv0GGJWzgdbRhNLFjsEr+DsPgtlo1AHKwIxq6gTU6c04tA+Q3fds3bIaDC
gwe4qLXEwDn63cgIXXMlIV4pnDm8x/hEQ/HJtBA8VBPK6g6gtnVtAeJw5ytjOe0bqiwKppKFE/V+
eHt/rqs/eCGs912LCI8HWDCN1A0Vq9Hs8jesOkQsuq88eAYT/Ng6e8UZH1izpEnQXm4TNyPNvxfi
3AwGswJ+RKgR0rGsd11Z22GRuSx6VRWkg5qSs6KS4v4ZWG4RRlEyelmBU4g/UjZ02Etw33FZzic0
wU1uJ/K75tf7UicUC0Ex40eg9EXR51j7aTdYBt++yA6tFA3grG1BdZAs4fcOBgto5sUVYJ/qJSHi
LOlMXnN2nZ1Z2rJYkTf9iP1GW4OmRApaR5U9Z1MOUosn2f4EX361Kmo4Jwvf6FfqyP80SMde2tc3
An3Rq+gzh+AbvdtjmY2hPsH3ORsAVOUm7O90ewoOnTPmVWKWtC1AP6uvT+2uI9g7EIrIegBzfgJE
8cEu1/VZOA1ckvDfjsbwFhCkMRBaqz9lr942UiTClg95U7M5lF4MYe13msYP/9Zw3llNDZLSjQCt
7YEfVDVGrPDYpMrEB25OxdZOeOE9agTsbHCB/VKuzCPimYUjQZoGPfgUz0Nil+9lDgVOmZt7isQS
8mwbpOJV+JCTD3OUZnz5cMl0iBb8RqvnMXFsXXJeKC2/NvwUuxGVQWY2rlWokdxUZerCGqUQxamY
otdP4D6lyVRCgqWSGuE4cNY+9P+DBrqBSOwgq6ciuitOZ6O1FRFB8qfD07QOTQ1DKk/zljUPva2q
6Gaz+H1Qw9KPL6nAAvbK9+53U8gOWUXlsqRcUt2fPilLF/Op9j8TBfFeopPmdaiVhW47e9PKd4+A
QYd87r4AuwZTKXpqUDIuxj+kZ2hzUJitmNBF3ZBqTF2Yr0eSfgEg3ZJM8WtfwAkKu7UhEIxFeXLr
s3n/VX55TSvoWpVkF+Pw3+EryIDmrTYCtv+n4DmYf8bVhUdtCDuot9AoarwUVY7HPKGE2He9q5cr
9+6m8+0yy3NJevavmtBpropYksxFrBXpvJ5B8inoIO4agOTdlhZnoqnU01XGOKTrFI5wqesRPYzQ
DllxYksXMoM4XrEZfEgiceQSbg8KvU5CJ6EHDZ0vush3X1mCl7EMzE4eFwRgIqRp/2z7usGOXbQw
k0Or92JaREt4eCTFYwCoZhkKE9EJqjFbBh15+4Iddeoar3jM46fjobCbJ+FJh3lRsU+5I0djDzck
d/ue6PYtr3JK2w2GYkLHMk5DbparVxdOyJaHv24utDiZoZbOP0I3N5YfBIinxrd1p2s9b9LlOyXD
jFJbhCAx+eYHC3cZRqJZnjEJ1T/bPWRzF0g/tqUh66TnTs2bu+hKgLmqkQsL3D4Lrt5SY6yN4La4
b4V+pFx79ZQd970VQMpQOgILiSzIlqchNWt5VoW7gpNfTzin7gVH6GSBR65bUEVmQGZE/5HCH2kM
2RRqBm59ccJ57bB2babe6uhPzZzxh3y756U272PqeiODvqciVZALMECJbDLyRyPbUD07KZ0HzlmZ
1yZ3W8nGhnbj+CpFlCeUgNhlUOojaJItLJkh4CHkFUDSSTlxUmi/Xju55PoU2YEoyxiC61liS8Bv
JO048cgYKNmJjQQRF+C503qwHPtufiaouePhCnJoNv7nkH2rWyZEIp9olS2I9SrfeFbhIq+yV9uE
Ztq0Uy7r49E04i5BRIp38Ny8WU1DSEugKrJfzH7obHPd68OnEVXFf4rB1M0HOVqQsuwYN5RcEkov
svUGbhHNINLiMJSUoyFFVOpfHvECm6/VOm7KLKOrG3cMziyxirplnX39+dj1SwQxmFUwfcXeplxV
H0BfGyfX2p/Bd8JgdCzlchvKkUGHibnP32txbhye5QJviSy8zaS9hapHOfN0nOdh0LUJAhzfmrcm
MsIeaOCjjr1BOJwCpXqlQt0Ejrvxz0xPbv6oaEFg/pp1EuwOnXG2r0Y9yvF9dW5On7uosmGEfZK8
+QHXowS+GGc0639kfSGW8nT4/UKmpLEDRmsnAslsN2w7gag+7IV+pC/KEQfnah8/Y6X04WKgbqgp
BVhVszdIQvcpfl/gYxmPCxgn1LANOSCMXMNCVH4UvUEzAo06EZEGwc0bQ0XZOjn8fxz1tcMt4SzY
x1prbnO0/1UVI7mcKcvk9nzxTgRstV2xzpyGCLcqlwXtCTR63iRENK4QuFqKvuc3RHyJDyO/9ao2
8sh02L5Mp4NW1/X/C3Z0LyKFAngBZaDtpq4+fOG2fmBeUFcem25xKPSCqA6KZ/6N85m/Jm5Mqduk
2RLtu8m7UWVzlPOBDe6b+YbJxsOK7hNQHj766j5PwE5fsbeKs4xabN0ts8lCwJquJPHxfsMigIEi
SZ9+1msCJXcPMxj2cuGUp94gZ03cG757rOIKY62suyU9h/GfBPRPO4K2Nm4wttoGs5SqPV3u7Sv1
mYfGmEBrETlSDpHeT/ehMDqdjs6j0Ou3f4AHzmnzjWoYM0mknwLIuWkxgNfdDkcm+7kq0xEgq5/H
g+I0x/TmLJfw17/P+YSIR0rq0AzfE7ajZe051ZZabmkS9EnjYZjZz8JWtbNN/kNSmqgmW2g12RIo
EyoDj6ii/hBxlwPv/uV48DM+pN+vtt/D/AUBnXQM9K+QKdhUqQnIKRVTJOCs0oLW+cNOOuba4BZv
ktPNQ9O2xzZE7mpCDx979kzL8BIlUXbXo6SeHD2JiOFzr41qVKme4FiLKZrgU6vCF/Pwnx00Rejy
0YPjqu5co1yM7OFfveNRPeA1xTN4ZhxG6q63SHpTfGa3L6BXP2jcl5Ok4kDQvCKXb8OrxWCeyKa9
uWQLnmO6j6+5mRBb9u62LE5AI52m0FChA9pYiLbPikFamfqSclZ314BBW5FKS1XWevXlF40xlTgm
7KMhist/EFP2mv5XGsv5JeN63mT5EiEFXLWojYVWS7aMzEtNbmUf6Epl6eRIX8mbIYn8/UO2xdHM
+hP3rk+mRWA4HvmjceoeAqP2rGzSlNpra6WCdCAOqKo09HbL8MLYxhXv4GGAtm9QP6Zzp7wiM1Yb
O22dF7KK3+oavTHHVbO1Vz7tXjoP2Id/wsom795KpEameWMjRA53MRDPi1VGkylIi9s9GY2NNwai
qWYmFw0LC3U8PAMSFv9pKOwGcta3qgo9YLiwJmSSlVfNaz+DY/yG5RVR2PwL27WWpg3ZEUFtRM9g
GT1OC7BSdBSzTWrHfJwO0tlblX2aYZvXGdefggkAFVFPGrLeLyqqQDITaY/im1IjsiNRXqWsyl60
YfFoUF6cpocyK6Qofo3l2xYZteZi9wye+GRUANthkSmD30Iw1Z6YPuPzEDoabemKn7c2tZ+Kq/OZ
FgubPvMnCPp+4NXNor02HL446FMG7NR8EkM+8l99UUQOtjEV/4QD09Wumy6KsQlUmSWeEAWLZAGt
UbwkdsnUCR/7QdaarrAJRZnSd+RcDd57CiJi1Xrppoe4C1OTZJBWitMIO7Q33Xun9tMPCi4ta31/
bt8vwLmrmtqt9PPuyTS+oMyThYOPlG36QSWJUOjwIl7M3n3LiJ2F4ojLicKTngKt4FAXSj++TtVe
CyzReTKbvFakxO5dUzzWCs7NJe7i7wlIBOjeXPZIHQTYCvpxldpzJd7Lz7aiA3bG5YLwQXQfGp2M
INs0qQ2uSDem26eUuO49xu9tQg8qHAL4g80aypEiTOzNZrHuRekDiCEgAu6M56RXXQhwRDPxpC95
9Y6NMjDutiLG8bReZjQfl5D2N7JNX/l0r9LaU6n69aLVVbzi0NwGQDnW35FK8pFv54DixjrHiGQY
hFMJlGLcSrURlB8BCQKaaEORAwQdNyGH58aKt9ih3VcAVmSDwcmXRnQtsuDgG1pH2s1w748paAkG
89eVWinftPfgfOOrxYQxNBz65+U1F5Mw6iKZHi+6QA3F3Y5LDHkJDfWqrtsQREpYHFo9+tUPsOho
kicAnlVERBTWg6oM3yHTlDjhZIiKa2S34i8Vfqqtyzwryn3fbsnmTQsTPB5pmyrMT7gcqX8aQ/oY
g6Y8ivljJmYManXYuvLk3EKaFVjA1qNRu5DZpHK6n++8BhiuwP0JLxsCKLMhpBkCDO/4bRsrZc2R
9FlFsH5Rq7ElFMXBQw3WwfOOwbDbNpAtT/VydVCQ93kWkxwQIzIWjYpb28KOvFqbFXuZo9ZNjoTd
KaUS9qHngakNXQ0dERXpAAh3bPPFJzhwWaqfRr2rWxMqVRHEv9v8VbNFuUgBPsSOv9hiqzY2V/JQ
pZ8q18Z4ym3MCW/3u+qCRUXlqdgU80MFi0edhEenDG/MW8Y2nWTfVYpiKO8Hd7Uk8OAHOpCiI9eY
rfWnp6plXfFG4OU9wyOoVmS0FIR6eDPX4+CPYQT3jZz1mTT7uooyjvOKdnRbWAFPPOXYDjBaayiH
ayX3uErNVPCJ1IpWY6m3YFxQoPATePgr4NXLhof9qUJitKTWKApUCgI8u5+A3L14Ce8mktzp9S1j
S47BEe89F9eNKBw2DJfWwKH85n+oQ1IlY5jy6aclorJ2h/6PGYFwqFSLIL933E+qJ2NRqQtxzfxt
I4JG/8j87pAT9pXLL6Sk45v2dFURhwxWGdoQj66FQK87UFdjEeEbPBAvppRiwB/q1Xv4n+zu0y3L
6lyhrEUh/gsQcAm4ve/HIY4pal82og/6LJUMV7xTop7gl9K7DbA/RM7fF15Dt/4aC3r59EIcig9R
jS2zaIHNaUkggqqDtUTVFGyWqEkFL7OL0b132K83yO6Lt7I2ZckZ+XNCka7BuxG3h5nyH4xZwRA3
353KaOGgphtjh/5Ysf0ukQwzR4D9yPH6GDLZ6oVuyOW5TW9qtqU2bflB5zPq7QG1wxzqy0yky1ou
IzbArrnmTERFRB+supvJoUkvRMpUdgt9XCKIMFN5IakEGU5mhDyQ/WwAxD6ccVxxXsYz/SCH5Zd/
uPysVaeSEcoifIJXCnr1YSpfYZ6BQrjm85gLCkrvBl0lWCayXQ5tRi+zGYKpbsh1pVUH2gY1HW4B
4HzsO9L3Rfk57BKf2AqLZ01CuCUd/BCD6ktkGAxyvW4Lod6GBasoH4swJRRBed6uNODAtfUywHBr
HSU4AV4PU8fJQRI1W1fuFR+qLNrEBiIRJc6HIYtsf1VB8FpsQCwlYFMr9eQFHWecRZX0IJSgwUgV
r4H0QOfuYjqqBNPn70oT1YjmV6vhDasZ011YItzXyHhv9/4WGtDTi6sRFrTiJZuoRReQgbaJXRqW
pluDYwjBhWHzlnEbAF1Lb4CXnLB1ZTHx5MY6P0KJ0VvbF+YwchU2/YWO2XfrnTq9/djcvn8tLB06
OU+Ua1mVgPy+g8k7VuYyAH6IQ5A8/oRmEgqrznlMEjkSBeg034FZevasK6stVledgvga8AdoIe1Q
DDeFy05ygjksnMojwFGUpUA/FipDER+6D0mQezqk9lIVaPZmd9jgDJBYHDpEhAzGd7Om9XtkGLTc
NTNIciYI7iZnEYeE2yDzIelO1te0H27zC1SqGd1YHKINcvusIdkFHD3iOO6Rw5bGHtkZjZY/GFYx
pO/764fPwFR+rWt3m41lgyNpWs81rwffV1TXf/vjsWdz/XjNgMScEWuOpB5rhmAqhSD/rc63yqq8
FdSoir8b0ZhhJsFnI6w9VtgrEORZwYYVEMZWccnfcwZx0kW+cZIGO41ACctKsFuXYh/NE8WYAoXD
zeFqn35p/7GAxw9Hi7Pr1iqA2FCxQtFPDPNy2qwVylP3MblMr3gasfPbcUPZIgucjRLTj88mCI2x
UW1ktbiIWLxlCXs7K2qhsZPdhWtFczxmQgWcOc6tnBq1sKpkSxRKAUSErkat+9AckCMrw8RzzMfE
PXCDeuDQavib4kh520tmn6uspGrJjgsX/71QmG/5qHPuhaoH4Zr//ciBUalj4zSS5HTA9WSxgWqc
fM1hVYImAuVaJqjklISo0UsRtkSXBsCMf52e+c2w0alr4a9UDBtWwegZSNj3Pdbk0B+UZFc2dfvI
hSFuIbRvIjeQ7zNJw1HgTAJ6aI9rysPL1qAdc8HGsCzvCOYnOIFjbIbHPgZOvmlLNys01V2f3sGz
RiNZCypcyrCONb3DAhF/V+MBeTewJfupm9E/3GsWfyPE5ShOQKPP9xqkaHZG5fTyknNEZX+H5sJW
W/9RTCuIzYyzv0K2PGN8zu7rqeOPda8Xk7/lvbntstVMgbz6N6xkKo2Myulo3yP0DZ1qU01/H5or
BUsYzsIM0Y9pMdO8ddn472vlkS0Zn+q34o/mE5oKMovcSwsYFbOirKSH1Nhum4kDFPPgqjuRqpqm
W7qM8EQPVSCVdClzY8Nai7n7Kyxt21ZVI8yHuiMukY1IKqGOO3bZ126bBy/cOmT9i/wgazx7hFXX
16kOXPoccTwdHplcXrSUJVflxaYf6lJhqTqIZFyIZLKBZkQISsOBmVHRTkqLold5AQDVPiwdGuoe
vbJ9RUTKJ2spnnRFuAD/Gijn4AjB/eY8MBdt+4blQQH1lKHE7BhNknTrpVNnQwwnwnmxRzbUkqXz
MAkGJJdljQDOx4bj+Nz7DL/oimxN4n4MBouRDw83+v4l9nL/dMblSclz5AufR5Y25dbh0IovpBO7
N3HE7WZkCAQiLX4/WFnI88vMkORzpSXPskjSshI7gIrBP02+Pbx3m5aUTPgGGzGOSsXptY7ChEws
0CFjtCKvS8kqNKgry3sjR9kV++L6GVTFdkPMZ3sdZ5Q7tzHBfuv+E0J6mZGThnraalFcOpvo+L3O
Vg88WbW4PSfJ2m/i9Rpbg9TUp8mEhrSPSrm8oZGtTdwuqI1nNTn+rxembuuMeB0oKhXpU0f1ORyJ
ci1VlVhUN+E+6b1MfynAZ2nH24r/GH6DivqYlE/1qGnYgbiUEarVGsUulAPyIwKt1PyAD1D5dZsN
RpTL6XxuOl9w/iQVTn3b/f+VYQa4ecJaHWTuEhohZ/mlM6jtKmNxeBfuvtxmgi2N4CRaDSWBJWys
UWWmZivKQJVRtWTnvBdrbcI+Np5cUmtfapYtZWnZRJmsTwY2BB3nmMuisrggBfpumLsV+G9ZkdBK
BCVCC3FjzHBE4gIaC2rg2iOMLmSx3QPaVNeHdaNe2NpxZhNj0j2DBWOpEYCjAXQzyi0AYXoFI/J2
SzJ2sfmVyvPnd/mJD0rbaiYgrNQVwCu/qGrq73pdSmN6RQXEE8owXRbe0h1FhDQlzQMQOCeMcKOz
16XlLHmCiaP0BisDQKpiAzNmTFjHF6vyXh/bgx1peN6dWTPvh/P462HPYW+7+gHGBGbwwj9/J45Y
cOTNS3WEw6N1N4O0olqCfJA1Miq5xueiubBrB5dE1k0iU1ayEkVvpg71p4AsNwQPYbpM+Qk2fw3Q
aJvSCGE8iADc4P1ZIFq0Ht8FeuD080qoLP0vbCQnZzIn36PK+oFzIcKTSu1hZutwuAG/X7uAq+31
t2GsvXZvmn5m/AQzmua/9d26RZFLmvaAFzZRBv7pCzg0Juv28vQdJINOPY2nwEu91d0yMYXya28s
ztEsyCYpVnJism7nPr66n4WXr3+7S2MS4fpGL6b6wVRwFf1L9qBIFA/gAJk7S0ml978NbJUYED1t
stz9HPnpQQ8T55diwU6SnnrCEe5KiqBpNswsUkuZ1ZNqgSaZmZF43WX0S8sziOfjjeTivCyBVf6u
ElXIJsKr5ZFJoUiVOYO+bzZQt8JGJd0fHZpouf9TBqr1CVaKwJU6CRElvLrSY3CO8TMlIkcJmTLF
ZVeJSZs9d5IhvkoL7DouTAB+0BlCe+4mCKHK0YZ/pS41x+dGjfRIs9D/LapgiXxPE+nMqHsZC4GM
H6LSSFOLyIRIW+m1PjlwtBYSYBTGpiCEL9RISEtx7vgZnmnYNlBddIYH+pjpBQopW4WOXayBeP7v
yVsr69pz5OUYlLqBlZdgDNCxGgUBf9fv6+K2n6UP52cnXKB9d2RPj2FQqvnGsNoOj6vLVjmdhNCs
Tr0UhadvnlCZuaPxdmlL2Fn9hciWtAs8lfgtzQC7qhXCoXDpUtBX4KT7axPt2MbIcHglGc7XBW/K
QlhJA0BoFeoolP0TCJKUKltsHzAk3iWv2B2r5Bzo5zTkR1sYcBZbXS11UCmP0cjMKNp0AHpjslUs
fiITj3Cyg+IKYWhmqwaCDgG4NnTbWu+Fa9Afb4DvCkI2rr0ODoSpMknwq7RPmE7I833cSzdAOS2t
uoIB+LrhWZcG8d4W7++p2/p8KpZr5r6mi5DgKM+I/wd3bKIOm412Coyp4WdL1W7MEzWZ+A0EeLWF
L5aAKuPphhTBzDWCxfulDK9WaZG0SlLMBqI6fRmHVFj8moSw1O7FcuEJxMgEd2uDonpO9Oqkx2nb
zLi77y/Vg6ZeqepyBsP1ifTXORal2rsnJzcxa2nEW+f8eFKR4D1tya+ulPeCRfMXJnPAA01g7FiQ
4tN9+otHmVEh0Ab7ZFZ+LGzu/0Zl0K4MYR9moQ6yK7mY7HqYN6yoqjPoDip/0os+ylNzIpI16zN0
wK9R3X3kzVB9FMjVICN9m/XCSwyJGvrvxZ8y0Mg+QqSC3VnX+Z61oz3w8r7J8cu+H5SQfoBtcv+z
bsevfIQ+ByJum6NAynd8Fvzy664mytNvm+0NU3mGc1US0cVmENV4mHB5VlLY0LdJb2lQdbqbnKyb
amQBTyirTfunbZ4Gw12P1SjzgrAW4GMc2Gggmlsly37KB0AltSGdwJaPSkhmuprIa3zpTEwt07YF
oQ22wwHLPzU1Ua/FIOV0StjbvkRHD4+C8nbnLeZAGNJio1vCAFkOuQqUj06t0QpaD9ZI7tk8/QYG
D2BGZQg507U1XeDSRgV7As4LuHMV9c0VAVALj8hSeXY8rR2ObEUZG9h3tRsGieUoc29wdliNoz13
57CV7m0GeZGjjjW9MCdH8eTx7tIGkEIjrTwdIp87C3dbfiGypu/MSTdPXt8yGwQRuZUydpVhpqgq
xqe11olotFaygDq+ArlpUZSPJLslPtydDYvqnveZi1VROtP6y7GhuX/3BSvhC9MWFHuZOw74jQ3b
j/ANgfyzUF3xU8XDZzhVIBrkwVJo8UokzHQOoFWv7j8PUNNGIBZVfiHJdNk2fCI03ruPJkLBiehK
QRYQ53oVTgg9G9JyKm0Fa9o8xuKJ+oFZjD+1ed/3hG7jlTcwu46IPg7sMQoLRXBSzLF1ipXhNQ1A
vqgbFj6rkqxfvZdOBt+BlAADrehrPWFDR5BNmwu3iuNX7HmQVClAY2y0+gTxoRwZbJq/KoWFS4Tv
5PjlrwUlwRTbPEz/bVKdXuov1ck/ZUGyHOfYeg8FIKAEtICF02Tyooopo7DZZuonawhb6m73xlO8
hkNrvsZvaHCdNz/xzC+CSHSmAWsnepdWpawINiwBSDL/mnJ78q2lPWsU1gUDAVnoIgY9CGHQ6adZ
g+G+aZkhJpmRdgERkIPxt8uPcZ2rd+V7VHfY00GBNTW+g9Y9hTSu9V2dp/23ojeepXauL6svnReP
uMwI5SujsGgybBke2wsg8UG15M1ybY//tmAOTF3UQlCKGrJshWxe1oPUpNlDOjoK8oOLleIUKTeS
U9rdN24j5Jbw5eVOH7XbbZetuFRucifjX+11aJeK0scxGseuTg+Hi0bxt0QDqghJWET6LORWFBzP
40Iv69Gz2+H1VUnvgCx5OHumBd8KQ/952hJVsK7YD4UOxQuYi1btAEcvn8LhADsv4RIspRLcAuLD
1Vm2iewPbGL80CybHwWA74XJjLZoAPvhUo4ZH3u74HDnXj/JhXS0KbQSM3IEdD2Aqwg8F6Rat3X2
0bAFw1sO+PAk/dgO+RM2uciI8ufHsOwhJdsCKZ8eueYFFZLm89p5NsaAK5i2FHjaEUhetxgbx8hH
PD4xOI+8Q/gBCjqgfcQVzkyoFjCLbLR0pkWNjO4OJyTSXPxWvfvi3UmfBVwiHco5YCoG+HRq2MgG
AyQkCogL3+ztk0Jp0eWdjmBnKfX2WnQRyGT1DhPFwSOXvfYVnACzINcOVvfunWh6NlLNp98m3FLy
ddOhmdkaHGcEX0O6LaaKOjHo/+i9I/lXDqvRgawWv+oYXstmVJj5TuXF03xtVSyvs1cS587LIy07
GqlfPtKvDkUwQMLIbrUYtNncrUva/9wTiE6a9KOhTgX65E9z4BsbCycTG/gjdln80PZTXpfgbbaC
yx7nuU4b7Ffp1rkDl9x3tv+0w5neAJ7UeUzjSe5kJrjpXjXtGhbJ5BxTEVy0mce1zrJXOC7p2LGH
3Ci7p2+tpEheXF7fXrdZqmuDLqMw5pETWgiWl4y6UBIR2xdxUNLlr+1j+A1UIH725XpgkIvQ4hOC
sy80xQ24/yPdx1MU3ae7SxnCPM0DeXlm6tx3fa3rOPH0Ef5dOLXUbMmD5dLDm1p3frRfJ/P7Hy/8
ijG5AkrFE6lnIXC2EOrjYL8y2TuyNnMs8tOmkKz7XxG2tGG6WUkl4dqL+GEfGJ09RbANIBGk8YAU
hESv82Dhp8mpsJxUWxpFiTdHFCb3NjB0mnwkyOKPYKi13PFKbOiRfR589XbEub2ouyhVn6ScKcrz
tq0ZRQTUB64YFOxTI6KXdr8LxQ51RRliBG8Trj/ytDZ/LnZCoV+GlBD8fqEd//2mZBW349q6BOk+
wF61Zxc4lu4jg8olcmYj8f1pXUrOFeUCuUH6yOMKKkBfLGE4ix7FsC71fskRwDzTkEzQpOuGDcFI
UMdQdUqu0wdWRapTL4LK0lqKZHQmPpjVJOr9iswuQ1k9F2UyBK1X13WFatpYdBrL8ktmgA0p8uA+
hbqTpHXz19FBxO9LyWi00aw66wrseh0ltb2X0qhhwkAi1WVteaGn8Fjdf3vFVokapeOBp1oGbWUT
vdgA78Qd161ThH3zgWC2vS4Vs06jKqGjXbGKrDQNcJbBhL9WyP67YP2AIY2aliIww3/PgZxROV5A
BNdLSU2j5w9hmRdOnfrT+axIb1++YWWc4LbltEpZ6lQea9avY6yyEDBZppxne9QnShpfA9uAOIJH
Vf9rSqdMd60NtUkkOFaHkY5v9e5cPfR3MffBgmmRgh1q0bDZR/uexPATpepkoiPHSkgumOCp/ZMU
WQKeaUsxlfIqpFd5m9j1LCelsiBBp34VrjI9TjTAHywMFIM9zYhjue+HEUHt2372/h3EYsRmQA7B
lgVYs6vZMllnHofY2/neXSYGhiw2hfbPfkrD4eF2dsEYbiQz5ofIxuDYYSsbzO4sHsoKSHzjymeu
mQO1z/P5pSw0sdTGJqpQChtVPOzPLhb37KfWx7zTyVzexhFMjGJxrMepJXL/FyLmzN2Xws4zqfZw
ZaiwBfTdnquWsMJbMDuQy8ZRJQEmu9pQq5fS3CyaC/zkZV9ySGGkW+gMayWBbH8JtcYdIDiDk53U
J8xQhQtrFeCZXNOVHKANmz0F5O/sMI3bjb6bm9f+07cACBswwkv3FJDhZ2i+SKBkP6r6+fIwQthq
tUXhhGUBo5HjIRbH8aaGr968zqqP4sWYWJ7K8DlU00ZvWIf33AIac6hC19pnMLaw28fW4VudoMyt
h6k+d/+6ofwFsQJA5Rm8ymJ/q2hujYf9fDZU9ga3T/SBb2FDZNZh7R0jLqLcPJv3q8nGD+Ifa97z
6H4ddcPFcSeGPFkZMekRXhf68CN5FNdPU3/ZC6B3WVjaq3XFbjOwCKoIqrtVAJxm8Ffn8rvKqNuw
346ikSLC/MvvKwXPc8QXONKf9I61ADoabP+vMtE41+CnvyJ0h5oxHWErN12VXP4wKjKiNfw44Owx
zZRUn1VI9RXQN+etz+JseW4in5KYzynlmt+YIC4azF2MOJMUCwYIfXqkpckEaO5+RonKZjA6Fasp
pVbW3JkxyHqJ8VaQfaFpWO0Nl13vEz54o8IEU+AW2E8+WG2p5YuXI7QeQNWJSjftUCf2otByTGsh
jjO8rC5EsDhYlJ4RKE8UHAbiXWzXrUAgUzeq69R2c/XoVhPxRR7nScU+9qf8Tky3Z0G8YrAYpH4D
xK1yNtpCUnpECDL4iFoEL0kjoscTMfXpQlB5weALOlPoSnC8Dgh/Szx0MYxdML7JfjdK91ouA3pi
bJcIff1FCMtVjKo9a3HuHpjFIQIS3RnifXclDOQf2ZDXdl9UizhKzG2g70nDPyUm2p9VpuekZ2B5
Af0dmhSks+bYHL1aYHjy6KjQSFWPBObYIIVMdRYymqkE1+sa6+56B0K4waDWbKUTNSGs01T+xNg+
Aq652ts6SrJuQHWGmr8GqUaBiXshSQjFo+FTF5hwVZ0a+sX3GtrxgZEmuLk8wZzQ7/F+o6UYKQ2c
fFp6dJIN3Qp8UlZ7aJ/pc7Tc4q7bb83Tm7+WlufzYZGt5mTc6TeQqqz3+vLcHaBleyQVVr34e/jC
8OxTeJtImLYgKCGagQjIePj02UP2DPjIIaIy1xCcvy4T8b9+67ky6nHiQxPTxeRk+CfLT43hUbTs
07sCiE9QqpTm/L7O3lCIeHilrj8MVouA4IhPB6rz21qQHr1zTJFz3vcTHiO/N8Bwhk/cDkD9GvBP
Eoy23f7Qiab0+fmY/6EeIh9W1YFLki2xI9gD6VynX6t1r+Goe/IHRDOqRwhtmiteYzk8AAWZcvBO
jPeamz0s1S/FaKyB5d5ujM58f7hi83gUPGx35UURmBHkBvX6AVvU+deIFEKffbVFqey0SnBEFA9g
Wdx9d1o6S0jTSWu3b4ed1Q1UNDGywLO059xKNHNcPvEGGft1nyeSU/F9G+vtIq9nDFTZ39wwW/va
pnOlqNmVV8aCUzQo41a3JVb8ST96JDJNKSHvx1CmS/4p3udxoYcHqV1/Xc3yJX4jE+/ddznAxaOE
CpiM347Dv8y6PxXcHWw5oOCJL7CDf1+FNHXQhUlkn9tsMgVo7TJKtO1CeZ2Dy8ZOS2BEWFQ+wsuZ
ArDgf24N1BMYuj9z1InFnuIhpMYFSaMFO3h9VRr6nayWskt+MwXwWc2vLi8bCVsHh0mnUdZArKv5
WSin5j3Ckj3ViCOpnxlzByYsSROqJMB/GSM0Ryt4qVjQed3SOmWabd6gbZFCR/3hIqNOSlTHYJsp
bUbWYZTHc7vrYm+iehL9rpVafoUhr0+OGk8wpOO9S9xsBcPv4crdcS62tHd+uC8DZuLZ3ZyWk938
4JRbb8ZjfkSrGg+qPE13xFhgDIg+tC1AVULDLq+tV++pJ19QtRbz3yxgLgsiCLdTkiFo7NY3jtpO
sJZphGa2PZCU8CWCHY6U/Vh2MpehAhsh9qfRqooRj29o6MEYN+9nXjKXRxXHl99/wjphutXEtElS
k3EoEuV0dvcGywnTTjG4CsEo0iR2BVR6S0ATTuZjzdDwmpm/EPhlGttFg9KRmt4bsQnWQOOZuXeK
3RPipprY1Ijg8uYZ6fMAOLxZlPN3h/E2zujYeSx81r4+nLShu9nvf8egXeDQx1E9mw0BI89TjIfq
6/YXfUv023SmgnEeBZHs3kbi+M0AlilXC8+nvjS2tZN5a4UAVm9x1T5h7X/IpZsDLTrMjHRLYOus
K6rUZ7uAct0bn0r0YjYqHIljhH2+1Dl7cj+RBjm8gnM2uXgLpUCiZwkHjU/Kd9G7WH2qypfWKISv
I5VRCIL0DUsOxPcSCMSRlJ7GZHPrupoRnzNr9hevrKGmXqFndD3pZD7HzMDxYl21ZOYtIQJY5LXA
Ij78wiJd1X8Cfl/0IaDTu7Pb/+qXKiza2/bfKIjkH12AT6a3wzijDFLefn49X1vnbUYcekcb+CRz
2Y6AAjsJIpc6RhYDq+jzUf90lXkkS1PDBuFFuEA8sHqvx0RkqiJECi4G7UyacTUAm8B7+kE+L0Op
Ekh+yO+ERB52TTolwGp6WTbkEJLH6HhPxPt7w6z+eDdQ/qU6fAHMivqPZcygRJGkRE+ELh5cLr6j
qcpOpNTyTwUxQ5b7uT2iXd4j0jvF9RDnMa1ljiSApM/OTB6bTe4f31Hev1MLY/sIWj/3gjghm7SA
WSpdZTz5i2L7gNRDGMTdvRtnSbcRVcYO3lmDekI1XoWZ8KPALyx90KXgszltojZEQczHGbu0G0ws
bNVrZPmGl2KHsW0G/snKDqpA2XJCrqKtuICov4vvDmDa4Q0LM/ovCc3/FyQshDJHXzuEqz2tV6nq
GlwKf9q5god60KOLpqCWO9JEvqKk8+y0UxtP1vnf9qaj3tslCFZKO9OOgU8s1l/Ws5/r4W84ojs9
TI6H+f3Dlzh6J88+quts/mgTXu9pK4K/AqwU8nTVa904wCKsmEb9iBXLyMPT0YgVfDBMw4UYnRnk
9tWp0GVub55Q4Qv9Apw+8sfhkKLsvcSHhj/FjQaek42A/8oRygGHitAfX6sXMy/4UEPLc2FnYnb+
dFLZLnguOPANtF3lxZCawZi46Pg7eDKUN3v/xzhwWwXIBfzQK2S2IJMUrJtM4G6fHDIUgaO3sFka
yyAJanW0QqCOCXLouGlVxc2egDVmal9i5609VNiWNt8lbL2xcK0EAmaz3pJQwN8FZAPZvQKuCCgB
1QP3qeogmIVOfIERQQ8j7DVO9LFaP0lIdq2Fs7fme3UoRHqFJBNgbzO43DNEUYc2hzzSE7rTDzsL
SLxcplfyRr/QL99rh92ah0bg7x3YNWlp873sy7AggqdVNGYNruX0DCtxm2sjlWv1LiX45yM8Y7Jo
nVY6d7Q3lPP2Zp3lWxE30iEgdryuThm76vlduk41yN+aluxSdptBygzO4SRaSEed/A5BgR2ofMGz
4gWg36+OjP+e+WMlBGl/CSuvoXn4eGZ17b8QPi2w9tKilCWKuTMehCGFEUyfxJD0GJBgdOerovgE
coOpDLLOZsjrKQu3HF6tma1/PqTfp1oKrZjCXJHJLeJFfSDJxsPlUILYaQ3obiTB0XMC9FoQGTwE
p+69VzxVgVVazbST3iY5TwF9VTuGAPw9oIXaJlhxuc7V+5L4J9dqVbL8nqFINh13clPEIZc2moyW
3sKgQILiDa2xEhv5P1l4gwM1GAVmRhLDBl7isd56hW3bx6ZDscFePhbovb4a5rzo3zrxfqpRaPzB
UGtzNlxqVCs63HE+ZmVL55lyleTxrX+fgdz/fx/BNlYOvAcLdslFMPk7gm4rlAm2jQvI0jynn3kW
FD8jdFDnsH+w2t7ARKH2L45U41WyurfcXP19lydHFrdw67xZwm+1cClOINfNEY7jeNWPYLHorpoQ
AqmnQqwNCjzKUBs/71i7ej2GPtpUbsgFB78O652pxyAw0VnDkljxqDrVKUDiqOcLMpxfnfcApAo/
KMJEsrL4PYg81sGr8IF2aF7Y2fpX/MWCgF/0UqJh6yfGHiR1KUEL+oAmknqJG0nB2r7l8XLeSDtc
5sDu8PB+rGenp+XHYWPeE9dYHnlYLPedmBgLWoVOtlGWgKhuftAyrR+DZtVdnWVHKZC/4hovNHSc
TOWZGBk1/1p8lS/K5qjyEVN58tl2n6LYLB0kKChmf6m8LioTzjsdC7eVRRmEumHf9jGIOlehKWzB
rBthD7N6rrxSTAixy1XTQZRfDBVU4/FqbC6INhuGdncTl71sI1z1Ub60WvmyhdGc+JEcdyDZVteZ
Lz0lkN2HB1pHpQxCMELQG5x7U7st7Exh7jFwlMLRcLySqA+GXVR3edlCyl3kqOHg589Y/h5m0Vbj
f2QFMzfajlkMAC+HT3T84j82/UpgmgVgLWhYsLZNkfPTdimXwKzbKuvu6IAAmpf1cJXyovr5DAV7
jFbJ528MjwmdDUQy6thOrgnDBnvcyLAQFEnfheZSeF7lg9AFiKwzfPbGdHg0eIsdm8PT/zWLzZQG
kmrjKkSsC5Qw5AchyEBURCJWGpSHhp5HEqRWIWzPvu9+N3YnGskGXLdPfBQopToXFYvy/3u2fhJJ
zrhOkH2Vdmc1Ikavb9pDlYYsTGzmXCo5JJyY1VihglVz533zbNnQTePI0OjAwQc9VdMTQHNOwuS5
Qf71fsaKvfHWOAvu/beZHama2cQU+Dn1p/fEHasELanXHQCbaJX9tgr9nVmj+tdBZtLsA42q1Xnb
J59s1mg+T8eKainK6kcKg70HTdrrXjhNnys4IN9hSuak1cQSAqIYfhof15x6JbkIYjLFNAUAG1JZ
bZLp/7MhSLe+gh8C0xBsjRXoUDN5E/ZMP0eEPvHAhgpKMSpsQzzmUN3i/sWEfGXjBc9RRsO3GMBY
wET0r0WSOUGDhvh3MNuAy4ln186hQrLn4Ue06EFJyhmahGBqXFnAU0Jh6DHuwB7veYBCf39kuC+Q
kn3FzZ/eDRgeePLRsLExCJM13KgFV5Mz3/wqt17W4UEqLQK0MNOJ2tzvsHEZDIVR6ablmpxLBJVZ
udAkjjbcQf8FRZEKwZ9YMdeNVgjLaVeKJbFPdX+X5NORQBB6u/4fcMNdoBz5QaVLaIkIivrDWblA
5TurBhWJikRFecPA2X0Xgdsb4n8VpXCcwJkkXH5jvCgBYI9M6Gorxt8xWbrnqyGz04Sbi5+EPSXp
kpVWbIKr1RbhFoGJ0TL0KJWsGYFq86k9aG4v9Hi4lBnFtHODuAwnBrRBCh/LUsJe4xB45jFxQy9r
PF2EnHRqvWjwQZaVVWhEAbEYpWZRX/WVY4W6GDS5mrKfS3CStuIKQMUOX/rZ4vbb+ZIT4y59n9Pc
oY/8no4YBSWwUSxCQKu5v0Gp6VJgbOnf4KxjXBba/P0o4dVk1AcNWerhphpomAVK249tSwIlMaC0
V/FIN+7YN9Znent0cMif3wR6SW82UYzXJJPFmW+QISpgNoF11qgnUat9y9xWglmejEODFwkioq7l
laWiiKJupm9oeN885wQHFLeMXCgpGC063CDOoTZq5o3mXQazoi/ttR0tzebODXA9hsjpocyR3OhR
6h80W/6x+ZcWtP61S+cUGr2T6J9Zr5tJmwNmlMMlKSpoYYh8oLzvmD9VahOtmwnxbfVpOJEPNpCM
S99WVWD9lvMwGV/ei4mr3zp8xiNgti4QCPAN0z7Ss7NRKIE+NAYBJZjp1GJApwT8kcaPbgjrPwRX
uGPYTFKY4Z5a7ijsUsKxHzwDVRlr00vzQtsaWpuqNov3gHCMMaaF9+JasFIY9r9a1qJVH8wwYE7Q
mav4KMjmwOhGnWQnyrkiqbyA3Pns99++5aoqV7JikWy85bz0inVO0lMsBTtoT1zIcOZu6H6DO0BG
NPpi8rIdzbg2cbARy3Jt85scAV0x/B879g/TpECLPDBPk9sfssT3EtAX7cwHAYWy7QtCmEs2J/sb
AvmIoQfFFytKlFOS+YxCK0ZG4IqwZa4QFfNe6uMYWV9Dsu79d+XyqDrLorCUj1ua1dDYgkjj85Nz
i8Qq87Gsx9yiE0LjOiTd8qu6jTC2DNqnPDZXxd5AIgO0TVL6QWZB2iOnc26PcCTJeZHOz0TEhQbq
0+fsha8VUvwKUwJc1z8UGPOXI+9MbDtHJhvLn1cnjVD1JpGHbIAs/yH11pyLG8BHrwPj4A/UaELQ
OJemHIsY2uG13R/J9mzL+A6rfUTusj9eGGfGSInvaf9gXDCkrwtXN/N9VPALil1G9dIHnBmwGRZS
7mRaSJYDQDAT58fneoBwwEOIUW+FgfYOI9cBDR5/PmDkciPEm3WlVXCjm+pKhP+f+H1oe2Rkq/X4
+q4yFH2scS+6G7ZYlpoIMZxR6HY8blB4ikKXAVOh5Ri7tkWaSlBoYaJm1Cf/zUsVErs1NcnUn6+v
xTBRR5Mv7bFKKy3yI0bB8ZHp/1czmUYVfwXU1NAXh9qdlCzAfGNRcoSly65xLRm7Ou3103EutlSc
ajk1Cn9t25Veg3h2vHlz+5fieBhb7Vmhm1dyBjJZvIfyhxUJ3/+WgG9ghONbI6pxxKzUdWdsKziF
eUy2WUhxnS6jtMcNg4T2209Oe2fd5VJfnxVQpdqwvwAvx6bm2ApmdGWIKj/ph9TvzjqgNJyH2YJo
yAeUMkx0dc9OU3yx6sikOX3kHhJB71OQ9OQzn6kgTxfvVuchc4p1C9P9ESeiFqsQLDPUOcYG2Ynv
hxUje/cEb4lMFXKNE+WxAyAYt4wWIN2qQM+W0pwtUcrzwBQlUps7rlu+Okl9xgyQzXW8JZnKWRp6
FzDUlU1xVSIbuSqXgocgknCzlwfiE9WhslS2iOSBz8TKInTFxxFd/TulEuhLZ7YVz/NiovW09kO4
qji/+LA3YxZf498xgztZo5+yoaQ9JFX/fc2Wz3HDuM5dZiQz3rsoLLDfDkWLhTU/v7vzh6J+4qdy
hd4pHtxl0pcBhYM9gpyVPCmrCGWZNhanNCe2F3GV7jF/YX3xj0YZdu323DIk598faRKYKBAuU36P
PcEtIY2/cKVtjjHhob8mmWAtIqMyR6tHhmY2lvcWYyZpmhS+DfMbtc4MqytZPQU2ZEqs18WeMuu4
8cDgnavZdmrx5aHrE9qg5tlZsZ7dHFY+NwuhNrux5ZKas9n3WCuseEu77TDDo34XPKs6gRsz3635
pmB3++mRzYG2onp0hR72wuRfIfgxB3F+yics3T8jaUWEsVjQ8nSK+qiQj7zKNt9SgYQF8894QqoX
jUG+nyUux6RBQD1IV+cRhtnrJIQ4YqXSJjNmDVl4mPHMQHGCNQ1WYoYDNMLJz32kljTm4ADChJ1n
JtRBPTrqw//W0NZuWx2bczyDJkbH9unaFxKYPtdjtGz4w/Zjs4fGEY4xrnml308hdta8ecoUtr3P
GwGDnDdcj/kVSrwHiDLm7CK61543sglPgv8aWPuHoKP/vY+IZKL73A+VrIFzumkzahkzX+mSwqqe
GW47vWl4Z/TBt7fWaLUNhsFSxyAtaRA2MegW2TQk4x2+1Z4+NNzBS2KZGT/YL6X+PHT1RptitLdu
2toi/8pm6+SXSBUT3nwEJ9SET+vA9Aww+jKvLlXae0gVhxwfmfnAh7qJUOeub121fgZevHOLe5QF
knaZ9xvhXZUD/7eT3zKXxcFQxpy67fNEKsGgGAvhYsOjnf46v8+Rnb+q45c6hmFnAdidxpnuGt0a
UegvfvPbP1lA60hJZ40PO3Ne7KMMkXPKZnk5MTFJZVXkFLPWGNzWut9qhArzwqC26F9X1fZKHnxI
0FnKzmqe4oy/fOTo9IllfiGAIrB/HOUcAGHtOB+9xF5FeuV5fJ0vChxZGfZqyoOc5vueHJ8JN2Dm
xqa2/V7IIHnXeEIZgPH0D+ALVeGlLnXdruUix9T60O7VeJLJoAehGnT11tpx8+DDrUvE8UgiByrC
Wbu2ArEeurQdlINVcNvYWPZfR//TUaHUnjkX+bAoqiF3ES8NGJlseFNrb7AnGTlaro1DaNqThdq1
AaawWk3j5hVMRzITRPcEjvnRehO2i+3Oh9XWaa98I/ofeIOflsP04ya0KzhqLEm/VV8dIFJoxJjf
FsnI5ikiGhuHh5CGKjz0u85wRrL43C8q4u6GF1NXu+jeDPq/HITXCF3DubnKIw9/vImV6kkJKAGi
QWXPSnsiARMpB/WLUimji9c4fMutOGzd3ImW/B/ucOlOiKbR0Woo00jhTWE9ZOq3FQsAQBoXl3JS
dQ9PD4JzN8db/nHJagnXvjke5lK095z+ys8qbg5JjAHVAPgCHJfA8kwfuiqElUo5jVIgGmKg6Klc
Z4E5fJ7SF2SkHiVzHlFzBp9wTjV7hYry+SlmXFM6mz4nj8G9IO+dU2Q2g1NIsQNVFtwl4HS/a/iH
bLzs6L4Y/lGZq3AyAFttbRiZvVwbNe199SbfDJ/u6oqDjpQrpQR7y136tuKyVZpDUT0Yf0Xath7N
cfbCx5/e/eLfQeQcWD1/CgFAZw3baBCo3mM3nFBrm0AxBrnk7KUeV8Mff3blKLDAOVam/IJ5wW1V
wXcBm8WB8pX003BpI36kyl7xhbg8nAgYpIKhIvHDcKbJcrHmyy20qQbrulTzStSFNffSIp1mDMkG
1UqzmUepR56hQtBdzIO1uHQM4rvtMwo9e8T5n4/2NMueZIATna4QqaWykczfpoWe0BAF4WJ1d0iH
Mcj0Z+JpEw9ZbDvfO5MJD3q3Vz3xshXooNZVv4Ld7x2aM2WtDLgXI5RA6py3kP1A+HdKpLUT7BfK
LpOlNYzlU2bP37nlXW5VD1XYrGan3jnSz2bI4Ugk7GwjJ9UjhlY5chqCQfnAyj5+0JuiIy6mEli4
41B2LYtqWnmY7YPWcAkioR+024ae9lEn7RufDV/6mvsz4M+Y5Qq7qCEeAIqT0hk/ud+0UcOYGmcl
txNpmB3NgwjPcuvXKfuQ9DbDZ+5fQdDJLZ+dmr3l9Khpb5dH0TEafrKazD9cmGaekDfDZPPW2yi5
b4JoWAiYnFWxmOfCt0Nj4NqwRSZqeeGhVt/Ih9YB4wCNDXld3XKihpr3qdBjbznx9BRLisi0rcpX
JULvslCCUbx8zSJfKbmr91I7AD7TyDakjdfVpAhsk7wh3SJmytAw9IVQW9+KnjYSzTVWbaBYUlaT
L2IVEH+bNjhmAeH5tWihTRkTuD8IqhULAgIFY15e9kj8dwczybYL33rlDj1Dje+uNaXbWiKLC7XS
T2hG3qdad60q6YBjJFUrtxlcEXc/AOaduJCrBFfXos7cMYYd+LI9IwH0RMX5k6XWtFaeGNAwGn4K
s9omBlzZH2tzNujGGVEhlqtLtmx9//SkuyAGRoMbvtXG6V8fbJWm2jZRBx1XDiomTDznOO4IFMOZ
oCnvOxISLQCyd3c1+WYgtMukTM51OxyxbthUVRUaw56HNPDchQmiB5b3ADlLqfBmYDAmMn0vqPTs
a+LEjfq7ZOryeq5ZpayzWN5IjA+2pa8NL6NbwS0Igu2Fwoasq66afDVaHq5x26hfUQOmjzGg4lzT
zHsfa06IlnqJuGnmHZiNphvAsyi26ZVVaz0pP9vpBgWRiKjsn6ACgPUzcoko6lx54sClPlD/5LxA
NwtOzifk/pyT5tzXk0kaXXUN9HK3lXOPJFjilI+mOxkQeCbJn3pm8g/tXdoxa8ZAwHmLqRI+OzCv
0hVRsh7Ja9bBZxXYYzY8J+XQoyP3CZbSZyjAUqkPoKT1zAYO1nYEoNOtRZf+HK8zrVfDV15vOTrU
CHDIcI+d+EMAzy6w7HtR623kulzq/nK+CIudT8bi4fTEMNaOtn+//VkZR5IDPZwGx4jnPf6xjrYZ
gLJXbPAyxQxWSLRzUAWulsrqjYIYTwEUjVwL9arPCyZ6Tecd9VBfFOjMuqYgbIvU8LhF9eOU9XtM
YbnhP/j5ciP9CDBmvmVvkskPj/HUgyB1pTTG48ITAcw6QP9Fse9Di8DGO2/xNY35o+iAkxSIv8a5
/RM/5I+IHaehWMMGwcaCYwe0oj/z4NAuYNtwJSbQLbtBXaRT8LeST80rIJ9GS8ajxR1bzSbtjPyX
9LETaZEYkejQ8RXZLzWm/g3f4wx/+GeldO2gRpGf+0ylgRw+JUDmGyq2VPmUESBcJOTGt2MHkClX
3uMRAQEM90re2YzEZ0gujNwzbc/uWlFZSuE0AMO25RjXK23akjq9u2cd7Hg/cVkSjQmPoeF77HPd
EESzl7mZjc+orsXOR1hiDWYEInNVtXo7QDiF45n1UwqGE4EJuffBrGuWFLsXyMpYWPRsFsslmhi0
rRBFe9TGiExD4rl+PzXIaEgVk2fd3kB0Sukld2we86BwuFjOX0WM2okIuCYRztuhLWT9PI8bTDjN
EMfIjskBC9CJzBlmqePjkJOZI7O5fOApICJVTN6aSDpmXm4VMNkXQkC5+Z0r4WK6Qg8pzOJtkzRr
+28UUFyDxvGaWeIzu9SPjGo7NrUalWy9dG7KPm7fX41dBuastfaJPPoYNoVyHBi9dBTLWHNYtsMY
jsZJTWNmF+6ueSbfavnbaZjFXku8JlQTvmtqCX5JeCfTo5T0gsxfZykkAOZtsSuUKGk4xntbzj66
oxPHggR/YIno5WAVYd+07wsln5tXs1yDJA99iEZnvr4pbU6yJPQB9pf1YLqXLvbgpTi5WJxSStSf
aGecyMRmCcPjE0DLIKxbtJeN1o2u+3naCPyq65OwGO6gHIgJZ+Hb4dShPtvOD3Q+uJt/gsfAGY5W
hw3+vzWJQgLvIoO72jV2VC3C86FKsLK7zU0WJVhFGVAzdVzVYVD4xzQbk31jISJgsh7YERE8gDct
BPArhxsvXJ5CEwdrT46UKBpThWGgz3+MxB2zpIVc8tx7mtA1hbp1dfg5hDVaDcnJbn93jow+MbEz
cWCdU8T+sTNW1b4OqA6UM8cefTiiSaadzZrR878UuKso/YGpWMzZZcOFMhQ3R618D7xc+pUtGPve
g3UBuzSgMAAOLfefo5IA0YtRRLWH42QgplWnfBbv6VAAAaopbDs/yw8XRhgAFmROZEDUXfpUA3BS
z8A+2Dz92rBYIPdcPeX3Mwx8xXB3BHgpLhaLKy2qkNHnIrO7Sx0oFeKu3FoK3iLi+ONZ6w6riy5U
uaNxcJ6XIbHx7bZV7cQRo8sIm/0UlNj96Mw29tmuntShlVkBGr8/5PK+eR4vtyaMNkbwTaqCWRlK
emAF449rUiw/V1eIxt99EKOe6ScCucX3Y8Mvt7NTzs+o3EjzAnr3cpZEDQ/JjtnzS987DurfwTkY
9v/gv1c05F9Rm3iY1J7mNvDhZBfMrN8Mmw34BR2rUKMohHdgkgc0G99uNxrhY0kEguhZtR9gCe1n
dU86Wfjozs+q4gmXmiFIA9Hi4G8069NFRXCXOEeAH5AlyC4F1tNJC9V7lfxhAv9NcBWCZqdO/9Ur
yv7Nf2Ii6MVF2WNtYUn5Hbv9ZCraCDH8YBMsKHUhChxEjdAYuOa6/L0Uu+4xgRxhI0UKa+PVxo3h
HLH3+GIK0udzvpye2LopC3gWr9KYs3Yp9r9ckHZGxoVAZpkup3hLqZP2i/bpXMN4CgqDWQwba1gU
10ZMav1vDmy+Y2vNrL47bXXr3hLQtP9deuQZ1kdIH7p5WwzewjdbMSCyPMf1ragU66+HaApQ1+pl
/ZeJ8CJpm92U2oBoIKhbqGWPOg8c3u92dN+oJ68sqmCrbejUI2zANa2WJEUXPuRIlwkAsbIBIdDG
SN1onAB4CYXV3bfMSTbParKEF0DIlMuAEBl0BMaJnuR21brVYzx4cYCIARbfmW6BxT8LiawTca+S
iToWZsfuZpFOsClkA7pEQQkpea2XB/HFE/X+puGL4igWpnDWXbEIOigp9Wc04mRS88MMcKtUTPBh
fFyBLXnRzGjwAD6O2UIRqq0VAFTw7FHgxxx544lxTBwJe/NEqTLuyislc7V3jp3boLE9xVVyD9Oe
ISp6aN48iFF47dq0UpocC84zPdGSnbU8Ov0FSArYzPGLhD9O+oCsQNxS6C8U/AlB73kR6QZB25KH
SweloOOkVFvpoyE8TThZy/sYjWvmwLPijXkhFl0/JGLyumWwPzEVmeIrbwW659soUD9GBsDD8ez2
jEAUeTJ6F83MnoMYbAHgjKgW1dTr0c5HT92v99rJy/p++GPwsBm1lM1NRpmda5ddqQ9CQ3mClOad
ralifAdTVWCvnC7eDAoX2NrkljbeLTP2xnb8daKtxFBOjA2nHsvg/KTGUng8YdCqj6/UfSwzxJXN
zFGDsMdv8RjUmWYQwe5Aan8sWPVAqo7Vi8t5rgcfwq0t5TzSwa4G1ium6QUR/qK5c654+gDvVsmh
d0eNc7cXE3LE4/e7xLD6yUs5pFjb5KOy9UfbDjgEHw8JNUdjOp6kGCBhK+2WA66g5qHWnAHwl6MU
ASCs8yBRJhtowy/dHNLWCrm4sbbGCR2Lw0lHvjEV/mEB9vsd19jitkl8azN5F3TOIXlZLnsBtqR7
TQazW2IdR9oX1q7P6WGbu0GhTtK8kgsqNI4kPcORgrwvhn58mRZSJVtRdSiVlPm6tkLHy67VztFX
P1aWDTFQn+8kmijlWZzVmEfM2faGXSFQxoX3WB4qJifa0Bwt4eJYWm5OrP4hoVYBKHLCtrFFZ9io
toxHCGwQvYrCrpkGhYa4WSyZE0u+cJwJs5IUIteq+R7Sw00F9EHuf9BVUsLSfNaxfkhybOGdWPF6
hgFP2upmtBO9mZGva5rkdPB1wNKE/v0T27vG7iOEExMd0VHjSNDjKVz0fYfF7bEMBV+ta/kmir2+
4qPNP9IsZgI4p3CTQ4xZ0QjoWo6wpSrv5O9JacKM38ZlSvjExG4vKqgocyMM40dvBOj08HAaiUZ+
qsXcZ5wiH0pgFs38HFXip+Dtz9bRcNUTz1vDDym18+YInGHRdICUb0+o1iMVXYcnwAQja5cuVoCN
uYXD4vzcINobwqHrQRPCesCR6SxeLD3pKHFpvQV0cefJlHrtI57vyQ6ef88A43uVn2VKuSigoBtN
ncaS663iaWaS69vq1zXrAA2H0kXu/FLGhnPicudF/BA5yCCgwmUlYymNm1vvcKWtR5o/mJXqFBS8
T/fL+K8+x+dhdnePerkGm/YhuJyEg4CxmdQaMDayDCMjtkVtpd1FnX9yMB9NqOiYpXi+JhC0xacx
iYscO0FOuSEu3LcNd8qhpI1H3mRjocOBjQ7ju9YN9p2ajZm5P8BNGVgdubFg0G0m9SuPMu0mYivE
jktn9U5yBM9zfqyJ+NCu7LyeQR55SB0vMGueQ2zAd4vOhx+yaLbWLDgnFQl9osrU+94GJdc24EGs
wcWorbP1HjSHSt8wNhfXI/umZ9ymG5vDQdL2L1E/yhSL1xD+OPPPYEWCp93lBWnz63dh3uGaT+pi
hWNwc6G3+zZftx4cw45w8xMBQkJnGARhJn0SpqXRqX4ClMqCB0BKseKRJa75yCL0DAVIqZbCtRPB
W2Zu/S+xD9OuTWpkwVHgd8ZmE4k4Tvha7yy8Li3mk4ykx5en065/XZldGzkOU5VGjFQWM1is3rql
8l4IUShW/keaVMb/CZrmzLZJ0xuXwUKMIYJqBqMD/p8lTzMdW3nc9tbYUWZxVl3z1Z9lehb6mFPa
xM2LjOD65jA+/4ndac2h/qIPdnhQR1x3Mb6zTbuVNXop+afDjI/Lu3ooVRIKuC++NnfLMAVlH6Jz
aJkd+CaFKYI6giRFoOUyJ2pla6uG+fKHSPL7gXpS+KUmVuHtunKMHIZVTWTX5/oNU/45ZheESK4g
NHuPI9MtVA3JG2Kdp0Z/QTZWcPGKRSxYbAhM3G36uYoPl/HJ59cNrXuMmmZCWKB+a8V2lTmxKl76
ollj00zSmm7dqufTdmMH8DO3fYwFKKVxgv7l309boEo7iDiY4tWn0Ltx9f/NazaZAkvNhJwcm6/I
59CRwauCwvjACUsaGJsKIK5mJRuYupGwAZ7eS3Ol2uBkFqeEQ2rH9Y8RqAQvfP/2H7Js5eQKnZng
wvHlXvu1S59tSljHXU91RHpIIb84Vo2oOzCc99r77Z7DfTq/7hk5HdGS5tkWKUoMrt9vHIDrMRJh
XRnXNQ9EFKQmd37ahmLi0sVGEJMXOJDxot7p1Td23CFWj5BNHFy0A1z94xoZq7Hq0wctgfycYV6h
toFpRQ8ymgMlmfNQw+heereq35JBSk8PToUQnbdiL9/4wgUA99W9nT9EKEygHJ8yIPRZFNkoxhkS
IasXyUjJcNotvf1UHlb6PPl7D71/TPzZj33PMcazEdw7mSWdaXLynYpNPNZ0BgscdoBBdMRN37cv
CGR8uI6OJQ1tYEg50HXYEpO5vYYgeb4e2qVUNvupeD3m/HTTKXEK06jX6rTF8dsm8zUXigYY2HJI
mgVVucUl5vPnZAfWi3lqhjHNydaqv68r195JRqH/CN1c+acFfxPQ5Ba3m2Lq7FHdmYrIS1I5nsEP
HGyWpGywUec53m6Hx2DzKPq+97sWXFsBhFC1TAHy4eATTBfZzRIWg+CZLvvNVjCs9qldm1KlALVN
39FcYduu/fWxtCBgnqvgzp4mWs6xSPl6Pr7Vke38aY8J1QhdejQepds0ZShCdL7h67u1mHGyJflt
F5AFGegDDc7765Ga6W3zt1V1fMY9NRFOg09CfqEit4zKBlbbtR5ff1HaTmYww/mKGqQvn/27x4WI
hXr8IU290x4WcA5nx5jgioSq0euKRESoAuMzAgZRhjae2AbIzc7b0USuWCuwCmtsPtj7s+HAAWU1
cd+b3Ol3qdDAWtkyhu8RykOaGNvMmzzSZ2MaM2pluTKkoFG0Xo7d3aCZx8dlX4SLzVlLChMyqua7
wI1GXjkUHbJDecvfkjlE3c/HPgmZJcZvLtC06bg0l4nu6Itn7svg1407zNPJMxTBXydyC6tsoikU
648v6C8TkhWZKTrmHZblagwNCYTWcQBinXyu1lqacfOfy0BHT5hF6X3TA2OLZ9J4Fv5coyP7Ns6w
JBzzH7MJ2ch6UsTxk8x05E4b7BoQ6IRtfKaCnLw5zhn2MsOb8083bWK7TXWpRDS4S/ohdP44LUAX
8kfk0p6M3BMBVibNOd3dN38wP/Pco/M0ked85rSRGoDeoOjNK/N9vt3bKYhV3GT5+G1KjQit3rWZ
L0KGvYBTJ65tT+oM79SPGEt5jnzxOF+OMlXoCAF1wf5z7jH3l8ASrH3Za/Prh7toZZy2u9nNVaaR
Pe5wTvlNVFr/koHjKnlbZCR/rtYquOR2hf/E7peO67HrkiJYg6s5Q25paMJsthKm3FCo51/NfYde
k0TeiKHvd2spXqcWnVIOmPq3wUnoeYhTJlA+2gATcj+ACtQO0LUJu1vGfgXNOofrMXoZmD/NcWwG
Q+CbbJuQDfXGJXsvKbUHR7uP4f4rqV2O37AZCH8oevksgfeyHEHQTFYJmnwOW5ar0LrOG54vk7fp
gRdAM2xl3hkDCHUeV2EyPK1cvArXueD6NCNKqnvva18ptlhYdZLvJRsMR4AUfmGXgLBJf80nhT0s
qytxJiORdtAXRDFucq9frR5HMTlUAGDRWgBM9B00Oc70kbYLksOGpP2ZVHMaQq2BqG843vLmmOKB
IXzYPvWDD3qpDlz+8Rzn1bB3fUNXqMb3f5vGgOOgpXbUTkqXH1S+11QsxzOzLUhvjObvRzSFrrb3
0iNx+OvstQeCDM2SubukNKvgRmiWPatJ7ZZQnW2oUfR0e4G9V2aCHCVfwrrE4Ydl8Jo3OkI0yCzo
6xkZTgp1RRvA4YXxeSQAdFJ2IvtHUw8o2z4amWN8zYB8Q5zpMo/uk2MsMQRoKSliwzIzoyvdZl58
3ubwZBHEpVF3DleMIP1oo5e3sS5tfTbZYHhxq5g41zZ+lAXVh4U07hLP+3qM7Zw/9kw1oCACTwmp
5YXBipckTnR0RL47O5FDfhJRxJvu7zQeZUujopHXnWWUTRhFQTajMXxn8Q4Wh32btzBlANdwqzty
gFgPlhZyvDcim6ekCpak1sR2MDlOnOC4aPsJaBNYLVk7Upcj8lNJv7AcupGCAP0j1Uy1CNs1f1tl
+GrAr42qGTyFudq4v0YfCrRC/P2RnSuypkhAxBNrBh5pLk617eKbGh1TzHx6d/fMLU3AWddeotAi
d9zITar/jSN4HR2sG/b8neRt1FxMXmAi78hvifZQhaOAHJ47rR2t6iCiVOwnRV5gb/8y3Wc7oOf2
nR90xm0GbzOchaW4RI7wShRBbNqsOHZHFe2vKOwtGlAdkEg44R4xxRV7ZoNSpvX9TcB+BB41f02K
AJ98m4joxKxAkE8/u125G4yRfeAM1K5ssmT7lGzCMzVzoEaBPhUrr3QJoNEW71JJeGcnfdre67Uu
L6qG3vG1zfIHIc/qUGCWWd+xb/fFw7sRSjFFGDy8e66v0AO3Q4A2WA5f+DO7bfeWL8DUccwobgyk
lLUOHbOfuRq5L1/Iu6JVvXWlb6Lv+U2r62wrLCGc8doecgS5PrLFqwVLA5QeXepzDvY3e9Dk/twf
v8soDn0nE0hdGumInhLBP+2qOc9ju15YamEWMUYoDL85zyRBVEHJguEX2PXS5BZPviJGD2Tj5IjY
ZES4MLX1A7a6nBUcRRZbE6yJF/Lp/idkTwzOpix+mXsitIu/5m5QgBLR2KcvP8mZmOg5ve5h8MYl
UdFcrWANH2S90Iv0xjfpq3DWKAtf72SAl71x2xqTxSCzrGGexcfpve5d0+3fvdR85nX3DmN4oPAW
5yqbW+J0QPhbiUXHhA83/5Ebsgi0xDN3OKtbOOztpnhTGliDbof6gBRwsG20e84L3plIsft9HUML
Xi6FjD0uYcA1Cr/14xlXwVbZW93UaQzLvaL3jnjanZ7dKr2cKFzB+19K03hamGl2OhCLI1HD6L/p
NIRqCiDMeUjRGYieMBR1rYeZY3AOla0MnLQplWS6kPOlgtikZpXt7/7TieQkSYpaMnblrtVEM2Jq
BTAqQn/FCwY9Yg9Yf1yKfnNt4BRBm/mQH92akWzY8oyxeZaRlbQG915uXTspDpu1+4S8b8sfbbkQ
3jK4dDMUmq94b0purpLzwn7AcCcxGcKvUBUxu+7apGoBABprYhkPQNBcXYz8L5ozctLJavIJIuOM
snCtDw34xdTfMbFlnD1fh7Pe+KFGIQQlFOeSTiDu8yCVGJr3bk1zwwiMKGHmuAha7EtlD2m7izrS
ym4FtiiPB3ZYabgu0ozKKk1c97drvyH5qF7NA+RTgaKmB8Bq7B0RtXw8T+kjpyq1Of1e2fbDOtXi
uxAwZYgnzz2sjFfb5wqdBdhCfzFpUyeZvHSQpBhHnxtf5KUbyy4MXx90hdQJegQtwBgcstDEx+5n
lsWJLzN33/2a+Z3WZNOBS4pLKWM6MvBMBa4ixjHV5nXH0/lxSjENGZw3WUdm/kZItpB489P0C8uD
oG8nI49a/R7XbdeDPWXLMXJ3ysaJway9BJoPUKjHPn2zWs0MFxyW2CWBEgcOoVC+o+q+bSdEreCL
yLCzpPV8CxpF2zwpAbId6r+NJsKiobx076QTIlaixG10nWBVTn//VFmLPuXxzh+veIVmIO8l61hB
UO2RpX4RbUF1I6GclTMHpVt95AuIb1qa4UOu8qxlFnCnr75htXv2WOKXGIPQApbSWK5cIEKXk3vg
ZfllI1FRkzlHsEB6rP4YF7pfLQAfKKJroHLtIWDR7+xhlnl6eO7FYaRuFZdALy7j6kK9Y+LjMSt5
g1WSJ49m9QWiL8nw5ih4hESLTRIsubYyvs+DWBI1EWFRO31r4ProdD2LTPMe4kPs3ROwkm4VZUgI
zbxDvXtqdhTLtbQ4xY0y/a1UT6weRGQlcbPS/dA9Dru5Sc/e5Fj/QqWrR8I0UA+ddK0VPACHAgMC
EhDrOCle+NWNQZRkZveuYjqLKYCk70Vd3XM3WCwGVZFrLaY/AdMVOmKc4gidXRH/hc/Q/SsIK0F2
DCTWxRdWRUKfrUlyFwMJ+lgkOEYMyMrl6QF0NjRmFItAICDQAmmDWygmHAr5sJ7t0mzfCIxda4AB
j4ULhTaAuxQjRh8HlEnglw4/uf9o2SciF1rSTT1AsaIu4PFfuHrfJKWeTd6JrmgNga2G86YaNT9r
fPPA4T60i9v0U0dAWYrjHK4rsi5nbcnyqnUJzVUMBkOWjFgjJV5ANXbsa2ydX3yr2AxWzGhI6pLD
cP1YbtkAxPRumOt2gImMXeDkzaJy/WrRqcEj3IFte4TqGtceUXy4f1gN3P4VuQtLi/ed4evIUsNx
C4U448cx/X5AN2Rs7nWd8Xp0YO0vrfMHlDOt4HOD/FEKTuV4wh4wHeN0sVZb297he4y6rsMiItiF
sRGYAQoqHohay01vS4a4+mmWmpxhoNEklbCov/AYXJ8rn21pvAsIIgxtJlhK1eOfQFx2xDB7AyAa
4Cu8SbYaN83sT2r4JYKT0PBqdwuQ5DnBXYoxz1/fAS2pDLO7cq8ekmta/Ca4gd+Ipo4sJ6JftQfJ
qduVm43E2DSrbFYAg/nC37pbiy7MmBMb8Wl7dr170tbtV79MT6cg4YnjpENQJdBVCH56pRjAcPls
XdN7SzTDo7SSuv5Oafl4RW6pUi7nMt3dholaRU2Gi5a0JL+X0zSwiQkwicAJEbhmGpj07695dGaz
ZuIsPW4/LTdur4AiKbeZ9bMKX9VwJT+VlCZBfs/3b+zy0gh0gMuXiLRYPx0aRvDK3Fbj1bvpoj1B
M5ebnlk8HFjtxfoyTgWCFuN6IaCvX9LG+nXym83SEHUETRzK04qN7wuNDTtMckXKivw2nHG1Oj0X
G36uFWrPG3r9x92yhLtiIy24guNjSDGk51bpk3DJgtAEfE3K35kZ1wNpBcvr0yfPq5aPnnVcagO8
SK5XRIm8FIivEygNWHPcMS18+SGDFoq2bGjTwL1dJFwYlESJfzx9J2FYnOFO4ZeYkVSK9jg4mBWj
vkGpeZoeaHdcc1tU7bJcUUxJTqGAxL9vSIQ608mKGpVsyfn09ltvJElV9v61UgsHcAsWUZUxAiEz
2z5jn02CLyYbuN2rJspKW+Y/jPdHLJgxsARBlkpvpo9b3zvsIQ9IDpCPxpRvNUO2Wv/nzotK2PLV
n818OjBr4lWLvsNUCpewGbUduAdMU3At+51eFBJr/JZsjkl8K1SnRiW6H+IVCtQDBWKHM/y+XT1o
0dE/FkB8tW4ZTs33MxhQU9li8ZXnm4pBRRtwcnlT+tzvGzt6TdgDjriTOBrrDYThtoOqjPDXEr/e
6DR86HsP/RySrcMaqpqIQoqjDhmQ8q56m2y1RLHse6hOrWiF21tBlEzrXtKCnY9yziuQwqzOZyB7
wTIV2VKOa4SdK6KX2zGYgq1ZrqADxdeQMrRXn4mgWLr/89DJKmFiojH4MsBqVCZvoK2ZCTrRBtrh
BcIdxtJ3GoxadtpaxFZex+Q5p4NSoysl4ap6HkSxdEq1U1x/8NbtGm0sWEdWyFMug95i080oeYeM
xDGHzKlCQgxFUq2ykGGVFlPusn0X7zwVmXOERoJfTeuI3p9tYz5zKVrCNObCL6YbxBUZAHbiWDho
FjHjnkne1Y7GEaxw/w1uaNGyPj3HZjaoveRy+5zCb9n27zvqvbTxOuoPL+f2b/CuQA4uTy2JNUcY
bpsBXPAoh0nfJyriltDMCkiew4IPCzg4IJcZsP2VzaEeK4W1bqKCuOXAZcX3dbLN0Fp8L7JHWKvA
THpCmc0F5twycjFDvYgSEtO6vxCBxt9g5tSg8PLBjwYFr7bt4tOnACzetFf2vUgkmTU82xLm6PQR
QZ+CfnnAbjtwYVMn78/CLs5wdk6TKUJ+15pFMZ8I2etz0qCEalqANcEXqWPuhsCBtG6haqVbDOty
JcqgNfscGg7jkUGaquqEw7NzQUqZfdbLLXLyLKjo1ZGeWEld9lTItPsrGPkzdxjofxv1yCX5/H7c
zlVYYbs+pIowS4JDZXBw8NEqtkf4ucV1CFiYIgSfs+cB6KcmzAzMXvDp3KkQ+clCewuYoZmd0sP3
DTKdGGa6oUb04nWNFxyizdA5PElcpAaL8dFeRLeWwiloqiYSBT8pl2h551oss8J3c0OtfKyRE/uj
91i4i2PREHLnFa7M1aAqSOTO4EIckulyXWFqpOZ53djVlFNseL9J1lR9VDj69IDWPl7NTYOU+XW4
vVXEGh4HLNqXp97Px6gW4WF3WSLsXCzUPmBBNr/4Sq62XAMGyliroLVtZYtIT+p7rKOUDGaR6pWz
+bOk2MeowABZzABJETn6uBRmXuENb9v4ZOMsGQxMbyPnZwNk01ForlBOrVGFFwbxCAY7U5TjbZGV
kUA++8iHVOK1x8mRIimVuZOwofcQ72IT78CCb4R4MA01QM2NNrtx/Yr8BWOfEB26R9JDa570LulM
M49Wnn3j32tBSESGnnQcCNg2izWXzC1vMBmJ5qd9wxzpYLeycC6Bm46fVL/lQQMpCkAH1VfLp71O
CLpkOv/rXPpU9nOGRq8m+rxf5Gko78AZy3fV2n0s18ZpALwxZoYoead97FKvOKBXy1uC+xwNVANM
sfA5vdHJzDHsEOek4iJnQjE28pDilMh3dr8O2XC+1+KmNqx1SZ6djRpsedPWAPseDX6+NesRF0eO
6MzdDELGfJfIONxFKHX0p3wKid3RpG4RIIlrpvP68t3rJLIfkuNZHffZ6KESJC6m6PgYgYQHZQ6B
++fpIMllgKu+D3adj7UkmH3EycENlojZvDVNd1Q8j1XoUOZOdm2AI6TWnVH4p9HRTWKaFHv8GQxx
Wo+FWGMy4KPbPinOdaeZ1PSSwjnr4kv/dvctpBAtKpQk3deMftiIkXULcgxAhuKA4u+7oXO9O/3R
7apodO+wuxNE/hYhGagyR4goKR8TWDkE5Kh/Ynnb5ezfX0PDb2N+GjIJ+rV0anLs0MtiymNXgINK
ttBMtyk28G/ATWF0RrvNviKrJlt9bnL1lxHbPuWje695f0cP9r1zGgoTzFRJhwIk9zYMDX/YaD29
amBKqv1stGb2jhaFfgy+kcfx/0gsJcr+X4ZY/Mm28DgzVYnWmWUWrpLQ6M5h6PLIme+hgOGutaOB
IcF/3sTeVZ9S8lFnG1rgLrIuUO9Vt9RVttELzxNh0xXBIbPPfBStl6nMS38e+IE4YsAoa//mLp0X
GjBP9iE3ZHMZ8MznyWyRL/mcQjIk2WTHEd/niAf4zZlAqG57u+zxCTpIAc/TA6p5fD5ePBAUrNy+
/PsEAQU/D8xlpwuP9AvekYFOT9yj7HNFETOH4WExDc/6mUgqHxiraUkJP+xw8EHKHFperWBMEfhv
cInGaiYevb9WzwdsUogb8ZqBt4qq9N+O8Bo9zsPVLxhYRr5o5ZO/RBg43OElSVPfQnhasv40N/Sm
dXknuWIPBSpTcZ/rjCVf8JTO7pimnC2ntjyhMPYApgehz33KIPwr4rnZ4hrjXCP7EXz7q7csMffH
puzusV7k/jXdFRvqnq35ZPlFtGWjF1bokBXVA6hcSGppFzlcKVzDySjSPHyc9zXzdO5chx2iOZjH
V31m3S9UDufHM1rySg5djcMyuRTKaL7IWbQ0W9Y0O+gLBmrRtzsm9udEcWuqH9d9hnfYjN42r1LL
I5TCemZ1/br5gvwqQZhVt4Ln4G3G+oNsSSdpy+4Wx0Iuu+oqiIiImID3GohzOrF3vld9cq/wGA55
4SaPIV7RAuWm/nMeSYNOOA3JcoRPSZ/+o2lmSXln0cGBep1hA/ei6k8RaakzlqBTV9fZaC41SJNF
1LZIuFFezDHixqZH6lyUmWaDVjEo1yozWV0nnAFPApYG46g1txXGLiG9Ecgq5z5D/E5fJFNB32hB
nkinc0EJZOplOSwk07YX50OWyvPOYMnYMA+PBP1vpMe3KLfkg18R33PUtLaKaiKJTrdkv4hZEWxC
4lnazP0RZxpyeK67ONyXSzdTXhlmAKY2rA/wlslQc+2UrRoiRbjLZk7aaKP4PZjq35qDUlkK/7+g
zIX+phjkc8UNZRiHb0UI1cXSz9nFeFCvszHtLVkp0OPV0zFoU+llwWa0MATdd6mmSh+nAcmxG5xR
c+iU6arFuWcllHQDcOqpGtw21aFlgUSl4cJO6ZAJtU2tKFtxIBYNEU2FSD+OZdJIfn4kxdBM91HC
AFvg0tEOQ2RI1ldsMaokRmW+A3Ltsg2cOQxDG7/md/3TqFE7j4dRZ+QoyvlT6TcwAoWzlxPT1pLI
vlqGBlMO5REicvevmVWZMAzEnHkQrmTGPypOEvBZczPWyTFqNspM+nFvbx2eCTPH9pHEHrP0gzYA
X4IN9lzaauPloiuJhNiVQYgfx61FPEvMb2dVJDwgzIokimDcH9eYKGNMmBV8t130486RA0HYP1AU
FIM39YPcISXHP10VTZ+CDuASkwoS/VAQ+S71Y7+1BolSm/IYLIMN6QjNuTeazeCkWfYZ3bAqLsMB
FS0+lcfNtkbA20oFttigZ4qp4a8pLYsoApaU76DXK4iJbE1sOFLLsngihkuzmOjgkN1JDRz54KdT
0Y9t2RBzQj0sPd2tWn0FTWn44Y6y7MZ5S1b6qABuY05b0ajDaENBhq+evHXgpWK+1hCI5UmvOlbp
Yn+hk8dsaBIpn7auvB9AWgAV9T0RA4BSEAL6zckUvKF0DTMwfAcUtYZ4DU6sm3yY0NXUVSfB29UJ
MsyAK1fXt608DQ1pb0dLFHBiMdcY2Sfb5PF9dig7WplXKLTY3hJjVJ6vAQRYNRw9MJSI5p6FL/2Q
mpNsV+vL8AFarFV2EWMFduY1KXX7nO+9o2VgYdNuqikA47byCU1Zu5/OUkN6pmalri+HZpHOQKHL
DK5sVOZrW44i1N7bVcyOI5WYutHwAMQ+FIdPFcSN8EQsMmQxx40yb6BdnoBb6v5JHZWRU6KTtJTu
0THn2lHBkDBHaqOQQVuzGJ2WIoPexIfIW2qY1qGKIEUZcyTwJi8qZXO69QbAZXhzM0gvPz2E7SNP
enlyg9V5sgwReo2wXCSwRnM4grOx4KhvvpXtT4GgOdDe0dWZ3xJCk3FmA+bZ2xQV9ALJS12grIBM
LiNMGpSbQjsDxSZSpygv7cjmz8ECa97kyG+YtdFbte4RnV85rC7xQDBYLpAG4zU8lcg2/gQXcZDs
kCwjO9SBmwnYGjAAjN93joZ6ytZFXmoptBloII89n7ga/7lPnXMmUovW6HSYrueR6LMV8JIAkpd0
FjX8bbE2+dsIj8r0pvulE3ntn8xoLevfwTVb8LxC1uMCVS6zWc9cAsHedliWPyfCQks7iogqQJMw
nBmYm36UQ71G2hT/7qP6b6WyPmpRFo0rujmF0vTA3Sn75kSZlOZ9HfP5iQAFTBc/+PcN2hEE7ljL
wSk5xKdtVuUI5xMjGHrkp30FxMd7K8f9A/JZkYkHl2D3hECBqppPIcYe+Ag34neTP88K/Qi8djbA
IXlBSRzVOuoD7AJMR365Rk7srKHBNIh4BZmOZGSn2QFgOqzZrsckCBY84l/LWjH9BMRsJF4g1brO
DUnK2jhAO69gDJHdNdmS9QkYh3EpcDmh2/hHhE7IrOLkSebBThb83Z4rVrYXQjpDlxmej+qv8+/v
FcGm+x/CDFY0vKtpwYC3Qa9qstC9RXgDsK5iAlRxn5dxYGXaVidtF6P58CnT0MwfxMfaO9Dayb5x
gYYi6WXWKkDaR4XrkMagub6dd1FH5dAl1+F/oBwOMPl0+oID9/xHlqpy7RQwe1YIHsx8isDNXKdc
y5vQfYVWy9MFwOoknVIOzcubEjkXaj0a3tI7FT38ahZqvSGg75p3K2AnJsdjW8hdcs1Go/wD8vPQ
GerzSDYIK1QMLV8Krf+at3OSX3cxUeiydQ7EcH/g6cpvkMnc66R5s7rNjbDvpL7uLA0fyUF1pDTg
Fg5Y9qRT4eaAG66szegVIn4SUuGx0ZsMV3ZPhrRiQqAr6Jsbfg2iR/3l4wNtyW3HTZTHk7sU8XLs
7esaVyb1UGcUUj4JMnw89tRQJJflo6gMY/trHFgpjNke0m3auIpnrWU/hT5DF7pwClFEP0rEwbNE
gEXahENJaEbqbSt0NB2Q583zO/PSMYK2OomUjxzwkRifHE0YGCxelFrXpedLbrwjX+btPhQEsl8q
2xkI0KXcCN4ezRcyjO24TCY1OCEttgmWcI7DANZQRHXg19Y20YBeO9MuxGqEjAZ8heZAWKc9DHFU
W9WVKCNdzRBQqWUpHSxpTBDuY0/BdwKpNsywzccdYkOhXjH8Cyrf5P7/ZugpCmAzihKzDXi025ml
JVwzNT4CClyHhc3LS8fZJzAq5CKaXlj80te3SCV3+3S7cgIrEDIlHtV1RTz0H7WhAzHhPw0uxGYa
A3xZ6y9/eIcP7eTdBBKLfe9wjhuPVuawcj/S7ouuhIFCLO1xdyUzxF/EfUOmsantU2j3uNKuKAdY
p1nvqyOX3dciIIF1lFySZyKCn5EAsDzhIVGmtwLNG56aI+W4FMit7NVrRjayHRwV/MNjr3EHKXvm
coNOvQX1VBX4k6bhUGizZCuKTf64tFf8JwskBK8OZ3JvvJCu9y3ykTk1XzH2KaceAE6qQt5BQCMl
hLQa5fsX8uRWUH25tb3jeNfmNLirfTGgJwPDKm0MdyiJMdYTDDgWIo6FvzSJ19Nejlu809Oqy0Ob
SFdynX9xlkbLRpOHa9xgBFvD27+9gs+y4xo2pAt32bryzCTAYkG8sS5AJH6zGRz73VAmjLUfMGTp
yoTx9SO70tLSsZkYc9hfJqu+4cYuwA+BoVbdV51D8f9Y9jKI6x5I+HdbGvRjDkIosBa3amFLM4eT
kXp0azIXXEtgGglWuuqdkYXl6Ac+3EiOkJswUHGVT6GmDYWaSpwIbe6U3wqgDkOtfhN6gxnNgvs8
Dx04wRL4Idwk0aoiUBchAeLQmwpGXO1bsHKdPil/kWTa4abAJRj+Qk+ccobkzpoEcwR+wfoXwBJf
7gqH5m+M0bgaSc50F4gd20bPNIbGZnN95IA+nLyr4i/BSQ1tMkIa4sOtOuJYIHMWCGs6B6/sN/ML
hioM2ttc7LPB3xa6DW+6Qo/KoekUjb8//zHsBmQBZv9Kz9rzWQWvuDyv2hUhpnzbdfYIibvma6ac
06YA9u1pOBRksBCP07437giEBROera1yZ7nwNi8fVLsmGXLV7XKLPQkpeDQqono3xJfqGFxIv/v6
JFC0pChdQ8xa2Z56/wkOC48QQzbY1KI+bfAhGusdRh9GWmkpaX3bBnplotmY8XHICyqsrvOcsarg
D+DGa6TGKXTzajlH8xA/23CniicvP7YAygIWNcRqOZ+E0ThCA7gvjpSoVKm1iWZJRsqzfWtFwctz
kNJuYieJgtCcqCC8nqQcs8td9el8nls8aMz7wMsAoVouA+SsqoYq0ROiTNy0GS6rZykXubbaaZ7I
QpS1IiKK+P5/8X89DjQRu6SVkZAV/NJ7MVrc/J+3l6vEqPy3yahkQFe10EHLPRulCjaJdXhLpidi
qZRHLv5mn4vEC09PsoKj3JVCYa7l4NwvP3cieXzHtrOhK2Jz2Tg9hRvYmljzNXcLZcj5JQwFafCy
0n96+4d/2QtT81zvU0Y38tUH2iHZg1eovqmQN38ghoI3oLE1ijO+3lLblF1thSWXDo4NDP8cB5oj
vAyehZCJY5nXJyn3WF5KdGccR8/bu+hxpCk4iSoBziM+fTl79rcXEel3+TOYtcnC2odNKtPmTO1n
JdZ1+127Lw795eyNq3jqQTnjtJ0rYfhOyHY4X85ICJJV8F5sRFLvvX0QVfZHcHmHz4dX6AO6eMzo
pa5MDKb/5SzKnpbzZO+IeouRJSJG/nbcLgjbh3XD6Sd7NNW1GX8VrtlDM3Vbdc5UL9GSX1qcr29m
/ezUZ/0TjAtcHWmDOKAgglCuvETYKH/BWG7j2ciFzrEDC/R18fBOfis0tE8C+wKPU98/OMiypgOH
+Qt6h2zpLqCYRvwBGxrqnjTlJo18XC0xLKZB3xQ0MVEcrBmNXvl4fmiHyDBxBoQZVfM3pdpUdqus
Xc91o/sYPuSUzQzNQTTZB0UbvC1gwFh+KyiQQ9wuwTwiO2Bn+o+WfdMlr8BN9QsmxczY/2lv6TuE
ye78HZIfiMU7g1HmRO93p6Ky7epDJcNWW0Un8aHi3z6hVrQjSBZFiP4aIknDjiYmB6uWnU1JCtYD
X9g5HtVYA8aNC/ge7l3pfSTVfzAsutg4fvyGrFOHqYTw2KpzS0pusOOI9VCVMkIuq84vrV2zLedd
z0pQ50cvgjfMhnabvjHffolfhH4F9VBFEApvbdOwMU+YMa6ggmYCj0GKV2aKXlbRw/mQje36M4cF
EzQjuc3F2GN5/WpujsAhLLQY8JF4RCDo0zskli6JwtwtZ+NtWPt6rI7SKPQL6Tvi7GQlt6/S4f44
+a83lgrJ9OH0248WR4owzdb0x9jw3QMHYXifGhrBmhZu3/7+pBXcG2lh7jpQsxCNeCplTexNQlZJ
qKlRMpIKNl9PFHyYKzpKRINsm7U7CIrQHihPguLcxRjpkBfoOEbPuPL1hu/LCwIc2Cw7LT4CIken
vNjmARcF5LD4eXHWbr4xKwAc+KMlXM5DRdShyQQahe2ncmzooT+lX7a/qSBeXPjllo7a7dXvewb8
EvsAo4SAh/ZcFKNL2AYT00EUtN1X1TmDp/3HrBB3HmjhxOh1iJPIzagw2Mgm1tj7z7MCuYRccH4Q
6e2Z8ST94s9Lnk1QQEtqxMtUHomo16BUdZkoh9NGMkCt4+nb+pnKfRjmraQXYyuG92DKsLaNz1LQ
LwKf5zhsse+3zRLGMV5uXpBsFIWV5cBHoqnWnzkQuLnRQPoxBbcxQgs4eV93mXCb3zie/nTZpLTe
vH+GLjz5W/arIbxMOHR5+kqALO9stZDQ3aq6MwAfWi/aFexJwkJ8jAsjucaWwmoslB9zLEfbPQ2p
/bXXwo7bdY9YAET+ur0XeF0P/cAuYm2FocAI0I47EM9uV4N9Lk4wynFeDlSI4w7U5+I6ckYGnfkz
dPHKRP04UJRUgYDt64twEnKa5pWgwfQ5JUd1VlhxY3Y3MZmwgC8QODyLY74KFyUqYgLPqEdfEj8S
N9VtzCI17XBrsGd9PpQIY+oEwODHX9E4uY9hoA2txKGQBR8PYqaqAiy7k3TTGwUfQxS1q17sqZJH
Xo1HLtwmZNmdW8PF/f0qd8ymhA1yeod55ZQO70b4raAsH7dxJoXRaFRrtN9c9aG2HGE7fo/jw+Sw
9HDIeQlP+wAKuNqc8+uhosrLVohjDWvbqJV4Jt+wTmUekT0bgT/U0q+wTrgcUle0F30Dd48L2qmm
ko0PzAUB9ENgnlyYbJNm/S/lPyTFaljLP+FFRS+cKUCokmrDrv4OKExHgNYmk89oYoo7/1R6NC7i
rfLS3H5DgoK1oaig2WXz9VMSrhMDazi+YXRkNqt1Yy1fpvxkvpn5V8gzdoabmGKJlzHjBVJ2o9AD
5X99i5u6wIIEr56o5RuUSX1GpfOK3km+6NbJ+UCS1qdrq13qCVzoB5GrjL0Gj6LVmXyKw8JT40zS
vMEttZxVIM0o20f2qvQxn9fE40SUNhqGBr2TPpa1IYXXSHiKDgxCIQv53JzEc446YrKuQoYv6WkK
/Wk+LH5Ei+stGq4X8UnxUusirSoeG3Z+IWxw7iMDrJANto3HoZaF05JJsUINRoQPEJmZj2YJhdqV
qwyjF+28uJslOQSD4Da9beMrDZm7WZOhclOCA72vD2ER3Ykw5xn8Lfkqh3XBKowHqDYzjPUaRu9N
Xyp6j1Z0mn+tbGAXIwOqbHED2nzauwAaK3p9p9/JmbBppRdAAQ/5m2kegqWOAbTR5k3XCoxlfrJD
VmdXroncQxhACh7dVmq65DMnX42hG8PjlP/oUc5ejHH+dgoX09WEfTxs2qJaPqwC/w3f/4Z31FSN
+Bqcm26awGHBc5QKLuPhhkzDGrW7Up6eNZTZxCIMJzp3HRXn192IBJD9rs4DIU/YIMU4sjGdaixM
OrWHuc1v1Sd1rMVdNJ9h3l/nM4klOUBtPnR5XazFIy455gXhREBlCa8dDmhd5kB3NLzyazZP8oS7
oKOkhtJthcroRXkJR/AwyqJfQichrHc7J/+JLMfVOL/FdPHbvlYoPFiP3IONEmlAKgzSjCwj+SZ9
BGkgNPhqlt59JDP0J9j1hPxMBIl6p2qbVpFV6Pj6BufK4x3DCUFFFd1GH8W9qvg4lmC/z8zrL40f
B02Rh7K8NdjrlAdMNNDpWLZNqCQ61LDryyyHHnXNQHxkSSUIiqgK997MItktMhjswvduNcncteVR
iRQjBBKeEGTbOpxKrfdV7tnJCYsVgc/FCK3RNTl7hW5qSTWZCWmgtrtk3HV569w21jAyW3g1S6AP
z5ktSKcskVk2syXEItww+52Z31zHFanBOp+wTnseHvMuO2c6sq4vilQ81Ek+YzzFvflQwDO1t84p
Inzs5pMpaOqaU463iE2etugJfCOa55yU3wTLd48HuSGMjWNwGUNaQUv021tPS8thed1QEdjf+D39
12nd42xr7EG8YBr+rWFdVP91ID8TM9xG/kA3bRS4KySVCspaEJCPi1sr9ZbRb71clN8qwSWDN2tm
gIhuOD2wxgrBKoJ1QIMoVENrAmdQL1rHfFqt5umUw+s7uUthJyyvBhsi3qZVKuzI8c3QwvNwEO2f
/K0zyqCQYg4HGTw3PccjLQ07Ci5dbNym8r33mqce1KhpObpkm/+p6lb2Z/DH8O6aiJl/SBCMrXUu
W8maAXI6GVKefc6Hh7w2Pyj/zELWLkbnFI/VhZTTaBF+W+Vg0s9YJeApeJXq+iuomIz6yYWcCS4C
YIc92Am4mF1ssMYMB0WO6OuomXJcB8KvurCZDkMFRmdAj0L3JIIV5p6d1wLtTgi4TowztKFppRXi
wWuDMPoOSnhW86vlDYzxdx07rfQ6tWJdMN0ByLKxfI7dwMibRvlDNSUDneeGHz+t/BYGbjNBhdv4
1XGpAVkCH+niM8CSdwwofBsrQcONt1FrhYullGDAByeehgwAw+yhIVCRjqXfIfC1HnMnqmQJ1Y5r
7F85h4NPUKld+hV998sOPcJ4vkJ4pam44YC3jCXt0v7UDluJRAzbNAD/AwKD1MuFfn9P2WOogEqb
eJHbpVhBnnaf+sbZNNnC3MmAeuyry+9d/zITEiE+AbiIySwf/aiJhNSLY14oqitycgWJOMGf8HmA
CZXSThE2cNnIXY3AV+/N+3zQwSfEt+PpV1WmjtjWv/3+Z1tmgGuMaMW0LA48MXlFL1fhPvEzjViH
1wybTMEuWe1GlBsv83S4xoZIS5B3r+yJnZ52KnWJEQJqpY0EeWMb6AyJfS0jHYdCXeYgILj6iEaV
pQ0xmGS2blY4H+0iBa+p9ccLlb8w0I5ol0ZBRSumEKMMSqYS2tM5f/yC/sy5OS+Wu1Js4pTyaYl8
A0oQM+Cp0+6hcSKUZyH60c9bx4K9Uchj+ZuRUcaOp283kAq6wKGdoTyCuxa0/UTUgUGBP7C9qqmg
MZ/eppFJfsWkN8c2OCXvRwN8jfkRpxSjonfGhmUC+uMPidPpcJu/GDHXb92n/GJzKUDsLo6I0Cz3
PjkWbbxwuLrFVg+TSQMp+d4TIzYmfH/fQD2x3mlZyh/VelUNoao1KTqVkquV0k+47nlio8ddjjSs
9kDySc7lbEExkhxl6qhNkgb8+LSk08LGwZ7Wj1LeECoSFJ0v0Lwe22EcqaM0LFLJ0suRDhX+yEKm
KqAzQOA+lOlYNk7Fh8YvXCPtL+6acGxb+iMngBjkNwRfuvDK4Ifj6qedHpd62C9B/0mis2cny5BZ
ecrdbf/kiMX327oi/oI/kJNJnDZr1n+ZbMCaEg2+HSBT+STRIRF+gr6J/esLkFMLnS7fLrGzBYWa
dqWFJ2Fo8uMDzt3jYpmj0GK+jR2FYv/9po2BepFFwf0Cngj140n82KzMr4akp9+SZWg/5bRc5ibx
uUjQzcTWFFfH7wPox38NoGdHEEfwuCGOQeCtuPWY4PqTbC/7ITE0L4ExUEDlY8W4sean2E+vsJaK
wXt1V3RnR/DoZup5GAglDmw1zaRcRQWJ2RP2Q6JFVaNZC/H04MhvQaVzX/2t42LndSVPIkqlTE3G
bEF9+6KEE4TudBXnygwOWuQOSUKkZijBrk077O53nYTo7jSiwy9UHAe1PLm+vRV8NC6AK+keI55s
3LMQqZoV8bMEMRZXkHicgapPIHRyFLYZPI6amk+Z1Wu5LhnG81buvDpklYXaTLD2FEMyr/HCyprD
1+bdNgjC4JwXChFCNxyBxkR3HVAbZz62I+fWbDw0RURn77M/LafbWF8p2AdAQ9MyIlUP/oCH1nIc
nCi/Q8AX9s+QkjIP2FuTyqXosCyHIz/kwfS+QpNuv6A4CqEQiVGRCOZ0R8KIuzEnFYAxN1JzPSJV
SpBpyU6f5LC1PxlUCsgk27nYGAykaB9yMfPYHtvGyn2iRxMR54AcTopwlZYJ61SbkJz/NMMBii9w
ljf54S12Wj+DdATfTRQNRNeaTArYoCyziaOQo+vk1UAALDQaBSmBYaOSEU8SIMDMaY7QX1Qg4gdj
m62y/ycVRBtTIaqBiKfNeeb+dQKMPZKbY+NFlDu+otnBm14fzsWsVkr/PTY/UT1hI8bMlmOkk3g1
pwD855uLiDFptWtlgyXdG1OuOT/FObcHGarD14kKiqOQ4TTx9JRJhr181fIpR6pMpDUCLKdVvbGG
6ez41izaLgx0PTHWevzaCQiEJs+feF8FhfuaUVyyStQHBKmX2P3pfJ0QUNX5ZWaiQsi3mU/FTyxw
s9RaR4vS10JVfujIAk4EwWDrxrCKKPPgi63d/3PrOgnF9Mi8ijBx4NYXfllV3JtsYGtSU4Oz96lF
J4SYU7sOP1c7fkvwrR5jRR5JfbHbK+bnzxDZcx7O2bMdpRiFzH/mmrEgPBnlJ1T4kifsNAcfOYKs
shiWuRQt1MoU5ueSUjTAxTrCzlIA/ub527YARmjbrtZyRnvmn9jNNJhn8lyOhXvPLil1QFg2EEua
cBYtSMBA8kDzOOSK69nq0tocsq7vBIIV/iY9Dlo0fIkWt5+MGKUtDvcacbtCI40LO8GPxQC7VtTU
p8EpzxiTS2PyLdau5ymSczCCXThLRxo6DsW1s3emZfuBvtXoG3E2QxYrDr35XTwXRuYWKLVbrdHx
Q3KyjlFiva+Z4Wa2x7YmnqN2Rnpl7TJyhNoKCxJJncAEXmON6HmX93n5L+9UTtU9A2VVGy4uo+HB
fIQhFHJ3n8K8xkZVrZ91zAs/HkC0xAvAV/TURNfB+g6l37MdH+gKVjFlGFpp4zgx2+I4M64TtLqq
SXtJNoTTPtgurgTo5cYwsVK0JCDKrKwKA1VOISkD6roXYO5i+lGrRT9k/AZe9GaExvJN0sFn7f/w
HL95c6lekKNAlNpT9wrwCBuTzF9rtRrpQ/sAQ8+cefpdKs7uEiTQdfuRVinU2T5m7t0/lQOCE2fL
Q69QbVxUfG14WY9xz7r9HGV6JI508fMPSZn0IdWXprQEeGdjv93diNgBpN0B3F2JSukXiTb++J5K
Jp14JtcrIEp9NshsFiN9RFrcFN7JzQH/LbKPlN8OCAu5qfwidcS6zYFHvf6FK0qVohFW1PLkCbda
TeABLiz9ZELF+9G8R7pSEPbMs9jXIJDffcz8A6iO00b08DobJ9bRgMrbf6oIAdAGK21ouASBjYGi
NJEI60MHLd949+ld+xM+c5TlrdUTLwigaPa4V5y1nljuy5SOMShYCXTUGeDLhQZdzgSSs9yOxGpD
/CClLlKCchYEq3IEZj7mRUL6o+k0j5QqGHK1kbwI/iAGJ89HG/Uu+BrwAue1S5ikSBpDZAh8/MLM
WyDjXApQYRuYc/TiDckUzuyVUGdo6tjmz9vQBiRRgHtPMfkqCV87UgurVALiO3barLRFnyPpfRWg
t3uGaDT5Lorzpiy6soFPWPAlXTmRoQix1FwpV154lAfPGYqfFAFQeY02b4kHL/rv81nFFZENcgRs
U5l0zAF/7AMPnNuUMM+l0rk//+3OKWvoEXLj9kMBW2KfRw77we0l2Xk8qrGp+z6mp6uYdSrKebLl
rCTygmllIEImk/JpGUcycjPawRs0Kft4svTPF6RiNvZ6vHURQpLtSKkn2lC6e5AXoVuoZwSztoEC
+BLLVPPGwh3PJNx+ruV4C4PFvMV7Ihid81XLEWIP6REudiKuiWngU5reS8UBKmwbSgSxNdSx+3Ed
AJBiGYlL7/r2+GMUyaO034vgSbDx2hP06l4W5jKDuMmAtetzHtsJ7/+D2FUtaVnq8sbv3N9QBVbP
DTIrGIH6LeOqEK0Mnpy/V2MkhGifA+/DvozIMfwAPvUFfG9Ld0RQ0lsRNKhL5hzY7snU+FimqaHa
+IZO6oVMU0LavSwwRAzNantPxfRtO15y5gAICiAZNotbKrLxYl9nUTVntEYIbOT5ApThuSuES8u6
UNvCT3tWk5m73TlNHHygDjX27NPtReS+vXfCks8XbGNogYB6lHRsSu4Ua+IyLg62eWOhefj2aw5Z
8raU+kO7uBz3frum4Bv3fGGwvBoPm07LkxllOVeZJ5McAwppPcs1z2lyoMCOBIuTevM4yE6HOD0P
kaOvqj120pIGqHQwV5u7EsDUDwCYyoO/b38sUr/fDbyOBtg4TNtwtME2JY1cJuYt92by0Y2ozv0d
wosp3NHr9ajo3qWofXHNwVc5620J4fezuhD3d+EizkE1Eo/4gmxA3d5qPOH1hdQBLYscAMtx79C6
jE/+IEDCsB3dDdKXG0sXr6mPMcPi2pqiI728JWcSsji03q3CQB5+A0qGl8iSxrkT0NwHYVHhj2hG
5jP2vGxyu1C36OUW1oiyXUKYWNTZ0dGdUtmPwlXg0u712PCmtKfojLFQ0+475i1sRUUIt+fqK0/v
0dKOabScEYPYDJyCgaNEPUX4cow7fSnK89ySZas+2YLOJzHtvLBE+7Wpz/Ue0g8fCpH5XclXj20I
sSyCKytuRKhf8/yLBZoNsfuvnViIXRlH2IQpByoPbMtIK7ln3cFYBJIhf47BTlecmIu51UkBequu
ZvqJJ5/IZe3ds/pzAX0zQfBRDW3wmy0UzHQdanHVYquZgOu3jNmPZVX6muhLE/jW6xY8/N8Je8iZ
x7nUzVhgaxgqLjs1IUQmfTjhc/4o0r0xDOMX4qSM2AyMYTt+oY3Y/4q6MDm02rdw+kULIc7oaMBF
jdklxVYGFPv+irQDwC4OY/3bfiJUrfXvMi7nRZXb7epoTYDG0b96Rhhk903CQV+jajXBhFsCRZ8b
ARdMW3d0GMKKzdi269nEr3ZPWmp/mY+3OT7JnBFMfpDBpXwCUL040a2BGWYUzkZllZmx4oWbxz85
SIg5doyZYw8/WYnsm+I7rneNuacWJjGBnKnMXyQVvP4mwrIXcz21dQLCwP9Ct6KT6NTegWhjvaIs
6cyv8rI1XWfk5Ql+wFrtTWiXLUOYZqbRx47TKTalXfcZzd/caBgBnb9aAPVTNZc/D+OAKSEt9+4C
JtcBV9KEEkBX+MArfWzjozKjvalGRAPxKCAkNheI9aXdBaUbfoE5pyTYvn0mhY8TZArYzzhLreo4
K0cgDUdT3xyh3XRES1XeYdUpBvYrBUNhU26bz2PZ3VaS/6dWwQ7MHsATalxPOiG820JPxXwwBUVP
sBwevzRnL/CbCcyV4XcqTrSU3+/wIyN0FmrB+Qud3ZljNnPM1zPrOd46EnbJ8806B7egSHy9WNyJ
4it7062/aNRv1IOhPTK4jSQpwz4scGonHSSV+8qXbtAesnWsP2+g3VYW5NazkCqM3vlpzZyZCyRo
rt94HPmdW/d2YMBCI964Z3iIZdKT8qiFYvlVb0q8e7voWwOLBqKkrg2UfbB9/eUTVZddqfh90fDf
S/NjhS17Ouv3VvoBXCu+IFv+JBciL60mIwNgEZtOBInZKhCZaO79S1YN6pKo212j3sM8qldCDIVa
z6uuX1/oarAf9ePrMFLr413ThGtpGvxsQa2+VXRyeana+MdhrYU1y5dt5ujkZeKQHhQDCsGObfjg
ZgZDGJ+uA95oLcwa9Alx1j/Jv9aJk1276eyZavqbk/nRmQSDgZUOfEcUXr0ge/HiTqM9h67j5SGX
uVGJznmqjojB1yPiIzwdPa9abSJfQimsCVFOSSigOmCXSHpQ11YTzvI6TwkGZ1vxyLGrAYTkdsZH
YRQLIHLUKrkdKR1mny0w6Mge1AW/wXO2dofcS38QZ9JSICZJOYJi7UsZSdveuEMbJ6a9IKeUNDVh
RIEWITzOjfXb1iuczgFJQ71L1BPM4F7Vmfs/pqb9gOsEfuwBc0c1FutMS18Lvu41xvcq/aw6B5wo
DJsXwaj4j8zL32kuvL8fgPnPFFhytPc8DTIqCMBRUHAqy+2P5NwPoNu9yZFQ7eu/0QPqrn17LQeB
+8Fos11A7pMtV2B2cw3y9p9N3I+wSm+KhrEvdqKphmkvMmWjfg/SE2FQUdiFJCRSMMkeCM6vfPe4
XZsBxA7+Kiw/Iql/sAWU1EQxaNHps4RDzlINhdctD2QfkWn/OhwPP39n9gWaPkresA6BzjHglxBH
rLMqYvPiiKkutJf5SaNy0RUJTJK9GW0UBfdd6p8eHuqu2bb2RqdJuiFVbGOcxfZfF0uA12lRhgUI
uHP/kav3gjpXXeyiRZ5TFM4DEFQUKdVsuhMumaM8WZtxccSmtA1rFbJf+4Jvp/DLo6W6xdDMw97J
IbVg1Xsvxb4f1NmCKwFBd7nT17BaSOfHtM2l3JylOyPW4PfpVmloIlpYxBOzrMGApFhQf8UkxbQp
tOP4xZM9eoBa+uazCgnHnGQORRKJQZmkcFSxRQ3BDFynRlesjOYulBxehHZ4eQN5x/HqyuzL+H59
WsI41SRn2FFoSbxdcbHTM6t7EfI5c7E2Cw6L/sFibu4zr7pw+kE1Rmq6oJl++wj0xhh4adE9Xugt
bdEckF8QpTLFUyORV3vgZ3grUZqHU6yj/sJlR9JUWhSJ/FdqN+t8Ycqf8AUIPD+BqA10hjbl9wVZ
PWhPI4UHaVFcl3zBTcXScwbgVGC3bvynxEhHe6GHbquV0MgSsFuTr6NLaOgtq8Si00FJVxxvrYJ7
UqZWBPeFB1y+3ZE84SuZXAx8zwIitlf43R7wVw6Utj2tizYwQ5iGEXwMMC+fGsHc87VG3J4uxses
byfiqN74odHKVNQARCaHUxm+uq/pDKKkUoq5surUOBTHxmARhYxpo9r9SAjbnQyz7A7k1yDrPiiT
TWc0fK9M39VLlYKuS7/u8qjmogrieQ7MblVV0R8GfRcxfsa0NiEKykP2gg9u0RRsd9yieqW0EhWB
fiShSLJKPAKrx/2q+Fqjt5X4JYTM8G4rBgoneOqfxwhOsJC8N2IWzVYknS050OqrRUz8IC2DUuty
YHKxunUHTHmZuJmm7K+iqp3vmH5uzmiwVVGSYpxK2KY6IlC2C/aIJyDbN4/n9FqdxpbiY2FKRAD3
WxWl+by5zQn+3YkND9TItSbPmA4CugRlO+nZQEha7/jMIusHAu1QDPLtSTNkIGiwFnfCg5VFcJCl
VbOH33G2mr7kFHHF6E9I3l2axcVSm3x+EFfQzYPnVWgLrMT1bOAjYPdH/FK8AHft2K2nIdcEnsVg
7WTaaIycHCI4jWAmNYCgp6AXTARxAODj7hRdjiT7IriUCJoysJaMa1ZyEOX0FdSJEkjSlyv9FaQV
6CITx/bb1yXc19YCITBskp81mwSzbTy4HZWhSVA8YtFmjsYYNSuLnHN9trMAOeKFZg7Hn8rZIECY
Ly8wbBjydA4qGlUYLncSWaNjeeSefTPE7TJhYirwpJiZnUae2Wt7vxsY8R/SEqwhIehwfTMnqCIz
byfY3CRdcwyYRe7YDSUhnAm+AY/isxy9Zu88I8n4zWkULdONDlfU5XTqC7np0eGa5lJwKonG/gl0
fxRK+niQCjyc7XjD2hwXl2XzgUBeqLvspkTFNA3bE/Ifa4in79uJlXhDCOZTisILyC2HaVjtSw7Y
PCwIA3pBVMlHBdeUa0ErxbDwkX0chODGfuknyHDsLs+MrIt4lAb5y77E0WL1Dgc8hVyuMJFQl55y
uw2YswGkRlQkl4cS8pxEjDh9dXRjEiieAAySQMe25JLj4a2THR4ZtFvmEUFFrN273vp1JpQQ3u9q
PoE4CxyRJDyxSVuX0Z6CASENTj16H8Vvau+KLmP8V/N/V/JPlInX82BbIoKvwDpWFjaMkPdotsxY
yxRRWM3UUOHnh/eZcdyo/WTXtwYDRfZsVfSrRzZdmaDT+8mL+Jr61D8cbvyR+RkPIHEPEvS2uK0f
frckBLdHnLoiDIw8t5KXiiefipYKevXrV0Fp+dLImU7ckxZdD2RLp+OMCZrHFkYYDMsH39RWMHL1
fBTD/JoHu1BylheDuDdfQW+eLTZp/XDLlNOmCu2CFW3nlW5sliM2Q1ijtfVG0z3+nM8YtcesdHZ6
NJ/ehfmiaIAae+k8W3tvtKNyamKTcljQet6JenYE7jmUxcpp+3GCRbUuqzYWF2zLzmHZFcGPJDix
eD7wTbG7/iOC9TUL2bx5iwGHPoooN2/PxuB0/OWI2noAbIpPT4+PN8o7QEOO0sib/avJVTrD6TWI
Z9ufqQs5Caz1bDAL6tRwv+t17eUeOotG2U8NrspkD1ce7O4enJzTA5sIJRbZa8ruOvJggyjdwxIv
F9D1v22Ryt4Hsh4WSSBOCqHN1JzxPAqeaKjbDkUu3YCJcj7QRC0NLcimw20fS/2Fu/adEbHQgILj
N+a7Cf3/bMAzaoYKQg2Cyq1kZhtWvQmhmBBfOwSvWA3RvDvcD4JS63QVSNAO9KEfQVpwK+L+ILFm
CJTGwlR5fJTnYdgCazq6lrIUWl7SaCglLPO7hmjS9mgJ6WKmoBnG144S9RrIwWrGYcQZKQK4CdKK
2Bqw7cnTMsg8+eB/K06+Pdn152GLZA2DLxro4dGa7NRoFTnZwAhstit4SpVsmqVEGQAQe4BNC4l+
U+R5whNmFWresL8Vdwr6kCFcKisuc4FBYjlEJQGuSJ+nmmse6NheNjbq5WYjjTVhqhrPx36Y4tsM
xfkbVo/f5ujBr72eNt77j5YL+c0vyp5JauNFMj82TDIDK8F4P/b5HxQ0wLT7LLPcMIN4fqd3eCCl
/6AhV0OmVEIT4V8TS0bnvD+cMYw0LkRyOZkW6uKY24ClTDHmPqGietmPuzMo1chrklSVVKYhapKs
bIM3ylFafdoXkteBDjMQHqkTqLn3Dt3N6Cd7CZt13JY/uTjiqz05gor71vS8ldae8n77mWQBuqTC
2pesRlYrqQGAjaXdl5NiAI4aMu6vXqke6wsYk7Mz9gzu85ETC2Cv/0bdox4WZ6o2Zig8GBea4hf+
M0KhkP8PSOkisltJ4IQdgo+W31QLPMrvLPv3pB6T4yQyG76Ph4bffvxyytDxQtaYdvP3NJ30xR8B
dReJHEROykRnl1lIbUsFKSByO2SM7ShEfxgIafgh5j/zIJe+cUe53kIjs0AZDH8A79GwM8m/TU+8
BcsQNPHAnsna7BYEvYR6TLvmS3b5wz+P1rlYFgkUW2kl44WfmaB4clTvfiN4iKTcZxhHaNuSlS1x
kyHYWoVap5TYgeQ795DYhP3uxggLXKgBjJBhU0O6ycqT7rRUkYy19sy4k4TcJoTMpkx3hqohHgtJ
LmeH4kbJJROBoxSsLYDS0IsQgNCrmA/bkZy+EI3wac6zNzVDkHfSAZPH6RNP7nee263B4pQo/UTC
4HLIPNlMWe/yXFYIN5l+LKXdM5HKRD8RQtNazBBmqZJwSYtLeH1CFz46n+U7Pzz9/abu8gL35QR3
FV1k/hMxM2gJhFyTqRkbWJ4do5KNiNgwXar5lR8S21qKW2pKeRhv5UT9LRHe11Kjj3rm5QKVlXCh
04P31OQYOl6OkaPhaNeo/YUsoR0jnHqUyXAo4xtonQYjxi0LOXQnKg3Oknja+GkyAPSM0mL/ejn5
nPYrOweccVvoj6dhNpWuZbWo1yujfktAbrNXEoLGNFXfGDt1vabI6S36VtXpdmdh153HksWH5SDL
KuiUVA/elLsWQ+nQQ5jVLWQyRWgbBnDKpygHnjlFedNcPWWiDVwtiIFc+1DxVdXnhM7vLXkCRqyg
YJQbDaWr4kg2CK9cZfbFcOgWTS0tXjgfqIRRRLtNgkkfJ9h0T1nsIkUwRyPgV5YfuhcEez2HD9wg
HnO7FRDMBa8E7Y+MiF0Jmx4+OLkwjLXgqWL1SkoT8thnzPK+owAfQGP14U1AUtQnxwYH32oSTRXf
za2JQQuUHkxrvay7x80ovZkjWupHymuhhOutkbyBvVLbcf+h4IpKJi81R3DDLvaUJCPstOqabDlh
pUWBTI7aw8xSnH1gWdSST2KJnpOyC/s02aRvvmdHG043yzLx8dPiKMLFAxu/472Y8r0ulQ8tFl2e
VnLI5QpZGLtYvZeQJeT2/mxk5siVxNYTWd+IKp7Mv5jr0ZAF2UEI+Zi4zOYw9Q2kxSCG/VOtWb0I
STwqMirKDKiwWExCXRxIRIuzmg3QLFljwpXJK37TqsodKXG7eNSZb8jiv9l8jx6+aTmz5Ye4okS0
c9/0rO3HZf+4YtyXiStxTg/hHlqrJNEJzcwMT1Gp9Qe4v5wnPp30UdlDIrE1XkmR7lUQFzNY374O
xTlAWlsclfer0BMfUIlHefRjASJR+BLopNaCHcHbAIgO/2IKKtSQXQRigVgqXGs0i5M4BN+W9qmy
kycttZEPScxAymZAKrPyexm9pl29LgvRfkrYXfQltVnpHBRgBuTJTcLXTn0F87mAlkHnlrZDq7lE
Jlp/z0KMFoAYMWS4/BCxvmO8WCA683GZCuDre2VA/Er+DGmIdn0rw7JfSb9gefGMsCz6ukZqOmkC
fEb9nAPvyfTkEdl8Xw3quprByVqZLaUtEld52xRlqsNzdpcpLYEZtaulFKguLpED/hIO25sN28yL
Q8iEAhvv1q5xwXRKqfHk/s+jIHWAW2NyAgOrwo+eePH6hh+CfueqQUBJoehx0gdUS0mtn2gk3gJj
gfEVM1s7NqcOvLeN/kByl3iF3ESaL7la67r1F74+ewbT0QucApEETTbTmVq0BvuqIBLlq3Urhiwq
GX9Fs2uHULzlqjhdA0uGJrTb5OQ6kwNgvemp5VmeE7ylLcI+23SdFpBuLVbJSbHhBTQHmSr1K4ty
CDkwTnMYd+E5MjKsUH1mGWlS5mXOOVc9E3noEij8OZWTn4YtJOeG2NLPfhZbrtFnukyqBL+yr4yQ
JeuyQ3aLFjRYU/Z4j0G5vudjTsiOnIooSQxx8j8aXN9otaZ6l8JGlLv36Vvnyj3J0galbzp2OifV
02bze2IrQAMcN3jx2a+LpdG6EGSEYzEuze4J9G/cMxXvL6599EE6MYQ1/wjrAiFiDOIAhqa49FfY
/0R6xmCjQ0U30Jk+7JZhTkZBVCD8JR1Mc9+1e/qp3Sf/m5EX0d7PzZ1Juy3L6Tq3u3fFPPlnltyy
Sb5t3jQM70ku1B7utW4n0zJT5SqBWOyiAljlp7WnMKpZs4TzssJQKKq1qnT0GvxXfOTqPS5ljLFq
OyP9+Er7zuGCAZsONh+DBDxioYmfmhwjxJ5yHX37z52wHbFFH7zKUWQGo644aNaIMf4OmaTEddqM
r7pysnYqJ6GfkBHeDFl1cQ3hAQkyP9fNjhut5Jsq3YhcxXpFwLYmht/L6Kn2KbkQGqbzuEvYWTQi
Jwvxd7UrqoHPZov06r8Sq+I6yrYjNhUpHLB8LwwipkJXzk8iy65S3xO4wnbyTMbhCuvEs4TBPIaM
jxgbKbL2PCvoY0AfDT2TPYB21IHYs8EamUcJLrfdk8wve/IBP9AvKfJ1umELepj1wG67lwJRu0VX
nEz0b8Yo2Po+XCIMLuVUGopP0kPpmovMDshC7jdhWLtUjlHE7EZV+CdLzXpnCEKF3MSWmt9SYeDE
g3R4OR+j3zkBxx9fe+m2y5k0oCsX8Jc5xVtfTiGSfn6hyg/fONgfeZPAkFZ/MIt4l+9gDMhrS/kf
QWRaCyXfDXZiY7SYVqbseTncb1FMyInE2CgG8vMZxX6GbgWom4uqAQHlkB4NxxPFdH5mnaSYAmzg
bFDT6cgvaNCAHFUw7YRXJ9onu9Lpu00alxNP3x07xz9A/vNeJHQIA+Zp1aEjsmu7eROUIosOuUl8
LjoV69A36U7Miz7VWah6eHB3XPaTPbzM6FwTNVrnZgbxX7OfKywg+ciyqC2tZ0xdl9bgOV2zZUx+
u7BPWwn9f63z1kKo/zwJ8ybUeRTFT1muQL+GsODHX6/476IUwyqNm4NMENi+6KFOWs+PJjW3yalX
xwSU2FasaZUjg8mhi1lJ2Ax7IUDBpVQRz/GAE2YYqKBi7hjSluuPZmU/hfmqWjNvL7hpb9KE5XOU
W1eyTRfkpERkS1Iza1uP7I1FZ2aopUOEoitneUGJtBqcwTyjq//A6PkatdzeLGQ3m0DOLHcT08AI
09QFq5fSRyu068rpleCvpPWMwXFFWqOOVb7vnSGaOIht/H+791mjJmK+PW26wBlKc5E12j8PaKA7
EPyeh/xgOuiWvyT4vRa16Orhrj7Uk0crP1kzA12PU9UNr69NVeS+ieXpxBjFL74V3DXsmZJ6JHqz
gZ0MflCueSuJCE8wqA35I4ulkph/GYfK/atUfaUPkhZLANSG/FIXe+zIsH5XYSlycSS5GxJvfAde
5fBugMBvA8CMusxW4nhTHv8P94244xLJcS/PTSE37x1l6/4AEE95lCbFk0g8IZWHc9VA0IWpUE1z
WUIl3NIAlTgn7ZWYW4OWWQGF4Bp+B79+ReQgaeP2ZWT4JN6xbJz3e1yD/uDxLmr0Q66OpRxFyz5E
DQQN11TB/FBqXcdQLIGNNmoVskGGFBN4qMEfeCOzEnCXcVlJ2ldcTDB/qsnrd86BVF3j53kQ4q7f
wBdxQKmPsx4NDVGqDmkM6tg+0LONW+g0blrsGB0VbbL3et+/+avMK3RGALRSKttVrdQCNpkJa14o
ePi6LzRPI9qMki9RyEI3kv8gi7yyHDruyAjyIuAEMIW/TbjCr0UWmWdpusIuEb2m2e0rhg7K7DKE
QbQ/YohKsasO+xae9jjxPlQEMBE7G8DK3I70+ym7VbX6x+ykxadBjAgTS4EI1G75VBd2J4R0KbIo
F1CI57DRTlVEiSAagqY5x8Fp2GNVnfAdD9TzmBNmqtoTEvDu1w+9Ck/c8DwQnLgynrDrILBiS1rH
MdP2rTWlC2KQjyFodp72QJzFB6e+omIbIpjiO+4Q2GKfvLFi+2C9GMXuNtjgjmn86v626h/+onU7
e/LrrBnj3em+E09yN8OFufFsztTdD3848l9BgbHYaTKK8SPjFsTVdxBU1Z0hLkLk450n9c/wHmZv
o1BlAaBfgqz4pi7vfSs84snUG6V7TKLIIMwhvHSi6MHueH8Ejuj7KsjWto6/TBG3dkS74rmHIxO7
t9WGjrS9WVKZq2KfaAAIGWSl3Vk3I2X0FBAJeE8XGXR+4qMlH2hgg8C296qleHXizxGKvUbIV3oH
xfSg+OAMeX5U+ddx8SrXdeo/+68UzQUCXIrsdrxKc5hz3vAr4ysYWDOM2ppEglzK/HiL0taMg7JQ
OEjif5LsgdQMw2PJ6Vl/nAWPjcCZ3f4rX40JkVczTbonwGDvP6Tm+ATWvpnOOyFMI/bHT98j0ZWi
SMLt6pyYLo/7h01Uv39+flhMhhKIjNIVEv3sCmI1BCHc7HMJbMBGQDZOMaeSpbNf2poNkW7cKxV9
5QqAD3SmQEyNU7hkRkvmRc5AlzGOpfvJvdXjvc1GTIHLJvQyR4J+0OAS4tEgelEwlB5aJ5olBMVz
mV8tURTKnXcTB/sMwo1fKFp5maplrRhrrcNcCk+lQ/ABZqA+R9bwIfFELC4OrRUGyZC7kTG7c9tn
qM+hjpu3VscUOTP9ii6bcFrPsjq0im/wrZotLQG2++9qlDlORH9cx9y6f1eDTunqplLjD5bej6Pk
kKt+YHEDB+/fqjq31DbWyZDx48mRfmbIxZ8YlW0nilK61xKB5h1eC5V3CnIerKs+xSzp5oknfWZd
CRMYez8HJnUdTcJ4zoCGaar/YrXlnupO7HJYXkcIORZ7MyrdFkK7xwTvDgron2Hmtrrb0hcZiViY
0ISYd+kaE2GQMXDv6+FDjmQb261r/y+iPHFGrfLPSErVQpYWSXalk8vp8VUf5kGrFcc81iOkG2oL
c6TXh1FYC4+dv/oU+WIB6zwSf015G7tr1eTPMKBycx4rPgxccS+NfDrGLVAnDU+HCutIa5CCZj5i
aLwv//zZewQPdjThjUcIQTL32UAEQenCV9eLWq6LvtE/EnVQyUTlYy7GZcofmdmd5urwpqNQxj+7
IvkVmArd9YzdYhd4J8hS4bJnr0pQHV7fxA3o5DTJGZIwa7oWOF1zTEy38ZLROi+boVyWIvk0+3N3
oUsMr4JJ7ad8Lsu52doayGJ3EpRHnpTlZ7oBmKopon0SjY1MhOJQkLFdbOcfh3kpItRL1JCJJuNu
XIMLHSwBS6fNRxUVHGe82nVqYxk7Q+HGjCtA6i3DuRZxnMjI2nK3/UBBnQHj+WikmtrbUZdexM7C
GgX+8sLGt3Y4jH7oSzEckYe+1cKLXPh/FeEU5c2Sfmp1Co2fywkBNWvbhZkPGwJmBgfOBtn853Nu
6GsBUrIHWFUIfNkp9MJiZAmyZTQYDQYyvPJXQg+24n6KC24PDU0/yOSfGgMWFmTZ5HuJbcXWrbrk
e4izGViPIH5EPQ95tAKKaSdDWhI2W0DmHSjJWalV8nta6zfBdheatP7e3Mwz9ilHoJJjcJzz5G8i
rC9IDbRyTjy36nkR8o7+dWMiVAYLQdY8bCkPmAsg1w7d3tRvNihfejBnOAQGwJOVmpgxDzhgtGNu
L6Nkwp+I/GikwPdDBupraRbe+ZqWKu0vlj/Jn0Bzv7ZgW2AEUdtfDB5x4Gv958OOQp1iwglM8Ocd
qftJlfYVbHWhcQoz18kdgx7Kb/IPMqVqO/0suXDRVs0dfv8ONo3zn62QA3WSGV3GjYVyseozCRbt
AwZB+/m8hSvCzihyCPCwg2niAJda2YY8IWpPvliiepjs00TycR96721Ak/ih834H2q+V1xS0MwKm
SDZVpF1pS9SAKxDyzfn/gHrNOoKgdCQxl0KqBDG3Myk3G1tNMfTfyko19YTOgDtT5bTeBjRe7u6l
AgIQtM4ZJKzQHgrUiPl4umAITBxDIbzD7KN0xxEF9Cze8n5xTs6ZBKSsDFwMoK7Zr2WiNXglZh7X
jnetdJNpknJfmqqF1rGDZptJ7JD2TRHmOdgHFcqdU8alqOLbuubAT/k5x5/r2CPUVIf78+ptCM/I
3nwLvq+O3bufrednYxwYLAmEWmGxSVpS6tMorrvuQu7mNl0WihR7ymZrYg//ga3s+3Cb2WawSGmc
CXgbKYEsrJBz7GlBf8DIhwmnMYHHp71doPI/Mcc9vCCCf8ux7SLEX44w+viuVtqmE+y7SvIfzrpp
IjIFNoMRdzzs1YWrmtD2UI1MVnRWMYkgsMOcElkNlnA8Vs7z/NKSoIR01/CFEcilBe6czTsrkJUN
BHa5hSV0rZJ0VyeMgpKlDkdugoNZcYWHS0Nt/DsMQ85ogSbokH0A8Qfm6QUDQtrT1ovUWdH4kMze
WJqImFsL67jTas2jKywF8Q9WWPmTYMn95YeMLa+yiey13EsbvI+Iay3+E56KfutNOn4ULQZ3wWee
2baBwQu/VyJ2UZ3LHZ2k9bZIYwtiCAkj0AJXmxk5zeAyOyfDCKyhOU99TAMc4V/r5KksQLkDc+UX
CzEWGH0AZ4J0un8FW1SCJNlBMOnom2p95ICZdu125veIhw+ke5udQGPg9wilxWC0s4BH3Et0cQt4
Oyiqvs/qlRc3D8H4yo6lfxMXH8M3/oHgiEULfcjmGBHLT+czkcnrxz/oLOAkJC+gQ//B5viqnrbn
z9d5Z61LQ5MQ5wpXL7VltoMjNd4hGIp37FMGGqFE+qpT/oZBmzMysrtqYVaK3lnOWfukO8+v+jrc
XF9wQp2krtm0TlDMGy2AXZjGdMGC9DJPwnSUadsVfhwHumJg7hdP4xIF574etwK5WNQktKT8rXkF
H5x+gjhvu9Q1G3t6uQpjZ2PS5vGh8tJLFTXk6BJu9uIMZc5wE0yC0ODOPJU7GMliD7+YbXXJjQZN
bXhBUKUsX3HLCS7mdsvLH65RRYJALeYil4SpiCSqv5WfZxGk6oNlLnfya5YQgrdfSsMaGHrBBBau
Z0X5EFGJiXjTESirB2LP2lO4qG/9nr0Z1QVf4q2Gi+vmB6kdO24gzwOTQbJVxEZz4pjhtPdTLZ4b
KU4xmoUUQa280NHw0Oc+Z+e4wxMt8RKsVH5iJZ6RW4qBge8DXJ4OlE2fqmFrmbppdM1Kt7KJ2sca
U/zsE1LjRrNHu0hqd3LABXYhtmcoIoaPaGUzdCSu2Ow+meZlmUEki5zK8G7xgEVEe7LV3SSXM/8e
Dy+ucGaJllvnLVvRf1kMkqkBnD8Mp899uKGrOheem4FpvkGhgCIqDcE4pz00XtogqEhcpkzUDxP8
ZTXIPgLwqKqHZBWJcXG3p8Qm44sDSjKUPPdIXWOMDJ4hYHesaiWbbUScvZFrShSVBMioyxp3eyR3
DgwklH1cyj4Z9MwpCye1kBGGyA0Sb0pNd2hBTvCUGs5hVoMwavy/E97ss+OXDQzUPyaCNqiNeA+m
fFQQH+UDQc4yRUyQAgW0OgtYsZ/4HcytQ706VKDepuz21eMvQhMK0PairNG7TmRyVI505aFhCAzQ
urQ+ANfjNYrVOae4Knd/D+5XVb68cRo6/Ahb9Zbt9OkwlLhA/VBBvkWKMfJdMefxAuq3ljY2L5h4
ADzD8UwhKmxmcuLncfQlT2yFoIF3Mk3yDZL79b9umgMMX4H147jRlunOP8zVGsVVZPjwv/q3ehvu
2exegOJiPqPmhjJUJqLTeSFdApgC6hWpl16vdazGr24uoYDUtptnj8jr+HU1CIF/FKSUiduhRMe3
RQInJyUb1YytCliTGoqZaEgS6CBikNmAF+nn0WE7qy2cxTdTBzuxGEcOw4WO89XdAyGcTEFCCsEo
zV9pVTl3hk4f+ON9Y3W7xUPQVuYi9ZdPOi5iFab/GS0Y1rOR7qv2+h1QPexCL3ccelY603e+elNn
EbtzDpL/vm2YPD+Lt+RjiUHD9JvTIkD829qY+9a69RxQBRAnJDE9ScYCR2IBmxyGNJ1ZZ2x+K5+6
Bvt3oguYRKgBdEJBxrBDcoeLcBintmIzan7yHyOWuFoQdw6U4priEFeyGqK+3K4Cnm9m8bmql3eH
3sDjKxy9EQ7rp+mdlrR/XyueKWp4mr/Wp+2bagYjmTiTMHjPmLi84JFzhWCdNfG5o6EgpEu56tVC
oto8l1BRJ1bfU7oIkMSIzcPi5tW0a5v8KmUijNkWphfO2FMVKKon4DpwX+qI5dbqjkuii14P3YIG
3J6AtmbRE/CuLsNr57Wxw+gTa3q3SqrOQMUGFuCLqbnZgpYR427GeAaiEJxB3nVMQ2bJLWdqN/jc
CmY95SI/nIdhbFi9ERIz2RCBSMQzW7V7EVxK7VybQ3CxjVShAFi5ffG0HQMG33e+odPaR4fQuPoa
UKxhNhHn4bPBxSlrRnyR48lSmuKS2WGiRQIMbC1Orax4E9Yl70wsUUM4UUFGXbyh+54/LjxhAKAo
ocLN9k+MKctoyuVK45S10p05/SQFV1cymGMDhgYpnPU1pfLYLBgJgzl0pt/682ZlqOHL67wK1Rmn
FLB6QGlhgL7vYqmswOrq4y+VFB8S2v8YL09jUx8yqG39OESeO8XLuI9kgsXDQ+wY7HElzq5You8o
RzmVqXKtlAnlz5iikrjFB4rA34iyZUZgLKF1L6LAsfMeOHVTBdL7AWf17A06I5EfgVXNeVqjHhtY
j3pgXqKCB5GQbvFbwbAAGQ7obL4VsMouNuc3PHzg7fl0tWgOtZydwcGU5DAgLBg+E9Y1VlHxLhq6
dnBtb4Y+k6sJlC+CfY+mUBa5RKtz9QQF4xsPlCOdCC2+ehEwVLvNvmhbgM6YboOLksrQTN3AhsOT
mioRUbIQ9Rb3Q2mh7YYSEmRbTozZReTNsbSmj9Qyrc/PkmYD98nhpeL6N7dDqSMmX2454Uyo+pfy
tDo1Og6y9qBuK6b1PXTrH/JnbKbsuOEJ3n2MxUkheFeUBH0P97AIhw2tg14kbIQ2DWEQcQJ60DJe
4e7iijpBjE4J/dqLbhAWOC9fB51mf74C3pSDqP7KyROicfbKEWIW3oBlpJANXS/2JoAPhCAd0O29
iLXS4J/OBau4PTDMs5CKJacVt8x0RXFF/RRfXHoPCWSeBlQzQwxwb+BahF3FDQcJW9hIWYbTmteW
IiIrZE5HmGDKp1DgnKty0i5feEU07ZeRM0ERoy8QjCwvx8tE+ZEqFyHJmbx5q7BDVVVjDxqoqe31
zZFaxzLm+A93mL9ZqYUqR51dSsytexZ5CJXdwccPzLzwwE3UbrBdWerLuRmSkML32USkkNBZ6khh
uO6vwhowNlQ2npqB27sqJvVSKQ7FdLxOO7X3rAqowDFBwBkKkaGINf4C14QUYgcGTU715wMa7egB
n1kIMC4s+ERpz/1GGr6WP7yAZxIcw/rAd4rLJUIwNE8ryvZfKs7mzAO24o8uqBYJmgHT+2rG5rOy
Md6qLeMjkBpTn0JxZKqLzlL19lauB7YR3c3fk3jmVpugFtkuZR1rJqBr93gKlyymvUkAXl63w7pE
/hBK7IQzPV+1elrg2mDmpzWPZfRZ1Ls6npudPX1KKKDDm/kVinzpWDTEf8hqYudrY1FcPSMDFxKg
SSKuzsCFa8Y4t37nWkvv01J1gEaRnwEe/gT/QJiwB/mzZzvGfHmbROud27SfBSI3M3LqepCckYi9
S+xbRKEmvjqOplKNr3bT4ctxwveHjczcomOmd6ZknDySZrSYxgtr+n4S3GsW13O0hcx0K49wcr+n
OjEORW9wH8mFIpCbfroBVE3rHdtOLO7zPuGn0/Qbtez1C38LmBJSJ6ua6iGj5I4YuUV/YizKP/cw
j85NTDkJw5zmpsdxBFws6OtKTUxWnGytOF0iH65i2BR9Sik1MRs7ok1g85mJteJJd8wrVfW0FW8/
nUzsx7pXRFh62RTxZPHPj04dSgr0WAZ3oBII2WK9i8FTgsKJyIrworo9RbDGF94j2M/fTDHYmqFZ
eLkUXDxSksIlrIaGC8NGe++HyJ9dIEpZv26KH/7rOntQetMWEIgf0Um/M9/y/eAt0bih8DPjuoFy
E+FcpVNVbJdWfHfizNHGigpzv4bQT3oig1JYmkB9xBQYQeUGNNvJvRUh2Vz+1zv1B2Kcx5o3s+Iv
GsYpX8yGD+KE0mTh0YqhccFEF+t6wP6NCTJmMauIIug224/v/AhkloL9hyOF4zX286jgP0fnaZPi
QT3c06lvCwcXjgn1a12mciibl5kQpVUDatUxuXgqSvns7hZlgI00QBD2MoEv7Uxn2yOQxeeIDXC7
pw/lx2quAAQ4Q+tLFNObOuOey9ymmEufOSDVr4UXVTSqpU/MX2QtyvWL93c8Aw8te50vm9YJIn94
ukaIt9w5hyZBv9E0EZa9UJRRjuiwQJxUmry5hByCjH7r1osauZpBJkeoM8FXlYEL1FyPBfh095g3
/K4PUv+a/+venRwEW5d9D+m+Osxpvf2hdwxtA7FlmKlizXWrAP9NLWFhmxAcI3LMcEIYmROHfAOC
0K7irwMxkEQnNafZgfNov4HxWX1FLQprldLf8VFISvOOI90GGwYabgUEsWpMCA0Du90o1G3JPFg6
8leCJ3PGCe5CARBVMPycOQyxMmsOiZyq0agXs+3XUYlwxcfNYSeJviC81pBxZcmHsrMlq2d6xKhZ
b5JNdydeTMGfBSX2/MJ3XPNCwoZV7pqyS6GYQkW21nDtJrR2zyx3HLpd964xhqYkNtFfi5wEMvgv
tMdktIBFQPs610ys0U1HHnbjYQxQyW7JD+dHmeO+Rr2I3wqaBJO0Qxrhcw5xN65pvqeMA4Z7XvS/
rR+wnEU9dNkVrGzz/9ETLivVUyf5yxwYs1qB5r7G32tFZQOW0o0Br6R8pefBuq7BKK0kz11v0SFq
aA/pwbrteT6X/pyEtp2H+N/8P4afRSuwVQfMlYtLf53/W7h5lw0YkPQju7gQrwLCE7jNrBajXWke
an7OffpUZn496kMk+gGNeFmZShxOGAxRyJ1g5X7CM6+XwQdW5rOA3JUVZ9E5TwimqAAEJcl9VnXs
46b71JdSMY+6zL4Aue/Fgq0vztxk0udsh/x3DLt+9aQSduI6DeGo2V2OheBi+lAPvJzvSYdhs7NK
9R9yVLtT/UNe1beq/9v5uxAok7MI5HV+ekOfgOIQZPmkJ5TLKbLW0h2vnM24P4rAasIoGA2/XUc6
ebzhKPdcP48X/41WOUc69rVbQ9ANfHtJ9i2SdOzi+Blf7vEqHRx87FxtOUZ9O258oxCfuHVDxY8d
yu4goygsBdMji+t40FpB1JAiOPDv4cnTq0O0q+u+z2ozLrnN7T491Uo2tlkPLbPFLtuxwDA1hnaJ
1o8F8zv4QmKBNMn+XJziZId/4qFPzgFjVIA69+um3astPtqg2EfNjlauqj2eafXm/GKWKEt4isrz
aZs7gC4Zs5U1iPK3PaYmWrtDKfC1e9GJ9iSLMYT+4LocMHGw1QFq8tj8xf+OcLeXO7xpDrLCyc+E
slRvevH5GsthicYFFK2vsj792pJpJeI9qKCo0d72YqArZef3ekmLdUE/cQS105aFuznRhZBsf1qQ
Wz7EnJTlEjV7ZYuheKM2cOS8LEiiVKGbGPApWIT80XmBTn9MOtz+Cd/bZzsBlGY5HIpaeRTwdPCz
j7/SA4lXiKoKagSNmsCaJbFqL6Qs5FibAgawK3TTifyWjoC4OOoE0O8A/LfXWHpUlbm5rc99naZZ
5FCuxVhxSYxdV6dUxsasgWFUC53qDmJUWaiUuh0a3MxoZ8VxoRyGUdAfni2+1HCwCog6SIazcIxL
mxktYnaPuvJ3UMNiN05G66r0ig2KD2vHb+EG1pFgpPr9GPjWwc75Qm8UNQyGLjcfaGMLV4hCmz33
ALGyw01eQ4bbQbDPcfLHJPPNaOl3CfAf8yK6tdJXJ8r6ROP8XGfubOsaTzENEHOzX45nj9lNoGYt
xqJFS6ZuhKFCN+vMncm3kJCw1RYZ4zqbElaqtQi1K/VHlgcP3ruFwhg/i2DlWgr+GxbpqSSguSKy
ZL9cc4ne2XQR6Y97iiDFujaVgaCW2U4+MPbjJF/j8EOuqpou827Q1ijQGUv59ARahVgcRraExw2m
R0z9gLokmL/x7UzV+sloO3UY3d97wkDl8IH9BlpjwXSHFgMBZYgdT7ICkWjeSCTP00WtMTlTAs7v
viZ9+tLv1T3V3QUY/AGuf7fZS+MVEM1ZgkytaZiR05sZBVOms/r4pLxszmHVaxwzlEuDWNbeI4qQ
FdsLKdG2OepEjyvGKRK24tNmG0D8FvR56Nt0La/uLYByLGsbZz9pYyQEa6/pYoAUernxT0nXmIMr
rwaGP3Cv0bfbCNRgK+A2x/27vKsvYzERu0FJcSEnD8J4e8qllHYFj8ffZtsCZKefH14X0vsuFdiI
JmvGQSBPUgUguINHGUcapjSa+kjr33bhwdIDOads6WR/vOIKfkDwfqVaZFqlHnj9XPuP/GkUq8Om
hu9PGdaId4Y8E+yX/T8YJJA7ByG5h8525QKslvvOGWWhw331l4/HH53RqirO4Ag2ZPxqzXcyWdh2
aXL/15zTEoxdOSGnVb92jdUeTe3HUTMoZ/EbCQX0H34vqHkp0yiodcTZQl1bGvql6L4H3RfxIroq
L/YuFMb43dLaGnb9wdrt7YcStbMf2c5su9UtXxKUv4IW29PH+v4y1ZLtyDeVY1Qwew3SklVvcuUV
dNoy7mOKt939kW/5/TtBogowkqOCCJjhKW0rmZWAyu76u8ljDhUuUD/xK2iI3SEp30vPuI1pFwTC
2MRfX5vZoJ1Js0CrRKVP67xutHD6Tv/15mae20VeId7fplFu95qPRAsLfH68X4Um59tkdTCMwqjK
H8Wis8phgapiUslgzxW37jM6CJ4uGAp0nsERuI+xNyHHGLIjq90W4mdovuykNib/mIER/f/DJOQD
a+NEWju4hN9S8NvIy7nCklgfQr1czdptidt/u6y4pcgKQs/LHx7J7AA6AkX6Tm+i8l3Ieuo7Sz3D
TYOZEtfNo4Ui6laRxuszvs+otLDBLuZ2N/1oyz5t01ap2KXYJwjlEedoCuF9XHkLSCNMInWgx3uW
+Js2lzFQifRGvmoji4aByvNhRT3m13P8QZlOjRULjskyyfLQdXEuKfF+60CTtjr/SNzRC7vEFRji
DlVM4tw14tVEa1rUi9PQL3gtjHmfcvfRJLVXvX4mpihkFkkciIIbzfSJg3xgx8C9Pq+G2k3EvdcP
GVDvrTwCWP/iDWKUxkwSTwX4fsdmnrtSlwac3LCXdw+NvdKXHLJJnfPbZex/QWTkPyofku2iP55B
eovobxXh+PWfWOpiu3h6VXqShpFXkujj9SkBwL518zBODdKFlZvqMQMrCa/kOO+A7WYXkJRhgTRl
LqYGnh6CBISCFgOAxrVpQbp29hBkgtCXVnzhFJBgjPoN9Nl+GZOeGw67mCsF4T0O8Qh4g9NZXJF2
uVjgbdgMtcjFkPiVahyC9duratPwmY2ofE+KTnspZoSYgwQLtC+lt9D8OAyMSSUrzHydnv8OQzkO
TJYPb8ILu9RcmeloY6PSZhMWSmyM3TKm0tBDgfeHg3UdAXEvnuTOo8Pie+5m/FJB021kBcqrBOxS
YfRofpG2cShTYPPLoPR1cWrMnYRfjwawHZ9t7pc2703KiSYJPoff7Vv5IKypn8vGQKBJq7Pi5/E7
nOEa0wm3aLz24Mc4JR6vK842bmXfrmMEyg82v97rdyzUm3l31lbkMvmDFy+WXkthZFXaNAPbvQ+v
ChQNAfBucwKAse1J3eNLSZ1Z+dLyP/i3hLwshBy8Lr/8OfToELu+y+EyPJDqCekLm/C6iNzxe6LS
3tzbtJCexL+0CjgsJrr8lDYGW6XdUxZiMT9n+OebNBlnXt3GRKiNNx2XfP0GE+hU/Z5onTaUuLrM
PmPdNfaoOObaUOUdrWx5+VCfpF/41NFGddfQ6NYRsYSEZDdQrE+E1T0gE2KdSkzLhFkSXLe6TUXN
hCefl1T8bledpn8w+p/Is5EcrVDEbyAKNN14oAdkafakJ7cPbOk5YQ6LQ+v5QbCyoKX4DOFmlLjO
SHKFkJCBGY5ok26M8dVJrFL54B9jELSnispPELbtZtEZkjGbMmX6KZYrsMozNCdnrPQV7whf5l/N
u7O1quR6GGC6PBrz4XBRnUdDhxuf52WP4G/1ke+afa5JotC7Lw4HuOqFRHbsWUEq8qMxsyG58hOD
eehvCarmbPW94uWtCJo2D4yBv/g3LeHOgvJt3rh9kUFpvYr9LyKjKaxZWV9yUjlg/ha+Kcg7klzX
c6f41KxDOy2fzZAVODQ83MkyWUeo+X+RS+8jz3A80PCMjP4DGV1F8hRAf3+XzZVFYtjc0A7SMlQ5
tkVvNWsbzRG27wyB1cUFWsN3F9Q7hFhZSjkJVps2uk4MGrMN9KyuU/M5944IOVH0uGZMr5k51T2s
M0zlyjdvx/sUwL6z+QeVGzIKQo3LNwdsvNVhqXddQHSFKhy3mSCYHJv2hQKjYfAn102zgwqHiLff
SM7Fqug8S/EENeg3fZh597pS0CDq2eDlXpoSqO0JmsKzB1DCNJ4iYvqHdk31I91FNnkACLBpQF2h
rChDcFQAww/Brs/0MjFUSmAoT3l89nQ2j4W9yCCRReCAIKm74/Xq8yswtaRHwYTVKtnTafJBWmWw
yAnTi5W/oz8M4LDRqtfBADQHxl+mhzSjrTxdsX6Bq3CeLG34cbLIm+O6ruVhp6UNhw7QsOgWlc/9
eGP9e9tx/Qnjv581aLTvDPjtiiPjq19KDe5cfs4ih93tnIaphu/ZaB/AVtq11RLywi15mwWDACMf
AsNzcfeC0ryWd9YkBWwzeHqai5uelNJw95KAtmjwfSzU12FuJ5GX9m83CciB1zvLepKW1Ja1OV6i
yRC2RzoVnZGWRhA52gThfPMj0rzdTzga5UoE/RrGDjYpa6kMYk5Vil96I4BTNLeyvPHQR/iR/7/s
Cznr/p5TG4DshuF+mzRY4XweFlJHWizfnSvNFPC/9a/Iev0o539KKy6rBxLWqLoz493ynTCajA4U
wUKXqXd+YCoJaFanGmSN/i1pYCHVDRR7u/2fya7In9OAh/qetsjc1s13uwZm/QYWZ5gm3D7V2pVD
AHRYMRXsUAWXolGPpYubNQsJkaW32PxX5YrDOwRcKdMqfDXUGDo6MF90Tl8VpGcbQmB0dUKiRRHh
RBM78WZDclYOsckjmpe0bG9AHSBjkUOGC1/pa1OJG18u0iuS7ks9ZcHJvwizamkQ/LvZtf2zUnhV
U4eh0x84B9qqcuy+YCaHbtQTAXjO1f0NoxCk+wTDrVRBck20ljFKi9qdn3/gjcU3ysewdDGzre4a
khtcWCvX21EsJPbGkC4APipfvmlPjRk7SF+0fnfg2kilC78vBpm8c5DzbP3jnQf2gaw23orveyqP
4b7x/thkjOOR78O9onOU4EEtRFBg4f76xSlN+LAUtsBeINg8P99FjdZtIlcSYtSIwmZ14FzkhMFY
1K7fZao3WmkEKpahrdYgDexYbsxyvBdvui8zdOKJH19RJtebDBo0/BEp97VfEIDDXZPerXKBxutb
pHHfsEP3DXJn8iADa9U4lv4bXyrVuxjkP3lwIaukqlukWaxXe6A7+TahqOiE+jIMc4nRogsEQziZ
YcHlzy8tm1v0WwuRX0Z9WIbXCJNlCuzpp4FZnG2e7S2rpjsF1xRhEh/wCx9KVkKWWrbDHGBMYPvf
XZNGZO2d91XFrvrh4u1lUv1Kgg6Kc51kIR/ar9l/Cmarhrd24MpHE4G+2kgbQ1mWrs/Mvl2LwOxG
Bdvp/VOR1tY9knIIlDZ6ngpBkbWqPLWYztUk+3UswRoyjPHKto6ZIz5Icino5O/tfS7Bk3aeB6bM
Q5Jh/w2GWGW7gSxsU4RTx4Gmf3PeEyTWNYum3XNm6zwEY2XUTQ+4F8HBFttAE63jk7cv/nTBlq+e
0vN/DTh5rpItOeGJJmna+PyKuHVmGRRmXLkzt9vonLIji+tg+ZZb6o3wbNWVCFocP0HFtxXV4+ly
qXww+Aqsbdkid5VL+CvCp8AO2daJvQkys8WBDCdioW0mSLAh0WZPGnCTKiBVsYkqQVk0CcS8PhCJ
0JvbTvnIR8vbEthwdorNkf55Q/XxFfMciQoY5h+7HuKAHnAye/QT+O/CsDdxidTSrK6GISt+4rZZ
TxzhzO8gKxkXDemyx1FRgMKXGKD8MKnFmxGejlW9ieK217uTkfqoKdBRBRCdyiFCmrTN09sIzWQq
UL477mvlJ0xvHkZJnKXAuv3TobxDg7Cfxs1932uD9Fsu6zaRE5/My27Yji/dKWwab8SckjxbbQKC
Q4FQ1zvBiHKcaIwB8liKBBmOpHlkvlczNXxANF7w8n87PhdFmU1Oia9q5466tAmmNyc37wz7HmYx
HKKvh2zPo1bkfCC3aD9eLPiVoStLMcaXjb8jPceBjCcYcM2O6qDyhCYCtV8g8uTJlgs7ABlg2dQk
HKQaLsiKhQM614jac0UL3moccxT9mTayiIt5Zc8FoEZuk8FCzG8vZf8CFk6cVkC3nX0ZlZcbN8//
8sgya9qpbHT0M/J12Hiyw5dPYSh7OZlEtNOvYq3x9Od8IQ3oLEz4vBC99EPlWi6nDdJ+rUftNwxF
is/s8+plSfK5aQU0GKxqZsbYs1DK8XP4mIUNajIIPpEJZ3gwgCBJw0kCXG7LQRYR+4950ms05upJ
J3Ur++C4WYq3U7twR6qxT70kt2YOJsltDu3AXqtpMN7ih6Lk5pTtaS15Ct3rmO0cbLFO/vP/Ww13
q69TV3+OJaOxwPDyJP9WKuX8ZfHaVU4DcEjzRmUrqNbVvboNz7TRidypB9un0X6G/1yYfdtZlSHI
4SUdEn4pGXJ4eXpCU64/R8rgE77o9zHPmvOahkRz/B5ykF093RshtytyKSn5U4DYCEqoYFuUZpsH
hgRKCNJYe05b2h+aFAYZEeY66mOdLtp0WmgZFu6vDUr/A2We/g7sptJyfCHpqpyAi8gsMJNoCaYO
lcEJYIPW8Hb22rgYYFQfyMbuOejYob8q6J3KKnvJs9w1MdAg/nBfIb+5jGkw5Dhu4qfaj1gxYo70
aSj9t8a38+iQ4PHcf/1zQApFkCmDzBw6jGNHiXvHzDGP5cERaGDJzGj4k2tv57LBImPi9acIba6F
ltQAfABjWiY+vnOxxcN4PnDkvDg7yVVFI4teMSniIrvLwpGE5FkrD/TqMAkHHa0IhycIPSJtOIxA
/Zi/VP2Kd1aJi2yg3Y2Ht4Cg13Ddw+3BIBt40nQN5g1wjekR6jdmRymYy4IkWn/pycuHHJ2rKmFC
zJ/WPw8YyXWYy06pt8P3iEoCB/oNCy8e0CT4OuxP9+y6pCaRPwC8MtUoW9QRE31+McKVklrYzyl6
v/+NEOhfZsbuS8FuAnrefkTGZUOhCLw9Mq8U2UiXSFpNV8tvFFRYWR2BQ8qYWlNQ9ZBEBkuzktAB
K325rFE5LxuHbov3MMoJ8RLiwasVzWxUV0ujsiK67Xk1zcJhAFLz/wtJoxA30mrqlAD9Pngj2FyT
KRqfhGEioi/rwPamsfCtn6WZOyTY9k6UYTDvQfHSkqyy1yIk79TXbnnOYXL0hWgkrCmDJwWmQfF6
syOa5fPb7k9in6GrwRKpSgGPaCIbDFjwaWcL/N9HT2fZjvz6eNIkM+FlVRw6lpMGBE203uQ5kQGr
4vf/mu1VmxPtHDrblkXFteSX8vPw0IYPArmGw5gFADhAvHE0xALRMvTRV/SfB1bx+f4x1+u8W6IN
roMTMkj1ZicAGas+rM/zrydffpKsSaiF24sICkbi/zb/Uag9d0ir5hMyZNYuDqzV65Szf6YWMIDG
0Rmqg39pzecjjjEEUewQrQdVQnA7SmlQtEHmgRWz6vv648BlwJp3H3rRczLPFNCiFRTYQyned8O9
8cX9x7v4IPyfJmDkLo7fJOxzbXyULDwO6M1Ab3nHLtPihmv/axICZuwx8I0bgyeO0Q4bUsTR77mz
zPrDQT3g2eyMBPziVqdE7ErIWN2FjIbt6WqpBmWe5pB4DHZU2EsgCRHNtvRFcsG3k/JRumTpSGlr
U4S/9EloxI1wYytMfgBu3H8tk3yPO/1DZ7ZGawXrRd3zfCjw++O75fIkV6MnU3RCc+/8tzVw40M4
JOH7u+UqhGUpjRdyrNwiG1ctTi9lAKGL3XQ1QpB7PvHFgQKDnp0EQf5r1jqKCPOZ2/1a85jL67+X
PI3+jmc0TP5U5btz9SifFBfs2YkedLh69/9TLtpDmpBwQMBftqA3Cc2BZPHnHj1NzWVncBQ8n611
zWUqol40o5qczajWn8SKIQMP281T/qFasqCCfusPfAGES8Qi7wycTi1d/6PaZOljV+43k5JV5lUi
4iMT+rDqbvm/1UgMGsIqk7y+uGISUjNKKMPOq6WFDF1euz0XZQoxPSDq9kMdmaCZR4i+ouwFpYtR
ofCNxI3uOdgRUwNiXUPoR048V0/F5rnOn87OGke4kPFU8V+6mFOhvWeu6HUH5G3vrB3joXQZ/fH+
jNl1OSktQ5jZ//1PTBG2gDEM8n9tdEv+ju2GkVW8H9s6SFWh3E7XongHQK/smZrSi8N31JW2xaTZ
wFtG/3vhjW6EYovqvzDSNDqLYihV+lrXlDyr4ClFCWAgQM9b+CDGyPDQg4B1ljK/T4CY2fn1RKqt
hxIw3JHrgs1pEs67q8ptUGWz92cTIcJslEMWykwXutRZ2Z97AcQxhllNGsnxErft9IdbzsHZC5aJ
Xd68U5Lrxmfl4P0GcgjBOG2xsNKKf75Jl9kBRGBmyEqWxutvCk/vwBqEmTyQl22Taqs8iDFrvkGT
DxDEQCVMs7xpHib/Gk6RPiFC85Gf2H5MaBnc85cuGQ3kIC/sBD/RrnH79TEaGElcI4EI9vL0aghJ
8pQxSUGnk+O7ArSXITZuWZ6KZf5QFddlIfWI9YnNrvCGYrwvUkc7k2Qw5okBeaQu9lQC4pdKliPf
Bq2kqRL+0Y289YJrVmbgZEOKOOQ/aQ+SutP7zYjUFFrQ7Xtja13MLcU+lA1WQImXk2bOw5qqLVyO
1xIOsF2d6B/xubPlIAU2X8vf3pLyX0aC9MzWJIECrxVsHg/i/wUO3ridM/tVpoWC1hwdVJmq+pZr
QEzJEmU4SDdE191jGO5iXIDgBotxMkbPTOqt9Bv4VaIpY/MS3UFIU7vd+lZO55wAZra3VmnMoYX9
b1FCzQmQy22OBlR1uuLtqFUszIyWrja44jH3ceU74dB/U8f1dCcMBIlPXJ5rprLrB4qphSyASAmQ
4rv6YAW+Y8S4Urvc1urXimSPROdcNPb/j5Ejb+mp06tuOy9MTUOza9ALvy5VQzeVHRkqhOn/ESs5
Dy+7A7yXF5BvOg7Rt7hPh0uoqqMfAXwG8tyiEs8s3cpix7wZR8yofDwy0f9I0U2zsDcMrh8+/iYn
BWbHS2F+G8BuzrwiAopkYV9w9upH/Jq8ccr0WFkU7r+nNT/tKG45RMiBoik4jRPNDSh/Oho+j9Pi
IH8OCDyVrnVSxk2/jfRxo7s5hVjcgTIFzr7XYvQNErpIKb0YNF8c4/u9Fanvya/iZEYLnz0Hg6Sd
1DtHSnhp4nc8CYNtzWjB640hWUPJqq1AbvXw3KiHh4vA3npUOB9L0362FFUobaibGAtEi8+rHj7z
M2qkGNutqUw171L7CN+p8zO4ylnlKddn3daoBiF754IJqeBxSsq2LCFj4mC/pjPfihBTbj7N/giC
pTMrwJDhHREiFKjONEDzdws/crKWqQ2uw7CZBeIgwHx6joCoMsIDKXu67PLURaUZUKt46w/QIBWJ
ZLAtnG7+6U9B8D7+pEmQWy0jiAh1noAF7fvf5cdqZgg+U4563rpqDuzJwVqr2AzE9YY56n/ohmQY
LIoCtN7qHy4mqCV8NgX1bzGvKVH9InYuuC8gvRONZRGSLGmT+mD8UWlZZSnmbNhbIGU+mQHX42KA
Gj6ngofaZuAhkR9IqL7TlhBiTfIkDy5f0TnmrYL6ypeOcFnte5OE+i7oJ62wQ+Gsb2dMsGs01v2f
Pnv01s6Btd/3c6UsxIjpF06H9OXl28SiilkQyIykaoOk7a4eD2ikAdNNSKTeehiamwAPnUiN+GN7
Mrm7ms2x5+BNqo/GiBspm/KY7eBMteBPHRw64Eey08TH/SaeeR9Kr3wBNScVOn/kg7AcPfAp2eTP
DRdo24Bx1etqHscYz8aXafkxknEPeD/kiIwGjf3M0bKOQ8ecnYx+8f/xZPGNOv3d/PlSoJBeWzPR
u6fPlcLpXnK/EM+0qYVZJyt9qRTf6kel31P45tGLB4mjHY85s3S84Wr7yJt2Kf3QgkgT+Cuq6btH
iu1UcYWkrtu1EsQrDHLDsPK67QZDvtKJrENkNVZz9TdFGMdk9aNFN4LAdC6P7hlWft0ek7ZIopTl
2vnm0Hke++Gu3HG+v3q7J/vaD0sIq84I3MbpOL5VlK7c0H130TP551U67KPZ0Wib/9q+b/L8nxSl
ZWPuY6EYcoWm2G1DX/q+GxpPj8IQ5n02G6noepMXOT63eXvMCH74qBZsRVl0nXyCeFwNUho4z49h
U+Fl8PQVvwVYKrxTFMiItdrn5CD4CnnCM6uXSh6d7/fn8qiyNXtufPoLo/dg0WVX04T0ZYj36jsv
e72xzOZ5otD9/8urjBZub15ySRU1uimMFVFAhs70j6rdltMHcCI0kdSDngNhnCdkiHBVFtkwPlr6
TWeKQHPSSyNW5246Kq7Pf6Lp1E4YWG5Y5B1c8T7OlbNhUNPFpsya6DQ+Ls6SFGbSSlqe4yvvJDZ1
rmRqxDZ5BY8JnO5UKNTrmgFrx7xKmfiyjW9ewNs8IbfI0WBFdLEvZYEeb4tgA7OtjxNcxdkR8ce1
7A4u/nFb2W4GV9jzkeasY99oijS73shphaHnvNcJVI8gZxxIKCKZVefrBOP2GlJbmWQokH2FSl+I
8l29gOXJwV8wDFospmFii5iT7HiN3EGgea1kSl+C93eiBPtFu/LL9uNApohw0av3kc99Ql7uryEq
ns1bONoFBErPiDDvRlYFlpglg5ZFOYIon+tFRU2Rma2BJdY9Eo5JpFPjMU73ENoqFkN7/fSTcR7C
E7d9tSntsjLlfjcOcv3GhJ8sMNU/TK8KbBeXhwU+T6m3vnTUEnXfOa6v82ykaSpS/TVmP7SPCm4O
i7pWLqGhDkkxYwiL4a/Cj+hOaxPnR5PfE6LKqEORkK/PHUUQ+y6zaHMlP1dSnNNAzuhHyUM1reNy
7PQ/8u3URT4+dQKpqhA/1aTMjvL624lyuKk2VnsZrE1F4MghQkNMnzfcoed8eL7mquxQscfQIKFr
cSIQqkoiwY/+JjLX6nTeXs+qbk1pg01g+C8/fqjGk93ftUVjzUtgf5luAcPa7GKyZx4Gl7gNslwP
bSVpWmQWrjnpxcjUA8bpBLGvasQML4Cd/f+jwnSj8tMdHKmxcOfaQL0O76USSsZufF2IcD2n/eJ/
5EWvSADV6TaEVAsAhkYc3HrAll9ZU4riQJLERsbVKEzO+7YtcKfH/Iem2gGnKU1PWwbuqXPgVmoR
muF7GuAyL5jI8VkoSDutImrPCkMs6I/4UyS21XugYBA6ltkdBayQrntSxBbuv3Aex6SvZEDyNBUR
2AzIh3v8Ed5WkUFUx0qvuhfQEhB8WFiNr9D7R42EuqFBRgIIR3Ze2w/nw55xezjCKZbYI97hx57D
DBFdzLnkOaElLxR1SBakRUTLusMUUBljPu9ipN+1rXhS75qXbUsESqIfVY8UAH2J0Ld1KGdDOe0G
wtPK9qh5CSRSlzvFPRRX+xaqwFDFI7Oh+mvUQdo5EPoAKx05CUMdaVZ4fUFt4ItCIsrX1JP+Ytec
1ezQJTBGDaqViLHQlmTCGkKgRx5N0JvO4kB67575Cw6MPJyMciZysvDdz47NdS4FNIPWNZ3jsMvh
TFptD/O3d2DPMyBGgsENIxGNJQTijxho+vDkzSF5AcVsDVCYHPswE4iKG3ACgHgmd6msR9aXoRXN
C6YjUmjkHYdvbs3JyVQYBQ++eWNicd1bOrlB0FIQrmH2YyoxCEPXa7fL5W/VmTH5lgYfIc+GwVFY
UQSVpDRV7ul6xIPVQQK8aoRcjmmq9aTPEAxHrOaCdlIxXXb3+uww/KutPrGggjIkGKtAnywrXMZh
iKgQXli2jQ3RMzZpcxkLQ3W/udvX8W3DKNTazJ9PjUWA8JEWRkJp9slMoi9a70wx0Ikys39oCH/O
O6YtBC6YY2c4uPMO5nQnFlKjfwnh1uqsgoSB3t+sp551gsy8QSi6VywvObi/9r9YfJEg2FXMcIIb
gd50rL5YXOzK+aK1krBYvirZe9QeLlQFyeINWfywVfTK9zf0d7ip1MnI0AJ9Mex0WWUONZ9rPBDO
leYVsBJ7fmV/uxobxUp0gT5fubspL9ersQ/GiWpcfgCyqBBHqmDckqUN2FN17I9ZsIeoYUV7YwRR
bVgA/ao6gnXJ3sqerYZRc7Vv3J9AONcUwqi9ddAATqgwpsPDzu9NsoKcW6x6f+ylPuqRMFQIYYcU
371fFg1I2dPdfN0g0Q+FgGUfWZEjlwaJBGTxMuowh59br4l7AkonaSAlL8fRvl1kbnEQu19l1f8k
gPVWvPLoc4ZFjJBKedUS1Znl28bcjLlhCiSK/qBMVvVJPLA8CbKX2p12wq+Aj2HwUv0oxetL2KEG
yDKtom57RALrvbK4GIHziDcjFXCxAT8CSRzaPXi/1QlC8+o5n4KmdxQfkGEo3Hh5Ufb1rDRKEIbG
vT2/iJNdWLPaRB+OQb8Vuw5k5Qw/361WuQspuEq5uP22BlFQuJKE5z01bxMRA7p/5ku2qIA6L1me
48fJZp1CWJQFTXIUxAwh1HBUOS2wS90B2/Ag6EW9Qp7sT7QwCr1OJjNr5FO4BFlwZi6T++GnQQuO
zjiOiRsQ8wuZbANL7b/Rj7wkX6CDNtwjyf2FIhgxZEPKfuyLhOJ4bbXszimFh4Zx7YUfHw64DGXN
BTNYeF8QwYaj7kSy1jqIuQyu0zFMVWS+aSAn7brn1VrdHX4It53/7Zua6VV6hvutVREulN89GDFm
UDoNJE6Q//2q92oSfbrvC2PY+9E7UXwh25McejXDWN7tBjqnS5AAebfaPWnCrjkjwVwdzpHnAuo8
Kj5wVA2OaVUswCzXvSzzd70B+iUwXRLLHWfwwOXEjIweoOmNyCdjhPqOiz2/OPhJ/bIZXHwhCb24
vPH7C+t4kacSDifxDfijohC0CtNFxiFfpePoT/JYzwd+aeBDEizdCIYm4axU5AWn4Jkm6XpbUrUI
gaT3YwmJdSlCko3KiRSuLh/OkqAq1ABITQzKntyTDrlQBkMPCYf8TNLnIWwaQTE04TGu2If7n3oe
qUjiKPWOiOw63bIqZW9qOZna6DvRIa97CsWJ4RUexA/lYA6+hs9FOmKt6GMBNzRmagn9I2maC1W4
WcsVoqI0i/icN5CdRj8wzf3OWcHtDtzeEZkfaPRK2cKHKQxHGddmEFeRN4e38f1/X/T02mxVJbs1
ajWMvDvf2mgbitTcTRgCHAQyy7l79O9YHYa1ITGQZFjHt04Cz72d2Zd6wJk1KF/Gx4+uNEnUuuq9
qFq0WRc6jRwyHdbyiPHAnUvc3gwBVOpcj20tcmnNW+VmVDmr78KCRQ8JwJjfkdf5/ECwqJOQ2X+/
QkIznEr1nUkYgKBw6rKofX9h1zs2bUfqBUIbw6khJL3WtZKFMRxNiskoP/tGlY0G3+PDInBPDP6A
6kHCP87sOHh1sq4vakvXN936BckUecU97CLWcpht1MQgnDwnTchB0S+CMwxV0r/1x9MWvJDTBqEp
E3vBdoX4ALN5Drp/Dxi+kdRCIbsGM9i1Oat1QifDro4lZ6B3EoJJ9Hm28rqlB7v0lknEGDrGCMYk
a7xgaW7/1JkAANowM07qeC/etvb8hdvOn/OuEKXGdg3byzUrkW+jy7QtzMqxvMXbue86Fk0HFBkG
y8uhl8kXsNbIjvfnKzIEc3DMmsg4aAg3vn+KfJdbxS2fYiMbLAFB9dZYJuw81qCvPOEvwyZHaEea
74qv+CQBg7iqR7v/exzHgxVymxwc9YmyAW6ttQFbjIZyOhNF+5r3XRNVTPzKo8kiX6VW8vDHUDuT
wOkTRPv78ec0SldMXx9MQ+6FKvRGzPi5ET2+5YveLyY8yG7wg7hM2FmoLBuRzjAPurcUIiGqc4Ux
2TadinfGXwEy6JNc31g+y+uY+ANF/9Cnonp6mryOkQi8f8OZUszXKfEFN+mBXMyy5aBpIjCQc/ia
MjMxyaimWBiCUB/HUT87gdmAEdtNrE+m2PqscwQtlCciR4pjOTe4NTNtTvSmdG5+7Gq7u/y6z5h6
vwZ1ecE7gm/VJHEOdm/iymllAFAKh3j9kKXnTzAzE69ZjgmZZGswh8Q9LjaLNsYKdYxslCxFuNyf
YOPmw61XQPrbJCq2jM242FdMJKYg3NJQcd/XPeNUksUuApTqYuul8AfP2WCf+RyeYW0h0ZV51lB2
MssSzBLkPYikhrAvu2R0P9KqQ5WR/hQCeTbO/FNJHSrjiunxAfRVS6gk3qEIgN0amoPJ28xelHqO
dFbpdFXo5alB59TV9iibshbV5OP92BxO5WLAyqesjniJbWvKQj67d0yNQGaOwnSVg4XoWXKV1mGi
DjROG7YaayoZjYn+6vGE7Z5rW2Aorj6r8ArgpHk9hOW5RaPX5OXCMbrDayInsS4+hrNgulXXCkuA
Il8Y3uUYcHjBzctTnakw5Qn1E+GJNjizrvefOkhcRbpyBPN8N+JxGLYucq0lJQwz4u6DQ8ysnbwf
AFJkF1+2g2rl+DxueYDmMAAPZttkfOGO8iKoBKbcTLNDv7B/uA+qfSdozp2HqBMuOOctejmAKiH7
tCz4cQ65cZkGa7DwGo/6t31MzUgTiBKgMXdCNsp98zAtkJaIaGe0AvE9nL1d19weX5EAmHrwfKdf
ErGdwouoqNyTliboSBUci7f0c0Okb8KzjPWTZujZSU5r6VnrzfyDb8eBvDImWCX24SRgeG92sFOs
5Ahulq2sDPWYarpelJcpYk80oM9hzDyjvFvL9uRlh8cuRXiRxFoS/lVzeVyaASGEkCDPPKj6zg0V
r21KoB3d7ehPe8PR/DxkJV0U+ychGjh8ac04BPm+pnp/qVGeTxclHfk+Saolko7dDg8CpQN49XGr
vHrdJqg6rqXfeE5LzQsVyTcBMFXoPiKBMLWSKUpteYBvleFWg9BbYfDf8aLTmSdVvaPu2EkWgT/r
mG+S0J0+nH57q64A2ianVWXGhB2/IGEyTZWZjj2I1DekVRjZ3lOenecAMTbvUSYIcVWiwvyIs8SS
tKib4iVnxbc87f1V9wmolVeI/1xNvyum58ATG1FG0EYjEREob9O0RfYd5hsUhFcSEwgIFBFRp6kh
NNCqrq3heFdPwWYd6oiIh7rxRzhQ2A3w76o+g/CPVMCjuHtaEujvZYIfBqtCdjvR95iC7laPDA/C
KDc/8WEVbio8sICJu0+sWgfbq+JcqtYMeUFgbt33+v/iwWvn69MYcAs6w5CcX32szuLVUyv1nol4
4kd+MOOeXQptI1LVgg03HX93P92a+yvi8eJPNabSkExZBEMbHCtndE6Odr/Un+GQA/+umLo5a8ck
bexHS7kgQZHSGRJJXC/HQEglO6IDz1AO2Ew6GZU/nDVldTjvjJRnitn0ULI559I2XjO91LAxiW87
7Os+wAqpGyvoBDOzapEFJWgy7AKrDe8Bd4uyIDt/hrLVkcXQ8xxuCFQwsDh2MDRc2FknOOOL8Fi3
lZmRiuoc2ZDADKzjyyN1SewhlXnqdC/S3Tl5LQSiTDT6B0SqzkGecX82Q/y7BqUyq0r7TNP6Hs3N
xOu68YAn9JBzWtqVZlJtVF43tkMKiscWNN3EkjzxFbxz8GMp6jHWRQSED9fZJyVEY/Edn3B5rHfV
/sxM8K4WBJApmDEDo79ndnnOj7V4ql8zGhFfj5EJuUy59Tj+Hf9EFh1tEzoM7speF9IVyzeEEVOJ
0NngLymx8iBgitWz0KvY2mRPKeTjUTVs9l836kBvNwW7cTiZl4OQ9VRmRrdnLWfEP0f++q4iQeEY
De1GujcAuo4mpG/aeNnl+BZccu2XMzao63xRiIjK7DEAmn+5bfOnEG0z0fmfA6pELOF/v4Dws75d
jsaU7T6Syy5kSUj2dEu2/5brbm0ZDdH8A8+nYbRM/UnkhvLuG2VTcMx8UPgo57cCYR2W+W1IKJL3
QCsia5wvaTRgeHNvawiSctO7GmRWWAJpc1Nowbd7WOMExE3ry5VrkqKQ7+PFK9/61YnuZNSTvqkq
EpQ6srQHxhZjo7Mpx96ji/B64OmDMUcbaVNt393NnvHX0ukGIps+rWgRzfmXedqLJyz1/ntPSTem
jlHQbx4vy00rRIjZRV67gITRg8QdIazShtNXcq0x/1TZ2CmimvDT+2XHn5O9/pS+qonNRzS8FUaX
m0pPvC+f5di0Q1GcuiHufNOQ32ttmvgFjUwx1z9j/wh9kGgap633ndicoUJqFIJ1krfMaT3Da91b
A6NuPQP7uz+XLvUVXVRpJFeQvbd4XvQyn9lTvGA27SxB9iLpyyCA92PReCliroCsLrZzt4OFUjhi
GqeeRQgQFnFa4hpwBtZUNtcFwMVUV007nzevT1EZdk3pJIz3uUDSLBuH4WgBz8awo62njLIdj91m
+ApuuafMjs+/lS7r7LXUfUl5DDG8olboLlTDXJfpD9UZq7/NPOZGOCN5N1Y5gTkNIQ5u5Wjdttmz
wNW8inRNEKMocMg0ZOsnlg2pJML0R7+QPIs6BW/L6ddcSSCGdy3S8CL82oyjaxlTsZ7olIUppVRt
YIcZ7LaKZ5pI5wKXtTi9xyb400ymwwRHJ1tq8L0uINFB8AVQqwRQiISpTJ4R4c5E2Vbiis+A5IZW
56DMxvN7k6ToFkD6HnnAaCtIaupdLiupd1gaTvvdc7/AcwQ+bbwq207/T7p87ljHuBJs0iPzJT0x
H7psZ59k8NQ+NRdoM9pKk6S9HLg4L47mJ1uch3v9Su/U/IXsTQTGEoTDDS+LvUSxviIA32+kN2YO
lElVr+Lk25ZMceSbRId4IbhbJFIXbc8Jdsh2ZMKTa9Wb4nrKQEbxmTd6i4gn3TcyiXMO2BQsVOJN
5K8WPyuqtgVxTkS1r+oxTlr3R8pJ0cEOeWHBTy0ItFk8DQhrYqROyZUuP4uK1lop/L3G918iaRTm
NbCLH3p8cduOGC5tKJucWAVFGv9CT8BclmKMt0fpHmS5jXS33sUpG9+Bhe6J+ba68KGxINydcxlu
2q8J3U3FrPBNnn+btmzcWv5XHqf4k/43ecLzyEeAo/djrT4wPPgyREf87iBaHkCoH8/tDu2y91+G
2EGdSxp7IvJKkvwUl3UEwF7tTvJ9FeGJGAobhzpyF0gqWi9MIfKoQ3Quk5nc/PX887PlDCY7mUQV
z28rM4RkYrkmp1EA8vXEwan/FlMQIgaNif4pWdhpAfPm4Ep1EQmaEjbw92kb9ykUT2fNGJL0gp09
2FCq8MrSotmY41cx9Mn8AUMdTXhiLdEGMOevOW9qjJ1DDrTV9V9yPvwfwrsl+eYbSSfUy5sb0/sg
aWWYoNC0Nvblv96Tf5Rqxc0g+f59ozX5c2UrZWxXDdDJwuKkhXD1sC2EryrI5WTHi481hSmeTlB6
cON+/VqFvKT3f+bZqKws9lbSKBNpzJ+A7u3O8cothyKVtzs5Fzr1u0O4ZL8a4K1jOaP+MVm7Jhth
5s65VwuGVE/ic1lzWUzcVzLPwE2V0va3mUJc4DeEMPX0Oy9q0yVqFgmIYVa058r0iXOzu0GZT+aH
PnFzCg9UtQqe6Bfm3jmK4HhgcAw5UTF3BvXIMMjesxkDCrQqmFF0GTxEKP7hmJMWI7f+sfzs2rTN
q8BKE8uT/cnTEuvtdZERyh5BOtiDijngfCqpruBkHi20JgQHTiSOUOQ7y5u6eVmpTz4Sf5Co+Sew
TDHdmr86gqr8OUZtr3UZtHf597H0M68/b210Gc+RpdjKA0aq3CoS2XFnerMJBlQFxXxWzEigq2gx
HSBaXSyC285/NKJdef+HE5PDH7zCF9k9gtYhErL4VhAzb7kjTMM5A75d50O70OCKCkkaDINRoriP
Qkpmiw2Jx5SA1twoFlm+jQ80e4euGbr5g6+zfbP3qUxt68rDvmDBUQCnASiC+gBjLMKOEHDblbFS
rXSU+KPfJ9L0ODuG3viQ6+AcxDlJAqFITxu/Ga9Z/LodShHOpCHxWTezhpJxAMtjda1qvJ/rgWbV
dHUKDz5dThN/2qXEjRUYqQsHyh2IDk+B5SvwBxP6SEcRk16th60tY5OS7NFPR/bBcfiDOdMwgqAc
6L+sAnEtI2j7RzgeoiHMCwwnz0G+S1iFM7M1FXrFyGPeEBStXyviNqe9eTjxzwHns8V1iRf26tSw
K/3DUhcyAjPeu2anb6wbJowlg0upu9ehLQcY7Oxl30vaVPo4HINkgtflfzOW2ExNTg3vZJLNqH9g
ymaDzGscuQudqmgHa0XgGB9JXDEV1KknPFGZrkYsIe0gWLB3Dlaa5JhNb5WzLehumiKjR3Iu/g47
8AknvOJf+re+LNoieQCVYpPV++5mCdEKhSIHrDeWORiO68hmwaxacC0RjoiG9uhh7Ij8E1LdLGKk
xmgHw0Gd+4coc/XNNH9rbvKX0QDGAYDmxRqO1MTbttXYUMJrr5c4Y3276nN92X1wmKHBrUGLPxet
PGzE4WfuPRuExnHeedkhTVRTvnW8HQIIoj0VsrzzReh8Gk4HcAQn1pkcg1yIWY3tMb1g+s4D7n5y
XY0qTKBdyrOhePycJ0KULRo/K4WSL3Q/5uCX22VELFl39b1zmk0KqVVlY4EjIWFAbwxXFshzvqz1
Fnk/uytbYNtvGD04lhgB4Uy4SNE8QQyz7rxWMaqfJdrai6e3U5sZ2OD8na1yNLQcQ4ey3kbiaBit
lJ4rt8cVHkibs3sqBpiXwOroTmyjC68Wdx1IXdspZYDq0LQ1VRdinWA7gF83DlYpVWtnfCSVuvLE
p51uwedTBwiO3Og2LVR5lh7lpXpBGE1tpcB8+VLU/riWr/tSDm39f3EZc/3gCsuUPi4hta6UGp6d
PGY0gFs2Te5B46v9yMaqH4yLENghX6Bqg9Wqq7tzGy7OrShwdxJ2xxuFslEENI2DOhq6UlihMKQc
zhIzMvMLQENvVrx2hCCRcJNfTVdostFSVGJLAcwN0diJlytWc5HEs/2pFPPJOqr31Q3P4Fq9oH7D
FTijSVWdAWUVuK5JMsqKs/L5rGtadLJofTAEcvYbBWEXsr6A5M1Z6PXkiItYMdKecwbTq1IuGLjB
7BCL41NbBGhlkA6LGVBk8ApQGs2FFw1HR6+0tumRJy5wTn9ludZU0ArUtN9H7X5CC0AXmLS3HGLn
ngIGAqp+/gdMy5ottG91IOQUo4UeBresSRdbvkl/UcmrQfdya8mSCm8TTdxXmFk2gNxj84PzoyFB
N7xofJb8+KBYzqSnzhsnmqyL2KHEWIyXkqDfvF9dbIZ5xuvvxcsS4OoqllH9g8Qmv2n+z4irlJsC
EKWlAihooA+/99+sJDhtCBhvrnVWRDboWG53Co0frmY0VBcEMwTRZzKBHl7UNcCRuyknWG8N4Gtx
TPPTpK52vUpddCX0AMBTcje1gDPHolvVyANcAAsHiSQs3F1+J8+HSwfOsuUuvKp0cSPFsDlUEY4/
bEgqVc2hBrYzYev2NNnH49QQtjSCiAWzPz8IZS8ZK3O+cQnT4G0Xwf+uhceWIikOqookYSy85LeN
LJv7fWPUmnZTx5gqVGfe3WIFkkAROBDGWnqxc58dl1XhPoRAjZj84pVa0ekiBZ6+VTYXBsKdEEwg
ZS9HLWYEhaFp0/oRbx08edmVbxk0IG+Dqf4ZFmiX+8ffDLC3Lb2FdfCTYHcYR4BEUj6Efakr+kPh
udWLGAQqxS/s3xF+fsXnM7db3W+58uouSqTmM/6j8c6RIhDCtX79LdDrWRuUxA1gdDoJG4DyRW2q
LOU1Gm5fLkOgaO6plIAvlTReXWgFkY0TYtpJK72b0uq85y62q6j5Wlvmn7rNlPe/84Ddhjp3uVDk
dMKU2atW52jR1j70dToM5CYF8rG4SBo/YiTyyvn0UlsQ+eVgK6JAywzAkzbbyQa5sA48u7/dsAA8
y03r2sfQFEzsetAlVRrt/nScCzJyONl+JQu7oGWxB1Uqg4MwL9PU1qMPNCAoeq86p8m0GAuME9UB
T3ZQazSZwKUuY/bpcRM7Ebx48QKue4ber7Ee5PFOdD9R/3TcPl4wYNZ0PwZYjDbWj6wR8aBZqiq5
1mTbIL7RGV0rBoSupVzTUjcRYQCZBTQbRekqOdpKpeMT785DAA/JvD9tO2z5o7GIhQ3OJjljsDrB
Wu4piKhGO4Qjgt1APKF3Jyfa79c54R8hFaQ7W078J11N5CQEIrindoJUKtaMC4yEwVHX5pZZrJd4
K+Aw27hPyYqxYGvL3PrR8pzuiQFgyTnoAVKAp0FF6937Wwf3CedRLW5g1h3gn/QvFj/qyQV/S2yO
nAanuVinA0hf2tH7/d0s8T74Wa2odua7hHdiwcehRXp6uLr2UvOrgUXPUw7f5DV9qdkYV3GKWbV4
WPZIC7M+V1++GHPvIR6bWIgK2+CNJQYusXaiVqva3HSQ/7AV3i80cSRhDxuzeShlpC7QK4bLCyha
SEhhYttJKiOtojSvekAO6Lln1sKyzoeoyK34S/DvWqIaesTR1D+rMJf9zkltOJCLtG5F238lc35d
OtMwuqLp6EtP5WGSebbMX/tC1rlRbboG08oI9q6ncr1GbRnuQ2GdcV3ORA9fVTXUXQow1prS4bFU
xWlB5CwgLt3nVWcpvfFRYuIjshQnfeTpJFy0rOShKvj7dyqy/peUwKb+sCM6ct6qryHfUSAzli2j
T61rG8dis0LbcWyz9AQtc/unR0b5RsaSZuUrxDYK2jXBXi+AwVJd9zS1BR8LngymT0qgaCei/dr0
Uh/Y17l5SF5g4uLQ7LRRtzHOMNXkEujVfgyv3YaiUcanMQlw7SwxW3EC2T6F8iuF6x3Z59UXgU+E
BNNCe9PJFcK+XbsojluRvz3TQ22BVYcgA+CBsgn7Fikz61xHyrJp7CmIwOobDBOcUTM42Z+xCaWQ
Vuw7iwsCaHsris1b7GzuNSp9yNpSnHr0zsLOaHT4tNKL9WXCT68h8JHa1ne40vAL6hBr0m6vVUSS
Z3jQbd4n61Zfn7KwUmhRtYnhXZ688WljktPegennpPZv4ihVKQo136OkOyTwDo+uNsdG1+zCTBFg
GCJZrMLDUuTZDVpCDjE3WhEvz2eKkabgb297I4VYphtmSR2kwEyV8oqoPE1jIGBw2PwR2fO6jyFE
7O4/o3s1Wdir+i95SoiIKSygVnNN4v9CqwGwfFcufcPSLkXi4QpqxZnqUjVJl/U/ZYA/g12pEUAJ
cneCNGTJAdmQcjjj5z6IV563vAgc6uesaREuqWii2u1I1PvZZKs1pESB3mvGO8lQwgoez3qtLYJB
0l25obHd9tBOJdTPC3GWCXIgZyd8C7xyA3CuKZQZu4j8iwXx5m8XIbRGfSKb8Gw9EVCy3DIHCfb7
IUKEwDMt92f1PUpXR4ez8IlCqFdcZrBn+sXLn9vzF4mXO6NrebvDz6fiCBsoq5QHLpnrEkmfgEQf
7W0gsYVVKMv/VT165EHPgmNOqizsLkx71kvJcMXb7mICpWWkFziII2RntXdc1G2DDthOfH1Ogcfv
034T3ICI2fMVsbfS/3x1cfK/sqTyl5Hwx1nEbxbagtLtoHypugiLvqa8nXsKKnWIYpHBFxs5pBpr
S2oC47dZOfS2n2y+uzj9Qj9BwewYqdrzMh9q+3rmcpVTKShoobwWb3Z0fXGllPuqW0I/sqqByylq
7DjB4ChnsoDV+KqzNxkM6z1/ef5wmCDYzftxe5VArHjZmnOnElgaHab9ErgbKK2D7C8QjXB4zRSd
O5mcta9LCDZ+JNQzlCgTGBSGQww5y5Gi3q5TDNKL+b3Tse18GWPpQDvFkF26JvYorULGJZsj0vUx
ptcYMMMRkjFa1GMMtBRb79ImBmrPJFIt9+uhiTvZhlhj9F2B3swfXBItVkGvRFXu/t593RMnuDI0
kGyzbxL0jNM+BbqSI4cvQeBjdbUCqv9wbV4143Jr+Y04KFZfZH/2Q9QFLai27WC9fhOx9Hnvqtxh
3AFqfuvUcfovTLe7m2WBMd1QYyUhRPW0aO7NqefhAZQnJHHG9VzxH1rdi9dCmUZbZf9Bydp0mhb9
dO5QlqxhVBJmjxPzgIiEOqxhhqLkwq9mZptckAr7wIgftuH4YpLs6s7GZyVgR6cFG/s6canJwgOW
BXI6SrvTf99HvirnBaOUmMty/IaJt12cv9fl/yW3RiH5jg1zZEknNwZ4r+rjkwhqE0g9KYcCvaAO
F4Sr+30WseNfQRSgoNkVf6/XU6LSyfOX2iBBabdjRNhsJ9Lak9e5M+rIRtdxI/ogmvjWlrvbUbsq
8W2Js8eg3SlLPjGYvzvK+NVyB3mweLIxG+q/6ExCKK6gvz3HlprOEUShAhuoqqFRfpunsCFpDJOd
VX/51XOyKdeAoqSuKQJy/RR/lxXg/jzAzNfqxdRohmZnCpTOln7t1JfEFaGhWvQCraAcCA0C7aqU
wnlJKiZAVAUQjS20DUxRuCuyTrkyPScXMI6FbCoEOJF+8WnXQBY4/aEDu8t1HYS80Tdd1KTupOVY
XuL2lr/D3413sPn5YxX/m+un85fMvjKESqUf1YfY1OzxigzNZk19LLJshLrwyZp8jxs989b7plCO
l2tTlXCfdH+4ULfNXq8DTV7qcaPEiSSvPUV5UGQr2aLXjb/cJd75LzQPdeJIo7UFXkJo0PN11uAH
DWR2cbJ0/cC3Nc8hXVL+iiSLQK+gBbqOHSTeeE+wp0oYQa9rkhCUxkkoqOFyn13y5Kj7Nx68JcC3
X6Z7lqnVwpwpbxpVmWO7mBtalhOmcLf7qUpZCxMQ9E0epCFLTZQz/KKpnQZWQLJGQwdFw78W4QZa
FmkVZSlSnmy6rgvmw03xICnVFzeDxaMtTEVVflKV75kdzpTm9NQX+Onv/fWHISFfX54nYQIbnRDi
RUtKaRPcyfyjw9VxpqYD4npYQH574w8BfIHuh3yo6wNzXvHJoOBcH2H1tPkvfLrUtsdgiEULeYUO
GZ3GnuGr76PeElQo/jyzHpUqdKIjsM2vnttVwZP6Db47NAG5jo0RQ3CO3jHqMTk9cG75w0GLxvgu
CIdXePduwBt6I2s0R66U3Y65EiAVfRKPnltB6Gl5TenLZtTzygTTfw3nTWhHoBvfscPcdHwnZP7g
OjmTgB4VR1MJDge96Eis07zrzlggduF8uOu70tqwVd7HVzENKejy1sHLfi6SKqaCOXWdWmGQvvRj
ZZql46LD7+8jI6/N78CsPtxbLM7N71+NCfkVOc0qDWaxFMrZFcU2CvVxOS1mxj6bSlVuc3BQnU2b
FHxq+CF2y0+T4D1B2wgPNoqtUWsfzWVfAURwWpc00OPqwQD2Vja3OB6G15erxIazAhsV21eQaLhC
0cO8kZ1yJTE7bAUXnpKSmnHAxW/PbsbKvSbOlkzjXFO/z2d6XwWAAKx/tmJ5cljvthSPhzKfy0zn
CJV3hpniwIdTBmij0XrDxLZOCYzNok1GcH4rlNeTw6smCJjcMvtFckDROS4NQa+hbQOj60WcSB+p
1MkBdoXBVeySn1t0047p17PHqEzHqpV45vDbDTHrnNT+z5uNfqj7WlQKWWzqj9wH/1cRSKSs1p0f
w0eIY04oyacf0PnMiYG4XThwBgBiLe0O5nJIG7LqFiTkO86uAj8wON2twYBj9oIwr+oQ3nBhAfcR
oUlI4N3HVijSGdgwJWCDsUm7ilgjwrft6M8GoylfVFjOgEAX3NhEzWQkm/fGXyX3qZceFo0DOYcc
20GVvGJzVXrTXZPfKibW7JqtVfSZ/NRFQXohyQ3tv0hYq8g+amLVcqnkx+EwXS0zvp86+kPjMNUN
I9rkDhl9eSaPBaNIAbyb9Rj9CsFbuDioe7dWYOSXX0mNFmuRyWYR6crBpzgk4me4gApl5wEuLAO8
sG1yMkMvI8n0TJWYNgRHcWYpeVonl3W3Y/0qZPmgSHw0jRp1ZFsnenf9rmUcmI9+D3AH3CcGEbo7
aSs06ZwDM9th1D8FXBz2B/IVMo/0eG4/Uqq2hGZjw7BRbYD7VVgSR3Z9ghyiQ+R6VdhPkHiBPyC9
dOdZZLVMCHSNuQbCoT8tkxUzCe7/QaRdgdzFL5nTN0WC3SUMXSI3HsaywD4tyLVGiCVGhNNCC9oA
yNPOXAb1JyLEaHohL5hINjWiBKq/VVYn7DKw5t+giwrgPAauCScMe8c0B2fvSmZPLdG7x1l0R96H
mWxSB2pgsGjqXwmOjWATB3rXtY/4N9fQhnrwlxVmmXCHWqWdcNTXk2BOSpHdc2Kye6lUsEHQaxL1
t5LWkucT/dnGVmKodj2ncjLWlnKm28Uiq/eKFccs1kx/6F/zI0r9Xsb4M7aZSkg0mkkDYLt6LNFb
RUth76stzjJNYx87znA0tIlSpyRe6/IZJ+fX4nSjret6rYBsWIWHYx9rjQcpii/us5hoCENPbg90
uMf9xDRSlT8Dq8RrL3GQHHw4ZlP0kxJPcpl5LH7uargdGOaiBoaSy3vfU46C85K4ljQhjJVHFecN
MNhyxHJViQJBq+3Hf7zt3lHCuDvH4fd3lp+fKnfnpdQ+Pr7DunIM24uPNyldVJ+U46qGY6zmRreh
9uuSm7bR0BtR66msGoAoL+GHD5PCVB18sFKbnt9FlsnLrz9PzovI7tpbBrU9+6RLH7AH+oHHwDbM
IVUWcLEC6rZU/MQBjLGb2IDIHM6pvLLo9KU/LOOHEb0E2Uik+YFMv50dQF3khZ907VjoSnA8DbgN
xCo+rlrjGBFZEYo1bQW+5zoxV1mujTdsWLctBZH3dp27m3uiCIolsnJZJItlXbB0OtOL4pRHpzfk
qQZPqXaxgkMX7UE9Elzrwmz5h6WLNYKdCpE4J202+fJRPeSa+n3Ck5Rem2OYT274V9dX91WLOI2N
uhvM0SbVM9QX7a8cVzHAMCgpezPGlF/bG9TTR4JUCz4ghfEDinXEK6o8knOJ7hc6PCj00OCEg548
0vICotPmVn4joxFWFRH9q6S4GH8jiAtUTTsnT4FpG4V1nTISTYiffhrvDUlnW3dNIwtckZHp0juh
dhLPsaHPdv0wVVlT5ubtkN8mnjxr0RpHhz/41Y8sdPs3axzdsrF293J/hygFanEwz6OtPF/6rHYM
0ZTHHH726BHJgcF2up30IG+eCh/FcGkN3FU8Wo46kXlVtZnX1g9ltRcPYicP5IkHttaFhzv/8HIo
I0kDzZwIUPDZRYuCOFbWF4/j0msOcslHi6p/VhJ5mKSga9W0tSjTX0Qff5Ybwl/25yq1f3aHvXu2
VUr0EHoMtvS5FlJHOweGc2yKVcn80ipeO65bjqfTXN+3sOnbVY0pXuJgK6iVpdtISWGXmRKm+PrP
puRww5qhZHsprS617YTcIbwuMcKwhxHNmRT+j7ww8OLc4520TQMg65DlC4SnHkadSetefWuughr3
vuTv5YfKJYd7CvVcL+qna5Cq0AF/Ye3jkcMOV3IB18Clq8dEXy5A1FV7ondLceewFn7lWnCqMkEM
EWHkW+bui6OVDADc1SWMBFrYl43vWPtWApYGWJAeKFzGwz9fgJfbA6UqUukreYYtX6kD5QAiM/hx
CcAAA1ApaCCmPUyraClk56Svo23ogcETXOG0y6crbsLLogGRIyNdX0ZzuQorlcR0A9gZqcQYlTP5
1OB4eBKkychtQhnwfSwUi5Lu5yzw+CR5TtmqRLq4Rc2VTSRg4yUEA9dsnobyM5BpETuuDY2U/xe/
NYpaNnhi1qIW+SXVyFm8FxFyFu4K+euEPnt62943TR6VjNWSviglhzICt2eQggxvj59ycq157Ap/
JXjV5g7j7xGpRpg/U0KUxRZvRVwI+EfAHvf9ICiN9+k49XHqYH1LoYMZWt97r48dAM2z3ksxQhGe
RzoJfvnb6h+qEFgHnRVOCTtyVOM3gwe2eMuu1anwzesFJuLWv7jkTo8jEHuGO0C7KnlXa32psIzg
kJvDJqpB8c226Hyxy42uC9ZHCmKQRESG0ghlLN/LRcRkU2+VcQOqg7w+3YTBQ/mRbWb0k/Auz9TB
50Bjs0ZIB80Y9bN1BxMn8T+xJ3KdBxmWEkZZYYEr8FkUuknxsczgDVkrktVLvrgyoDOFXa9iKLFG
Y2igBGM1MtFa+l/Si55eK6y4PAIJzaG0G3GEgkV8qeCEdDES5nb22XTWqIlV05v/unNJGR2QSrVo
mHHDe4+PDWD5a6AAsPsa64L+deNYAMzDvDMDlCKnrneWdBOjvdmzBfHyx2hHJUy0C0sv5eNL9D7K
FV0ZRgwW42oxg5xxxYC3hzA6H2a8F7V536meJHOtdEddWRcysnez2J37ZD/9V4QFgjJkv79bO7EH
AE5sq5pFA3ryamKB4ydnsIiXYDw9tlBnOOuTbnXCZ87A5NGZ6scDtG0ooXE61ERU/pHsrP8LCEW+
p06C2lNTAxSEzkezEUvljS2loyCF4lqldrdZMswVtHAgkCcnZlZh9sPyx87xqyjFtPeT4N1X9+FL
tCZkKVh2vcCpr0oXTg9i96QRIUvklrPhO13E7D5vfsZc7OKYapHRClp+qZPZdD6Fg+JyL8z0ej//
cqfq5QBGuNoX34Vx0GJKD0/JhqMroUO9xFnpbSo8EY1+bV5H7ktLgeuhDSVDDko5QjfDr/ZP/oOQ
WkW2JGJwg7OAUpWSh2DWah4JcEB7VXHKXW5XMGT68VqsCeKnNa5Nun2wzkTJcR1jTUCu3jWQeQAc
+8zLg1atZWzspAYruWfgasj5gWRIvzV0fY7DhVcFEfPvSYWqrLdi7o6/So3iX/ukagCdGVKm5qDD
lrbnXnHjpCAgzG+hXrEaWtyhGugvNTjMznc7VhBuSr68/il9P72UZ1vISwO1rOD54zLjkxRC+43f
/XzzadTFHpA6+6P14ybKhDNHegZ8gnS3Vn+FfvgRfZpWkeNcQTxAxty5Dlb4r2ooUuQIdocxl7sP
+i9iIITipnpvecyHCdshaQ+N6LcElW5Z6i0JDBKwy5qwQcCbg6bA47wAL+rgKWnlto4QHf/AiusH
RWFoEo2bOH1/QCn4yFrzS7F0zIQfSktrKd5bx6NnX4km6liqb4G9OdZjwj843jlq2ITEggFiWRK+
+o72mR1KhSVLUJmmIMJz3fvwzMAOFJGvi5lA67mJbcwucUwqzB07l/DxpWZPu6QTVa2IBk2H3iyI
ny/J7eNo+/yqwMICb/DFxoPcgaouVnTRP6Sy0CD9/yPc48OW7ums5BNXeZhGoVtHIf1FgP0wwr8i
mW8GkYri2oz0898Gczv1EELKgjO6Axl5dlMKYXHCxVDuhsjowXxHQKiWvGVDH0uSiwvVdZxgCB/1
RtVpYgDEvEpgsFrqRDjxt0YM2q+VdBerWp3bGcUB03pz5cenF1Cr6z/oHbN0fFYRjSQr0rYE8nZx
6xaUZI/NpFY0KeyZKsCXE3DTfMBHtlaUgrF4I4uUBuuKWqNe2Y+CrXF9Yt8YizeQrtBGz4JDPNcR
PQZjWw1kmWsm/OXlTQxN9S64Ak8DvHt8cDCSG4a8mj81O5Hr3UjVWHR1kQmUxXN7prjlcFweCwfX
0tRSqsgLFEsE8tb/wJ6XZRoDImMhfTQ6EJL22NybQfkPrUklQXrSmsNPi7uP3KdlUyaEcv63Nh7R
AFbYDVhCAXj1AUFEmbyLgmz0rE37YzUB+KMcaeyemrVX+kC9Ybfx/jo91kyBJqu0Mx0xTEa7eKV9
Lp1ovNd2pv2bd24b90xEWCb0vIWbC5TDcSZZHFRbsugadtI7U8KCgUVpaXz8f3uXMQ5qwvvU/v5/
TYcqHjD3PybnEfu9hwQUTcaV3UzMPup/Sjgz3ZcXmP4Z3EXxVHSUoNuJEo1IS31gPOT5y3BmwsU6
A4i7W0PynCh34ZkMKUBArqbrQe2f6btosL0xzh8sH3h9fYIacebT3UDssWBj9Ipt1P7QaQAKVxT0
QccnadKMFiMO9elq8stC0wD/n+cbIhM9y73eXGWDMkzZesEQNXbXqC/DDfhtZcGA209Sd/n3X8R5
zl98BhxWuJ1j719A8wGKZ1fkVpFQDyngSAky4TFQ6q1kbsdF+NJKEH5OudYmDlJH3xATqBaCEdFf
zVuf2EuhYGZ+sZwYRW8OI7tTMhqjrYMLAnYHEHi+EKu2Ww/kpmsZqsE0QIKLEDZXIS3loZ4jBxgN
nh7HyG9oMAq6KtF/SsXWP4S55SvP4Jn4Q9sw6SyF2ggp85d1JzmvR8J7KaqVi9tsLRuI9Hf+wXve
qjqIA2VNjcdcGaYnZy1jE5RUN/Ip7Em3bHocsm5b5H69hGRBcDNJQYlqEWBKZKlK7n1Mh+DMISk3
Yre6F21Ce3PRMn3wmbBHE6541MF6ihdR46KAxJ9VNNw8C1U3vG4c1QmXsL52ORx0PSFpL5Fw+hFx
ClGPmy5j9xDyF7nHcIkFEvMbFAEOd7Pnr/ZaoqN3a7YIwr4ArSJjHQX7YUVMqelc4ZKP6cWNpwsu
btvzdgr499zKE2seDftPsz+YBmetDCUh2+3XfhYNB4MFv1ULBk83bg4x95uy9YhYUAq3mhp8zNxP
VkTz9yvDOZj9SsCws396a4txE7/rqA+iIdgfYDJ3xFuQSPOKLx51pz1BFqzWtCjFZDaVTM4qNMQK
TfEDSUQJzb5+KNp/eYgcj0UfvOWT6EoKyBBYO/Yt581jBA0Ot4ldSlU2njdJJ46BsUm3Q5GIJ/DZ
FcFCqAw+SaygFeoevZZYLU80MAjR6J3k9GgQ/lnuJaEDqq0sl5lz7UThnt1dAei/cpQ25SmnfzRV
2K8l+MtAcJol+qQk4DfWzrXcaVx1IBy6EKMJ5ex76loXph9V6bXPGJNwTfesSFItj7L0D3t99A27
/hvEN7/SgNDKZjoOhwrzJcdVRxNzkMoz4OJUYAEZ3TNNTWRVno4RN+rgSjFgh17oDxvs+eH0oLnF
q6I4k9Ehg2E4a69/1N0a7LX/CYQ72XGFEadsnvXNNqfed4C6w8hrRWiPCrkzyqSmj60VS4f8Dyue
HSJWP5BRRWBXJyoH2CfmrXTpLgjK4NbQBSg3TW0J9bsEAhOlblD+FxynSrl5gagAVHkg8/1OdUDi
GbAmLJy/ZFTW9VnrcB4bFTwKgirZK2rZsuQ9JfSyXjI+61FrzNxzbg1wLRFG80ls/TmIPsrbKgQ8
iSqlNuDAf4MKdB11oHniVGbSjYThdWBjawg4j9scTtsv7jHp4MjOo6z677pv0Fvueiqk5VssIlL4
xD78Osci/gClk+Bj3Jv61/1zQY/SkjkzO2KvVRzrCX0SOJumP9AjR+n/5/mWbkfC6Tnpw7Bo+P9B
dDBtzAotwWtunGknyJTNQh/C4ArZ5N7J6SaGwn5bfEEUveB9P5Cpo3s1kjHdn1Z1QHjELvyGYx1h
CvxRtu7XPFIsoaw/45T6nv2F7tL4f6DI+W0hU+7HgiATevihk7SPMXk8jHLusg4BSCS5ppJcd6uF
PzdfzqSkqaU3owkCR/i2hj12RHMrAi/6RWofS6GNWbHBi8pzK7SUAyAFhNcGlooNLhGTo5Gr73S6
nKam7siTxMGDwMITqMHjSDGgl9Csxg8ZrCQaxncZonN28HbWheufp8HMyBUZoLkr1VMIbu2gdtJy
sspzN2Okp6cWq3lNM4ggYLfimr0y8JQhWno45jE+y7+Nx5cvAkmPxubzA9L4Dfg3UjTYNHPaxda3
//OgtO8VgAYTdtAJLIIyGFZ+IJ6iyDB2QAEZ+xION2OQWhu5Sb6BuLEPbNlIGRPYZAqlzAneoLR9
zKZGsl+3Z5sypweBvq1441wqAEw4JS4hpRooQiCb7qNjwU1QlXZPGuEciNq98LFodOVcy1AjRy69
KFiCuZlJAbPan4GP5GVrZ613LhowFJA/98Bw3dFp57xQmi04tGAIBPErs8NELYBnYmNO0nPK9re3
AxtPtLi9vL5emErk3nyrZscu+WMUq2WKjHqBhEkeB97FYnNgPoxPzujRETjD9T+JIxAmef5jMKmE
cATb+fq+VtHZU5hRS2K1m8D1C58vIQf68luVp5c6tJN7JWIBKV94dZcYCczpIaGACgEOdSMjD29u
jC3k/eyFEstNn7sjG8mMCAMFQD7zhgKNgPRWiJGxBjYKGMa959VdNGVKx2A8m+h61N97JkSA6D1A
kpdsSHdtYUnIUtA9CRre+n9/ih0S2f+Rf8WuZr04UsDCPSEvVHc+EDqEYc4XzOGKEX4dlAxJ++Ci
aFKhgT4oik2eX75fJUmrCgtYwGY2vdabYhniHD8TpJsFcAX24HNQPnUR0tCrTWmzOLRIIiuyyWgo
i/p8JCKoonow9u/4iy1DQOoK0+Y7iZlWnBayRHqwft8WDOuLvCJGyMhQT5u7lhXSi2cKGgOqCnLE
+6Srq+atqszZEJHVks5OPrEJeQUylP9bdUm9BKeMMKo/kRyWagXYgoNKx7AHeNg3dK2AaGI5+LZb
kU0UWMBxEx9wSQpoZ7bmDtej7o+cPFNNi3sWZRLEbH1BRFz9SuA05hv4PwnoQkXpr/nHGosve/x3
L+5U4ZdN2IqQqvdTUJblAta9mHq5ss3Xih0MRDraHNQ1BZfUB7sSSGZydv5IAajC+days6xMnuyf
a7v8Bvov/7pVVOC4NL9QeeT/HrRoD/Baa0n58DuwOBN5jHJ/z9tQoxy/KA99FPJuMkoibDeDf0xb
h/h8yf5BQZIeGJ9NtgQCwB914f5XpeHBYo21PH9Y/bvstMr1OfjmdZegu+4NEwX9Dt1xzTGnKH2S
hqF0c9cTP7DdL7t+1ILl0rpHaQSk1pBvBoOLQXtcPOLpxq/x+bZlTan5ZHs8qJ5+/8yzhWQvIXaK
WYaLVqzMAFhHe8fZqeR8lb7jMde6jRSsDAXKrIhXYTEGho5krgV3QdlUpaVbwFoP1w9aKUa6BBJD
KXum4+rMqZnVICWN0ORuY/2vluPbJHj9e2HVrF9FvMq0iiAUjpqe2yRSWQag5Xl4QIqsp10Ydhh0
MFdTDtb9V6x9vXtH8XpcI7yMExKSYWmD5hjCriWZpfpO13/p61rArUyh/9Q/U/D8GjOGuCv5XNNA
GnIUpO1pL4Aan+C+e6I+LxUlejHZaHHiFdbUFrm3ArcAqpfNBp5heMDy/u55rWHGSDsnQ7wgykpJ
qqpr7t+R+/CKWzvGn0uCam3Em+TcQF26LPuctPkvmJ+FP60lMbPkUWqVWEJou4tSPx2OlADdbNRH
33n9l/VS9pXHfN8yedJLFuY3ja2mg7vz0Is7BYT2sZFMYG1iGuFLxXDXbKmCNHR/a2Z9q5QnOLwf
EUyim8MrODWc3EakW6QljsxXsJFO9lAC3tMU9ReTfPXDEYnaFVRCPGea0jLnqesjAQ+nAHxxPHkE
Sig+pAEteB9bvm8I+sCpWh1jPQZefbyxL/XqYgXQX8wcGqGp+JkjootnUXzjjROIO9zy77yN59oA
nLHs3Qnga5MOkL4B9fSq3wkI3aVBPJyTQIWHo87Jv9uqvqA0sG9shiJSSEmJUgnFVmpCXOp18DP7
/X4YDg8SKiw3Syty86cRVWg4z7SE4dISaWyM+ieiZLeGsKxOLoX44hhZHSEFWXrYdVL1/4/3GO8x
jbPtMzXyUhbMSApYRM7HPDNzru5Yr7SofVmLWRjCHgDsApW1I40ti1oqRP9RvrqXjT/SY/RGiqU9
bLuUwbZn+aOdUtfIMfThYmEnt//AKqRAj1TttQ+U2V1sL8t4iUEHKnQMHaB+dfa9j9ManpXZ/2Q+
Om2MB2hHsz7T7l8FhObNsP+2/prpTNNF5QLeRFmzJfL4zJqfHQmqqtQ5Q99GsbgK3lKt//sPL51T
BojmQsxnoPG9m8dbpP7B9hFpEFSOkpAhW44eO+LaMIjAd06VUAI2qYyEocfTnpQlXEwPWaBbDGm0
/MDvGRFwDyl29Fhh/22M4cNY7wB+NFUlQgtpsA92P0tb0z0E25jCLFJJQr9fDbUmTtDZSZ3R2kWi
NAT5aOL9jA+djKhQLtEQQ0nF0c+nxSdOo/Qzk838CYYx37gp+BB5gqO0JxQUY+xrMYftfjaWe5fs
80HCL1eaLG04qbArTinROHx35yk+BosziR0qe10rPJVgc6P7rcA1KMVLS7Xm/KI15TjhfWIP+Nyw
U4xKZt9KKV/4YQfnQk3VwILeZE937Y9vmhZ4caJQclNTX2isCL+w82X/jeXCS9q2tNH4QgA37q6P
wERClDcuG0VDSnzQsG8xlQjMEVB1G7Qhyf/Nbcdh054Vhi1qQMqajbEbFhCKoCxcoNw6v/c9wi0P
/rH/Fqs5uaQMxqlnr/W62HjElexPuSSMwSrtHsrCDSVpMfwRxQILwm6hP1g8rr9HYJUfBR8QJ//Q
8jtwuNgWNLr8iuuvYD36G6FBszt3vSs3Qle2Fott3clnF3hsvaWIDKkFu80p89khYJn6QUtbSnl/
YkabJzl6UMTmimM3oOFz/Y0Ixoc8NC4gRKK9UYIABox6hxZ3KMkGxKJV7ERxUst3QMhkT3zkcc8g
ZNa/sYiMBIh5R17CIiSTWngdBBWj7AkRHKV+ZWAnZYlJL6yQdDWENmFI7YYBitPkN3dB55J0qZgB
UlcLkJzWd/E/iPBxv1tBW0xFXQAElotgYPUyHZCnmrOcIUzXYRel100yexEdE5wZad63ALh46/yG
Pax9NXIgAyn+umWrOESLbNw7dGN5+ajswx67aEaWolFgYkF3fIgOKpYD8Gexn/ubFYK3JA6GI9E9
IAPgX+gJXfH5Q5MElgJ00hZCj2EgVS7xLj+o64nn4YuGRk6ewIagr0vepFWpfX9mT9TqGhdJvgUO
Zme+mBkJUSjiYxPZpfF3rnqee02My1nz00h8x5xpkEql8FjUKY6uejI/bTMiQc+VjydRKBkD5SNZ
ZNCODCWdXyGAdeNiVOkc5GG1v1ISNgCmvY7PHuqQJd0RV8Mp6zEr+CxvWwGYj3ZVeqVXiEqq5tdx
AIzaZf5MvAwz6qKK7ZNsQzAkp8NBVQw4huYOpaS1lKsC0s21W4NCc/YlnRKt4+83lO3KIKX7zVe7
sIsjHR/ZDyk597ExDvIKIOw2Gib/++SOz+tYJADhC/w5ThEniXVZbiRpTftAe5RgfKWBVgEGDvyd
1DazfqvxfRdTX1sG4OODBmRowZxCi//64yYPR8qwvTdhYjc9cVU/ZUC3ZJLv54syZbyW+V5FVBkI
/5KETToQQrZs0CjuwXlFTbTPo+K3LcxzSfre25n4ujUUPcUU1ObwUAKZmsqa+i+iRcbz+6824rCV
cO3Plhnwyacj9az1FQF89OiyczsX+SbswzeGsC2180RO9NMOvVcLRt4SjiyFOCCoVOEfmD1QZFvc
JHNMirt8aKZlalpJ3lW+u2/uL+m6Xr0YQWgWOJfSDCv7hpcyQgLz0+BsPAnEZT5+NZqxQJOEdG8d
DCz6lo3Ikxj13REalIiAod2GGWq13u2yyoh5OVL9Sp5pcW/9e38ZhB+TOrU1o5KrXFDuHwpuWm+i
vEcDafFAnwh6wg8ssRRMQIrduwm4OfTo0yaLyPFtGHswTWnhMKA/GILX2bPicaY944PXHO37jQub
8jiSy9GxabVzEOjktN22NDMChOd9LQlhQpSlmiD67b+ABTy4mtqZir3duJWjJjSzA6ekBse605mp
yzxQy7aoBy4mMeBWKOSpiIMwTuaEIImOXYcsnWMJn2UgTpEmOg9Fhwt7oNRqYiMTMP/83vRCIOQQ
PeBYSS8uTaAJtqGt8sB/K3jTEun60nCntqW3PDckv6lNTfe7Knb/nLqbfa4aRyVY/AH/yJVV3ssa
uZHH4xXrLSRjGAjwXdurY64F69WM4NVQ+RuaM48BTo0APecgYtIZEV1OitGWn91QSKZv43kbMsJr
D2jgIGuHB6jJotZZlNGhJwG5eqnwM5Kjgqu512jSgS1H0Oqceh4Afkict7d5I0LDojwWrmyHxYki
xgZWHFYWl7zVWUPvp6JwB+9USNxAudC1S8f838kt1iwvTWBy+95TZwCVfSTXb6nI33tojM4Tn6Ew
vMWq2IyV76ttTWSSOmXNf0xzNjChp0mULNmzjvcvDaJFi9rjdlPrX4FWIXPnj3rujRwlpRn1t9ri
S1EjTkz+Cy6GmVq+KedmUeEU+HPzInW+8w3+ovfRpWpVpnkUXjbQsTaj2tYbUNV8sfBzOnB2IviZ
WJrO+rl6zdH6KasViCT95j5O/96up1cqj1x3OTdlaxHZt39xX149AKGteOqfEfG/fIrHJt5P8ZXG
AjS8v7D0mBjaHrfSSWrWvCMPpVamqs9nroJ07ZX+XFCK/2KWXs8d1pmyZSOMsQiyGb2sQE+tti/0
5FQCzx1w3jkQpP2RQzRZvuVziVPgjlMX03AB5naIw1lv82OYbSzNPEWZkzWnjOF9sYIM1P6NoEhx
zr9s0BOth2WgaidAfhqxMxazsbi8l8dJt2LG23E6J3O2t0df4irmB5eMxF/6KBdIaFWCyv5SDbZ8
MEpixBlsDtHnzPxwjn+WnBc80fT5mgNNJPj/2X0NOqx6R6PNO0JfrCwuO4cfVrpTJ+G8Bj0v+2wp
w3FDFj7ojdqeksfsqbfEVta4hfwNUEu6N5KGOieUZb+3vt1wiAM9fUrZqUxXSSkZNqEB92oA9Ixw
ngQ9oD1Cr200rTSzFSu/eMnwIj8JBlN5VZKT0l5yr5txv8GZQ+GffyYr6fKex1ZMG5jZlRLr2m3N
jqKFvpbi36K5Hg0jB+w6p2Rt2XDQrV9sI8vMsQW6O1Tps+9z0krn7/23YqmXAc6/QOIlHE9EOt9Z
EZo1fnZljLGF2I6ONvTsmUQKZccNxnljCheM9u1R9U04k0nqRvyIGW7txPjCIpqtE0I7tDUw2RNn
Y7A6LVVTZaghndBdFWLW5+JRCNsnCYRebyo1ZAO2utvn0nzxEOA9t5gqHFQvA1hCnGksA+AbZAvv
jfNg4oNfH2ZYMbvPMrLnOKz6jE64/GEcDPBRrBuW5WIs2ThHTv/mMN5nWvS9kluFQYjoqoJ5IfHQ
TkKrLs5UV6E/eLuX+ZkQl3bl9rnjy5d+yQNEOnKAoNO1ZGcE/SHNoi5lVpNAvEFE3j2hVnuuB5EL
Qt5gaFQoGRDRnJuR9VBLs/fAZyi5VNPZGpPwjzkzsIwtNcEYAo29xRByUnGPfTgABpKBvl4SAm0T
+SIccUQ0yJEPdQ2LgNTeSKkpPHJpjgd/WF1VJLpuWGkVXf+omNvwYgznl7zjLtAGUDD4begd02dF
fBItJ5QM0sI2L7nwoqe/0vDiaPszVlwGnfj0+zvADecktx78Bi3hENgt4P0Kffwo99o+BtSnLCwp
mSZD5C9pPF39KztAOuj5o90kZ4O8+bVj4xCn2eU/JzY6Zs4h1Ou1y6gZA8YlbSoc8hTvE9UlaRf0
J3CqmEb7Sa8DzsfFmfAuUz+3we8HPrdqmeUJGApEV9O9ZR7ax1zdUfO52Uwg7diyGyyqYq0j0Nh3
DZ3MiuRpN5mV8xbADVQBlvsBCnspdCFIhWAxCRSMdNsP7F28SNcpu94bxdtCZGnhb5FRh3JjDInO
/6CvB83FkGGL2KT50DktBaxMzpXBBfN3HfFXVosCRmCGcufJ1vwgEw/N6wxb2tTlwR8BUmgxo7/C
z9oGfJSz7R5HBNotNajZhXx1ppvvEOkEnqn2AQxu9ccD65gEPxKEKF9NMmU1FVCzhk2Cs5uiPtXA
8ED2IgOWIVyKjrdNKbVHeUH2MA/XtAEzE3EOmU3+3mAR62CFq6UxwOPV5PRuMkYH/AgLqM+jJz3G
eAn4YDzLAZ1rsJlwskgt3PtGC/QDPjr6XfRcfp/k5tOe4a+zrJpP/7uJ3INzkYbjRV+Ed/wCe1zZ
nifQPu/CMs6dMHIt3YhMmdFhUwWttPvEGzgTwc9SHIb+FLi6208RdTb8UfeArePFgdeSOCS3AECm
uioiKSgJlcrvobRNv1KsIh31G5bqWiDVpo37u+rSkVbDC9gzUXR8V4z9aD36+R0V4wmT2M+Cga3r
uAvDM+laZ2u9KpFEZM+tyG6UgCyLFgHH+jSABlh5OnfQBiRRje0/zDXQIe/LajTDsh0s5mcMSfsL
pnEmjANv7LfUnl86rBR/5jgfh+TAAD8Q3B1eyY+mJy7X9NrERV3Pva0wiD4PA0jxvxhWbEK8U2qn
3HKL7lO9b6ZFXEqqjV/cNTj3KPGefgjK3fH6P1KjnIlbgR6wEJX5DW3qUctp1gaELqN/8baiT6oM
JKlUDi/bq34QQ2ITV67JmwzedYLyzzd+5uzp4VfLN2A5Mtn2TOjp2WAi3bkoO+5q2BBsK2A+nLsB
gKDCRKziwl0X9+Gx0EBHbruUccLAvkH+BJDi2RyJinjcMypD+8oEQb9HkjDdgqRNlVIAYRljIpq9
kvM+3J50PRZAVizPu/Frjb4F4pCBMNsbt/IxsW6r5mzRjpTdE4vzHLl2aJqr2ehpOexsLT2f4Dsl
aWIl+xxgvjhu8l3z1dizqBItHAN0y5Pqybw/1CbbsAxbgaibNTKpDg8yxyFmO7R/blY7EdaZo0m7
qataarA01yZ7nUlL3D2K/RiSSeHpAs9XCLg4ps0eh4CuHwFc4Gpq8L7MxTNy97B2PqhFMN5p3fq/
oCd/fOQcEbNi8IHbLM/XJnhlNXrVS3+Kk+yYIeZ1LCSPf7HYdbRKAvCTzFZJrhSJesfLtVPKsKBo
+YlDM03XESfhTqoYhHwE3cZW8VxrQtQDgKljd7LGQLtEW6fx6cCofp0AvvaElR2j6o0AHVnOCYbk
44AMPDErozdDrBI6IAelKsB1FhfI+I9eyUb6Rn0BBMpYfmCH+5n/74mMhONxvTtSWA+9dv7cpUVJ
G35NM202zR7ZzWkfBfyiSRmSonqTr/AdRPe6S3g/NXrsrbb6BlqqvXq3kmJt7xbdy0i1Jpndi18Y
WHlDnfqy5woQjEQHMREJniABDxzKb37iilEoYuQ58/SGpJd/jO52bSTToM3m1ES/CK+OKyQzBBBU
xqrWVXhJneNvSMT83yS3sXqUToS7OJMQf3DIRrs0eFvJtNYnZ0rqYsu+r/8xw3F8xq71tcXdajup
JYisQo7Mjxn2tdCq/k8m9+DJmroMqQQv6k4kuA+oFWks/njfzGl93etHwPXcwhC1Py6jU7g3nswT
aABfVGdCMmx6kIqCoIxtVnPP7D47pwhyv2Btyb9e6P56/jNKJiB0JlVaG/kTGl+0T7VzMQQeICEp
bK0WN4IcKe9xiA4ygvJeXbOOFgYyFxDG/HpUqo1zvDvHFw9q9fJP/w8DMPjdW7tQY6zCH0t8Qknr
OMRpfrdCcOlljOsxXrgMmnPMuEg8VY+l2ACNxsSuEQqdHawRrZbyv2NgR6eLVh9kpCtNk4W5hHan
JuLZXeisnivrSlOTQrZZiGx5yOY1nnif/M+wZm1uwhovLdGyGaqmaLtjzxNa/C6hn3s00tjqElji
YarWazoWczR8GgKOEQJfqjHs56Ma9TxZPjcmIsxUk22Pi0TTDBXYsfM5BoVij3JzenjsYN0ZysI0
LHu5euvLMYaSnkcdJv+tdDk1L1E/uXmwJ0BAoe/XyQ8R5Eflzpo3z0+DJ71gy8VppwcJ5lbBGzKU
oRVBv2/d/IZqsb8EjWixxQ5jZzPMmZeQ6UfI/AplPNVJd5W1S6U2YGaJWoenBgnJgRPaLbFSSneS
zja3SroCPJ/3mA6/gJkuSRfKSrFQ/OHMlAJBclkuGok3zJNEAf+fL1V5pe9x9hjWgLHpU45O64i/
zzkui+S9yocHj57m/C/II+pyQTVbGu84yA5qDtGQxjKnKWFvU5mLOztIbTAwCBtwpNze4JB4JUuX
c6R0rMGjFX7DNxmOV+rtWPVxGnpCEdgmyoAnNebixbXY0Vw4PYDW7aYXIhRGlUutkvwnnF2zYjX/
OHEmf275Wma8oDMekl1S9bLfzmjeXdfPF7QxibFzGLME3dnDPQ/lxOL2emNgh7ofXHLNwULWm8xg
v/oUbfqhCjnpNSNFeFYbCrzzGfahZPoqYE7Q3cz9H1CC04fVISFMkCNfg07RO/WrjK+HzdGfsvFI
ncQWVe3VLsxBZwQrnUguALDRa9+5qmvJFRnKjrvJuukRyQ09sMNnaUz6Ukj+Jh1jgxaYj6QQe3Vg
y53TZZZYdx0lNHXvmEALwjdzQUpGczOx9yFxDIlIMLgE/O7glZ7ablD8QZlHUWxX7mKfRWoUmQy6
2LVeMMuH0vtUJTVVke+NGuAWbgoxar2PBWE+JXEJ4SNZEHEasWTJlgI2HO7wDx/ACtprUs+IhpZ9
S3m08k98a4SgjIvFm40cinA/MLekD7AO5G8LDss/JGMMa2wrNZvCtKRZJXZSEN4Dv2PJ7gEC3He9
A3rHXOXHgORSABdCKxHq4airBj43wiYICEQ+qR8PrRzc23auFLliimVQVpn6j30mrkLfHXeSFjfo
4FrT5lcaADanIfmH4zv6iUPx0AlOiwpLgpZ5KErZHG9+3JD7lTqY2kMRMNIhE+z5a+S4OBw7CmwP
RzBGlZxrS/happhdYBYwkzi4K0Cy/Ce4+GH49CsSy0gCqV60B+MUZMJPCOxyWR+8RwF3BzOEif6L
5UFOKHeG6zT7C42ZVw2kb8J3jsR+8vNpc3bDbz4H2v2EliCs2hgDZfb3kYK06kXWj3+AEHBDPDje
U/0yj/DP6aXywm+nCOUAkpVy3tToiFYSRR3xGTI5evqHlMWCtcPSdXcqNAW4/nCQQBmgtbNzmmRm
p8Km+hCqflcZzZTrAr0xvx/uUKhCVZNtpLiebfsNszKTCdmSeesPwwhMi4U3nXVW6Z72PAW4ZuCQ
++EFCaxTnN0c7OfM+ni/tOAYyyFE3XXmXVqKkFlex6m/taCd1nFelDcnTaZBhmvwwQvulY7lg1MK
ppkYy+EnNkDhQQLvwAXwWoDYn85BpX7SwwsbiaoME6k4NteAwGzHfouFWptG+6npLPu/MUHKkDoY
VtFMnyZb/3KTL2HiRyO5bb7OA8kVm7s7mlgtpnbkH9l6VtQ6IhpNtd81WPB1dDujYEVS2Hd2JCUS
KgkXGmpVEoCCuBgtlKFX3nGM9KVImW/rAU+dTqq/f7ajVryX/rFY5vgt+E1N9qE3GnCPq8eJ1WCH
uTitiwQRDgkHvg9Z+KVYhwCDV0K0IfN4e3++YrzVZB7uepiYHwdiXWJf4WGb+p0jWNkRsHnqT7lr
TfcKUDTgF3OAQJqVxU4M4W5RaIc9vEQlqB/4CGVxf97lysmWWemsZsboT9uD8dRakK9EOvDi0gE+
upnghVyMD2xkQ2H29bAQDiOR02DxFjeI/V8thmYJPNRrdaRvVJU5Ee5D1FTM+01dm1VlpZsyOdyR
c5/29VA8dJhP4lHEHt5gyyNt0WsVEagiHtLb9qNGTwJlOvpTYilRUwST3KcgpMm1dK432Oi5YUeg
sXeJ8hfvx97SjMBcu5p3CowQN50Y7tZQ2Y3BUyWTX5CnqtJNRkd9du02LyE+chsjkeih6pP1XJiZ
oos7836c5OzICe5ZZTt1m6LLiqc/lrBykRDjZgfhj/46UBPB/d6K3G12JkRNizAEzNvewiuxN2Wm
8CXlAzQc0qxoXabWpfwryuOsdLwgp3baCwKQP7/Y8EfAamUiOwc/epZX+4iM4PUNhfqZmjHSfigC
lfWSg/TCFKsDJfileGCuQ9XW84aL/V0rwQaxC6ZDxSajhHBe4ZD9pL36bqKuZlMOiVKvFWMoEuqW
FFNPLcZnYLnVUei2Xalb4vx0G0iuc4B+CsGH1sVYjnCmYgii8EwfRaP+Sv/6O7no2EI8eveqlqdl
BOdwPazHYEQlIVJ5FGCtyvuoEa9s/N3Z9rhrIdkKI9jQg5RhJCflKLqulwVtdIkxSVRmPXuBAHUh
OGutbF7LpRNVHu7Ws+Z8hnjNb6rsbb67Fcr6d0v1Jkr3ktAh44T4cCRsZN91BGFc6UwtBkLQ0DaS
ZHcA1guSUeQydUKsIVpFMjTOCwiQ4cFthYSzcfjZQl0T6fg7puGZ+aro4k0mF2qjU9VY0yrxb+JD
TsWyiFNVy8pUO3PmlAgjuWvTznh7dkThA5ti7Aolb7EH1140zy0AF44hREYqJC+oMzvq3DHNBT4j
FZjiyr/XREphIbAL/NKNW02QDBaSO0L44BH655SVGHFUdg+LqynakbfFPdu4h+vlidNOo92UdOZC
+6WUErpPzVTZaFwoZjATDmTVC9jA0r3QKM5LqMevAQYDmIAIbxUhZ7Yvr5Gq1py41FEPzQQREqhy
E3d55FMwYvINOHTE4Q9k5FBg+bCkJfrkvPXeUAUIdbedxlUV7n9HCk473ugNGBg6y5ko3OcYw8t/
s66N9wWKkxtjUa7j/86gYgLYNZ3TLsEAo+QPL0Ctmz/hj3JWFTA3Dw44rczBBnu/A9q6DF6paZtK
ojcfTShfg98ibHMNRA8llEUpk9anbdcQWiUqtvyQQbW2ZYwhDnZTyor98LMI9WGZ4KEAzdyseOUT
ML6ynGUNiFxCi3vGkveAphF3LlW5mlbDCitVimBRnfKy3zey+EdSoJHD/K66VQ9izYrcIAaceN0w
O5LwtpbjQwkWJT50ztl6a8l9rjmdXtsySdOFHg/nRghmr9AEiFrWpoysA2uWcrJ4NiiCf0hp7Y5t
6a38o6k5nD+EIi+po3sq+G/Pfg6PSj59kmOD1gVNsFjV28FFEwuyvqxlBNEXDcGDBhpdRs0yCFCw
bNdeBVVRUqoMX2qzf7+K0fiw6KjWyj4XFx7bXJ0Q94y/bImVisPGq4udLDVo0yNDuYvn9wtaOSG/
072HtXWOr1xQdJXCVMLDLFy1thoAGlsBFuy79K9B3boSsie0DN6zMLCxv1KHVqRJv4X84ch6ayzC
HCIUKTXV2LRKQeUJDUvFhKwVH2pl8NgvLeCiVQKNlClelVD1WgBNpjkdYjQvF75fWGX+Ljq4N/U7
fUNVzqA0NGC6UNnaekgqDQvDr8U0RQ/k38gYHYJ6azqqrxo4iDhXXPF/Rm7N6bkYOClEuy6Kh1xv
fvkWIpi6qrBCkt5Ezlpr2zz2TagxMxrJCPlKu3bvyE8VBMgk0DO08L6tPmwGP3o5gIZkHnHy2xwh
jTzwpqxU/XD4Fio32XqxEuIc0QeYOaq6RAnXgGkbjOe/F3u75gxe4Q6GNjsQSFs3p7OTEIFtF/0E
/F5wLk221zPJJyCn7Q4MgMx+4/vf4ogIOX4y/0XlInQB5Dobr6LxFHbMB70yg74u2yX/smxV4yri
Kw+gMFNDVW/hAViYt84piw5mN2eY8gSnDn8ZjgxSFe/sGSB5J5hgSoiMTjC/Dsz/V+kwseM/f/L3
GVqqKBAyqs3d9yh85jQxSVWSZ6NOGM4qtcnIULo86UgAoPtSLmTxtd8Lk5Ks4i+fJkkuTm1JeBNT
hw7p+tLMIkC7HrU7JpMiUd2PMCw+Nz3y8AUhdrX77iUmjamOI+J7P/I1arJuMJ3tixzfOhlFlYCo
i4mhFZJuitZfD/9H+kewYe9wipw8JJdbse2OoPoEjx8cUUvlL1BQKOeyz5lW5xGDdOjMOPsRzPje
tAzsrQLDyNoZhH83a7kIjwFXlLAoWUQLoi+tICAP1R+NhqzJ7PEEbs5IpdWSytYA/w6XBG86nb7r
7krBQhRcplzFjf83nBKHeZ5XpwV480YsAGU60We3SNLQgsDT/IQaLq4SUxFi7JL6vckjMZOt8dUE
5wetJwq2A6m8+W6sJcf/I6IL2rtwT55JGhsKfuvw2X7uWJHVVp2rQX6rscjcr6XO5SPGsBMSsjCJ
UDUeYf5hFFvx7EkhabLpZRR/9gCwgfBnudG2LGXyNjo8PQqa6PJJwGPzXd9E59L74xK2cTU9KWhp
SpfQLM++0Qm+uc8FB1xKdMFzVCDsmJOgN9CZ2tihPAR0zwS8yV2gn5ubS3CrmMaFwBEKcvbNdKIp
rMReslTjzixZSMvX6gfHAKcXwUOsr9WiPRhSHcovzwPQ4TXb265Rc4gzka1uC8IEnrQ2gul4wHTH
2Xvc3mkiBrbyoJpcKj11C0yx3Twx9sIGCkKeo6lZdKcNra1+4WMwAkyrJZMGn3mGWecE4Ggo905w
4VQvPUAwZvBtykk+YhotQixYgl3UVWNvjdqegJeMsy7l8Z9q0rtMEG6aE51Uc/jQkJFJkUyWiQYu
TD8boK1tHzyQXVrq5US1WUCtYpVPMTFrfzW5j9ENe6DQ49JGOJdfP+NeKehiqASMtGaCaplNhJAd
gZ5Z/+VU4sNcTkxCubbduB6EkfBRpPSWVjjFvSqp7O87+4pR7NVg/XzDb4wdel/AuRC4YI7jj6AL
xlFuGSW8UVRpi4TAq61UeCvJnKpVt9Z3/a8BcviJPdWGvsAaR0abmnc63YdyKcPRdTMhw9TRDDyH
j5PZZ+z5XgEoxTZoBVf4C+ul4xo4jqma/AaRevatXrH4wNBm8kMWAksj7yCvhPsD+QRaqi+A1Rn5
ok8R3MNnSTihnkIRzCLOArvGo1/0OXATTIVnIqa5TuMTgBE9BBt+k4iZvJwxnStsiMSbYyyjQ0rW
D4VhfAN66lxRtD88EZ8WdIu4LFhxtUKzRZhsiotBCPI+QFQ4D8T6ZDybTaAY3+RNfjlS6mDZzdTa
dcz2gPSNFK/7cFUZ1XEBGTrbcj+D+FbFhpDZxm/layp6ge+2Bm7MctSOAz9jggKKKM7OYj0cb1uv
Ha4CvoiE2LQIID/mv/hld8PM2O4zvn1KUsKFQCaoGHo44LDt+R9g3VerBQN17w3XRJlPmEPv65tz
QreKDg3b2rpHuMZskwTnplu8g6xtdhHDrW8Njn3BB3mKlCdrmHOywNDqYgwOSbn6l5oqSwzfCtgE
xXqHv5O5uBMm/d3L+Nj4OBTK1P9j9h6KjXmKZXJL7wG+IXIRmFssXZnhu7IMk53cguDQE2bJZKmM
KX+0KrO8rW0NPJ5lvhRozAoBAOwxnyCew7Fq1drFqugb5ofjjHyJmwHdrqUeWMu2Sy8T9r3vxqNb
AfRngaDw8wcJ9ajvmxcpv7sbUjeKHXEw57xKMzKv+rqQjXshaQmx3eMlOzP90maCWDSTtE26Oq6n
PPRM9sJuNoEG7c+TrAlTr99+RIZJZZW7c00d1Hj4BvXb7GYgyvp5xG9PRfAq3J9tUy9ar4m/jkrl
YiRhruyE8px+8FwPf1yuUeWPr2HXBC8jU68pxH6n3o7UM6yrlLAdIL46/He7hkUzPqEwUVs21A/j
acaxTeffOeEYV2eFfWVPJGcGRIEgj4mjchNFtTZFbImn0UOLx+7P1BPwsQU4JPzRlnKJYsa49D3+
u3J4dmz77aQIAHP9aS0kYEboAetwY9dfmuoLCrNUiczBx3vJNBhMkzM9fY2Lf5BR2l7H45hMu3bh
cBj11Gutbdk3859nyr8Eny0TpbqxAHghCJUrd8JOx+hZ64FOfhvE1beoWths5hC8ThMQEWdmX+Ip
DgWZlBWkA/HkA+TH0OkOX/ebCF5f6MCvpovyXfwC0OresfW/kwxuwAn1qGfjkQobom4TdME4SGOw
gnpLn7BlVgxWU6PjAVQoCREGMS/mDMxBPlTz/y5/DXUIJn0j4jvY5nPa2b3i7W732jzf8oVAQ430
j3KAkN+8vrsQpCO1zcwabQCYG1G/jFjcMkoKLZ+Uq+lLWa/YzdEJxoG4ZNMMuAjNkGe3As/Ha+NV
ilxPU51++U2tOk4Y14AaNZYz6JPfxF04Dik9wJ33MneziifQXr2dIcbQwhzLyf+6k1uHvkZXIHuf
VD+SDCHnFOmBJAYB2AzhjdwwDK6k+5vv7eTUrxkyTNkfWgQyYGnzvKD3I2tpWZwdYZz72PERD3R2
a8V4oQlkgvMBf4zos77Ju/tXF/8hnfw1W0h4ATCydvpvV47MJoFAYOyUiBl22V8NMSK5J4x5qedt
Qv6PscxW2H8oJMWtmePnmoFsNaUEjbx1LXsxOUSS+NsNuHgPndRNiu+B2F0fCZ9RNIcOfR1MdtbP
e8iLjlxNX14Su1iG2bX+C56HlPfeXPh0xtF1DzUBRNoBtoYbL2ymz46nsAhB3Czfy62QjaxHj1tn
9OJalDUWfwfC4ZkFi2wjrNdfFRIU1mQ+jSybwjkXsChGnXDohjIsulcsIZti9YixgxqOVpzHYhea
nzd3GhG0iWsorf2m2Cv/2NmzgsMgyHILkGCrc+qCx2iSKU4GhRMa3qhToT2nD6gV+MLTvadGicLz
AyUwnA+X5vAtw+Kpv/FyBhKkn1mSe798OiLOF3uioZHPDeid8YqaGQdvg4CHvGpWdrxb60aP95zf
hIyx88s+BpZwHj/j1yvrpHjH3Y0clY9LX5E6ATNsx2kQdHR1HYI+5VuY1Tg2LXrUeKphm4P+YC7K
AVw89Seq3NeTLLXbTmLFNUubsx7BA3J/SG7dHPABwwMC692dQjDHKtgdQyxsaWjfBtDTOD8f394A
DjJ8fVGyFqgSIomTf/jz024sPZPy4hbUlN14g005N2uIi4xUxOOMabBf0QGUCyIZ49Fj0aX+xjq1
ugIV0chmQ8NGZBzlL/EI1iblQTw9dVy6SOppSqvxHy0qgglUP3jFOy4HC4p88hAHO+TQgLrLV13L
pc+rVE9CNNf+6wWAmSKUehXwYMTOSHIEhcqzRVKEqyOeq5o0Jj7SGI4CpkX1xxaJQp/M6Kc41Na/
zJLm+NtYr2cl6LnPbTe7wAqg/m5B8E2tViHEeDMlmyQT8EdJbP8AHvFyGxqmFqk5kGZYj4zK6o36
gtH6bJDyW/Hqu4EhiMT5U9tz9doLugctyiBTwSHCnpFHVeA5zH4VjNrQjywsvI+EOzorq2HdNtcx
6nFockzXxy/QK5/HScuVy7IxjETANq1hHgalmefTsMZVJ90FQsoXFNyh5vLG+im0n9zFwiiwRL4I
IgTU2TdZZZ2Lm14Hdpuglwk0CJ2k1nT3oGHi/T3P8PmJ+GXVjNJ4Le/q0KlU4e2rKay7zhN+07C0
FOCh8h0DBujBL6TwAnzd2qfGSravHMQPhIMaXSHiPVv7SZoFdeWUSV2HUh7tksjZws341EdLKpie
Y3nQeMGZJJusYc94n4mJe9W9UvgD/9txg5urprLq81fKIvPZbvpGGkPaZMNiDtpAoI6wzu4UrTYz
GEnbVG0FpFubDVIKRR5E4QnN+0VJOZ3+2EHTf9+a9g+lQtL8C6O6aaMlgx5PUwP/0Xa1gyXkYGtG
wpkmpFA2Gd6z3uXDm6UXmY5Y8m7+T8l31SEJSzIdst1m6dSCkBKYMQSdJcG8O7tb9pRaT20AKCnX
EXPyBYPJq7S8/Sqhl12dEittIQERef1Lu6IS3W2IS6k9/d2gMJqhu1PTCVzcORpCK+jCHNZgi0wt
vOYyeZXcqKbdEInVbCOIeA6L4lqRmMNymfdXr66JRgU5FRaHi8Wi9QxaZXem+KAMr/aNEVetC8Tz
/V1BLfX8VYVfrl8adDhgGhRbJU0zNlW2lBFBFF+HuK6IyrpOm+iGMqEeRAS4Q7rr52s2Nv/oXlAp
bitdywzx/uWo+zUonBa7XVGkHX6vjdniemLWZNa/3J0RLYuWylFWkfEldheIbhwS5MtBo8waK211
+GPvnIGTi9RMfR+zcOkfoICq7hUkiQRT1EjwmPQBdhLO4D32IL8Gbbc6o+mslORW3GO1p+3YHU5Y
CZmVrtIFTmwuVSQ8PE8Tl3HBP+Ce1slAwbLLlsBoiA2VTgdaijhKFN4yyVisLjisiYx9MN0M8lKm
FZdGm3Y3M6D+o7a1h09G9pnBGbfzCOZahSf6Aayr9wGOszgEJHh240loHKrzA+ceBbIdm7Yn0SIT
BsbIx4XVjkYyxxgroJHG81+07s1FreMo5lBcyUSoAhwX/RKiy8eb893MVPNuBEfcWp1b9JFWb0SF
l39m+yO7qqvVl0woRQQO0mbucq3rb6gnrNZPlkbVL/r5g012I657id1Uli6ejmwHeTWcaIKh1hWn
umRQJ0tNxs3EmGHIw8K8pGxN9NQEcnoE5rCFodmJNyp2uLhZUYJgMqGNkc4wIY2R08SqLtC51gaM
cEGI32Sqpd3TFGs/Huj2vbBzCbbYiUeBoYWOnbexflPbD1jy4w8EkGWS+WVwZNyWjR21lf40YRAC
djD52lz9SccNkJkj5BFgYevIC4US0xwSWfYmOAT3TTUCohtajCxPDCMZbRwuJdzVPzdTgceWqHaZ
s0qOUGNjPuGLNpFISHBxudSnOH+O/ectpLsH5OzxmK00+j2NqbFpKQip1JQnwbHQQm8GgcYuphri
H0dL1zPujG56FduUmsZY/UkjZICEj6RjjIRasXAQ6UaLrNsWgidnMpFlYRrTki2r+sN7tEMLcc7c
05UooyVmWFRSzBPUiooo/HXWyn2sM2aAm+jVI9w3xy87LB5A9LzBblis/Lwmktl+laLez1t49/uQ
35x3JVGVbeknl5/zi0roUetr/omffoxqkgjFR3FN2ax3+yPxnWCYtRG3Aw1cwHEEYILekV4E4rZV
JXX1Tvztk/+3YGE/kDisgneTN0LISBFK/O9D3rTJOGQsXDAe6yUMwrkBcqd6hvAIkKq5oND0WO7t
chnFCPlQelN4mu1Q9D0U6sETvrMxFgGmO+dvZuDMUjkayDhWRvIbE/8NElLMZNaaxyNlPGAjIgWn
JsthlvRbcX2VO4WDoUYMpFMyC+BbTNfghTyLBsm+tpG4D+QKNQ7ae0VOA/ph7G7hL8y+BCSwkybO
80moC0v6oZzMEecTrnyENIhOf/dYMaiEtZgDglbNc1+MYsi//kSVTaFa9Vebyls/E+F5AG5qwdB2
GSCJsVZ6bqorFEvMIGMIvI41I+xcIotLZ+WxRxpkT4nMhENXI9h3Ogo3xSm22v/CeVlenPDDk4Da
9oZ6y/a+IDEEIrwkCrTM9THDPeOzr8Vdhm2jeZM280LIU+ytzaUVVKae6Vzbt45+ssm9elCPIpjr
W4/nlcmn60MdVpPGv/5wLg+qKknhNZ7jbcxtnKoKhkZGKajEtjwsIFVRHHmwnK8bR/D1/LEVzqdE
3XDn1SX/fQCs17bDRwmyZ3FkD4yREakuapNNlH3zfcvesLq8dOTQ9YYHzg9Tud6dqNcn/ym26Pie
AomidwZXn3rlSqNSooThUHqqCO7e4et3uAWlpKHVoW8Df9HX1SAC07ZZdkn7T1PTh1/POyvb5Mu7
TOsW8I1WN1hbtzHnTFc1dXYBEKbmvumld1fobPrG74/mbSKmrH3tJe/n6wY419a9XN07IR9DUwgs
f7gx1vCX5RyXhNl9aJF7pf5BwE5ah9eK0szalt4cALNFBe6rPcs0K5IA58YEXPgaMylKMaFFN1Ys
hwh1eyu9NiAzfdep9Dp5gfNIx0+xITHtmiY15A8f+J6EOus4ZyHqQnovDKjKAxfLIjj+gUonnnk3
Uf074TIiWpBD9DRwkIhnvPOK0mzXPzGbefL3Y4hBhbjBLCnjBQE/h21XuaIpM1/MDvGLIJcXeL3I
GUr9Jq5eM5CRqhcN2BS7Ktx20yDQTK87p6in6hqDteRBRRNi8BldrsGcLr32bjyztJsEj3POgCqk
sPwNz6j2uxTR1KgW443Z4sfOoDt3RoQMRgJ16798vrrtQgRkf2WpiTQUYVt1rkxaEb1VOfi0CWnO
fo5WK125gSYraREFLP/cGpP6s5HNe1yFH6fsDCobZtuI9C+du3561busjNWZiXTdHqHaZFxl2dHE
g98+yranIAaoEZJTigUzh3v8pPaPIhfRA392Uk1Gk+La/zmbVG6QBWW6tBzKgKW/zatL671wd1Kb
9sFrnGtU49mui/y5Bm+EmZpmaXBwP9GkV/emJneF9ixdEIAn9XMu89UD+vq+/5c4g+Tzt65qpuy/
lZWjdHsLhC+ffM5O4T6mepAFc5PElapxXIDK0cjVTeWg5p0oL0Whlw1wl1hmv8kSugKkW7rXy70X
SC5dAnej/Dj2NbZlz3jsbEPjsXebEzoK/NjvPpAi84aoPhKEkVTTWVhINUk+f2Yf3Tg6jnnwamPS
rdU/mL2R9B/0Qphjcxpvo8EAnlkCayODb4dripRqDQS2ytLwalELAVkXhv53e+pH+bHDzAvP65dL
9oSJzls4sFlbva0BnBl6Eh6UJcuFZaA7emw9OyzrFCYTWPujnXioUHJIP1o63CJqoMu8FWbGlNJx
HBfChpr9AYZWbFUXPbClUwkhxkWxLlUvgMmDViYzzwfFtWfZ5kJNEoExQaehx8UjI2v5tvMC4dcR
qpSOUY2kbDMnuh6DR7LXyyHIpdzM9nTT4OTTxuCl9QHSvjMiXsBIydBFfQX0sfks21Uap2685nXn
GS1nse6hlY+Db19CEd526wpGZi6av6xEf5DZhcLnxh7sFsfgozRf6CE+zWN7YZGSTkApYQapwQLz
RWsai2dh1n1/T7wqw+gpG/rYJpIqUB58dx8LVIVFfqAZ50Vs1ZoE9OcR4tb6TPp5sx7MWkIm/mmD
/9Q2J9mRYk1c23y7ZUdwnrnHV4aibzaYdoNRcenfD0P82NkD0w1xVgS3OZHRGe2Q0FtQQp2tBY1i
d7S0ZcVdcQtFQpqn2npNrLtAcgc9rbv1bA7FYWkAXEnwt9iVcE1F+GjwtEsYObSijaVl4fyuX2lZ
MvRS7ZQ0YoVUriS5qicSQrKNu9TVu2IdpoxKDbWt/jOTieKGbG9mqX4/9aFwd7OcDErYNIv6IslS
okkQZupR1sW4cI9fCZXUOL3E3VM/33xlihqAQPteMDlhVWeaiZr7wLlGr98/Gh1iQ+uBDKMIwVqj
HWwEDsiaE6x2VONRN76+MRlb6cWJf/4uOUdOIJtcMAQGxvfnga5N2owauVGuHCGlDPCZSaPC7buN
b+syG9QFBLerT1J9QGZKt7YLGDow/FCbt20y6f1+cZBvMVr36oPiFL8YzW0i3fCSJ6vjzRbfHWr0
VnEblz0rnBqw8t2Zfl1hCrLpIPMpfmA/Tf6UdepQiSLCFm5y1+i8zO54gJLRLsR+vmLnZMi9r5Zr
ljOWesO6wcjjhXlbtEq9lIWQm2ZVTrIHwwzs1sVsjnnBddS3muvxIycwJ4q16+YSVG9yT77g/YkE
oBYJL8NqceLIhP0zKAKDDg/lWduPSnX6Ry6IvoQo/lGc06wp6bjehlE+HENn3vvU0vQvIpd08IkA
sIl837i7FwG9DVPMCb5jk6bwa/6+2BQMClr2+mzN3hucT6Mv7IXaRdja5j4ychH5o+hXrAk534mH
bw1RClzijoaA+R0XK+tIGeIWJ8lrH4gEm9ogIUughTTk21KhKzIuhkrgSVnLMJLyd75lVOZCXsgm
AP4tqCeC15TUjvl+CSPbrLhkqf+K5mux2v8qjbUCbY51304OW/30d9WWpj/tXEqt+5cfzJa4f+wR
C9/Q9FkZ8N0Fov3CFXRu8iD9qP6UZwCfMDOPbhtbt01H1Befph8D65GdC/++r5nugtMFVrxaEfIL
qayap6Z10q9l8nCidZ4coMdYHasRLnfANqtSdB2RcICT5i6hg5aOKviMhanfRt5FwrwOU04xs37g
0LAz6RkencWQaBpatBhY0ZkRljZnGi9kBVYwUUtMx2uTgx4If7H4X4ocJEodz6NNaIq0AOKXalQU
qD9jL+3YU40O6zcFyHZWy52JlG26ieCiorQHnUew0bxxq46HfhmSCXq/KkYZqgBihmjF6n8/6cn1
2CueAl35F+a5qyQr0da2o7uwhkUsKL4qmnQ1nriLoOUDbCceRJ/cZjwjEdMcbd2PppUBL7fKXf1D
62VbiDK0VZz5dE1a07l5pmxZGsutmSbsNcfzd7XqXYzy6ZYmzFeHULgu4zS4zuQCtFcehR8r8ipY
QM66pGaWJZO1IT6gAHk7BbL6FNfSoXJer/d9c0paQsiSKPjBDJV9DDacilgT0Nr1H0+Fc9qKYdZJ
3dgGxHqwiP0oa6aHv3hD4nQry9HTcxhomSD6b5F6IZcaDqyKnMwSsajruFL+VAQ6LyTxqdfYNIMG
fpbQe22xmpZomUsG+hV6uKBfBsIhZA7eRkBuFWrpWQJ8IAwqI2fZ63YueFb8uJPwB3dBGmuI6Xw1
xeWY1EE7ce6oFmGPfw+HSj3b/C2wQTQkNaZj+30vbfNL9UJM54HsvNhbou0+/yEsgF/q98634gPD
GGjQ17ZhE5m12sbIXuvHc9e0YKviBC7uoP8KOkFoNI8mIWtboLViKfopOL0KaA1FV7tVfoW6ufWC
aDawS/+fJEFGJGEkKR/tu8RDM+4mp1TkriYPHpbFckfqB95xUKp9TdU7Lu2BcW9DCBEnszG5qvzt
m5YHGoGapjheAj2yi222aMTyD6HRrk+sD3ZO+hGl2qVNpz+Sop2Ud4d5I/1M3SeFYIpjbK1M7mB5
1HNQjLVLBwRabcUCagJDptgPzkRfmv7u0lEqspmqz2CBzize5pR1p3DdDEjBJk9rLPoH4e+98J5q
W2kMnXDMn+XXDD+eLx0PTh7IJHxNG0R64r7bpwwb76N5MZi8qfT7lGPdcxKu8oHlk8Tt1bnxRNsZ
P2qXX06fNCGezKoVW5i4BOHYRlpsj8OlxmEc15ZZdapnzCQ2S6rN1zXIuQVFXym+wGr3MYBq/dWl
ZbcJg2k6XPxYOYeiQfiG6nVc+WJl6sfG5+BUH8vjb0AKikg3EfJUira18dlBka0MoRjs38pmDRhn
Jz60+rAPzGs8puJScSfLC/upyLqUa8BBSRGvSWnBr28wtOLWfIMKDliLfF5hVzZOnF8esEk7jhM9
0o1n9LwJ7JnFP5dBFQtSEUVZagxITVSyhKhEob7mO4B4DtA+t02mPFLtTmVpQy8LOnKyAXiIyVkf
2KSeNULy0JkRoigTB/pCxmFCvbAhnxn2EFSuJRNOSWh/NeUodYgLNvxRU7odUzwkUmQPiFmvaD4O
Vd3zdmIFnox2z3UBkIaghxntf0tjoPL+lS/ku3qdEpeBQ7/zKmrQFnGRV1jJbaMdpuQ9ZMBwKcO5
35kVTKlbIq98xy0FepxPFEAyVKfbDK4xXFqz5PurCcxQ+ErZXhAU8dJnMRYhLaA1QncL0hX+a46f
bDC7/0necSX2lOfQrbLHbitLgOQcSuJwRldGHJsEM1Ppvv5Zy2xucsq8rvhhJn3Gc/3T/TYS/SiA
EuMvbgW99ByWZ7K5tv+erUreDl5tpLW+SvY7K/RpIMaQVoj8xyhv+h2SZBwfpA/gartU2Mjv0WoO
iM7RteMfEVJ0slzXAuPYqpYJN+YQN3xWvHEvXc/XNsmuxgxqlzOOhHEE50cyibDpOG9m5sxPNwGp
JwnfscQahAT3loHzKHt/nbXIVBMe4ycajHhEACooTbloLMomImjBDWZoZlThgAMjYv2mugF2lkRP
T7nNnmHOv9A5YanyB68JNowaABDadR83Z4zwbjVhNS4rEBTqBr9t9bjOZ3QgDZy4FAYOs/q+hID0
CWhqtWPCeMQ/UOU761isPsSTV8EvO2wYH6xVW/zLjJ2Tq44Kz3FDy6xdd9IQuMX2ol9fdb7myGo5
hem24gR1EC5ATmI5LJylgvpnMpTud7XtR8FcX5TmHmbOqvAU/uKM7FGtMpmNJPW7FRcE+B0iZg0T
hfLdNRqVCWV+CCwaAYTk9d/CyCUQnhbQHtz7kX5W3coL7hrwVgVHk07JAtJSKvzlPpdwc4Gnmuhw
x4KMsJr1l8/wA6SjvsR+wMEdn/UzAm6Q+d8lL0HRgMkLHCOHt4iAK8msxMfeO/8uaA4TV/F5qcj7
dt69nNLsLVBmkv/HQdUTzh9Wh4Qjg9gWX62A8k9rNa1NJ5UXfhoEimSnnr6E6ujDinPL773QfEmE
hbtjjZ06ljZEMCyLgGiNCrG7sVgRtjtBIbdjZCmmkAYSBsp7cNl0fPzbiVt807IT6AbhqC3kJSka
WWdWF9I6ht2ltLl2FZEw07szDrpUG4awmRJTvuoUFR6HgzbmmWYVDZkq3CyLo4cy6RbHJHITOhHJ
804+hNpa4m86scJTB2bxT9iz9sAYpF0VzvhQYIw2AhSBTf6CxdTTtHpHF1MaZL/gXf3YIZsGsbMx
0DUCfvUNXjezQWPGGYiI0JoB2m6K44ACxgGNNUmWUoYykgwNO0s08rgYafoIChuiRYZph5SK072k
Ugx3sv4kfULlvPytTS8Qn6tcRBn7o4GNH5gK8G5oL0b1lxuAAeX7HV5eTVOYiKZLf8dU7aWZ8sF/
TbHxwFiXY40G1GsAQ00fXt0rW/5Ve/Yf4arsfXuoZ3FqRoKWK8kyi+XGeus0FqANW90JjqG+JKI/
fDG2WyiezzbqlGNFEqleREhfrGPNEaF2W7tgtc4e97Ad7o+2tJm5vow988bQpaRHDoU142DPqEVK
+0bAC4CeRUi/arD3Bdrd10jG5qzBy0DMhXYyOUhutnxmpcruuJwu0tTcwtK37U+jSVBHaMDtlkxI
vV02YxrnUfeO+m3gD4/zjL9EBCppemJO+IaQr6HiFwG+4FPmqi3z6HsuBFKP5WQP9nBF0ONVvxBZ
0gs+x2/Zk+YhUkCeF5L4AT3TzRgyX0UriQGVN4/2NL6+DB07xXEhodLiJ2uWn13xMdtv1VZaIrwa
inhfRY7ha2UzLCigwmOPW/uuZ29yzXDSQQzZhSCnTvoSkrAJ6JTjZHUeq2AVELwXK6O8A/Ums086
FuRiFCOvG/66PQP9vhnp82dTyOkNtw95kB91qvysofc/6TXlpGP1aeO+/8/hChYJTJ9T+7N204kf
5JgpJ7TAHKql7S7OWjbC3NQiheq1ffT2aYjJVR+RkEZIIAPFya8txWC2vBxOmtfKUysNQABXAaVX
D5MkcWehm6CNTT9Lw5uWUF9DJM3RbeBeY01gtpDxOXFe9pVigYny4F7C7BSojkAPjAkn9S+v/+WI
NIJGcRLqjjsby+blX+SUuYfLm6QAsnuwAO1FFOBV+QMiwhyja1tq3rXX40hb55HCapT7QqOXyubc
BJi20zwBLW0go74GC5gUJkhxB01fRZBP3DL6UZQevxw1n4COw6JCLRDcHl4Qcm+7PVOpJbThKYiw
hA9tQVb8Qfsbb0gwEtZ7JTC7gSKRLqZwXSANzpS0DJ0t7yrq6StwTOlXhZFK9C+pcXnl13RhjXq5
6Kj2X77glQFi9w1wXRF2dFwvPVcE8IGzqniJ+TkeMk7n3Nx5UDwmxYkgqGKU3kQrgsIm20gky1QK
LvITt2J2XqzbXMi7lu02B/CZp21p/oTpXCdlGSa2N0AOW7zD1c3FX2vdW7WVXcd5VJoBF/nmfKPW
XWRNkHHRaYIT7lXbhlNGi/rEauxyGkuYjBUZ3p+R4Dq6gxJrUhYirQ/eq6lkHqIae23bHKE7ueDg
2FIqU0ng4KobP5XjF2kFtTzZAeESoxCsIDyGogWeRzfC54zoXtPOAP5bWULs8kHVqvipd/Rq69Fn
tqafzmaOlJZlp3T+3wXL9RM+c74fpEXTGCelon8HGWEKRqrPxEx+IDxhVoTo1sn3sc+OaYOqGJZf
EC+KqtawHJQ4xeJy4wPJSe6LCd7esARDNoXkCR6L6pP7VCVWctbxwUmA0pKWOCVZhQ37SBqLblmz
+YvrmrWV0RPSkP/0VbewLRaCfaByTLqD61DFh659SIReL3Pkz3GRtg1xghcCV4g2fvvbIvjout0A
L5/eluCQqfpCnpUpR9SJmGjUVgbMFEMMfHlpVpauzDefDslJLZFaRgZpCydxApUQuEHG71VRSlY/
Y/pXkSHAjiyVyXqC7UhazfSqvJ+ActTTcbTXoDMZvlpR29LMenKoq0IwZzPGlhbzFZ7lzVy/cUY5
VC51GtSKfsA8eyV42NOGWtxLM1/y8yaQ8Jen1X2rwjXmlP7XswSmeWMSz9WPC62SuF9XvFICDL7O
QNqsRoQALio9lFhZ3qYJOI4xL3eZFlP+NAbZmeYtGyDQnBh2vH8TCVXU1WAApJSdtJx4Qe8Fy+tt
Xhn1y9OP5KjScxRwRL9hiItgLZRHCLPblyZCWg0vMhHT/PmgcIdRh94O1/F2FhpsrhgtOJDzUqGh
MDCd6gdr4lGfo6jWGceur0Ii1YJbovtZ2etMsrW8n8tZWaHdemy36gvDyB+z+G8pT/Zcyqv0pxL4
JmDoJwBTahOQ4B/E9fMFIa4fvcBx//wDFrIJVSijJx0l7U3RufGHONr4C86ZO/IdxmoWf8Af2vjl
Uecxo/lghJBIArfScFwHFerP4nWKddG+j+7yE+k6u4WEQMVi6QMlz6DRz6eTm1y/qrX2KVPgCzbU
SmUHt3+qfO3/FXEQRy9/S4NxsUsaGSzU0bRE3CqBGRMbpo/IBuOrlbnhbDUN1lNsBzRUPkySO6Ry
89lR+6k04bFvkBTJFPeq94XUFsieYrZ/XvYDIHTHkhA0Zjw9X+l7ATl0XF7K+5fB5BPX+neKAFCq
uep1dSYS1PPB+wLMpYtbdkCcaplf9U6ej8q66SFGiXoeBT6W9VrDlfpQ8v12CXA22oSK9RJZVKAx
Q2fAJ79HgXmalBYG4ONUT81Hou7wg5eIpzEUVYqpUtkxDbAeXrm5YbvtINFfEDsG0PzrjUgTpw/y
gAPJHDOQhjFxPkjeOOXpGdj0dNk7lfuGPNecJkky5ei8UsmBlzleT7riKK+uX+8w6+6G43D8gjYh
3lzfY36OXw209oEsnU+KLvX9OfM+tSjskii44RzBsZSLs+dfzVel2noZ0iVUz+PPxxh+C6dKJ9d7
jittvbKf2km98/zyqKKItfASzdwLqTBwdJEyL2CbHfjlLU3OEK/ss1iWoScRe1lNYwlenBVqRls/
ButL0B44rH04tUfs6DW71n0aHDm6Pl5ZQ1uEdG4INkZkyAxQ+Q3U5RJbfG+hkVqKQzIbK3Jukf8C
avUzRZU+7OR/Hv8P5fkWT3pW+C1O094/CEG0jr7LO/xsGKWgJiwQ57eeWGbsMMyLj07dn+gq1+9w
5KhYDBWkvIM19D6Af7miC9O2DMfHAPdZ4FEWl4keryxVwBvDcmSsnh/ncBdLFMGbhRFp+q3NLajI
7Cwx+qqnGO5U5u8MLoVfNUVpyeMzTO6Xj1XBopnC3H23i9cTxkMtM3Qh92lBVH+svN1lidH5g8No
BMAK7bV2PyEshq9RpE5wnr9GnvD+fEp7G0F6dcE4f4kn5PSLjs3GBDHy8DIwRlbuIBiURhQRK/0G
uJ5VduXUiM5lUhho0XH9EsT70vIVIBY9sISE2XyO38w6903cTdDy3DaeCW0HhTrvVHb7tLbycTiD
LbOWPqfhRpjvqNVbu86+IVqGPaZvFVbd5PTXmPPGo/24pr9dZevFFiuK0NurKfSRHp5jvBYAmngP
o5VIE9T/SlrtYgT64WxJURAfbMzMtKMpHk4CJMbvPc5OReu/zxIWjwRLahavlbv1IDx3hPPQHNbe
bAx9GKxBNP5ezXHf71UNcyMF+ajFuDqlJmqMmKYCmXQ2DM8drh8jlvSXpgrJMrgSrDYeU6oCDZGU
pI+PPfFUFVu5rzP3ZX/wo/umaHQXd30hpJguxcdeTGAddD4cMP4Nwor0i+t8LoE3YM+xb1NliGXM
8idpRD+bAIgt6KSRWP6lKERnk3E33uVPy3eqZz7EQwnxIS+r7sH9XttoHyCSvXx4owJRTeu5frR3
ZKtqBxWyAP4zLt8jfm1Mrq6ZlUFAbEG8sPrXLO3R24IV0jKTZqjzWqdQcz96T/plBaIm7xdNltWr
GgQSAujDFlFfA1Wk8DNRsYmoewPb5nliiLAkPbM+RQrbJDsFjDs4iPL3x0zPGLLb+21RkPoSqYSX
yjB7ajbE7IoRNRHluvFyL254RwL4FRV7nigVVk2fg7supl80Q1TXDy71jHZtDXh5zm3LJ3H1KEmj
0fY1RQ26xFj2j4lzo/IX2v/UeZ/U/9X/Rkdj0s+RTio6O/4PMmHouh2sQnBVqIrYb6aSTE6Mc3j3
PxdiyDVAfaMSMv082YDPU5kN3kmjpOZrvglrlMLXgPhjse/C8DkYBdT8C4IU1kPVCZmEJ8fK8cBg
QVj+TlusoZVC83773dcod8n4aS5+JRcFkrnhsZp8YNQgWcWsioiFGWa2aO+t0LZBnTW8difCYSfm
u7qIp90Rul731GZAV3m/tZii3zXDYSH5cD3n0NIA20apPNKiznyBkP+7n2jAmQ3srKXUzhhisWpK
uv9M8TKI3NkOMB9kJ5P/QaKtU2HtpS81qMMiuNipzqkYFLTlrT3ZAynjFhJWqLNo6UgrG1GTY4hY
VHSN11Ir7wA2yBaIzFbnDYyULNMAsbkGdN9ZZVq319pnZTdKRMUo1feqEmuSBtRkDVPry5MlghzH
uJEUKH76MwWMjF5pgseEUnJGRAU0tK4wVKoo6MNFLAYZd9dpq0Q6ryw2uQb5wblERjCFpSsDx8zC
2Fv8i1vs44/kqwapC+NqB96IaCtdxTipK3vpcBABjDDcHrfeh80wKnZ+vfOSAltVz8DWd2GfS48R
In/rQ7af8l7x6u0AyZs5vh3QnfYrnUsxG1psH5Y6lKJC4mxHr4Fai9p/MNAp7NxC9OCDirVjH5xm
1+TkzMXbtjjcMI6OyOjpvejVV2Yz3Q/+qKMAR80deqB96/j5aQ0qK7HeJuoYG4U0k89rJu2ppkm7
wdkHcRo1cEYqEemizPxAooK+kfcJIFx5JtueLxBv5v4TDwK8JZ6tzSu5vFMegiVYtUrISFqmhWZV
JxQd/f+dcd3gNX8az+QtAZ/VOid0b7h4eCOI9iH4o2qciXvvK52AiWSytPXswgd8GfC6aRSnOXkW
MCdncbNDmnnNp82G1JCfWLe9KDY44tL7Pqv1xzeijPHj0p7y7eDXcawRXs4UvPcLN2lmFOWQoWHz
xyk+JewQIrJq6C9JBMuRoFr+cL0VTeE2kuE/LkarbBXdSnNzckS2G/pQESdhk8Zysk53V1BtNkjs
1svputAkNoeLeLo6AAgl+mXihdLMpuMl35bJoH+3pIBz5YVFl/rO4muUTSV34Uo+cwl/AcW3N+qn
77XdgK9Q3UCsDMYUKWd4k8qAY12z3ywlmgRDs9Dtm2JN4VR2XsM3z+RHlF3FxTNDeLdYJzjR2t6K
uq75pn5VUbfxfQhRSsPu/JE+ICFDt3PSMYvCC21u3T1UphqO6PKIH/BY4Zkr4wkC7Y7+vIHss1zv
KO+WHujk2bFxdwfHbLpXF4UxEyL5mKOVebSJ9E5csyfBrwhelOMPkw3RqICEy5eLa7dpqhOJJ4Lt
HcyxJ9SPzZRcmPfKXChZChPM7mkQiXqkbdsLygVINEbiOk3n2xmeQUWCwl808XfrajVNtHC8qVVl
Vrv9gk+sgNBrMDD/DdYpt3uxl0ohEmWZxb0OwvFtH8UIHWkIZ++PmF+7gOvIDhUuvhkyY/PLGLkM
ILDaB5Tvkwgf3Btct0t6PHC3y1fSNQiZFlp4B3kwzjdc0/iYDi/DboqPGE5qWDRgRHaddU/eRiyt
azroTMKCAmaDu8rQpliWtIh48Ux2A/bcVRg9dcNqGdDFhS8naGs5orGySHWv2Y7ZoRWWPsZMLl9T
GFJpHpPZMIb4BlX02y0XB88wYneif4jYClyKO7h+r/RVurcDB+BIPuLtS8e+HMm0MyBMDfzUUGql
ERlUWVBx9n1cCAQq/+UlycLisUvHSq+LUWuRj2rZaSMx5AOvxd7dppHkXvfaJh9BEB4V1buiI9Y5
Nw+tDJ28fVQOeQtD/PdQ9NKL2O933cx9G1RNSMmU0huQj3ifKfAf9Ztrr1qpaDmLr/UAbB8yGhT6
V9lfKONjTQUTGeeWxpOCXCwKMjm0t21lBzNS3456773PiUvotVQ8rOw0Ky0qSodTv5S2vJcp6NmR
wFHlcy00FAgib5bHpwoCskO6IAHosXtLigU3ejkFHthTdDHVtT8iwVUk80KKxaIW9+m+XXRB+xF+
pSUz9aRQeh15bj3ftmtjMKCqRVYCSHS71NiKOE9oCj6/DLPgJwXn57uOzj6ZqRq/uq/UnNRGR+dV
7O6NmXRSvuRjwnk/soOxmxuKJ4TAIVCMWCeSsvYZJOxcB/cenTf1tvazchI7ZMo8t0YGlkdfSWjF
v9ASYeAqmnWV7pEcmZ/BKf0MBhxGtAcrAJ8lHS5Ws0r+LKIpRzVkO/V/D3HHIcUuW3k0kGBITH16
IoqLCf3wEhh2LzGBlc2U07O9vQUFT/DOXhe0yVcB7yLPtqbUsVaKQ5BL4FdL9ndB37SPCwYi/lgG
UZJKBE4mVlVzouS1YeQVabEMbhCJnq4fCmRUojkpWKtcbMMU8YnWGmj1FlrEcrtccViOaaiI+lxI
hqJkDspneXeTx4jBsuo2rKECfYvDu2ibt987TFfJ79IwXcUg4kUum1uY3rce+8ZWShEwKEOpehxI
ZXZ/D6IELs0ZRlSZCYp00Eq+eVEJZVdnt7hEb4rutHbV3FDNjZSHRd9UiYohfChQud2gV8fV/juw
1gm9X/oZf+zrPHESIqGnyhfORAdAOwSc2S7Du8afYUIPq57IQjd+tPPVtFKEVWO3VDqCqO8VFCwL
r3GZlmmqfQmEt2MOq058vfeuemz85EL7Adm5pkltO2vr70/LhFpzoapHbXJCrQVI8Ra37k0Em9Aq
/70q39pP+MoJiPGvTMIssyIqA6eDaxeVmJaiha5hpD8XlNjWuosYT5hC2I3VfKAm+2U/c5HKxXQW
Uy0H3PDBRYQa7w8aen5Q0Uds9xzgy54wpeFLJhs76p2xe7sdO23fzB2cHiecI56dM0BtUWmwZJOT
dxgEFlo6jcSLNQfsHMbbAczgPBx1Pu7EZBiZCZmQ00S0pUTdL8U85ta7+JHJjnfgy92Bc20SJ6OW
MfDOkCA6pZ0KTTN2bFHQIMbWJIpgbwBCAij8MePbnc+zV9qBO2ixPUYmdrrQhMP2vG7Rb/59D7sz
5f72sFKjbBT8j7gdFkkGU2z+5UyjMLEyYT+SfWMd3aznREYgHHOllULYVy8KGorQKwzzgCFatgwE
PBNm5GFJKRI2AS466btGdWlXFGeaBD2jw20X4vE8vh/qXZrkq8WT6gPV04y3GFrBailW2piqy5iw
xFQ572JUS8o/Q/HG0jA3Edc8hDhrTdJluD/EAgUS9cichhJ5WnPxknS5KlG2beLzrZ0mbd/zk/6y
oqGOeVGFGysckSVKAYbf3PFVVziJoy29/4PHoJZdOfu2+JL3EKC19/na0Yocg+j0txkDIS7XAdPJ
gmzCOCrj1wh0vCcJaQJFmbVBWd835ls/vM8N+rf7xDwWLiqc9O2FHbFd2aKi/7StJZDamZZWw9HG
6osOAU5axWvX8OLeoxML8XrxTMiHqLPz09vXzAUS8h9vtsJP+v+OoGpjQOHvMNN6SttAXDll2HKI
w6EW93SGLg07UARCPwazXY1aRHEvrE8YmguSm+QSAN6mAHi+hCNeuqotn9jtHBqIeHZax1J48IrS
YkBg0VDVQ6hVAF1g5qUNE1mWq43vmt9nEAAxLpv4NWtXfrsMu9LAlQRhaXLbkQcRBNpA/IAJp2EZ
X6pdZPZyVxvMg2qlLaN+v0hJNhTBggwZq7w9KS2isoLYnm3BZ//wY68/T2LezvRgohq7OoIM7FUp
3oDO45MuP2y39xTC4KC0WEvNsKkHum5cglikQP0gi4pBPIMi5V3mSp9axLfi1BP+nrpYe7FX0ZL2
K8Fl/JE8TSvTUZFUVhOB0fsZ1EOptHxT36ypMemno/bgI98fkJbtFi8ASR1wyO3yyGq09ZDFvyVu
FbrhAeOapSBZIMPcfENidEugc9DnjWn0w2TEn0X6z0RwXqrSo3zb/yhoUS5fETWHa93bBgXRA8SU
9CX9AV+VD66GLyZVwdTUZmwQlQ/0X6GtpRlKPnhs1KjQZ6lwk8i9c+iu3s3294oVFy19sSzMvEhL
TQX4HNMkjDnAc4sQXSNnUHm2sR/rCC9un9f4lj14/6QDg/C9f53Ax7YpbLW9L1lW5nOfQ9NRria3
0tCXcl1roCZMj237tLJPOh30DyYrbfBS5c0hZlJIrrlhCOxC62lftsyVOLDMyBbN4y4Krl/AnFLY
QjsYfQ+eKU6L1+SWIRc63KJH4gjEy9Lcu+5dHw2LxZMhQg3wZsoxiXIro6OQ145FqKEYDLi6CNQs
/hZJkrooK57UZ4YrtOycEvaQTOk7mokoTodHpTnv3ilVAu2olrZ3r9Bn0kY07R2/Dj+fCEneuDh4
kvZKyGeVM8thLD8om5oCOXdlnlMrWeofUHw12DlyZQeZSQncLck0Z09aRlV3WWZ+zS+bg5q6du5z
SPA4whPodkgSFZ2QoX5WuwfJpKrH7gY+gEJaXdYWGDNQx8e+Yqik7OBoUxmhvJG3K0ECjD9lv4sH
gMHXuNzuU69cBbIpKc6iBuxFkIZvGMpQ5sxKkT8l8Uq4sI2jv5+KaA7Nw93/d/dWQqlTF2laQNKq
DQqnPNyyp8nfirp7Qfl9fTCJuf42UpNHbcDkP+jUPClmpXt5ywMRe/DmjMxUMyj+sNZ6FmKs/mz8
7sr5KZBkJ/rm5iJ9x2yihlNS2fO+De4ItsWHrNuPBO32ctvPbL3IbtTumQbYZxfeemab7q1fuFqn
YfXSBYqAoMWSXOQcsQpkNGKKBWoianRnNU4Rqtsy6yci0lVV4dWixb4oaNEkm91c0nO1xxKBMrdu
pDL5LkghUsvzPvQv6/BU6vzVfOHhPJDmYJwLgbBauBM+QUjYCKxpR9Ov8h5HNU0KXSRok8tx6CtS
vb0Nf38NTgj2V7gHghEz/pRMy/cNL/KwTcim4Q7gHkwqtiRvK3IiBjk8LzHwUbbPyUs2Uv1UfLIz
/atbrVoG0oUhzhiHRIhpdjvv20hBMmVR+NdLCgxeTNhDk27q8c4Ah60xZKG+laKoqEA91LcbbAE1
hIoM1k+fMQcvvxkPh0Ttl1cN7Zvjx7HeG2PXC1/SYM1oAUC5O9J7uZMc17xAPuBGk1p0Y3g54S++
fgz3JIZalVcipjTEdT5zVAWw43hNWf9EJC8TXXay+49ZfwyiOZPm6Gnx3RrosrtCL1X9oy8EQKpg
y9GJ63Zb3zs9UOc4cUYWXhxKA9v/LsEyBKk4VHU95ZPd5LAofWjEYgfF8fb9QlQzQbCsNKTQRj1u
feOg4udxOiYPsQdKroFab91V8y3RpURjTeNZDTwTsEEjcgwollla/t3fH8KfPFtZgxJiaY0tP237
xgTWrT3xIJDDBMbk0hGUEGBB9KsltY9pLwAZCQpXu+7X6jnwCYuwrog3jF0IyIcncqWIcZdqcNtI
jpar9hny37Q8HlmUxVWneugYhtWvD4715oQBT3RTetvIAZjXGNnurbt4B/l2GD9zHOom4OBDDSMH
jx4BUqy4lEGRSbo0fyBFOwUvdrj46NjuJ8hYC35ovdETrECfs4MIVngMZBzKkqssalCRbji63fTF
47kGFDo/Y+2tzD3BC4jglEaLiPFkAAdxbSW2erD1c2BYFlR+dLXKRS1/pGOMFKkNypwVSqHHjImh
68bH6pMFh7tDj1+QLFfwTfbMnDBi40UMRDZg+Oc/IyRre6vb6yQ2Znab1CYAv6k2kclA9q7cnFOR
SPVVi1oxGYjfe9tJHQYVbpSUydw5XL5xW9Qrg2DCDOkFmec+Tv6g3mQG6mVdSvLrM/0MYOwF6RWm
mPo3+gf1TMUM3NS8lhrqZwC76BZMyQ/pPdiyKf/UP34tK+LE/PqWJEhNjPPwnf5D5oIQbLtF7Vz7
KAX83iSwm3I9qeXapQi4qdJbefnFs3kozdDGVCCnodEkDPTXb0nMMGphoW8ExowmTqWoRbOioGIw
vXO5+HGxbf894qqGuwcmGHnkMWOpmLlNTk8MCCQG+tOQn6FAcsHABjoEg2EMj5/8mqXF2MZcgwgQ
/o5dH/HacPkllHR8gs6XD55V7dIRoxR4pWfAqUFDk3fhjrx3NkgdZVn7KhXXCMiqVvkYG7bhH1b4
RS73Nwze/A3z1TL7fNjg2EhjcxtTZDxvL4qjFzRE9JPVUbk9yxTjI7fDS8qmiEO61h+wKis9yEzI
5ub7bkYGxJH3ik1S3kfmZAZCRLGukYmqh7vP4JQc3VVQxJa8Tu6liYJNOanfapKMb1yutrtxlkAw
pbHyU9kOrN3j8APB0RFafqVqSk+p91W+tXXUinxc7biGsS3VfHXqSvp5ONSj+1MSX++JwMReVReN
wxtAHqSo/ksmXzYHyOOKWdJhspWmpDEYUL0etuh+6X65rQ3H/bf+GIRk1RJTpCDpuwIwJVCn4g/h
tnTD/+pp8VF4KiHk1flPHWz0/OFp6ZGw97AjpCis2tQOapntFhrItjwABg0rlV0XEMn5Wv5CICI1
5IRToUB4WrNDd2QxAlObz+kox3YYGnb06asSGRrY4jM6Zg+iT29NLaqhqg7Tb+B/n1SC7WueX/uR
fGWM+IdhckaH3TrO9O7sMZi1czLO3WXVZylgYvv1OQ71tlPKnCY1L7U/5UilJBKoBcW27H+gSfkM
Z9GEfp7/1maYGAonf3vwLcF6vL/gU6XdbotzbpfcjtuUix5WMDqf7yYfpC+xjtj7mSTRmBkyfnBz
IFeaVs8uArcut1oNWIBE8Wy+94zqNu23sfKAxvLGHah3zCu05JoPLj08DvnNcg52AQJvek4hAGnf
li6DQFkP8Ioc85DAXTI90wkHokFgRPd5vuwoP4ztI03rJWqyut3zcg87mrmOhlUEjLPB/cKNb8WY
6H0v1Cui1LETOe8ESxBidCdnROpxbVTzg424WSxllxZMaQ/g/E3EzSoBysi9JBJ6mQMNxqbpHIm6
PBxL5Rg7NUrPlBcDjfvCSuhdZLfDctNmltqiXirEdiasUFQ6q66nXseLCEDy6vvQ/KdSn3IsHHG4
8ix6A3K6VwZmpDM0wHafG4gVFQG0q+H7Da2zdDuvWiBbbUxeTJRiw0C0wLJ/nUaLNaGWORZNSBij
SAjxSdfYRpFsqr1DHf2eQJc0AuenxhBA2pBpCYP9gCsGHov4dYQaqe2gmIol0FxcucoXpIlCb9z9
q4da7fPbjooY9mLCIEJkehnqqZhiRLv/SiuUfYUCwQZuMxsX9FVvANIKkamuB+9cDfMclXsUDvul
jEGzX+ZQrNmSfGn+cUDc5o/k6qFSvCJKZ4W5IqoEzpwGqjhQahDw7lx/tqfWFZyIN17XZ8+GPT3k
sDin5kGHRsxHscvthZ0xNWX2xB+ykGBY21JtEaoZ3b4t9DAzTLlZqLjtBqcAk8lsIX9OX7zBpKxJ
9xwNdc3lKtIpagvjZfzSy9jfvSLv4G2g+HgdTGy/mJXs3HUEfuz/1TSXkaZ/Ey4jNAImPgVxL/HY
rXrVAKHcwJ1Q7Cs/mZKowSO9loBJgyHBgtYDV/e08xfmkDNLP+HejefHbMfPxdA5vzJmBrpJpcWV
km+bx972y8fioJKF9/NcITroivmNAPPC6q7y9PNhIOXeKBZUZK5HMGOBasRib/AH9MpcrCa24zYI
0hzSFGd2DYI4lakNKVzjQIW36B/3vMdnAjAb8UcFkwlv8A4YfAlO5na0tI//hGFM5oPHin21kXN8
ke+3jWNIzFd5GRyzJaLDAhrefu1J3GOrtB2ElSoOrdxGzhmN70a3QCh8QMlwHYiqZBpEG6C5nxMf
tPDnjeNROYSq11K4R/jk+P0Ar18KLtjqFTeXS2HhFtcyXTmsNbUDwONXlmvK1m7KVswhhslkDf0P
oFxAuPya00Ufx16JcJ3ts2NaR0fYcVOX3p9AAynvmb3jQiDRBzMmu8S82Zs2aRXxJ2LGzl57gU15
PHlO9+hxflerlvgrc54vAgOQGhqvwg5Kyh7fCb7JfeVsHotUpBBgW/hjnPbrf1NY1BRQM8wn9b1r
Y8J/WuiHiqf4wrZPU8E37sr/OclLgflDWnoPUk5fBJVHjvcPTLJ7Hf0mP+oqlDxDtj8FO+rqZ8zT
BJb+F+86RcoEpY2MTUgSNw7JUSrI1BprwpejaZjkeWQvZyeIcNEFX1TmrDgv+sewaY2reL8dpZWV
rPTh1u5PlsTtgf33/jZ3zcSANvziB20lNBbjcUsnPpCA7VeErI+6u8EZqEBD2DTVAThrvYR6iXXh
OSCBykVrsUYRENpcZFdj+3AxcIfUKthZfJ1z29kM64uIHJSuzcNO72s0YUNIbAh0IpIt1xatTiha
XH5VOYO3/brMO9QpsOiojHFYu4n93ctUx+E1vSQ8+B/ZmZWphgDuDu13nlbtgynPzpzl4P+9gIlB
QP+DJPwAyQVBkvrd73FiHymdKsGFN8d0SNaYBX0M06X25/B/PEAnCON5YnHyvbUxIVNIpQZN3s+z
Bn9eWu4knD/+KbY2p7DgYEjaYpldbLvQIpRaeyWj1B6m2Bg7YJB6hGFuXmH4DPs+8fTg+Pkz2J82
MrFq73heblKq8b2+HQmekkA7uhx3qMn8kThDKiYl6hCl/SFQWq5Jwd/gsUeuyd2Nz2Bk3jsrVob/
77qh0G96UIpFXgkM0qT2g/qd01TdZnofz31YNyUMWmeBdhU9klvCiYGlWkGh1jL1YEpHkBY3d6FA
wpmJ1GPzdye6Unn55zUnVECTfGqK46h6Dk+ktRjcYTHUaT6bCywS6jL7q2XEmQAYlDIW1i4Ohuc4
e22QCMWiP8MtuSqkqgY+81V9FKHBkqp6ME/Z/4Q6hqsF7y5b79/IbjpsnziUiRGeXboTEdMdo4d4
rp4Amx/G4G94Suwv/97GX72y1rhGEFlUDAXpeHw0jU9pgaJ4/YWj9h/lRY4ut5/MO0tbXR8LOwlj
/NhOqEM7kg2nSW/7JuRWffF1UYl+TDgs8sNJCT3ulXGme3FFM7dFb78BLikm8B11WCgKA+8Rn90Q
zac9hxZa+UCfZcueg0ZE0uXQPaSwWqS91x2+56FuzlUuqTDXabZpGsgQ7dxMj2xANNqtccqvFLqz
eVaJk9ipVXMMVN/4k83CitvwbhP7L8HX9zdopcL2s7JIYACNKqP0sndTkNpVqH8hmIWg5AucwHNg
gmf+PziPSaCNUroVGBpzPJhQZg2csYcjpW/8MtP56ARbbSuHgbwSmNGuZ3td9c+PTCD9eqQMKLLy
9C5P5WAAIN+u5s0w/jEx8HSW8BawvEAZbdC3y/kNJsEbQlbS9Uwig3k6pV09CPOeXmSn4GoitFo2
O7oAt+UZgtBtqyfdqLwd5UCuGlgG6tkUI7JNM92CxeRvPs0MQkogK4m5V0n96wgkB5gTNtu35TBC
DEf3JrDICPiKMcMVz78A+1WNUMmGCR1i+VPISI33vIb6bDhRqnzsaOEpBKO/nmMQh+IM5fY469MB
FAuTIrrxv65eeFdNYzhIGjmLHUHc/5Q8CbO/KmpGXNMlaZS1ooRiy1wYcZZjWtmFCcgmQAXrNRyk
QZJ610lg1dYGxBxZBB5h5rOCaVwkm8oBBmLXXlhjbV/dT80iJ9lSRSAw1ip23fNFOLh7Hkndsrcg
BqcelAmjLFOq5Ed4zt+YJ//0XRDdX64DO2l557+a6O2GBNUSrSfN84KEQhq8mdhYsbL14DC1RoSJ
HyQN/SzhgYyjfn4WuA82wuUa9vkQ1fBvC3j2VUKie0wTp4Uy0TAEEKXyvmcWDLQgU60kZvBJKEgR
2jDswhqZ4UEYzASDNPQW5/FvdKpcRUF54IFNu/3nG4c5k5quuN94+co0OCy4WvcU0+hGhYxZ/BfS
0Jb1RFDFGzGuMtPF0hNFw8jg51yAQzA7oPeUedmvCQ6YtKz2FfqYsB+oppDRFmpuLD725SLwn4xp
dmjWEda7tV9osZq9jOcZy+0XJ62l2/ElXGt3s7UTO9y0r9Q1xikye6db/lb5EIAze73LRQfQJtH7
lzL+bB+eK8WOkTNFXBY4m4xzT+sWsMHpCdbWegPo/tKFvNjkFASpnEgZ24ARnXwlO6edS7/3Hxzb
VmARY+U6ngw4yIYgUUPoTbh2QZUcWZlGlmEsfs3mnRP8QD/T1YNftDBMC0ALkfTP5Z8OxvXYRVpo
kICxZGP97eQehxknqXvbu0vj2O8bYkFRcl3pjknPEaGhRP+JlsjOaNTCzLQ/IHdhdUiwQbmTkuJR
tTrmo+CIMt0nWPaCDb4Dp0rt+2oRO3VM+UxSsjlQV3OdLkhK6Xm4/QZrz6CfkMN9zhhv5O1SfilV
qxbq0PQUL9zXSsJehN55+k7T6g1+tAg4fX4MmeF7DdsgmwZJxanB1K7a3DVmaZBtq+H9FxkQ39pt
/2WKNpyuR3dgJdmY5A1sV0PEYJ8Y/T6Z4cXjO4hSSN44m2Ak3XBdydETqRQ8xxCRgJckeeaqZwFq
Ruw0chVSnpyBHHFtZYSfxhpSMD8sJNNNWppK13AK0ngSuBqrEvmXUoJwTjxOnUh4JsKk98jevUcy
UKA8XGA6Fh3lf3UkhazZkPy0v5u7qSsx9mExJVXszVwp1nMTLulk7rHpO7UM7F6yFc2kX9dMn8pI
OA0re5nNvmFZfQY+RbzsRY5XevvkZ5PIcxJDclqgSnjRM/X2W1OSngptvycgWH0eL2uLP58QcHll
kFcHOmfE2SaZRW3DgP/LLPUfT6yvFIfoaNol4IFnUJUnViDakCUjZpCNsxnAx/FycfaIqgKhLJK2
GcuLxUFB+jmQCMz9J+NCuErmMkQeO6CfYt7aTrLi3w6jjYu0Nnr9uuixuhhfPsFmzYg6SgtVJe43
qjQ79sv+mMujgS85SepoQdXbUj86VjzVd8silXjvBxw5DtZOzNqp4g9V6PQzkDCtqKzb10KZ5y6x
JW99HTPfUMsiiINfr4e+Vk9UeTMcXuOMMJLNBP7X6na2MbU4rB/9IdEEi0X4yzajEYk2BXXUaigK
OVwT5qyqV6sds8N4Sarqe1UeDc2RCUyxO5M/XxulgE5yq7cUzyHqv4tEIl1jOwhxPu/A+HYReW89
8nVZRdpTZzyujE0zfuzlLSQkEAMbWtWuZjZ5i/ZbzhVQuHMRUFOZBkTdNhekEMHulNYdnVemTIZN
uE5nM0wcFI+qoaWsW6yFJc3VvdW5WQV+bDf+zKkQ3q3S9PYwTzZuSvLKRAP5A5EbK40UbdFKftBv
K49fVBkDaxwY0gQabplCmFk7KYnZUfJuED7ZEy7jBXEtQhpzNvtSSd5mB7l87mtaqWV1USxOhhUD
zJi58QdhyV2RC5ijK8Qqbh5AISuGk2vxeuJyr7tOPX71C4unqWlnKre77+eRd2WiZVUmqkFjQ28g
0/zidhuSbV7gmfl0fWoXYuLGU2NyxftuMxeyt9R18bBN+sONwYEc0Z3OKHmRnSh0GtNB2AmkQpYV
JXhZfrbm5Nr+obkIjMfCeLGPPxHyZ0CdYY9eH1jZ5VYbQqNIRxtCyYhqIfg8Yz1P4PRbdBL3U2HI
c/ORScYggXo0OPRo9HLmddomQ4Np7XcUptPn/1EpzFzoXcYx5hSq2QnLSve/sSIJMl7oxR9HYePa
Xe7MYsMhk+l6jzQeOqHMizUzW4q9gWhFUms+6JsiDhisgAiNM7Y8/unPTwOzooA53OOjgiNfeFD1
zpgh7006jjAP196x/MnWyMDshpGLPopJRtZW434SN+arLN4xYFgq7RrHnmQ1cHXbrTxdCDHClg+v
Pi9Op2huPWtkhtb/cbKowd2CEenf+KZM02+f9aG8UK+pCFIWuiwHGU38a3FVVhZx3rFccGEpESLR
pVArVtvWeW75GcXOy4m1eawc1veOBOHb+o5idU5ZVPRjmm6QTQuQ5jviymF8Xcyfp11hBJB2fA7H
afrQ3ddb7yA9lg1f255f69gNEZV7bmx74D2zobekL6ZCoTjzdgcMmyoSsaJn2/LhB7kSUVlCGc0o
nni5cCU+HzJ9Go9nLyYNFhpFRfLszAN4EFvLD61Ts+ej6Sa+tMCKkxQF3ryp9CsYhUC4juxtv58n
rEbdQhD5avmU1HQfSxvZrMfb/oeGt/QlPJbSVnKj1stJfpBfUbyNqy+eYZ4IHKae3UH8/T2JmOap
KhKuYUpFd6jueR76gr0n0SIGqPXcFaAn/kRlkW4vGy13BaA5ykALPXycIUnjtE0OHH/3ujDo/2cF
ofnSV2KM12ZsrEKGLX2OZrE0MWRp+eQ6AR0BsTKlo8yOqLxkbuXFkTOGfcr2+o1kmHWU75ZA/ppC
zEcU8OJzquz/uODAAiTg4eVGS1c47ZkEiuu0snxEG1ReU/vKaqrEmd1NJlo1RRgSRtAwfJtUw4y3
Dt3fKXtasXf/XMFn0Un8b7fDZPj7HVboRLPvxJ1rtmcrtyCEeL1O2oPjSfACle+IoRG61GCDz537
vEfePJ1brFPnOcnnbOYE186XLS+Y/J5ixt0CUVKlO3zqTG8sI0GBk6R4D4GWFXig3s9lgHMQwbSD
zrvlUOh5gMckhDuIszlYUA6F13K9dNiojvuZSkLu4hJo7hYhRnV8d6q9alyNKcvm9UzKy4tHeY5t
VgwvYWZoe4RzLPFfS4O+YUhNumpYwgo6CNucn0GBG33UFvrb2gH70ZdhljR9TbiGhs9G9REi/2DX
GlxMOWPzolPAuhGm0VefLoaB8fN07fwn1K7HDclvHMyasavSWcp8rBk7tKGS26zqsVMGZAWbVQ9c
aC/tOL0cCHcF6mEZ2jnfxSOuqzp5kkUKA4zvopIVlmOj3GPoDxjeNSVW+B4XoRonJdg9yajrSnn1
9mEhqOlKZrSn4EpRhPlGeRDjilxmi2c26pXCY+7eTWH0sUBFtcONuhe+0xgIKwhO6fLIhRXM68PF
Ax1vr0KY5vc3HGuu8TQ/fbyu0VLjHoJZrUBvtdxTY76ipsUTQZxEWTP76gHYi/XYzc/G8C2gyKNf
VhbNjWwND+o4vOrKErFs9pQRJsEeNoBUR16KJ7ikDzvkg2U/zzJFkrEBNPQGB1F8DJvo+KS2XsTe
76Bbl/nuVD2bCUN8iuRXRBobAkAVSwEFSV3RCjtM4Q6i3YXkh2Guzhd7FawiveZtnZBqtC8O+xTU
GLgbOTCC31lThdegUHlSvfeJXzv/Xjut+AghD1IfOEOEFoLpsHo4UFS0sKz7NBejGkMPxZdcSBdU
8fC6vxBa8WWXYFNToPZ9hrC6s7ByjIpbHf5MC8gb1YBn0FVoIZXZRR70S3YB7vVwgGekz9wg2hXh
VVcbdhaPe+aVXn8AS+wfVTnltp8BxY4uw3m3Zb0RZ38Gr4VZnLAgk1i7rUHDAhYMX3Z0shoq9z+5
vTxh5BS5yV1j7KCRn3y12io0J2st9+Xla1E22QUPEkXRyT7hltiLmSqHIn7BUH7V3P5pAdHp9oxq
/vEeGgzbpFOevEPM5nFPL4nl07XpjPyXIXurpvTw4MJsqAOtbbM5DflHA3A5EyNRHrjtsnvcx7q+
BeVCxh3zTRAZV7jtN9y8b2NdG1qhYwp8ZMssM7ny8cLVKXSVcut28V2PCPEgXP7jVZSwUwyRE/VB
cGjlkzmXYw/cRlsGGMNNgRSsxs295sLa2tIyTSFQ+d6SLxfli2MLdDY1hPyaX0+NBaRcrBxSoCJb
tqRcp+6DeQwZXvdp7E9R8BbQPJQOXWzll0Ye9PXWb427FwEr78i2WsvJSNZu+JhQXtJiuJ/UbobS
jpA/8RV3NY/RQRGi0m8awZxapcCD34Y/afuLI4F5wPAjURj4WbJhAxmP9xYw68M3VNaizdC3x0BV
3sv6RRbxkzt0xt39/CWcTqm1DAYifW6xzgeXfZeaoEjBl+er2z/Fg5HRDDmHGWO+JAiegxMty2NT
GC575Foq3NJX4wTzSOo69AAIFgxCXsuIkJZcW+Ud43epq++pSQZM/bEwMkzd9eJdj2DrJbhV9gj9
mqlNLXplR7kU6xauPwvgt+pr6RoQRXcruA5peXG85rZKWRXyjfYST8yaFosbDgqua+yRzijmOcWG
A8ZHoudNr2rDQg3uxUnzu+r9eq8lkNF6uAN07v+HtRI6U8Ct8c8lgx7lU9EZ1MCRyCRu969mXBYR
3YtrGldNleLkmX4hNsL8RPleqBdoMQxNrwtAbbDtWR2HOdAELneJ/sUhfPcT5WoyVenhxf8a3UWL
FI4OPMAAH4JJjsm3VAhp/wKPouWJghQjPlBsdSosiI62FujG0ovYzPD/YJKwL21Filv8U9HRHn8R
obYN0BOX7xOplEwmJoo/4EUlPS3R/hV2IgSi0HlL58lGLJV04fL8G/osbVruqVK4xcKbwvF0R2kc
VGZqWENbmc6EqNENuSoy/Mw4akq3vaclc3vaGew+FpIRwb/TRMWkD6+HTdrN50cwOjkKbb+o3f3q
dQ1f7I8zh+aSLXww+4+giktktj8wscXBTXGdvUBaR7C3b8KjSzHbmoup2g78wYIv56gLlIdc/kMP
1MICIi680DjNuY7rXbesQ2pqWbV4KHRjpbuHLGupfimwFEdokBGz04oOFtO6RZZ3shZKQjFydLtd
Ph8Nx/rGbsaZiwSgKm3wTPT25qF3Y/HEFarikX+F1rTWyavmNgzxtmPFzbQQGGyPl7QYecNqQzeS
vQRnIilV2fLNdEzCJODCH+O0ZgOrb4DBPbx8ZW+ewCA4SitLB9F32GXmszgNExCzQpEYOQ/itpr0
vI5HNE6oWVUayUh+NLIf50PWdnna+mvKUkKnjqyQnw5EWHoC8FKRRxOR+cVBDOcLgucWrtxNC7EL
w0FzmEeSAOJsDn8yknJs/t5c3r1bbnYwjd2A+1Z7hyAy1/Q7D7NkxtjsHinGR+wRH9hFpyCXTiBg
2wSRXvH0mtGFHgqhZvPJFlDvwu1QDm8Jps7oCFQP5xqeLrAUtZqJmzzyn/1LUPeYTwq5GvNsco96
mLplmb5/rknRQ25lFPpjqblzP0jQxl4puLZnTDwFPvNDpf8JARQwoSh179BbAwtHQIWsrBu6WTWS
AAZtnLcOmwggGDaSU6ds5ItHHeCIZdoHkFz4KV318GiO6Xe2fhzbqv9bBg7Ojep8fd/ZX49OXTwo
KuqH7IdDPy5/vgd0rcj2nnvPxHYcLC1SzhapE6+/ZfMCBM/nLADxeB/DKchY/cHqIGIhaGGkRNgI
/bgWIPCtHxnzMMieX+RULJPAbQWBPRgk6aHyEKbagIIucxgGKTZHU1Hg28PEQVwKjjL3qO/EKiVW
mZlKiUKcsyHLolUQrRlIrOPkt5leBomCqiHeNpQ0u4/nfxYZOgugi2oautdp4PSPU15x15RNWDUS
n7YraEI9Er1tIBdfr9bJI8gpetPXwI6vMSafagcHzPCeDVQBIWtIDplkADgJvjCMxoKDrKfBPOi2
SSnOj9RoM7S41+hRBhDaB6bNKPoTK3J7uuivwM1MCf9BJr29YKqOmehMPIpl9vbK1wGelP5vNvAR
wNxVKnE/hCmkTTQBQMknARg/nGn0elzQqwdRoJOuiE5SiH+PQwOp7GtgAZ25ytFJ/RLf2YPqmCr1
P2jG7QbPsQc/qCGjP/Mim1v/c2ZY31yMbEKoqePtW0bVSNmtibUHgWcf1DS7YzfPud4UNa/de1pC
NWh1RVD3hryfFYLvky+c5/1mLt2uCx3tqXjBGza9Tee3mxhGUed47buwe/aOuKaurqhcodouk+HA
TL8Ia9XBX//6HNdpVF52ly4qANhz7/h8AZwMOKYLIACfxXOYrx6A9FZ3b5Dw5pHYrFMxh8+KAxGC
B+nPZKD8dovBRsWATzd+4NtnJkVSMZibpps6CaZVdVUGzIR8gBgLw74NiemrtyAxvnbcr3OJYrMn
aBXhekd86o/gXCPfDw5GuAhLR7rl6dNZZJzHyQUt+opEiHIiVzIb0N8AaiSB6aSZkRvMnmCrq/wF
eI0CXu7/PeqY68nbFob0Xr29V9f+0nr/ilpnluzrQA7P7LsuKsj+SCYAwRxqEs33S/aFsybrhb7q
OSFV2Gf0Ze8YwB3IEDJpUqKay968nZrXaegz6pA6qcGRl1YDIyXR+ac/AzecqF9zx8z83vExcgZh
vO6N7dmBnMb34K5wBv20uPSYLlXBMV2bq2UuTpXXJ2n9agTT1dQUoiRooBedF99girj/biH6C2lY
ADk9x2KJa7hSYvfJQmK7opTf/7bc+mkM5thFOPlEQjkC5EmF7spUtvBQQGxbVURi+sluWFxsGzV1
O4ZApPCm3dQ4KQ0YphoIyCnwz6LSKDlbcnTQvygxFjuY1yR1ogBlndINw3FVVDGSKYU8WdMjH4mc
EerRi+o4akpeBTpQ5SzKaQXlCpNyqRJu24bjtM/o49kNGs4myC9205c0BCyC4cjxShWVBW4+ZDzf
LiXPNvVoCQHhSOXJUCRnFRSk5H7acTCYzNNVEWk+PSdkzkVwBpHLiNubSQV8z1iMK6+sw1HCkNY8
65bS0qXDDxzNJc/l6LnKIWmH7plPn8foClgz3HqI/w6WyC1GXoFTbMfSGQX5bUVviv5Hzjk7dt/R
qXeGFLXDeSlP/bCbac5C8JY9E57j6Ma/0ua+y41MaC9BVU85iD3MZ1EciRAGY8AJfe5+3Yusi7y8
okNG6cPC+NRCULCBzpvNFgiSc+oL6vzXDbTP3XkMZYjYu6CUWvR9O+GTFmYs8kOj2/zmnj2SGuDV
MgkGeoX+GQ0ZZk5zBc5tveeJiYGK0DyvthkD79uXjc9pYlwFSY2lbTgf6Kslf5ExrpaL9YKqo5fY
a2YZhEjNyPl7Ci8WftE6GNbyEsW1DQiY6qlMBvt/FvmKVbSH4LdavLphq7H4DnApBa2NcsQou//z
4u5Q/h1OqlKLQCoLHjwSxqfRrVMjAjgNAdbNXg8gcVoBg8C+6rlyAcoJTIRl5q3vEEvG/3FCI1kG
KPTg+vnOuTzZcEfGRX4mKW2BJ2LdX9Nks+DapLJX+SxOsO5CY8CXF6fogol6yy364Q+xY+TWgwEH
NDE+ixEiIspPAm6zX2Jve5DNr7JbPn1AuPJgWOKVXKKwC0xnKz3HpMfx9V+mH5Q2Gy+iLOMI/DIj
2GZ0jadqFuHZsL3h9GEl3s2HRTSnZJTg/MPwmbRJz1RbTlu2eqgPcTvJ2Dq/6C8bzk746nzPy7bL
zDVdLsmIUSLzTvOuomh3MwCzfJYcns89OklSfD9VHslQP3mMSW6SL1XLG28sA6NmCygy5m0BVMZQ
RaFd8M7NUlgGUs4DmSaYYyirGUXtRz6djPTSixVML9ulULQtPnJS15p86vWVwhZ+wXibTvgym6uq
0GroKvib55wwuv/xJSSOJiFemQSfhnEUlbAXOhpFJVFgJK7BQ/hucXm+kuJo8KqB6as1ZkWk2ddK
VZrP0Thn142Fvfwob0a0TrgdePL2yIJ4MKRWE3ETH6WjF9V2KTkJedY0+YFk70rQ+Vk3r74qH4Xs
akVOrARJtPayUhTilMKQ+ika3PAHPdnzK/I0aVjghSalHf45pgvz/fCPfr67nVqjERo34q9QPTr4
M9BbHlYRdjkodyBsxlOL+ccUnZi95kuo4IqR2L15nW9jZ9BiRH1MuANI+SyQiOq5deRti3bhTGU/
7inU/aeBxAIOk1SBRGS2tumNSO7W6uNmVTTX7ECXZT9pLCUpOz6D62G0ULj71dbfXj1kbwZ3gn9N
yjmmfkVLWBQhi3qxugWB4VWixuCkphMMuk5IfP3qkz1/Ad1TDWAKi3W+jQSmqpvaKNBehjnfDPaR
x2VQo+nuZF09nfLLPJx0KDRYIu30JP5Jti7dEm1q+rZFoYC8/VMVKpVajM24rsyq8lzQibrb6RDd
MWvaOUB8O1UNekGPXXaBQFk3gPy0pFKvKjB2G/o+eegL6TwuQhc4LjmXYgpAEiLAtCNTqDxv+mAU
FdNv1J9Siqcofqm3FW4JyCzXC6HRQDjTVHft3Epj8T+qOUzbzOntmdm+0lNU40Mgap4KCKmn7X3O
xc21MJTdFs5KlWgVolpxBnuSurUZoPyQqTspjxCWs2gWkCnzE/rM0Xz2xoe98qvrUI+xXyz8PKEA
k0ObiKalL18mvyFXGDQ9O+HJeJz49mO8DpIZZmKY6ipgzVRGwkxdK1SN9HHTNxIVMyZ6qhtNvjI8
QgzKeEEu3mTd1N9wPCZgt0qMkMPO1+EHuYYx9WM50dfyox/fKGCfXSTdMss5M/W42S0viC6+54sa
GetpPgbk35ombp8cjbjXS+ysC8C3HGFGSZ1vdoIsLPKFziAADW5LuxKtVE6mSHVFQ4MXxIOCW/9I
/8hRaDlQjZfb/4oLdM5sog9CCfZTHmj83SrDTghVVlPJoYYIVIwIqWnqNn1WQsyHkqFcDSGafBw0
Hgx5brWCzc44vF0KqNWtKr98It4HHRjyhX9YoMgLZ6O1iJC1GLffo0td5sAXkEvqLeKeos6nG5eN
GXX99cKdyi29E9a7SSRPPTXBuWaJCym02cUIk3tUJwgp9eyCkG+Dib5B18zTcidnMZVyxXR9TOTm
o4l8seYE9OVELyHsAVPcUl8yNAUTR/muA66BHye2F9qyRaN8fos6+znEVuTX+/kMaWrO2Vh6x7Nr
o3/9KJ/jqkGzwxnWl0fGBltZd/vu2ZSAWF05nACwXJxQqwJMRgtlioxj7c5g3cxmoSGWbHuIljPo
4Wj0jblX5CdAiqcuxhirYFP3HSgpexjTlWl6ESwuLfVe69CSYKpdSanRWCu/YiNc8YmXER7Ty/Vw
QnpfCNLT8oXWSm5c+kVP2kH3JN5etQpc0/ugVWKi9iXADASmhLPlfAfwSlQSg2iXEabnAc3zUrLB
ZgzaUJraGejQHODtJCHrwxC9a/W08RYGNqFU/Rt1ABa0rnH08cNcW9z4/+AZj5JQEJnedf5f7fbZ
f7dGTmvWZdEbzTYbXKWRtR6zOVBuNhPDcY68RayebX5Tc3Ce622fkQP3K/IDlb/fvKRA1it24QQU
l1SqTidCn5nGp8GlOBnhqUWR2vvy1kF8WqrwlITX6OPZUSiy+vLGu6P0HNN8PxidJOaJUHyaaY23
57IXdNjJlkql6x+kOwZmCt3k5aIzc6JlGm2TVSEBYUuanxMCJFHR+N6/dTS8UrK/qvsy8qUbLEb6
zn46jaSgdkuUCqO7bzcEP1ypQXY2Gtz186S6KeC/nrivBPOvatmTGsRCfbSO2rF3/2sDNNoq6uBs
kL/OwWQN4CBH1gQ/E7TfE+U7wLGKGeBPuejoimUTolyQ66OLe9HtPciEAMbGCCggnuc7RVZxgrVN
gYc7V4ZYXakvYNfcESns4b7P77v1CAWNRPQo6p8xtpu0PR1eEVmRDzzdYGOFcTI9ept7yN2gjO61
QehppdxXNXr3/yQKDkFM/EtfaBo9NtGp8l+37UE5kvSNJYijzYPAD5LRoSTyFmJguO+k9RW/L2gl
d7KWcnGP4cS759TDREtLEIO2LJ87SSwTtXBQ1mWpDyORE36whDoukMy5JPuLcCYWGnkqasqwuQ/D
odSHZtnws/Go4WSlvQNgyQS7UXXw7Q7QmjSPd99HCZ3N0qa7IOePUjkefdMy4I8j+ktqLcUNrOaX
YPG3HaHBfC638mGjASIe1m1CQlNcApT3P8arpoVj4LnK/FgbNWj11+cuw5scuSbDgCANp8p+IugM
2ZCnvQ4pdnd7BhZH9ax+GgSQ5CWCDNk+6PaCOc446SE43dgHo7f3EnEUE1VNncB4cWrBagtLtt04
n2D5oHDnfFmPEjhLKRzerjJaUTjWjvzaAOKvLH3DeazXtqQ7EuMw5quD28DXuUh01kQfIoJ4v12M
XIJNW//e8JzX2EwpsOf8YexIRJ0XkepEfXhUdOaZOFdkmekVGk2kusv/n2fbEf9tfMKFCPvX+MDK
oPXkvcYEZjNT6CjyObEcTDUsK3TnO1Z9T97Z9i/QOstIc6Th6K5CqNPQmHSXEd7w4qTJTIueIH4X
JeuT+sViI3sjPwzmzav9YqSZ9fDm9ZsMX8xqg6RNMyhzCDEJckGWgToBPrvQgowt003tTS/HQ9Q4
H3SzgBsl8CkDRHzF6l2F8YE5Z78rhfD5vql0Ur6f5EhhtJz8yMg6cozRVCDt/jXWsw50xxuPbiz1
Ye9K+2x1caIvv8hRi0pbdifoQ95ei1WluI+Z0NorG8bp/lTa4jWFZ/mQd10wapHN7SNlTapB0KWt
CvqOvOOYyfp7n4McX3wRZnMejLmI+ehjzI4/eylLlu3D9l6Diobu2W+uUTqHkM8nodYWr4hPXeB8
X8/ooCXAiF1dpKTSS6L8MDDGWJk9g9u1EEgOB4Flu2hwvPnZBijcOIkbbkP49krnSV39aGXIfuh1
B4tnJW5WlSnQbhph0zuF2fJSz9byaHoEsW5YDSwgPo5Y9EKfWohqHixwB+4oSivWNxPcnU2JYkCZ
+ZMdmBwbhyY4Y1BoSvubWRdPHm09Z3r/XM6F0t6607PTQIuuVwEPFPrAm3n1BV/j1GfMcyI2SPxk
yxo8shhhxNc0YQVMlTBzxb05F5uxFmloem0RkA8qb2RjnxNW+3mqwEfcBZlaBgAqO5FxNGj3rfLP
cQbLUjA9TcVhko+7i/NyFN48+fCQoHz2taGkxyESLT2mJ8ERvinG6DndHJ6gEqcQHE9E3N6d5irM
GRJdGRah9B3UO2L+koKTIiYwzxTf0sylKQhC1ZpLth0xZ+/2jOwtoDlI4xWrkYSBAd6Xj50sb1Ij
XUUwoQDfGOBymwEu0ZL4OvjukI60PbprntYBhwCw5HqFo4sIslSuHFN+v4oJJM93CRgRGXucjboS
EkD4MvmN/4uBrInC6kprnn6OBmqSUFnm6Yx70v1mNfoRSLsLa4mkUAveYIreZGXDkchJ0vTQhuXS
tueYnwo6tLIjNS+DUJ3CxBHwHTsNtN6Dr3ZzNNSwYdvx7L1eZCRS6DOgUngmhI04ZVDlGtdLiYxk
cpO/7J3haj2G5hQEU4F7DE6xaHw0BganR/eLH/3odKELVmpMofKvx6E07ePSuXvLeT4IhMKIgOHg
9ElHAvslKwmWI5w6zWT42GkxDIvuSIGCubc9tSS1EEKZBnAseSLUAks8k26fNwxbPbC/tkt+RW0T
jKnPxZ1zeSaD47vNDV5+00KtYzqSHm0WeYA9oHSlwEhqRtdUPJdTPZVXdx+WICDpflIW5rk0eALt
rWgLH5UAI9K3Z1yyNetY4XL4YFb+uNSnM6zL+gopsZNtqYajbYpsj+cQ8ZIbNOfjyFnvqa0HeIWa
AiWnFVG15xD9HAgHJz81ACu8IWT6qyUJFpW2xLIkE8t3/D42iBHkdrjGxYqzVRFKBkmcG9ABTWIZ
hOrrQ/6MXGoDptDBrWAw7Kbq4iifZSyb2z5sFe4qaj2rJfBumn6Ucd0CuponGIfZ/dCY5kZSouR5
a3irx6ZYYzljTrm6WoYSBUzm5t043CdAzchX6XjI2wIJeRTm8QbDMpfPMEg7VkZFVgVpyJpOipeb
q2UiUaWCMIEyyD2uy1nD8toQ8mDT5EAsBPJQera8auPmq0Dqk2QAWLlJgo2bxvbjnbaJ1vKYwro8
j/RLh2n+o4GV1fvT6vXGql6nGNxFszAPCptp6/DJgIAGUosP8sI0uYipO+KPwkxB0iobt4W7abUX
nbPaQQO2IgS9a9hD+PCcssIkJscC4LrHTcpFNcO1+QMEX3tou19GlZYg/9vpVoifnbHs8bvmZKRu
U1nsLi0wDojCA0MkxidfKip1Neict+SZCN1kXe+YQtGS/cqtWI2+bIseCjQ6M2POiV9FQlmNCZWK
pldShiOQnLrW2eb50Y52IwDcOtjPiMuB8jN4CmUrzfxwa5VZXWncvscF2gB9Q3C+T+1hLhG4adeS
r83CoeOE3tvgkTU5AMtJ2hASmF+k61lApzZlQZh5LCT1O9HVslSHryD1Utn9mcHuLCgZcDK/8m+U
dDWJxBLBB5ve8DtX3OxFwbQ8SvI87lxKeD0YbrOSy0SNClkLJHthQl8sey8GM1TZKTi5uOCNDgHH
R5sFT7RvZusz9smB8W2bcFrFfuruXKvmQmGsmKwVWVE2Ui2szBOS+E1vaai6oTk6eMUvvc4grM5R
zPGtDJMj9KJRtnGlJxVKl7jlfupCbyxmZWQLo4SlcWZIRRkpzWmxuvDiyvMZibJGDjdN7whGGN7a
cjzd/vf0PDBKJDzfo0pcW6NjowWHDvT9z/r2kEgQoAeJT3yDacb2+8sqr1uwBXBYXgFsvSwiFSc2
cJvtljJcUU7FjofpmZgEfpdejJuRfC14UFDk4ga5/quc+NJViNeLfya6YiMGh+9uJ5GMKqOGe7gD
F7fB9DVbuPSZ+K1EV1ftHRytGZpLTZtCkHt2wbHW1RnkqqX2M95SEECbt6KoTjM9XfVY9ZZpARs7
JL6bV7sAdzMGUtL+TIp435lGPOn9SrdqBLZ3K8DjuIuw8MTXmHWLGv/7dl2PwZzLoqIRwpX0Ee6Y
kM1xeaqiklHcPD3knR2QaEk+mQ7F+TpzNd0Yb1wwmdiiP1PDaJ6zc+SRwFdr/Wi1FAmhM4fqEvfe
EyykUVHXE/TFG/qqnV60siEjdl7OgdGizVDuzregLrBtuYmJnouAXhEXlBpinF1KBlJfHp7z+5Zu
jGTPEhPl0i8fdzIyQHSnucIUR0FNJrnC5QEM9lPA8GIFSGU+YzqzAvK6tBGwiR0P8tNOS8F/aQ2H
p5UqIEFnAU9e1aS/AdfOQq0E06voE8s1qe6+XQxypzJETz5R4AuDiwTDg5htUlgmQmrovoP5mXwW
gX2tBk5DQPILJpCo1sIpCCTsODrrnfTe+Z5K/xCjqC7//wuV+Rp1i0yXYmdM71JcuiMXcBnR0+hF
QPHSB8YQh+O7LFNuQ75EWowHT2KgmZtSc0949srnOM9r1P922k3Hpm5TQkkJxOevrsrZQ72tuXFl
C3DG/3vsidExzJDgECYXPIGtz7EqZKIIGk9pFHsEqUztzZjcFQW8GLN9m3WWgoFOux/kyA/4rrYR
H5nM6AvI1TtWCe0CBG6OTtIY4fCh8MlaCcv+EqhDuOelCqoZiOPKKrtFFp5I23RkQ/2siIZMQ5w5
mQy5CZNBC3M4zKdTQMMFeawuOyKkHAkkeXXEJWZR8DL5ka8rMbFDtVzEUREnagcQYc0RcMH/gf4X
Fj6v1K7rjV5iNQgpPXIi03JglPfJlqB9GDRZ2W6KNCQXcueeDlcFk4+MINPq24uJjMx6vKH8Tsjy
4swsY60CjY3vxxR4a1x/aw3/+MceR/A3SRwF8jG4IueGL/nOcWY+lZfF4xg3WSsgNBefpdGLhT13
QmqDokuXXnWE1ALRc6fvGYaOHomXBOocVKd4o9+6cjckRKR5c6R7HW/I+1rJnY3w2irI3608Vfsh
hnifVRX+CLy6aaz5+iyDrJmISQHmh4/zt/XYL8j0kL0I5Sr33nZyBebIhTN1G4QoTfGT82hRtktI
43EfSqV0+oys1NFgQcVk/acUppXuhYW+WR1cbrJS+kj5sgvwhd3iX71NipbqKYL1cr3iAqh952NW
9k/WlL4dw6qlCv3IDaKL21Tt6GUNPLqtm62Q3Zn6/RWdh1RDJYUzybhpjb6cWyMIIWYRTinwa3MN
3P0zqG9tial1FWRfDUxB7zS7o7wP836zkbosjeKiYDZaeHrJY0IW/ynpleNXGImIjuVzZ0yq09r5
ztKkT69aL3na/nnc4JrrqwNQPdv+48Gydcvb98W1b+vzKNpMKsoFhwyIScI10dQU9pg+CH4sfXD3
mcMrum81dogBmeiWkcobCmZYHFqyo7RXM7uE8XjVL4jaoRTtUxLbGUSL5vgfMjyqbSVCKXRAWBo3
/nhagbEl+pehk+NNQc8EOm+lmWQtXS85E5PbWSfm2rCShf3kxM7gj/Q+/HDWYwnZwXYb0HlLxAEi
dbP/0IariYIhEdPJiB7C904p/zsV7ShujR9uyJdWFLRKLym7R2Ko+MyBdcViOSOeWSEUClQm1AY4
zf66Vx1EowI4OrQNiIxUNv6wLqEH9nH5XxtzSadpRJNYdicfL9DwDoOKV0bsxbBWoQSwt4fCMUax
sdzjYWw2arc1Wmr37nrqrlP7POuqYYKOcMaGNakX8E6Plgyehf8J/un/p0qFhbdZEV+xNIvZiU2y
Mrarjk8atbl9/OcX9WcutLAne8HXIoRDkl3s/4n9cMhLnaA59R5mkXqm+CzmiDmPjiDNyvN7N/bP
Q7IOlDXgo0DB2JNV1EGJthk5owiP+hq0CHRJYX4e4dyDKmva3lttbTb92SxmouBIH+dCnH3/QQj3
pLWPZgOi1Nv/6z6ODQVa/aEipWfObGZFsxI+cArT3FDZboS6nxcClNVKbmz501uSIII5HERGeHfW
ba8bD3z8sP8U41GMRBoVH4uUt3G3XEFm5ZqIMDiIEdppA0LtiZpJBkpml+ouUdG3+4sTjnw18WM8
00wGIUYvYkfcGPGcWWJ3JQIdOSNApEIcAK+7pZz0wVE9fdV7FDc3jIcBKhyyhxwKmz7o+8p9g/Cw
1/u73CnqnuMCYvTBf6WIDE3gYxyQmO8PDTt0DH3A4z9rQlksqHbUnLQCevbLIi10n1w5glOrpz5Y
0afhQAg58CJO9OUQkEq0R7KXTVF/MIPDiyvk0y0NOuqjfxhJ5rmjIBh7kB2Jv46Qv6Pm1q1C5GSf
lxlJq2ORqLy3FQLyGD+ve2cqo2bs4nXOeLI8G4RsaAaLTxWe9ZbsqJjOOnztM0kxzdpNaIo9Lse3
2A6xOdbf1F1COCL3jggQDh57K7UnZLUbv17HxZloJQHqoe5qHlv62n0HZIIgSeLCTdP4PoxhQ8u0
Xs57rryugVOU/NkewfN7Ddrl6LesExm15rB/dc3OJofnK9sua/N6M5GTwz2/9TatZboG0mG5fcxE
a1f50JzTpKX7u/k2+DaYKETtAtUYTsu9TmOr/HHaPyTsKRscdbqcoYGh6zUx70+ROWc8vf1othIg
zSjeJ92jpWGRigYwwbpJf69TYzclO6+gtZFM+T2hk/XkjgNsV8Xy0we3UQjxM06O8pLFwK76mbJm
WUsloj1Qum6DqQHk45sxhqjK1U43kK/6ytsyDYWGV0ZNc5Rv8oICJU5pMOGB6ibgea2+wPtVJU9l
VufvbS8lfcsa3/Tqu9L3b16k6X9xNtNmEMfyZ9ZlDL0UJ2K4gMVlb6wITrNhVGHnCPQYRmu+o8Ng
SkN+MedUAksL+1ZQ85SM/fhaiezl5q4aTtTqbdX0C9H9Qi2WMds5U8c9HqY2SDVwVdnP2Md7pnBZ
A1nMBETMv/bZvIhIV2KCj0doLz+4LqNhiqoKVJo6ESA14iSi+GDa6VwDiXp/U9xPRq0gWzMQljlK
NDwc4IZUan/4r9Gt6edPcgoKnd77WaDlEbcqDvxChOnfey/+7DX+0JHsU1V8tu+OXldb1q4j4F1k
S08wS2UjdTZqmaCnuLwxWKENibKthpHd33XEKDRNT5tkhnq8z8JLhxKFFytaEDj1nAbm3EK0dX6J
i16tmFwHIoOo6NN/IjrEZ/BHcJ7r8pw2i6PgxFSzg6ycXuMdtx2Yh+dF0LuSFaqMPDMEC3nzYKej
29ZrjGR6ws6Al55nLt2xyypJ7VhzC4agk9FTDh82a7/L4vqEjnlzlNaftwO8mEWDIdh2idkLrx4z
biiwsYqkc+2txlLnlN/RxVusDhJ71liBi11WEUXiYx4HKnW0Tv/VoUQ0CzOY6TIaSIZK4Z3yD4z5
i4kj2BayM5B09dD/0ru8tiCnEG2rLEkpMB8JgF42UeuLycmKws6jEy77O99dvODsn0nrN3GevGE9
EOVIREn/L1uwm9JR0T4ATO7O3cDv/T4rzQEGcf+3tLjseB9MdvVNpgJYJzTlHoUphUJwvT9TSssj
brwbux6gePoQd97KdUJMKbubYLplsjKbbJGB7Bnyk86Bxbj5VSc3b1EpZKOFi7SRED13hjHNuQsS
M3Co6oBEOBRRrJEXLH5OvQufzKhtHKXyDN9E0ns+Clpxl7oXvruYy9mx/3m9YMdkinUrmC+dw4FA
CyL5XJMTqVwBn0Xq2QktPZnWBSKrqnSkRAIUcWzjL0QVbPjuW2zh5qNjmzSRIUURkv0PAaQ7L/Aa
WeaX9286kmyG/5Q9fkrtzA+ECJSqJE4xqjsvc3/TXF4tpQ6cGCnn9VzMZ7HdFCwEuktXWvPcoQir
K/LYgd2S2paczhFsh4bl5Kf5YoIsz5xZRZAk/UCjQ/M+AdRynxeSIRy7pZZxZPn3/eL+VkYT3pOw
PDhdHKb6Zss1M+wgbz3euIdbv31EbxXfsnRwXzD+FZqr+qJSWkK0yAIHEBmrooLi+f2zv0gXZD4d
B021azDEqG1DfkW0k1YoGsH2qY2ZE4imduvS3JeaLzHsIXXqAog+zBYL3EBezXE6bEi68m9GXQHK
QJJNsxuza+SOdeTR2zd1DA2tZeLsC+5qyB4D1pg26hXoOm2rlvqEHC5p0BSYvg4fAAEwVpDgp4jv
A0wX+xo/KV2/vvKbPmmTip2re6c+AyMNqY1dfU2AykGuCldSaSyZ3Uy94CA6V6SC2e7EPIVUcU1R
STTAkbht4hJxxnlE739+bCBnvGaq8ahDOgNUDEl3Ofdl9/wcrq6kXG8RSrHMWYIXgl8v4H4agXMi
cPWurAZVCEwJjLjqI9WkFIl7S/ysOerRzhIBdrE+ShSGH6hUEgNp48hPIoNc/hKtRFQeUrLsyPTU
0mEKUpW5UUxlkjWLhyRtqDOdoBeeVXDn7/3yUuLfFZsWcwAj1xtmMRWG5/ZROqzbLaJ2cx0IfBim
qDA/kWX4R1m0cg2H6/f1OV4SOUp4dNdiIPMXegJx9BVbtgxGuPthLeSk3xgr2zTKB1Sjc3Y+LroI
mma9YBkVTcTWYarB+vO2Gopu/oqhuMF9sCJOJAR8zr5+mJhyfttPzlsQV0RlqzgEXouffhI8hia1
kCnTAO8cTeQaHN5ogNcw797eS60WfLVQme1kOw/CyTNQn47lJLzDPLy+dtHzhOfyn2WmfZrrMmir
4r5gxPpNzsoaB71W0m6NWOxpzeK2bcRPz+X2vVvmbLNd8KbNBtePRT4H6QIIMe/opFPY/IUCBeh3
+9OwhnuUe0wdkArwtykuwNVDWGHJXIhdwVA3blP9Im02S2WU/GOjkyRKD1oriTHYWvmClHjSMe9K
KcYKtvJgY2eqXpXUu9pke14blNX58GO4W+5JOcmUwIcxr68pk9DlzifYeALGtLTqIoPfYQqdxOnG
KSFsIVfDSv591uVJ+Z9qMHX6ReXleD/llCT+o4eg5Rl8MkfqsOA7i4Re2yInVsxFw8DY3DZu0DFt
ZWJ9kj4L6oiV8nJ36eFXXoEUtknAoH0InZyCqZO/i4qGRpYX0FhSgZxU/wl1/aqkQuCTZaRsAyZI
n7teo6Ncv+/YsNE0CURQl/7jm9dVBFOaAQbP6RzdVxYYrcD+H8+xYB6kKkpfSUATC6A6ftAbD4pq
EOy9N4/HaR2qmm2JtQCVsvLW1H6x8Ks4sqzygdVkejAschn2XCEQS4cMJoUEshmVfBhv0WL35MUc
fgnSgP+5mVWTvkVzYg58r3UKyI56X07UXgH6I7YeE9laxVAngm4X0QBoA9ZReCeAIqDVaf9LnRhx
W3AIksvMOzrVF/J76LMvqTHrTW5+DNpIiwPuJe/x8NJ5MExfQhGQrjaXkdiewCkVdkj75RtPGoQZ
BLA7ETkeO5ha/JQXVDUtqw6d3xsgt8pjrEY23yPM17aUeT19H5B2Nu2z3fqVcI6h4EhZYPjDsEd3
f4qZHHBBl8QmzEgD+LnClhFVVdQ7Wt+IHHCj5RBBkYs8Fuobb69SQE2rqEEEOXJpq0uzFG2QrJUH
rMKyNVTqM/zjHgFBJyLyNkNSYg+zSeCOCQ5FwV+2b7SmRM5ERmwkw9upwTT+23gE0SP0wesHwItV
ip/0XXpl2uYKuXaCLzblM50qlwjOcbW6Cdfhgmd3IFvBIhv5c+kiKW/Tn0ZwSsfy/rzkDs7c4+al
ddtg9uGEA7fmEvAyrmKVQVuFII1bCxhgkzsO9mJtCP9zqrNQJnX9wZxkQLqWk/HxEl/272sKCvQw
j0K0rBnnUOuUS0AYB/B812IMzU03cHDQuOnxhbVa9NKVyjXYM1T1izapR9CwWWqxnIne04JXAivP
YHbBf3aXEeLGxoWWomMl0y4RQllFQ+WwGafEhlUhsXkLVV3Dd9dTJ/XXX4SM/SimS7jrImagrHuA
ioeid7AiBMkqFjVFomVdeuvsrwm3R/dFAx7nlXJM0ImibLCH629hYNh+RVMGIEUcwwc3aBfH8Hj9
tJ0KUFlgYPV/lvley7FqqeLkzc38Sb5LFJGQvyW5IBi9L5ZqdS/I70KirilVn5dQObS0Z/9rn8SE
nFuiNbIlJUNESFAFuqTMn2vs74I1fhHkdIRcLKLbCwtDoa2o3HiC2vwF2cCsTvLSakvL0skw4S0W
IT+asB/FV5kKWSCUOMiW812aGxhy5AigyjfwwsKj5Ca+mnjoKauKJ22SeNq6ERxM5x0OvMlAy5AE
ksmnxidecKDdcJTI9Uizd9RgjDkLT3qTZxIjYu5BXJpxV+ud53VzBwiwJbM2xqjzfffSFDBoPM6W
g9Qq3tsJvPHtmb4LyRjeRNM/BuezgOJMh1wJYy8YaN755Z/0pYEn0cmjr68rYztfK7f151JhT+dI
xtG8zKlmotSA9F7jIOlKPEgfEvy4Z+g4mecOs8SFpM6vj+HthK/2tW0Zf9gtv9PdursO0TSRySlU
Rf3CH7uK8qKHhVjoFRCoUCO8iUo7ht53zWQzsR/4DGAac2rX7ljmXLDZZmVW7Ev8+5LjpXSI1Xo/
uYgh7q5vUdHH2H7ME3eRtSOijHh6pJqVShr1b82VBuYxpzGMnaNWgsQMlsVjuJEXq7gynZLHhdrZ
QGotg8vTFFZDFOBgWEFAu5oB6+EJTD9DuhYDE07dM9UKIT5xKwKBLHj10lpMdPnUsgb36EmOkVKK
/XoDG59nGzvrJpMHx1EsuqP1l63HxldmptMU8adt8tl6NGIY+gVRXZv1qQLyFRuoOCpHFcvmlT/8
yrOPEBxQWI3IhOBLpVlJoio5+1I0XeLaqnhM2eLO+pgfiNAuNFnNP7jxS7kuD98ygxSPAE8jNw57
9koJDvzrAf3HQDfLSizyXofc3YKpz1Smma/XELxRM1QNqC9eFHc8g0xccpDRP2aI9kFVQfjOKMip
xGYp84Y/IPnRqBWCccRaC7YEB2Gz0uKyQNsAIIch7jcCZCftgc/JNApXZKVQTt0WgJMvjgbm96en
V05F075zjaljqwoOCg9FrCpfqoMNR7ef5wVidiRp4jgXMY+VMvWVkPRZ57g4meKB1SJ1CwCboS93
eWq6DnfC/oPaFIAG5IVP1CwyUMvgkmczSMtILpBwu4mTk+ijs+a8yf8UBXBFXIrwJ+2KvE92msNz
LJFQUDx3wnUaA5Cjkjenkz/bFFbtJ8NNdpQTAPCMb+e+GkBetl19N2NfVhVeKccRaLu5biH1LJBe
hxg7ZL1FCYOh9mt1wxkhZa2Zl7CDyPjG0qYlv327qpKDM4ysJCaPBckOrCuGr2smEgLOruutluWn
IYuUTL0S+xfBmZqULnMZTKSNEHD+DVYqCvtBluNrXPVazaLYfr66KJxTzsHxkYe9mhcsj+0EpoN2
WXfMx+KUgBZxqm7Z1UQInf9lWBLb5BvUjrVXfzDmXrtiVomYhZ3p8Xz16t03fMKdCkMVwM4K0njM
rkgOKsWO/ov3J8eOJhyaITQ3MzEXZ0Qpg8Mn0SBGc87n/lDIcd6KyiNqaI79lwnloTqsAgc8MWgX
8SNtpWjI66Raz4iPjU85dJwQRv0qxNDkimEK16+9qR8lW6wzkC/zWZXInYkwKBNgcjEjSTI7Rwer
fLnSCxXUf1ElBaWLB1bJH50OJv8ba19/Dz5WGqDt163u+mdgqInT819KXvhvbfN0h8UT4k43cudI
4Vyp5XZOn7oV9cXFa4uXAkO+B33GIPfn7qdDKWAXYb6nDm8kOqKNLzFxR/ocOQJl8yD1rhbsYr5m
AnON/uk5eH2fjog3uI9wChPfJ/DcTOSVsivTu6EqIPz4kzR0EQb23ZlVoo1Em9iQeoB7Nw8g3oxe
Zb9frHX79C8ZQlwp/wgODsZfO/ZskylYaLiyGqqm489qf1u1bwm/qCeuxWbE1gyLKiBl9ukekAA+
CCrWaLjp/OUZJ+MxmulYb7ZIwpHAbYlFs3Sqolv9yjAwJgdzPiEVxoRwnAFpoz4ZLhm/wst+xJ6w
zOCxOiXhDgWuHF/UK9XPFGAU4+e5WjHekdk2pgFwhHzRee3VihIyVfx7Rn46SFIrtMqHdCDvTf3c
zQoC6evQ5avlY50f+037CqzQQL4DowGkTHP3bom1E1znT1m5UccQloIBCdeIiOpSm0lhvnJHU2oN
4JtPJELpz8IEn6li+Txp/M/2auKBWfbbv6/sp1FDnzVBpfcpv8MWi1u4AI7AB8bELGnXphzYJQbV
OBSaJuacbHPm0w9AIxl5F0cCzF2IUnjWkdVWUpR4IMLa9pQjObTP/BqYhSeXV1jYV6+aLFVqmwW2
dP7eNw8w5EhlzycZa2svbFhjf9WPID23/8Jfx2Q72z/3Hp+4etvdxq31n912ZJcgdjyxloYeiTDw
bgVRHZHUKHVRW7ltwlAMEKzVzGcCJQIc//+BMBfT5nvbWoEJYsEBJ28P0vmMryklYc/Gybchighh
XFIKLM/wRTgws4LvuFJIy4iqSuRka3VYPRqkx/OrrYb7PSiZY2mjS6+2uQEXjtzeR3Xbu0zeeueA
JzIJkMrUSy3RfxMNqaCWepYmYVxmaCJ+xOReaZ2SKlTMyF//0BmGC9POp5549V2N0BOft8fS5R15
TL774/7c2dLX8idDXrsV5KJ3hOi3g602TpwbW7o7SgAMAW05WXgtkUvX8+graPg6FmIN40Kd/onA
O/MqlGKfdXAx9gSbTwW8949RY6/aelljbNM4UpHEpwBlbGptQQvzGU0+XO2aZv0QPiJiKYCsKjYr
VJA8lvpeEx9ZYbV2VK8AP/fPPxxSOwT4PG8rl1oq2FaeFZaDb90hjk1m6SZy/Kwank04R6ehosY+
XxmWIOP2O69EXOq15kEJU9goUgR3ZPH15jmP0xsYpSpExgLfL7ZgpA0Vv9Z6YY7gC1A8JnsohERf
vR5iljNLavyJgKcNZzWQftYfy+BDGw1NSOeaxxRtaAc6PcHkiqEn0xVgo7k7a0g3vdqnIKcBPHc2
DQ4O1icv3ltBpbTvdqTssbp9TqP/FF/kJiIySeFmLKICOE1pIbh9hqUmjlMo48QNg57vUfwTIXQz
M/91PtTrNxXZQ9j3BitMwOWN/r36FW7U08jPxgVJOsVdVFMOV8csNtoH6ztNqOf58lHwdnw8VFY0
GfDZ1HTsLFFrK9szhtrcepflgCsdGTD94YFiPUsSFV00pQDapIB2QOTrxZBv4nxRX/rp3usz9pSB
2o6nSEQYqqDFSupMs3y717546+WGoB+JdVv6U38dkgISfG6Yqjl5OEPamQvp3svRJpVGRMh0XEqh
BfAoJ+2NbFecljQgow6uINGBBGTArG0Dx04qWquSQXbrngosxcQgiyZMUJ/6m4HwhOyalO1/aDQU
IR5/Y2Z1hu1lLW38JwihhF5mYnGazW/RDZgdug4QmVQW32JaHL3Wqzz2E/PcdJ6XIos0KBsjxtpD
7VIquJL08YuMx3h6iJG3CoM/FsJ2S0+67FOr5cOn5N4VZ5YOe9YJs3tPtKQcdHvMj1QJHHTBg6vt
/ramlO8UKkHRLrwPUn5IfQXrk7D+zkRLUnwvIBsaS86MlOxlGxByyPixbeNeGQM3NVSG3icNTrWz
BmKHRF9rCpTj8LrcX6lPV6UfXp03brSHsqRUJ4aLI211fbgayrHfplF5Wvo19ANGMZvcmPMXr41d
hKWU8jxBMIx18xfBjfj854l/i4H8dhj+I1q/qJ6t+LAGPPBSoPJwKTGxGNNt+5VsffLHCrQGSsrY
egNaTRYKbsWLB7U7LjKAl3GXcDmYMWGTJyZ8yVF1XfeJcJgnkA3Lkhu7c2FnsegBgoaCMB6shUYX
hoK2vRPMihje1p4HiXRT5GypomX0ZB9uCcr59ShnxaUnHgNRV4p1OANo1Nl8IEqeCB6xTJRBxV8n
LOfDyDDP9wi+toXHfYx+D9NEFRsfiD40d+1l3NLMjpnNbb9i9RBWQkjxiTMeHcrHTiFrVsT1EuGW
s4caObRHYSdfgxa4NCgnFMUiQhWQxm2EHTXQ7m7czAH70dEnZ9DFZUESVxzTHjYUfIf1Jf8bkDZz
jJK2CRNAvRsueK61kbLVFDDJ92F8a1Eh9hzM81XTT6CCAM4I0pyRNWmAB94mfLWsT+FTNaay9w+k
ioKajG7nn0sZAOnDUhv38jigsGL0h/R3KeoHXHOkYFbA56jkuRmIqVvMprJd5qr+GvTfw30c7ReZ
HZntRu9/0uhCP+gLJYEulKaaD+QPyq1mO3n6y2HLQ1Psg6sIADyTBYKZIsiGb3ekvM1az1QdX15U
LiitchR4o8pykhniMMNPcINHhXPFMegE60+ZS5ZBLffTyPSe6zGum8KGdMPaAiXFOyGXGlL718TB
UaxNjynuyLxq+IvMDUt0c6jsP1AwZBvXCLWntEQfeRrMyhgD2dAI4gjxQ47MIOSxFNHuqTj4Vqbc
WbE/CGucDzmr1cUok3ZkPmloqXF8QqtG5qDBn/A+3DH6+QlPuSvuLKgyoEvDmNH6BnbKMbSXzoJz
p49pNxnYyzFkuRzgloiyh6BgiiHy/DTRqFcgq3mISBd/Yp+nb9wGjybnQJfdrNV7cxFYvzWabQMT
uzo4xmzrbYiiU3/Q7TXvieYRvfC0+7VKsxCstTTRkgKbfPwnrOow/knID6lCF+4NHfx/U+0FF4jM
Fhsq02soF/0eP63H4DKYUVc9Xy1lXr4F2gfMbVqa5WqX+4AoNmcciXXjZMnNiXPLzAimWyI831l0
1w+4DfKJ3lPAv9bcjl6Tg6NMLJpluwcb8s/rz8METy6VpkadfygQ1uNsEKIigheVBYo2tPg4oM+S
BjK5BkvePkXswgWqTLuKOh5VnGQ12fHhxjW3Dvhbls5L5omzbr7Aylx/o9uOc05F9Xr4pkDckJcf
JPXDm3E0LHyWXgq98PvluSZx35wt2sxaF6wQziLrGREVmaGgGqNJwUgD0yaz9/rez4148gKKHjZ5
z/dObiIq8doc8oIqzKyJQ+tLDpGPutftw14+2DmXO67TOCz0By+slusDHb+JkQOZd7tyhgg8e9yJ
FEFKGmCHv4K8hwE3NOlnt7k1IUgidAEyncI6jwJz3DXg+r7kEi+TskwNxSHxZbgdjqXENKEMVjUW
Uh7WBEM9hkbwGyNy7vcxcp0C/J2wvtVRSTzWZyQmiAU8okDU47hkXov/PdLVjyYNSHPf4xBX1OsG
jlJrG0Z3BoZPpkPNJ+hxUrJWv1DDzExXL+ugDzX+scOySs5PlPLKwodCR62fuHxWHstmT95lGDJ+
I+U8N+JCgUMhPQQqhvrXXERgk8gn4TNShgvhZednhV8XqSdBgWUSucD5wQjH/VfthXGvAT/PK0le
OqeoTli6DYMbLUwzTV6HoyzF8fMVfn6ve73cW3dID76jVMMRsN5uzrRSv1i1k9FPk8qVSVNzhnLm
5otX7hPyXR49rtFYg3AI9uS12UIqJPeLzSzNVDt1Xf9AEbu6tLgRSbog4l44d0XAlMylCmo+e08c
rVCsyhwdSe8CJrqRvqdrnJi7Ywnl8q6yUCs1GcIZnRifClisqGdK+1HN/Uh6r939M3YpQzrQ9sCs
KOUZhKaE5vusK5xWNUAcrjGsJ89Ik4qXxXiVuofOQSdWGt06Vv/aw7C6EWlHHUPmSx9UQAyPV+W1
1qwKwk26dt63WAe7pUisJmBvxxR17zF60qGG5LvU7cSxJbmQ4EAwfe8aTpGZTyqWq3ICjynHjWKX
JjnQ3yGOzovG3YruPnWagG32XvmDVdIZuWlmV66U/YGPqNP9ZRmjzdtfHRJ05BhAzldky8+EliV6
Z+ZU0Zvf5UBZYev/b6ykDixYjOjDapQO7QCYE5Nw71CnX5jCSkBC+GvAVgubEKSIOqx5YO6bBHJF
7MP7GtStm1/hAYRPR49Wm3oArrAdMqw/5X70u9Avf44hsfvYsj+JGFrfcTTo+dgKQo0FD4A3F0ae
7+LN9KlWQdCh3SPmuOjza/GM8HySYcA5LhR99wT/X/OYg1VgINXPwzygxIR4rUBr7MsxKCpJGwHD
CSEVfxvFPKEFmtHlcxw9ALhrGkvwXJo03noCjmR7JZ1/SbPXs1N2mVxc1o9zDo5GCFyq3BQ8be+9
fgRLWAfjVpOYEj5W7IUnKUgqfjbsN2XVcPGBeibwp2kZ9AqolAlq3pxfU1tixgCvYLwocc7pgdop
IztP4Gf4SYab3gWpZHJIRODU5vCYCDSNUvEj2jBvME6hAdmByueWMR9EgetuY+gMoaElsf0lQHZU
0qpOafJPuV1uUOB8Rtxq0TDlqce7H8zMrLOkC0nHvnk+j7h4D5SSL6cptWOt1FOceDUZ9VA2OzWO
Z/TAoKAl5udZtWMb11hw/3fGcvPD6NLblC/eLR/LUpVxzh4sYHCRcjd+kiOI/4shlCMgyqDmMtCq
JlpLdFRJ8vy9KBd/W3UiVWBWaQkcdm9k4hth1gFf6zz6Tly8KI2Jkr3BI6xdAsXu3SqDpybcbVMd
3plRIqSlh6r+T2EKnfIo28KIFzujue8ypv8Q9DStap0j4K5ICP+OYpQ9UELBr1nJk+HnFpviS4eH
LNz0kJl8vdVn40WsMPkOf+ry4yGHNjT3S+13MW6Q2/ppTcKU1yRfBiF/2E++bs6XpAFT/cTC4YCQ
Rt0wU85oBvOahaUXTODghKhvsAirJpHsa0OpuS5OGTYxhOTQF7+aNeU6BCdd/4+9Cqil7TU2HCig
x386a4/2gWbilotFWQLeqQekrkukUm3q0ehOgpVdSeTvpTFYw09g7dKT8GCp13DXV+I3jBiQ+DE5
b5QEKoxVtzNItXJlILALBO9/WqWUElltGQBLKInBjzN8wAJiAcRCJzR/HZGlPORYC3PDQPEctvIm
CS7FOp63zuPVzigHxFrPzrUAW/JQYPrTU8Acw1nYGZIO5juQX87bYBSGs221LyarbDm308Gc7EAR
8eUQf+rG+WTH+E6PxH2NKHynDG0QTAK9gJkmqCptQWy3drVYFuOdmOVocNpVbIBizXd04DWhm6jT
vhNabGl17LJFmoOGSEZsG9N54xffyHezx9X5EakBoS1/3OPbzhsMF874rSLY8a+OQwzcmashDbBw
Q2AjRSZVydwao3y46+MbFzpLbknail654lxQSITJro0q198URv6Layxl4AKfty1kBkBoEIgNvIyj
Ywrvn5N3peCL4phJbdFxPIaVuQq3EEdBApJT9xzWH5b62Ct7oVrNJKeKMD/ycpARYCEbw6xl11sq
KNOgzc/oBtuYB/UxIgAXVIg3PQaGVuECEzoDYgIFvmawtxiWjxMRAJj3kHdQVoC8pjLCnVPgUOUe
7cMlE/qPEYP90iPPJKVBU1C2COvB9BTQb5OIsuihK11wiwrQImN7ajiPu7eJauyBbQAB+uogy/7D
t7oRpbYAqSScHuoxPw29c8q8bxMFXUHKKxkcKclAgTB+hM9TV8KIZir+0pWhf5HBy6NS+QS0mvGt
uh4VUJxMdzMACVaJLWh2W9QhtmOlAMEKj8KbHyTig/L7dBRyHvUltjE5Qa3CtFXJVKksGjt1io/2
g5cLB6XXLj6iUfVXc4+GxEH/6idf3mKLGZv9lYtj9IEoZFgYJhaP39yxTnZbX8z5A/g14iCwnu3Y
3CYI8rtMRX6xOeeKR/vTUTYmpMYwTA5wf1cWlQ6WTCksQXr6Bt3YL6mX3t9zW2hXWmzHHyLs1CGH
XvGPs7HMMMsNCLBiCFL9sYk4UFa6EaqIyfqxv1uKdGUoavpDaysNLHy+WUBnXkgwRgU8u8+ZM2Qg
Uyg2CWmGyU/ksbe/h+XWwvqxgTIIpaEFBjhOaE+lXntwF4DRydZqa52uXEvICrH0AiD0+rTtCJM5
QMgR3l9ZFJHRloKPXevZZGPhT1K2Mpf2J5rc+TeGUbkh63yDROB20PBtQiDxEF8qyPnH/7G+WRdo
ICNSnsjZnMXquccD+cwzD0Nv7tDV7+3D28M/5Bmfc66daP0lEblxUuZsx6gk+TmcBUDH/p5Q5TCA
/6/XrIkZvlNSILKZu3d2RWayFxj5MoeycY4wrkZdMZvFL/bZInQaA5IsNCD3oRZrKV8vG36mvcMe
DF03anFO2EP8UMXZVCz3H3T0U8/qPDGOGP+vVbnJH/bMBgqgPl6aYla1CvaGhJjz9tf6jfC1VAg0
Bd+8RvrqKkcJ4QcJVF6mI2M6h+TKwGZ9C8UDc/DLw9GXGK/L7CbLv07rtUTw7QP7c5eUj76sNKTL
gdlOYVUp5+6M0ZCvwko8Qr0M6G9rZT51eGMmfo9VmGWEycMVnLIibXJmFO7DtQnrGoacJ3q8P79I
JPJIm2ecrb2D+Et20MM8J6cHEYjH8vk8kRR7u/WG5t+x3NeLt9qIo10Ey5Lq+US+kuQg2x6VTPJs
OOtEwaTsWjiG28/5Icg8HzcuCMvULYgUk64zsmsvqSRQtoul/hW34vjLzv5JdOfFiJ7JapH6BnUp
ct/8ueArCOTNkcQshK4QAAXrigi5hn9YWbXiH/9RIzH4zv8UedYxogWJBBhRGMjvY4RGVq9a4LcT
NuZ2uVdlzrb4h3PjOYyaBSEULQRQg4nBPcj+sBm0sIT42gZQiFPA2QIh4wbiaB++lqvo057/NokZ
nqlrXbTzuTyui7uWl9NZNT5mlhVKTsBAHcTlkK1kxIZHndKXrrXKHi4Rai/OQks9rKl+nUUn6Nfo
cN50j/ffrFvT0lImKTOGskxD0LCpRtKcfj1Dm4M6HizQZ+22yk5Nl4Xb3RVNv/gRor0ergZm9eD0
UnDopG7Qohb8EbGdEAE56/jJ1KYeTBmQJRGnD+ublPkdB7dhwGVDiNe4SgbHQAx+5N88ddqoRmIH
qSA22tnmK/PGnYJbbpD/DuTwNsA/4dq56U3NLEHXPuB1WSuGfUOMO4nBtIhbQjn3Tss87fuRG1NY
B90nM8iK4XkU5s28AV0HD3B48vpp+/lmVFkByZ7PuFP+eB+d3loXaAwVh74aAzl4ZlYLnQbDcjNk
6Uw8R2eCEOZTG6AB5nh2WQGDEgUsRFNfel43lgE7Uigfw/nW9tR3uU2GuVdxjdnzwLVi7q+M77iJ
QznMiuIivZi/0w9RHYos7F/+s3dv0uW+CKFcRiNNR06Wysc54NjvbH7M0pEutr5scxv4Fl7Tl4T8
gs/B6yNJDcII/eLt2mzU9l6z1gBCYp1yF8DlXU0jj1EW44CziPbblSWdNOGCHJ3fyS9gkK6VZH/G
UfN1CDAuzIuc4Za2hJ+olbGW0NtsLVQId+GyLwg2yVQn+tMgSrk4kkVjEBoEyDajWjhqQZW63Kch
YwX19dpdktQheJD56ZwtwvfpKmvlCsVT70PI9p0Unx3oK+DUJHC6GhTjvIkozrxSv7ujkFGITLvx
YTAsd/d2Qh3l/RyryNu5yREXLgXuyh2X0j4Bst9ximMgapgVJgezf2MNz368hzh+ajsV9oRVv4Wn
oaop8f1WuovgP55DhlxsPmpMeG7dEW6PIB9e2KauMUq+C2iqd3NGURAyITfMI5cm1LCBcEgI23ul
cxaL2AXGkMPECK4DllYDj3qWE9JfH+MEHL2PGdMaiqMyZhnEq9AkRKGfaAMzXRGBPi1ZZzci22nU
4gH1MuVl6pwFNSCUs1MuR6Yh1humEsAm8UhfBNIqct7X0/LIbA2juJAq/ZgYAxND9z5R48c+cx1G
qNAug5q/tY6r2uniTGrfmFmcBAnISfTrKWZzLfkOqTmaVGZdqqPwaS5hfCFcun5ozndhDAwjqorY
y3pj5cyDFFcxxCNn2uBirMvjaM6jdv6XFrdINOQ9BFocD+NJrfipjL+3Or24R9ydSl0pZ1gvP7Dc
FtcC8h/3zFiKvmZBIEdHtLwBgV0mml0OUmreLquVa3NuDs65DPmp1FaSLs//LsDLMBxZvdzlSR3u
LxAPNQhEGndx5YHMFr90DbIIN2MumWTI3RUb6agRE1MfwTILKJL1xJqM/7WkB1aVfejU2LvDgIha
IaZIXA0mUeeZQQTDrtT9MB6Ljtf6JbqTzRPreQ/fUB9VM3+llx0NHiiJz69gY10F9kKTSgmPmYED
ZONTELqzkUQATdf7ue7ACBe9dryVpS+GBW2RQbBxYilkzeH29udjPabhCGPjUf0DfEwDG6jL4N+3
Jks0M1WNZYJP9whdUhjlzEf3RmHD+Im3bUe2Jq7wrrLPPN3pHbXXifPlap+T8ju9kH8YKjTx/Z7W
34mudL7pbp/XBoKl6bWkyKD/Ql8lUHYskoYsIDvxRhWH/CRocevyqti4tRMz3mwa+gx54mdJAUFU
JLI7IlNBLvMPy2BbvTu+gi8/D8xrMCPSHEWQiK7ezu60zjUkGp92WifnrMbr+ZOHbVMe/hkSygGb
am7RIM2bENCiG0a432WG4H95D/Xw1HCT3mwM4Y/yTzrfEEfxgquex9BPfhZ7rY4+jBidOvB2nXaO
kbU7YyGrr6Q1SEg94Nkn/OKLNkLA4pd5FDRejOHHwKv1ND6q4kEb+yVW74rkL9+fnC6nDZDcvCKP
r6ftpI+9A0UEwy0z4xSTxSfUEqt0427vR7q0T9oCDCKnKlwF1KlwqjIpgBV53Qc3KI+tyKo9m20Z
oNeuJ2ILdNhYQWwJEv2Pe1DU2sKkXzxyokdIqZS7roTomHbFOjHhthPc28xaheQyyC7nUa0eAfqX
LdVzZGspXoC2+gdqnb73gEcr4z02+BCyhUgNk632Afmb+sY3Ey/1fUl8s3w+hF4+ykRtlBf+exwV
oKqTp54uM9hVkQvs+EsDW0/GGKxSMCktktL7A7tqwuwDV2VrOQkQlAtJlP0uN4nSY1J1iX/PpfBk
UNDTdJerFnvZKPFtyv7RtUpHfMGAIgKfYIYKziAS/bmbvkekqQ0zjT4IhmchND5jzw2iStKs44TG
g9dirwSATxC/gythjKVmVOhsFt0u2oOCjv/gHhYQuDwztFJHwtVnnWkEgZWz0uu6KiCIyC6Q9qvf
nyh0UImtkMFqe4C9BI5lY3/Hsel7SuvH33qxJWhFDPHQ1maXiYDbE+6FSUVS309qCDBXup1BbILf
vyNzC1GyfzdMuMcNRKstNNztf+V1O40PZLqVz0gyPlXK9kvs6RcjLh1yRWhsKhSyvi7GHym09Cix
s/8fshE81jxVTW7/Xj9ngLMJXczOErXD8N4kGhf88NymLhzcZ0MB8XLz42hRHMPnGzynr3nvaWaS
pBxkjTAnI2HcbRl/MmHHAlJlSCQ744KGyCXVaxbEfbq1yntRw7wtWUgFgdhI2LG+9/wJzI+YEDD/
QC+uydvanaYNbCA8JTe7nlnHPfAW4Oc5qw4n+LXxR6NdAKqi9GKK+3m0ejgcwdzr7/lAWWEx59r+
vv0Xo3rE/bmN2gkoH8gsvmd5kjsjxmK0rkORunwUwWItiWEJ0SGvoMEl0WxzTZOQHFYbnI98tb9w
0HXc+jKzLGsnXbL8WffCzwL/JMG5OfNJs7FoR/CS5xk/uyJ4mNy4PkVmsgER3XGzcJiXieQLpNBs
HtR+Dv17tEjenNJ2wEvWj4eifUpYBhmApWNfJFJGOQTPFKbe5/4+xTJre6Y5sbbdRDhVPo4hJnbL
wZcBeJMwhZoVZx3Q3aOF3Wj9Hm/HOaN7vMFLd8jeAom8aZjV20O6TOzfmJyv7NLS2lgza+nd97SZ
kCRRo+fsTAlJ5/D91cRRb/nj9CJCTAubriSVRUkdyob3kRXLP1sBvk89jlm+yLPLMFAc2NwU9New
gR83Kgih4UZziubWrHG/XZ+KTdgHqJOyD1RXHvFTb8V6zG+kvVWy+cN5WMRXPEBCgEdg7MixOCN/
XgN9rXkT77jWghOX3/yfzy3mLn5UQ/8aeh7fC31DHbXdjYl8R0Jt6P3jtIfdlqFrQwh5WfrBUjMB
ssla04y7q/W1Pot7Q1Wy32qp3nroao/2SUogxxoCZQseMwNbZKYxrpsWxzIjPp12swBQPXzIV1yz
KsAypEQ8TQMDHaSj8Oro0Y1YCrIbL/5iWjcubFe/cx6r1y8cqa5ZfZJYwkZkBSZAT/gUdLY9Qwft
aI+JdrSKQdRS2DbeKnZVXiYQxKwz8u4NNyZzlBq+6HEgDC/VVUMoaUkUkx7Y7KKzz5bxxfnbM7A0
LaWTvUGYoqJj/Py60PYEJhSm2aTAf2t+Jgl5GysQT/bG3A1cLJISNFL58n3NWtQEqJj5mJpryuZz
EcqqOl7kfnOJXdX+/go82U4VfqFjfVFPCw8S23mbIjwk0Xnoj+Rgr7I+E+vSo5Co1trX93lOa6au
oy8GCWKxyRP2u3z1254MYXoGrXoLIUgHqkZwJXNyltzLpUXkkYjvOfNnDLeayrriAsg+/Vcm9sdy
44WNnpXd4AwLtmQMWbLHv84wQNCReZfQ5mN40y5LJJ2pUuVPBl7u1QVmj0PCsgEcWpfAp76rrbE3
KuOlWRl1t7+8SBcqFEn3EMTLfaiZnmawZ4f0voM1OKM93NAp0S2J1K5H4uztpIY17aKqmicDsUXH
G58IBj8qZwXQ+KLQzQEKUqouZmLw8PncLl/PmIjgbnflB9H8i9lRKPm0bNbyg1YiLtutJmyAM+tc
l5X2bxiXSlFu7f+s83ewCejrTgxlGAk6Il7cSK5E3xITPWfRb+1eHChTGOHF977QI3cyZXUe0ysh
nlVHxJtY82RX5BOXM+x5AYDlx0sXD8Au9DMDoOqqkNeKP+D7A23D4my6O1J9nNA7pHK9YQszPVk1
+2YlzLifC3Mp4Q5OGOXRRPDK9Oulk4yivHjgNN1gYqG0sM2Bo++45aw66l+5QHyuVTmyGWPNtZIW
4YxrSLAUelcOElzfDm78ny+B5RglNXH0CSjqqAGIAqv6PbC+lfDBWtdi/1HtZ7qts1jmwjkNmzmK
EeSX3tydLXLxWRnJD+1wazAXj4XEqssWyOh2WsyIW+Fp2FepJ1TFOY4SJ7ntnGXCmhh6laFeeO6I
nG9hWu67LYo2WtS6nCESszw2m9v02EDtmuNEdHpN7YCoTAE8mcSebYPac5fiOi7FZ61fH9TqjNeB
liZTchAZnbWf9h3VPUNbsutt9lqxILgp3t8eiO5MEMFQLs5sPatkOxa3zZ1H/+CReVuOZkt3yBBi
62b0SKuqwkEORFDebNQQ9C9eZN7vp3WNIDEELGTrtaK+8HcNGi75Fq0t6f0CXkMAioCJUeeiHq+2
hCunWwzTKlRIDIWj3K3htXf3odgdAkSgKQ8jiYj0z/MZ/m/0EDj+cphXiWRXGCN+YwZ8BM/3LT9O
iJ4gk/lAej9JWWxKz8oItI3u/JcHOE/GH0LFx7f38tI/fBFLvJhqSa1B9G0QzgvCoWIjaNcXrSaG
rADmU/POU9GpnmoPF5ghdH0qG/sFASE2X7FLdXmpOTegv4Fu+LjoBX9vsok0WNGvAdTLnKYZQFp5
eZ/+Cf+igEMq/KGPsitQP0UhmC8VE8Cyg1BBMXJFUWLPUW4i7HJmsKdeT9uTOpNXrZfGJ7sU8KSe
neTiAZBrDsSaa/iBkx9YL8cE4FCguZKS/MolKeZ70i+a/G6xtlcdi08RNe7AKiAr36FnhYsQ7KQ3
pd4DVdBS1/kV+Q3n1FCBGSDwGyp3KGiaYuyCUbqFX1ebRNWKiE2fzrQ4pRdrf6OFgwcoXRtk/Th7
QqDFNKn88dTaGvRLyoTKX0Lv/I8yrsWqn4DHRX7Lxba0IoqXpJojgist0re2djUfYPUtXWTfbdUv
UUHC1Ux9FOrSKluHcQM3HYhq1tibgTCvrUPWrxbrOBYmTggi9vTXqUUJ6qWF/AApcAQh/EkC2okc
YFDzDtZ2sOoRPA/8kolaAz9XgUeme5FreEUWyGJs8GuzMqtJ5zY1ohZeJHUXhGPYttuVe5GG3SeT
7n/GqztS5mF1U7RHbbSdf17WbHU3TYsjyOVBCFpEp65inaeIjetOvTUZLFW2U+ksz47y/XvoGS5+
+LnCPFLSpWjLvywXmfOBMwFx58f1ShKskqMcAdy0B2AzKtxtkJISK+2qQcFMJ36l6Zd9bVLMhDlY
UMV2r2Ho4VR4Vx2eIOOQZC7Rc0gtolLj5MDaBTDBhoBhuVFPxgK/qfbdnsY+pTQry0kHt6cYx0zm
wk2w6JxeCtKEGBXNT8KAc2YHKes9mY6YPnm2IhLjZ3FDRjtSNNg2yjXr3qwGD+ceKmT/yEmfMImN
s20DNlrxH2YrcsJ3zNcIXwsCuYjkNa9IUOMY2e1w8mU3Kear7kXDBwBfxqBDNYQCC+MSW2dBcq36
SqMHizVbqXZvNABRjjMMp5u2CgdqNcAGYreAtxdOsHR41HuKeSostUVnWuX/bjp2AdpJjNB9GyeY
JPi3gEIB+MWS1K6Cl9lH1nQisSbWdIQMVYkx8i4U9KxFsN084xH64iKYPXZal+UgBmNNvNpfQbgf
23lGTkCumlB8Jos/5eQKBzNHZZ+zpDvFUDG27DB19hLQ5C6Prue9Jw2oeOO/tDt86hrjio9JIfQo
Nv5YNCeSCdTT1fOFqFmVShTFGIDJN72MXO6znnuWbSOfEe3phiuIDz88eRTXqgkOXl3wBIJjRwWM
4kJYXrv2bdMJi0OIX677TVFWOID18cC4HeiCkrFl8QdODBnT3oID75Qvl5IZwPTsp4T9fTyXfTqm
NPI/30Pc4xXo9n2a1SbEb5jwpT5ALA9jlPL8POQ17vSYCBvryQtBk8lYWqgY6JiIE2JwRP/D8SLv
R6rQYR/sILCrFiHYFYORDiAC7dghCLpwNlvwPAhG7/8ws34NaRKZ76CMpEh52+ovMONYKf2yaJaG
OvivmQeohZnoFO+JYVA0q6bKoZcxn5p6sAAlwswwgsOF1TH7vShhn1jmVk3xdx5VT9j3jhCWOxm8
Ec9i0zvFxy03B0967GeLz4YWMf/QVyq25X7FY4aiOahlY9tgdQwJK/2rfb9PZ1yBYqw6CTdDddCQ
AhtGpw6sqU6j5txSutD9N4wjOGVwnaoa4pb+XGf+RC4re7W3l2hu3vshMJnfP+F82kmVvh+uMElk
18P7dnmR6dS4gV/wB7apvwI3JUv+nqz06Va2iSqmY7veDW/mCSccBswvbBgx+dDQWPU0NVN5MZtM
HZ/mTNRgLW9LeAIVTGfhjvE/THIUGLRGR52s/6XlBh4AhpV3noW1VmGBO/Y/8ngHvDD+dT0rgTXT
vjXwcb+ZJjm8BV47TciKnvcU4kq6kZSVwx/QywlG0mAoYHGPJtkcnDDCSFc/5Wgz4lGaJg7eBeNE
85SN6j8ViwYiWXdph71d0Hd2tdluQbsndVgiqWIYMTbsZyFpGlR4sV770yxOXWmwK9E6dvZo+mDg
FhEi4PJqoNd9RqqECLu510oddlMBtYgB2HD0idl6FH3YDHEy2pQIHS8Z+Lmli2cEIXqF35oSuVFZ
/ujWg7yJGq99GptNHB8kFUNTP5Fy3YKJ4IVwZ4kr9zqOtDQAj1uL3I/nSTTZUsoqT1jh8fSLYxkb
vBl7G7CJaVYLtqJtLRqQkIolvRjm0AZ+CM1yS4Z0uDPlYcHWDt6HLR0eAwHjao/EmqKLp01o44t9
QKzLEnmLQFB7aO/cV7YftWn1HOZvG1keXWY2B3lycOLodKpeooTWXqnnzkZUngzuM00qc4g2TUxx
+SJ6+9rRT+w2/7aggRUzehfo4UH/P2b+tm8y5R4+AXHiOrYp6fgtjpNCNPyMjIo3PzjWYD2QYHtH
oqX7bep6e4Eky0Ldo7TX/eouI0ildaXHt9AxBjJDSJeiXQmXtFfPXfLbr+r+3tO/dXLmoNJWB7o7
4xo68ehS4zi3aG6VuV2gwHnTpCyv+0JprmKVctlyfSXmwSW6+jV2jxFXHr04efEjlqG9yvtDuwBn
LXLhmrcuSFOiA8U2XNtyGANK7BK7BqapTHy5OO300rcnlX7Trg75AyFPCG3YECLwaZ/OaqUjW8I0
6Amx7EMdi83CfmvJG97s7K2zZUwCOYwM+janBN4LNsbRoRcqtUgxEWEgqNsFyvXYesAODFhdsWyR
8791rmpMFj0CvaqvkdQ8ONmA4jD5i08Y/G6nUmwhRb4RaAduwV79NbQ25Vqe28d5/ZMr5SlK2no0
gbCRVVLx4PgHZ0RzgBqt5NM0/9aISIcXJ/EvxGuTZygCiIz0dv6mXL+rVf9YL2Sd8Rw7QOMPm80r
XOyGGH6fAUOQ15GyGcEIq6LgCCTILaiLUaEsZFu0JUi9Fg8wltG1V8u00jG3x5rsL0eNhbPMdBSu
QnCgOUD32LU3VY1+lwvx+/E4AFsjMVmZtX3cGO5SxsvU54eImRCa6AfdmaR0j7bO5zo0hJXckkOk
PNRcVdPW97KTiISWe/zS2Sbs9GkdXoFanE/yOnXJXfuEsj57eBd1fMx+qJYzGflRjdM5xL6ZnEsJ
AFnM5FrmOE5njLK4LNFZqDkIaqFMJ6f8FJbGVPTtvsURJwezMLC6yksg0y2e7DoPUYSmNrhrn2e3
C+dcXmf96A9Y2T515r2HWuLRy2S6rdYLKqp7tepUxa1p4lOsvcsZRaY+PRvhY1nvyAJdrTVuUz7f
uObMZZPqNHo/+VdC1HeWlPHan8WXq+q0BwitMfO6fIEBFZBHbclGFlER2A5gg8sx0p7Gjb8fabPS
XPSGROe4EGEwpg1/zNeHpU19FRJ2hZNa8ARofXaKD93UCJ7AztZKeQjChhSG+NGDRCViI/phegWw
mEYRzhF9R1e2Fgfh9TZOQjVl5iiFER6C0dNSv+8iEx3U7xe+ErpW25lfCgDneg4ngs3VOPgr/Slc
iPQ+C1jq/EGVBK4n2NwhAGxaCpxGdCsblVpQD0tyqgTG6mG46Zt53WaU4LabE/oUwvI9VISM7XkA
F0idIOl3g4jd8C7001YrdcWKh7W4lUANSLO8CnIMICmI1JdjlzLVa3oVPMQOic0BOge24IVOuUZw
Q2mtKjSYClh/BlCO37MYq/6i6mhXnBsB496JoS3iu2Sdh6ArOZ73h846nTmNM2pkMZt1W1sjpVrK
XIs9VAEwYTtDNHy5fbQilZwo7PBIR0+viS4pln4MrwfUocN6cpQkXvYXyOK0hdb/brDT/1gfwYYE
km7+akvQxEV8MleYAXU+pu/ENfYIZ/ePAgkUNKhVYGW8emHDDEf5dtwR8z7Rq5DluYfyHJ2xiPOY
LlomxCyh48eme8iBR4hU6BJsJtLduE1oWznMNQSolV5WsHrsBmKJM/97kOKeC9bAnlzldzYdkT3n
MJQ9ozwGLuo/8wQhBsQW6XAJ381dWugwlCl5ifVQLrspOdckESd+57YLbM3AIHXt1LWv67NwtYIu
o+fBLFh8xjpG+n27mfYGnUJu2Mnli0+8pzeuosJq9/3g7HE1aHBVVG6NhqAonf7ednZUUAscWqOu
KNoC0qPWSvyqY2iSxUqaxc0uxDH25iLHdE3LkQXBd08u5boaHiEjzRYI7oXYWftj9KHwkK1F+vBv
55CfRZpt9Nl0r4GlsbO6WCrC7xbfdTh0vXfM6UQxPGPXhGa7UxV6RfBVdiznrAAV0X9braAMIlAi
kTY+iLn4MvvZCTHZeI48bZZ4ooO/0KMjLXsZ/zjubDs6h21FuxP7uXlZ5juJAyTnBMqKrQvo4vtI
FLJd21PJddu/Jupg94qwOThCWlrz14PZSqDD/phogJ/P3qR3uALW5CpenqmiDHWO7us6wAvIRvBq
SYLvm0QwaQAKY8iie4llWpTLb9/BuloaEjBQlF3z+icGoETvFvjoii7nJoxakmsgoBQIf+FK9GDQ
LHls6AIB4xwUWipMe7/C1R7HBJaZjE+3EtpVVOFcGQxKAJc6cGTWvZdQq5cxHwWm6ON3W4pM9tmh
oVm/GcWnmXwSFaidTaj5EnqWOXIzraiLxi2L2OCxtZWheFbNOKLvoTEsNLPXWwz67NhSXwIMaYvy
APGMIhJq9dqMoc5w3AvyDQGqvplKNz4x+qH0cJQvNShcLO5mnCEzl6XD7fOXsjmEIkiCb/GtEJBq
k6MCw2ipchP0yLVY8hE+CF6UiUljXJyJBRCmsK+KNNNSmv0YPwJ/li/hYXPfKwph3aME1K72pG4F
GyRuQY68J1SZ2XVV18Yxaij2G5c0TQ1MaBlGM6u/qKL9twC4C25LrCKnj5wN2g4EjE2v/iTCuv8/
VH2exA6RLVxqzBbbSCwPVvasEXVmXI2YHdgQPwkSbKwfcYCslqqNmUVDWhCYkmV6ruqZCVDPfuDF
azTAzKNzRafAHOqUvI+Iw0cnUv9Aqog1OgOg5Sqhq8L5r83iDqGkU3+u137LsiAEUyDs1ymBdVy+
OAuNZpagk+rtSGiMfNBK1+7exNMWu76u5x+W8rGkIBDUg8U1Y5MxVZtb1CyUPeMSUt4Es4DarVWC
uo5jsoTznx+j4RoWKvRZ4T8y60O9rAWxFnqUQr/JjC/jormTlYhCyIXQgfQkGwl1/+x6u92I3qqf
1Ob4rhkx4ex6orn34UJLzp18lUdfxRfaNuts5L4MVBom62aWB8czrzMF6+4pPgWX9DUvaLkVCPO3
1Dz8nzkHO4Mjr0lgiLkvnaXQybflRkz1yi/0RJKu46qN6eHfjDXho9U2yMvsSojTbm13rM+iU/3t
80iZ1P+IOKPE69Rj1UpoTMqNa0uDuZlL6ewHn0vv2DEJ7WiOxLF3woDvWhi9CZci0KW6PhAD56Ss
CNTr5UuHDMlglmsG7bLfXr0txHHdZ10nV8wnZQYaeV+VR6p60siJ4hSCHzVoAjvF2Dhy+BqGa/Uc
PZakFYLsgWgX9xXKs7LxPfhTuVlYleMp5pGiJ6r2cYtXR0oZscDZkkJLcdG4O/VMM3nfnSn1F90q
iEVwCIeDj+9pWW1k9IEiAD63b1pjgNwi3v/cwSpj9L4erx55dl5Rm/W58TIyc9OMvs9YI5B+ew25
zq0Z221HgR9aj32yyFdbh+QbAnuyJKIZBsB3Y7jg/ZcjEsI7PljJBMthO6ICa9lKOdCpeoMaLO9P
0YRMsmP94pkiv98jaBsCZ8ULpmoOsbCfzeWrNJlIrW9LNatyBGPsz8NGuEgXzkAMbeAEnH6gLrUE
ATybbbMLT/aO0ZPlWajS95ZOaqx0sb92NnwY/exbFzNCVcRfECCRt1QFCBsxIvb0b6H8M7PCn33s
2fNDEFuk5j3faLU2ANAhsyUASOj2hFQmG7MUdb/hyldN5Ju6an8yVzhwDYWPv+Me+9+6vMwYmaPL
/gvZgk/Iffh7hSEbvHhZuJ7Fs4UeLoTn+tX6CFEZ8OiVT05sxnFGNh31/ccTVVvQRKVQl9znZSh9
hiOIKurYKXDgaLUgJLKcmN3NQ0zvbjLu33p1H1nRTAhPRaz9bhsmvbeUau5Qx3c7xLE+XTr33hek
iwwVyQpxP+Nq6E0Nrhtku4E6Ws0jL+Im7DFaUspzvQAf3FGiML5YFX2kNq8dADb+ev+iLiLVHgTp
g/Tu6O/XobTrgs4apZb7tnBNREGzkM70+SCBTfttq4I6VIjwIG06OeO7FJmnparkzzNxzsoCIpGZ
2y6Bc0A2Zio584QJjkpJXVPYAKY9fKR9tMedXMUEaKuoR4IMnDSJ3VfUtdD1oedsihE4W81gdH8I
HE9VYzVFF1jhWeGeOd5RJHIo4B4TZ6CgS+DdkeqEOag+vFDRAKFbU66Kz0+YhCbty/w364JCH2P3
+1+uJghhC1VmEwycEm6M1QzOihApJjB5J+AtzcSMW9TqotyDs18wP0J6PLPwlCETmyVQ5t6oufdS
SOM17PuxX+a6kEIYDRGhclkc49ljwVVMVwiaAnFKJXaqpwNdR/W8DchAk1h6dobe3Ni6nKHGicKN
t+gA/4p9vFd3ChbZ50dwiQOVMn6zPwktGp1ilp2tIsgzuNlYBQWxy7JamyGJe3KPtFBgdL/X9Ws3
HePRYZJQR3Ja4n08vkWtV5jpXoCsJ7ENp2RCUPhjFqTF3gUUw8PTuB3e3Hx6q0hxC5801orir5jh
ks8inBzQ22YRAYpoWbRurIYjHsWqH41Hq1t9ipOptBIDM3Yw8KYUXf2O/M7p6oroU0Bn6xSX9hSf
lNZMKrBthcXkJuoLRA1qtqFcuwp3LvuT4gk9j0gRLMsKO32o+ipfG8JLGl9IA/6YN3hr8m87AiQW
xrKvOkYBa5oD48wdcyN2tIoQs8HdQRUvuDKSO2Dt1NM0hvIO7UOTmVVCsnJcRqPFkyQdHrkM2mql
QMFr+7nMOpPpVuBmyJWXN6xP9kSCw82msHHr+dsgBLYdQVf32Uh/cYBeTp1EMMzm4Z+7AOQ2WzVW
cajJks/7SFQfKoKUzqgVDlUbCgqNW5wUIyST3cMPCfGYlshSFJmKihxAs50LQr3vrWluCM7a80q6
9iSnY99arZPkZ4LNllAyZ+IwmN1AxldwI3T/OBZFTnYd5L2zB0zsUDOvIflffylHeDfjIHfiil1w
Kc/A5mxIBNXNDa4ATg2wdx2/FFsXjrPZlM9ggr0XfUUWjEEle7xg1NoGjusCqocxnj3P+IE1wZHH
f0fQqaQkmu5gDgbupANHHzmFbgCUTODB7c2E4VI5eh7RIapXUUQToVAIUMJoKeepyPyRGKMV0TzV
YYUKXXA/UStcidgoXOvvaC5QROQlMwYlr47XmAFzTUgsPWcL5AWPyJlbt9ThCeV2ScPFVCgJ3h8y
feJChq+2zgIPZb2LejGOwI8ChUgG1ssfbpO95FIZbSDLR97a1KsdskX0qu03i+OMQp9zJOyVcnaT
CfDp3i8l5nLnlgJUP6O1GFJca1wUFSTIAxMvWgB9Z1v5KxWZDDa3U6UEhsrE+mNaoAyo7pTtXGdb
3sic7gtBl4991n6fh1JeHigpsONBupzgIIMcl7dUaRR2BpqE/vS6TtQe6w5jYiC5/wPL22GNYeFU
QIFp5FUv7eyIuTKQmO1T4z0J8wvWlhixsTW/yJG8CuUJB297WEPemx3ogLWlnxk3d2NM2LtkhKB6
ZMQcPZqm4UsgznM53tRr1iosIL2CKJyPICrK8gpQJXcEk+esb0mGcstYp5oWJP+o3Ypg1SD0Rq4c
dY4OEb222vmOo5gHhBd1g8cojyZ3fXSQ0RXq3p+dso5PSWTUBlz1rEERobpM+O5XM7fMpxIi1Yu9
NJ30EBthWkT4knPUiDPRKk2oZOE0uShC3gHxyzDhs2W/AIW5N5AZihBoS+ywfGcbPWKdRwAxGWeX
DOR8sICg3MVUryu9OR1ndvJz7ElEFtedliVae9uh6G9OmH8UszoGO0QZxHKPkW8AgtwQroppknxv
DRCDyGhQ1ZrXYPclxZedNTuuKTMg3+kchACSynTMUhpL4hIhnA3doSGIolwT7XFFAspbsbesh1hc
3UcUl+Lo1FfQanhgC3uI3EgeGHT+jo8yofO7HTjcCsFObxSTdHHe/V2Xtqc9dW5g2dlPMV8l1kkP
R2bjEtbMHNoxlHfWRjG2gGOfZG49aW7HhOGyK9u0PSi803NHT0ZhbJvrIGR6Ntm44cJJKpO1UiIA
TfhZtln2GgOLzShQk2zCiv4wkjhUH9R6G0qRUYMoTZbx1O267Dba75nT6O6KGJ3sFyQdnCTtPr7J
1oCfYt4+nhOw4oUtPB2eEo9JkfmPfNDGy/HJpqx/h0UZCKQnB0ARcofmCuORjW15HJpcSpDjAyQ2
9CZVMGAHlDbW6eJ3Wd9rBrNZUcX4UqfzrlKZW6fuEDFtVP3PaJ3hbK6EHuooJoU4YAgYIspE+QO/
oOQQG/1Tn+TJ144Zd5ZwzJxwyE0lcClbJLA+jW4lWgkUxLM7vjofNr7PsJJxLdgWBFX8ZmNJ+UZ0
ZLWEoNozjeFtYtUSXDhOBKkPfaiWMcC2fc2TmHVaYNiVmM7rf9J+Kq5xspe4KHyXeYmgWa/SOD03
8oHCknWcK0wm7d4uz4WMT7FS7DoTjcUmGKLLqKBR7eHaxAPLPYCeNeyfvpaBCr/46a3MvO1AsTB8
v1TP/HPTE7535d05IukGVYiqnumYxW+c0+Zf0aNcMSEP48XRODK1ER9UO73whue+84sFb/Wj1DQb
JaGMf7myNLMd3WQpgPjveGm4CKzG9vGiR0nRyXw+tKSXXu9O6j9RGX7nxaPS3fiNC3l0cLS32p3j
efyZs2iU0GsV9q3SesUNcZaaE9rHxTewSF3/7gDnH31xKtWZg5aKgkhRohPVTQrwjPW3iOFm1y/O
iclMAN9br/IulNH4x2dDT5/MwdAsFisfybhISKAnUTwExkuNCd7S8yX03mNxuVrKahtgw1ts4g74
7VR1tVVf2O2mbmdc0SDQoNKkDXGUxL2ykx03EMygSXmyxRo0oVo7PnL5/pMMc3+zFNHDDmR9pOlD
ibgt+1HwrW9EIStqzVAs4JqEOqnhM1qPbEBRnSdAqMFrOmHNSk0VqS/BcFQpzvww74JlUDBrRbz+
7hkAKWuqNJCbfw3Fbf73mjHWsr0DDIC21ZR/Bxx8yS/SDcGdhdSd/UtSelLbqXdO91poHYd8kRPj
fPBJMdivkXskHyIfmlFx2upCu40ImVS0BTT7OJkukQdDybGW5qUDpSVGiHaomSr9OYxc2yAN34gw
K6t5a6uKFPDW69yiRYk253AfafWD4oXkfrRA9uFArneGisfeIWXhqIT3kGbQzKbirsrM8KAYYUD0
pDV6BpL2vN6amsYAKY8Jnqo+7RhDfrx/3OiB9V4QiwJVvZr9ZmbTevRpqZj3KZ076wbp/3nlP2A3
cAleZK8uILazU8MHUCOTXU6N2aDKvwGUpOw/JGnMc6QshEU9Z8csPJj/KNLbbXUJ13ycMiaUapim
lbo0+eMONOPmtNFrFaepyZ7QFZkNq2t5tgugN/BsCXIybfeWC6S6V9SlPYL6P2MosX0r/6BwytV8
xLxs11nOd3/VqC0OF61gROPaqP2CuVH+BrGJ7ynLaQKWMQhl5ydGJEblJzupuP7L77Tv85A7vz+J
f5HT6VWLtLeIVBOByfYxCx40qfv1nQVNIpDWYkZGZmWms4KYt2WV3Kn7TgyxZR28vsIUMIg5F6yV
H3dJilEmZDDn3hA0K6er45P+pWGRuTEpA19f+tqdfv37Gt6fZgH23tFacxtnj4GqafKhdgCDxXBZ
G0jFZcDSiQKr7mHwiye1TbyOQHx8MzZ3I4J1vUhv9bVzHAKEMFwema8VjFahJMFnpMYV/eA7tuZg
HGuPH+5Pg270sZIOPs2t9AyKfbrJHXpBZ2xe9rat1i94p+opMK25YGP5W9mXWkRTI5T9GHVO2mvf
PcijlEha06IO9zTMeyq7VAXrvvcJGb42ZzQkKdu1WwbiRDBQUoEuFGiUy7diOTRFGiIZE9huKXjQ
HuUL6J/MvTHldTFklV9Q+B527LpNpKeWK2qrj9nUV43isjcA8jq2JiqCwXwqhNVaSTJs013Phif6
CtmJzckHlomENYmdf/Y33YGdL36YXZ7xHEuWzhsB5vy9UBwwwp/lfBzTDtn8pNiHCam3aPzBgMKB
H0U/1RU1feNrG7ON0vZymE++LllgILhAC0FO/aw5WsNM7+iochMsC+l4yobcCL2k+6FMh+xw/BGn
E8ERpU4QLm19yhun/pzewlNU8DAkwV3+DmxCWCWRe2x2GW5nNQCMZbm4Ou5mQFAH6ARepLROC9dJ
/SRrDTPawLxMSdjogT1c+Bu4aG08hQeDmkw6G0//Iki8r0CVGYIKIaIIvZ82Q6dmMxcyWmBR/kC0
xf27oNlxO58+yh+iioG49o4FjEwZqc/5aER1ZjwDI8Fh1V81FvfMjl3Vze2qQuFpe9jlQ8Oq7P9g
hDWOWHbodJhwluIaE3ng43EhzsSnTth2ZwX0t9P8T5D6zM0n5A93WEsCrLfVlkd7bpinqYi5wsEO
ehWEwGMnWKeCmByUPkiCmNkIU4wAlD/TVjXp8+zosfhaXSd04cVs9PlT8gyjWU9Is2PfTtlTEs+C
lDkEh47UkcuIYvgG8ErJKMEY5bML1Mg/mzx/OV+MfS75UEFznwhB6/Bd0TkTwcE1U25emCmm+N3n
xQt5/vnR/znH17ZNsbmzfoYnrapNBkvkASIVzU2F0KyZKy/BvU54XHwwOgS0KzVMMPwMUbllSbAF
1KDdmYN+C7+ScyI+VvByJK6W1vazeVETUoppW3U5vJ78fd8GB1E/BWcxaOYKdsB0u38LU0YIUrXO
lV6RfL8Q48lz3cuBB3pfKuZ/JqsmS50VqHtC25u58h2Vaf5VAfgg1f2997MtDDdkZfbk7a2n7J6g
ktlZIxdqR1iieVxjhkCZ54QKHLZp2fDyqbUgmFgDIlm3PH9MJ1vesDuV1s13fZm5MDjt0Af1182t
6q29ZapGbJ/IIG636mbV/rN3IYiDvHElWRWr5qCP1pZSSj7zJALEVnGPrqAPFGYhNvHelD/PIXXW
AVhmNTBYFWMyFkTB7jkl7nh/JcnmEzwpfKgwX8oF1OUaUvTCFTIFXwwJCWptEeNFJjHEzu4UXpo9
XsyN8HC/ZE/oXwRU06e/xSr5T+nPfSK+Zm5sRiWflxhZPyhPXGPYocPdJ2hJ/pG95VO6Ps9KjEWR
1duUy2XWR27jb6bOOzoe21swJ3AAnoqhQ1gIamJ0pe/S7N60ilyhuvVqfgJmfpjMGRhK8ISBhaYb
pQyBxqLro4lqHa5Pz1nbrZ/udQKrodRAxhOfWHDIo4vHbpt1x9TXot9eKB+CgVi4qZz58HfGD7FY
jTSwd1k+5C0CB2K4TOxrtzg9HHrGj6V9mu5uQEojhahuQyZLt1nNYMmst4qTkJTEUUMSx6kkzQbI
o5yKRZsZ/u9m2OrBgyxIw8SscRSVboXMCM26roqxZNnToXTsyXks1/QrTuWh1NQRWWw4cJAavk8n
6+QnGCpaCpI2mjw+O2A7cORP3geR2qPTGrMx2LU8ErmcmA+DB7deXihv4gsqF/rHcDtL3B0kO/8d
2zlf4+TgXJJzHhChsaNZcei/rw8VrSFsXXkRN6M6KKywNCykCFlGkP/K9CU28LvQ9Zn/QafIJoNs
aZ/xmm6Wbn4GOVn/gbAXmr6aAo8GT7hocx8vYhEdXC2Ot2BxFAAatMs9c4OLqaJ2COXt+Q6t9J1Q
B4kNQUDUgA141wBQkysZoH7anb0FU4QXhMumd0Zah5xGsrqb8n4clF1gfPobmKRO0qwBUeseuFEC
f9sdJV+sRNb/pn52DEOVPBBbC37Kn2dCZapAp2R6uX8YgMLxUBEEHP5Gxgue73pbXvoq27ttnPYn
0Mx8LpdqXLCfRQWby2OkfkTkouVUnxhv8H5/xGD5invGNwwuO/uPpbA52CS6mxeAF4vn5OuPdQ6D
bWVUJ1X4OwkZU6Go6hxvLeKF+fG7xUMdqDFY033LhpOPbpLPlMYm7xH20Uena9GCGe+k3qLK65v+
yfOu/A1VhJqlpXSHkq8tlvxV0o9PgX3P0TOzc/IQzkgJVt30NRtRFZrvRzCEO2bie25Lxi9nyeMd
TzqBl5n+ygNY+cKxUTQb5jU7C6IcnYb0Ibtmo4RCTvx/co9ZtHbTcNMzeL7GtRq8LwNxeaNGIO5O
+sPiq7f0WAa2QmyJrkIeITycabdK79G+vDi3o/OJDwb708AULxCUQLu20s6K9atZocIxg5U+iaSW
dWTy9fWLoD8NVj1ah0q2aemXGouvPvmWmOW64odaaNIdTuHq2GZyT992GJDk4ltNwWZw/APOVIMG
uMcDyhozEzbrrjAv6hgcaDSOlKPjykAp7t2iNzs1Q0hblFnCdIX/MJ2xhEDhc6vPoFiDsA7VC24P
u2C+MynXfp2RqgWYVT8z99snKQt+gfZ1JVxMAYSDmJh//mlV1rJv1Zov0avDe/DGHYd+hKvjMVns
k2Ghq7oLQomidL4fTnG8Z5x+SS8VkQ15OfyUTMGLGIm4e//qJu0E081NPyz26cmtN9296S3t6LD8
onxH8O89BZ1+4qKzQSlXKi3/yDDhDQr+GSZcxOqGEgi6WU2FCx9n5+cFrJVY43658E1J+Our54Ku
W3GYUHHgpyKOmwYoxo7tFsTGBZ775s0GRlerjDEGbEo4TtaNHNX7dhBiFeXJWU2lHlmWBlcE5Ga0
KEvHAXl+CwgCuSoYX5qBfkBsZNUVYWYT/6Hs+YvVEGTEYGCg0XK7EzFcwEUbHyHJt27CtLaBQTvv
dEvv4GGnMnt00OQ9g+ftcZO/dJ+leaYHb/2umaSs0vUDBAoCHlS0huD7T9EE2QQslPLuknKiWCRB
RHL/kMBhBokiKqX9JTt9cT97ByUFSSPcD6CERvzXW9vlwQuY1ztFfsIQWy0lv3ezRejwvOTOWHS9
Tg+Aye4TKQyjRdRFnHDbOg0VZl71KkmGISNE1bSuMCZUlzYQA3WAC4O07MecYrNwgSnyoW5vjYtH
7z4V51JQli1ygzovIVBQ5hTdMR9qVJy+Zr1900X5FcKI845UGnhRnnn4wDbp6dKi1sQx7Fo8KsV5
/VSO8OldDKAIyw7x6huU5jfMXmIDg9wclUAWDS7H1Thy8oXgSIfUcdqoUufQuJGQF0E47kBH6E9s
OmumxZR+fxBpTHCL3VNV8bLXBr28Xms7h1Zgr1Pdv1xHpi+YlGKt8BevYJagtlIt9TspCmz2b4RB
+qTECiW9K/3XtbRUECqPRUbhdWGm/MP0JWosYtfRbNOUHJn2N454BRiT0vO5FiKx9kcWdhVhWVcK
UmiLkJwtfbtFqPEGkB0N+2yeE5/0fjQVXqhlYQXlCMQOjq5Pak13E4y0McsT8NPUf4vVPUMbJ5iX
QK6olsgk3YmPF/VqmGOhE5OBKTg9xwVfLYdsYKgxL825H0FCmT8WXduIZyTtKUmk/jMcRu9Ed3T7
8qQm91hgQYiTw13caibOuidnZ+ryMf/jnkmb01AWDo74hZeX5LcEwDwMpQd0LnBtmrozPLQ1/fUS
9atdcUemdYW3RH5JV+3hPH9M6vLzcshfnNNbeRw9HIHpEUhqVjCVGJvwVXKUW0FV0PU2g38PAAE9
X33YOi9KgjQWsTFXHfJ7Sl0Y3Q2mZJ7qkZfsuNkYzSQv45EhG4ANDmYVEa7s8mTywN14dClqdFpg
BUHaw31aWZJKqAeju0lGFhCy3ebfvi2tXIxr3RlJ/3C0n64Ykyj7taO03HFhEXbFMP/uO/ptRoaM
OAJeX33Zv3FigXijaiQGgA12RbSUY04Bhf+5KvmOxYAGvBVG9twDZCFYgD3Cns+42HjpO4NK3ZTD
dJVyQtHdsblnOnhDh6nFZAZnPQtE1GF4b56zlDzeDitXYIOS53MLUQLYVQRky46dmuMxVeZOo7B7
U5zr2egsfGVru988ThZ/ujOaa6i2egnBxgzkRcban8rVF3QKKYBimK2ksJVfKORy9jMp0HW9cAbY
wAfnWTEs62CYhSzs+5wFPD28IK7T6kD7cThzs6bpiKAVlhng+w98O3wfw9G/NKPuYS8CJn1Tqhos
yn0BKaCABDQyuqEy3GV3Q+rAu0NDwhKQxmKXdr64ZiXpoEH3I3aieY4m17AG9loTHTb/lUxpuX3S
2AsKCUdKwyfHjfQfhnWSo6kz+XrLV2LcXSnG0fDt2NDzvqQ3TYfCbv08kELAoCacJqANWN/n6HRw
khDbN/kZjtSJ1bod107PYI10PLjUXM3dIiUxFGdb65GiepOtnjCK5sMNnxU9MR25MJcdmSyiFTBR
XfIyJyTA+si9KjmIy00PS36X3yC8pEiy6mPLDkuncpFn5fRk8vTB28Xn5JIkvBdHyADL/AeMUP5d
+oFi2N82COmWDmeprVbd4HQVfDz8TMX6KTPs7vJAClgTH1AVxxQgWA5jBayLogd2fAWoGc/1btui
InoYh5JdzeQo//Cs/+zbtMV9xTtBleT7JS1LNCwcMiWJ9N9trtJv+WuRB/GUfmweC8rv/Sswh/2r
yZrMTPMDWaz0FT6su7CaYTo5nKgkdZOaGVVjWgdTjBs10D8JDbvGJ8Dki/d6Y8Quh2p5MhO7nakp
V3zL5x9j53HUSzqe5RpsGg6MdFHNcsg606RIj/kmRsahXi98zEsnEhxmfD5BGqeFwQdgDHT4okVF
CDrejEtmMefFf8o5/DnS3HeKhfDsD7jkF7RHt0Ra4lw8gDXUPEjZRFmIKgwxfF2A8R6bRY55M/8x
ph0PpHbCNnM8viQ6gyamzVl9Ptu7G2BGCtPH7USf8ijNW3TzPJiRv5m7dqa50hvx7FSZDNy1sWSJ
wqQ3RJbX9Y9HTQxZAvhqjYrS/yCafpgs0nybyQAZbeGGltB1DweK8UvUTy+7h7RvgxzPuxYuNCtm
L/zqtHUXe1zFDna6vXjPU+xqW2O0B3rt8XgBDG1Nk2t9abya3RXmWBbk/MQVh16DbTXCfBYPlMYs
slgNsCbxuBd9af9zR0oV39Gh3spgK/DcYvaWO6xXJbpGJ29hqpgMCv0+XNAxXtCeZNo1mbsFFOxf
CSzJyQJJJGNkZVQMy2OePu0PebxP5sLqAYa4NitoKsERZqQuzeM9CR2pW7+1gjMRcQ+wD0Bte29c
lps/BBy0YYeJ3HrRzp5g8I03VX73zHCoeyt0s/+nrk0esiYdWvG9+joostjyA7QAoBTqN6b+MGTt
7cd1nUAdUGOeZK9jgzCSQzJR9kgEfoy4PumymUv30bpnI+b3mQyDiY+J0lY7WKi4jvjRvqv4WWr9
t73suS9ceuoYSRNzYV7Ek6CH9bq1TIQ90SPtaIEytw8OpxuQIocNIRZN7MNxwW/awAg43eDWEp8c
nKKJBUdlpNc2Qpr/EGGJQsJxVggZjYvCG06KT3FjAPVRPoeSRWglwO1fnjL0BDScMYS9h7zgwOH8
4ZLpWauJMlsUcUjtjF1278ttGrewKFAFN7LfFYLUILTUTy8+XjEbES2RWIfK1BFyVTUOn8g+RnGI
FPckG/6bThLaCt7sV4Zve5rhlUljmiuqddSRfyKWKekzepO1h8QuV/pcdJefqg7SgJhxiNTXY0p8
2gBeBLI4CFeBk9JroN1YFrA1y2gtKb2mnuT9V2Aoov27UDbpWQI4USvMqxrY0gmnJ54cqTzNrG5F
b3KIFv9p5r232LY1YLTs9CZW6sg4vkCB3h98QAYxroApyk+GBsZnAJWeYGnk5Nqy6o39PNAIQaWC
w0NKCCdce0eZdjACiS27VNmJEn8kJEaM9/nFffCTOigk4c9defC64XgsiLQGko87qVXh80+a5kFr
onBKm1uORykuyQS5zLV8KbjYkmcHL3V74vRbhLmYteX1cm1TXKqK5dZuQrya6qeoX39c6T9EQf+j
ExZ92OSrc9N1NTA3qY3+3YexFDhnsAUN56v0m2egMNwU3Lp6wIbdTWh0wFGZwfUt3HefKurF9hnU
0qh80KWVWpBZDvTc/4DWX2Y/Zcw1TNj8yK+NY48OVQdQEkwHiOeyKLXH3Ifrf9xbqDPVZ+EG0Agg
rvQya4+uBCfXiHMzNGIScivtCAlHsdByCbFNZ0XmQGiJtch/lu/6Pp47vGI6MO7uakUzN75kBrPW
ERFhX14UHDw/s8A4PHJREfRn3YimkU8/7jEKgE26S43zGgoJrDeRHIikiUGND00sfcPWkTASEMEy
YD6Ik/QyQYbI7TTh8J65sNCUN5MZ6+eHLrfEbGcXu0AlCd0K0vsCOXBp/UW0BU9DWkXXliOigRF7
rVn3U//jPCrjTGSEpf4roBXkGXsq2VmWv6e7l5UhzAuQI5PidEEcCTU77MN7kGkb3NirwYyerd0D
OeDv/2Z2NHqpQlPSPOSJYJkrLfplXCe71V31PHSfal+gQG7TZt1ej/NPMH67Fe5TWl/Oqg2aco2U
AHCe/LSjPKWebG5PwDUEZ7UP2bnntljzJPhtMf/N0zhaovV59QUFYowSDAlN/T+mqNrkXN2qH4F7
BUg1hQZx86zNlU0cIhH5nJYMl8+FFuHqlNMoMX8zs0X6YiyNVz/qXMK8sIKUoqCBwXtZm0qBo1yE
KPZQEXufkfKNqCw7hfjDrOnLy6GRji5ppR8dVc07leJ5SfA4zVUbW5Rl3qkZqVhULIqkej6EdHmd
gKS4TlLyzqZNhQxuyWh4sOtELW+O/BQYciJoIka11DnuBDI9p8kIez6VrwwnKjZMa1CoK+sZrm9x
k1ZaCBMgSadY1IOF+9i1R+kVEBgAKXr4b4++ejUSXyAjXP55Ka6Cb7wdlBKNdvB6gTLYOkk8fjZ4
RhPZZGZHYwxFl4n/hr/cm9DAKW/R//G7BTy3yzG9mmqqfzC43mxAM1Ha+nyFGHDPv3l6zFOC5Z8+
r2Tc16meWh7KQPoJA/Sk4JVDRn0XyoRdrmrY03JJ9sc4uGPnIwBJHrH3Dzr596BSyvZX2WZZcb/m
V9QMU+CFkFKp+AYvl8InGHJ19q7e76btGtQ4gFlwm6xm+sBQR8i7PwPVVZehlK5SXVoKmheGrYEV
KB6QSjII/LIJRinElK6GXmvxhoMZhW7Kn3nrFMeTwUxUwH9loMJvXaNZXcG/WFePUgj0/9/HcTbM
X/g68xvr4Lfw1OCtUK1wEYu9ugeo50CbiH6PAOyNT5w0klZYPyQPJi88gfcAn9fLbehNenl4TmXT
XjQFiimuEbQVrVexesdcHmC8OCyPKYYoowkMWAPYCIfjKcJV5C8BI3pFQd6VAN9M/zbm1qoGVnQW
TiriN/rWPqzbt/Qef6CKBwxyPqKtzHon7CCJRLqFbvgRcUIqepHy2i2mLm4A+M3jI0UhZZSNvV4Y
svIfTWxkO+hG5aKlSNVpEEDrOOeEP74YL4CWxqPFYrZiRiw7ecqdVMXqaHn4JV1u/amA9uPILTzB
aTueoIg20NvlYYnuOatgbGW8Kwv9k1KEcoRj1j9mZSEonq6PruPZuF9Lz90CwXqEOcif4m0IFE3W
b0oC+zHihqRWxwEaqK6bNMnrsvHySrdnow/rXOA85QJIyYXOCnyotBmLJvIJsaT2DOAhiJdcyT7V
9Zc34AkOicpV/xD+ShOXndvIkBGMCjKWXvsUZ/s5NM0qI6tGTg51nKrvODWJvrrf/EtXxcu8JATx
AAA8Mvy3C2nc6uhAMWUboKN7KHBN/V2Nq69wnxt/6QhNrFbqEH75hiwIIpHSOd2gPm2jHRrpnNfM
0ucQCrfDx+h1J3vK2FcxrzjRqPL82ksqqmBYC5/TiaoprR90cU1ya+ZB3gV2V4r+W/PZMwYKAPQf
moeZ1+9U5N4wlg0VEZgNOjCfcgEa2MOhBtOY/wFyjiYvLqKOeobZCN3fCFzskE9Ul8SCGoQEphdH
XaM+oieuUO3bJh1dG820YusL578bgaAcypJRgfv8jZohibgYnXTlYmU7faQs5whdAS4Axo4tyHw+
y/bHH6oFB2OzcVRZgUfYr39UdFmw+NYhyTg/1G9ZgDleaOBsBGOT+cU146iuYxWRSK8xruiB953A
OjMJ+q7HjcNLPKZiswUHS9ofHyuK30GFWXXq2EzuNSA/wWOqFddvgYUoD0iotkuSpeGr9hYB0Kce
3eTPncpK0ApxCOtkFgYs/GQJQ4nyzO46ZwjiYfTlxlnJ2aZdm6MkrORQ1zllb+3b1og8N3/VhGlf
ViSNlWPR//nlZ7DwjCcj1EberhBpsXI38pgWv5+Jq4STCufItnHI+ioxuTkUreo5GHElHr+AWHXc
y3DV0YXvn3sUlO2Q/YblDPjIDx4RTYKvd6crjognCSftvX1AZW/38N3LX1CdHCfLfjmaEVg/B1yy
5u+cgVUmTgkoX5+eHDfgvUGKDKBpYMPJKd6vmZJrGWIsT0uRQR1puBHDoBDqhewbG1nUaxAnbZqh
qwIuoaJ6YyqpbcWs8tHQEeLH2cgf7GT0IIvE47r67kC5Wch3IjNitzBOzS9/G+1MskvlApVHijMT
J9tsM/Ixp/7mhytnvXTMckNvE8Z1qiH6YgM3Z0MKKxlv3gq4DZNT14DG6gcInFRSYEAn15oUU/rx
wjHYVMtrjTr561kF1PgEabxSySoNlDH0ddYAIeQ7FBWyYUD9MC8xCCKTuAttvEmSCvGHtbTpZH0l
6pKNLqMztr7mYydW6F3+GJZY7bOErSOd4z9Sp03hW4CYR/OhMOkcFwU6SppcJTAwE50DnI8qoZuj
SVVP9HnBZGZXOLDZNkuqsyvntwrTDq9dWJ/HFgiUkRVJyyYHSbLWLHXC4lYgV7XzEdPA+1W4mTll
xvTAsqNk41hL+soBTCE+iAOBTvR5iV6iB0L0wBg1Xyi06wXCve9/NOrzaeJEipnCzGqH/NM+HE3T
XH85Odfh+QblPaRs+RTEp46qbhVzSeOm8H1683JEp7MvZ+kOBh1verQYXkSr/5rZTNh3B4rNtTl1
bRKODRcPvrNFqKn3ztP91wSxoHb3WWGmBpER+q+agzhMW4IB4BwACjp8qWakvDI3Km6o29Qi7mj1
H+JRr9K5IrIBsC/KGBp45Z+4yewtSTq4qmeFVcvLxwnw21niIZg+xbjCQ+A5X7K684hKd4DwTUAU
3uy78MwcOCZMrXlqygzCgSi2e0x9RU5d0NdEtqlcf+oWQyvzXA+VzsOc6yEk1mfQDDXBnOVxXASO
0ZvYeQKIIg1yRuVy+MeU3wI9YRLTHURbzQZqL3gB7//Tm8MdFLWlk2rx1qWihmBgYZ8bVb9Vlx19
Jl79xsQhDjw4WKukJuLMTuhAvTDZuEUYLcEVuMuOVC9e/07AcBsveTw4wM6hd5bZjeH8gNRHrzec
tJPY1A0wIYaySoQ3XrMaJNvJuinN1SoPZsbtXdpxJMKOY2DCjv88x97NBPRoUZaKrdZO5SSduvOx
7TVgM9Pzh2X/DP9Q5bSGaxT7HGhBAk7Jrfx+uB23dbTPo+znujtNwE2nCqmbX2xQona2HOIFiP1N
cwFSaXeCDuu07G4BpNSAuZaa2eypIdYkx0o1/rtydFxypU5ChCnhnh21FQj6RwSmUL6XkfmTF90U
4/tpc6Kge7SqPOzcHiRxTkGq7ynfDPeHpaZ+3U6AO3Hr4Iqn/XaZZIoOS0oV8qGlxvpB8aAokg3H
yfxsxxTHN3CtpZZ8HjmyBQov+5Z7XPGR84paGx2GnW6ZwbVjZ60yCk5GdbFHmIP+ejKYJe8rgtIj
sLeh9vwVtteySHGnl4lqr3LYPj9gPfJLAYX+qRnHAVPhjPtg1pmVDeTbqXu+R4ZNcnl0zMEn4b0m
T2BcRmpAbKxiE/vbZUbSoZlT/PWxFNWsKnX58Z3Kb4P0P/SGkudKoF5tSVp3z0iI3WI5l7M2AFsj
T6l+31s8G48UneYjDsanMWy2KWhD3ePKA30z2Srpyl72ZOFj7Ub9lGZbDodMQlH/HV+hZ6JL0SYt
3zSbmUCqJY8ElqgGzgF91jCqeis5iLiPXWeq1t2GAxbXKqEqb7PwxgyIy6Rb5Mh/yYQp/Ko6Tpdl
iAWi/nLiJysswIgT166AJ+o+N7+wS9/X872ZLLzbPheKcwPuMUH2S4Vdr+W5eXXFr6vr60oA59xM
fn0D4UMUmWdBaG1eU83AlB+efT69RM/HZhWW1VNid8gSYIV7GJ3NLH00FzD3y3vjxxSP7Lfsv7iy
mndE6BBZ1He4Tl3Sigv+iA5AjJWjhIw6PmNTIQFfE/e3IH9mvuKAVBh6Wkco3u3/lWFLaCZrqhI3
7yhEI1tMhEoxtUbCaWevLGcS763c2E2pTEDjCt7zQeQZk9rzPhNIzAkOYo+w+VoK/fBc76vTBe9a
eyAJCG69UgA1xCFfJQFr1ayKnWfc/b9cUI3e3ubSZ1SzrXP+dZua5UeH5c8cTxGQIx4VJnCkvafz
fRPoNYRMDSIydebfMY5XTlp88YTRzBOs7d6uISIHuqpMMJjpCAjj0QBgzomVuf/BYQNQxAIZpKBN
PWuyE98T00Uiy/txsbtkfZkQuaK/v+/2y7sLExao+ttHCU+y+kasdHoNmjmVCjIUVyASVUzQ0Zkc
s7iAoNcqUvqwjvSvdNty8su8ZTnY3p2cEJFqR9kS0NW35y7yruhE0Bu7Dn2yreFN/SjmjkVHxa2N
yrxisFU2Mm2D5QrSCZtHR0zgEE1BMavkp5UxsCR26WsEoWhvq+sSVDQlylQjysDcDY80zkZ2HmC1
l/gdMTxk5pCPTVqgtWMCMaCEXYrMdZSceX5XWLScEeUkDciInvZZC5nN4ZOpFQJvJ27dy2brGSBG
6i7D7EQYZdBXBe8QJwj7lxDR5S+NizoxRC6/akAhaLTZKicWErLv2pUh/pwviY2+XSjlYNFdsh17
1B2JfzEjN+lK32p2ZOo02FURx1ZgBnKpdx9R6KTNqugr/begwDWsRv4DTgAl8fH+UWNOIGklCVCi
r5oYMiMH6cIJdqrGuZCpKUG3YdkGBavcoJCrv6I5dVZ2UYeIRHWJUtrHIWRKtBF3ljXs4PO0p24j
kI/HkycdHeUlyGlJAC8cdlQwID+EGaPImnKJKtzN1ZzSjsui1xHVn5YUAz+lpUlpMEBEgfB5wqJu
2Wg/9EPGsYQuBMXtFFHTtfUyvbvuXypf+l/XX1BuOeUL3bsHau1EjJ72eSoMyY4FcPiTIs+AolRZ
GEV+Noc2HuK+dsHF/n3QF39JDwbpEvIS4Aqknb/i3agh2LwkaLv8uu43i3aOEiXm/SxhmFcju+Z/
9yoZD3jxVINHrn3LDLP8QXgou7dS/AEaveiPgv9fpO+nkYe439e2z0TKI7iJxcZ10hZIwSs+MQyr
TZfnfL3dAw+VFZ/gzxRTs+fjp8bIOMLTeAYgqp1AxzrVBUOufSW+tUYLFKCmhUwqs8zXke6wg4H/
5Be7ZyXg9GCqoMKPmVFAZPidkB838/QBcFnzpcHHn4gK6TRDkA5Y8sHhGVmgV+sDMBVqfSAEY19O
LS2GjnO1OQmgeQV6f/3vY3IBq5GEHzIhYcCf59Qh3EGzs87aNiY3ik+1dMBI+jNBAmFs+o8gx5lJ
wnlrC/djbNSlJzYF/jqtorh/el8o3CzPUSYi1Oz4z8Url0U2cI46D0BQ2WBizfJTSpkQW/ufCWBn
qjF8J/GnaOQDhN0uzSRsu3j5vBnvGiCVbRQmoqWIWjzrCnYusndYwdrUdTl8Kq5B7pMi+sD93NlQ
fZfCPj+kNfFugjZy3VUDxKQapWO5rWX3I5lyl3gAuoY+vnN9yxQbjj2fDhwZG1MboY88Xs4U1WYZ
BsYmdtOI/+T2utd+8Ej4SBvq5bQT4RilLysWZbVUgLaDT2P5tEZ/EkXlRYPwncPLHxFf2PxEXh6v
CKhyD461WysICuRTkq64NpNF5MCcEZzL+SIogTLaAkt5+peazZWpqKTXG/vXwyoiAHwtDr2Rql4c
n7GR5FtTlcEyfiggk9jX/2167NEnFV1WUoMWIwKeuBh+1fGgm3Q0akpfgcG+QC4XHFdaC7E/J9C8
xg+xPtCeDfi6pK48K1y+xDKTbwSWF95TspitFUAQcyJwRZtZY0yub7ptdxkTfnR7vX5FPSEbYB5U
K6Dp1XH5+uw0ta82tpKsTpLy7tNFc4Q2iC7tRU0AbxkHs8q4vCDGiMSwLKpOVa+dDHD7pGhHS71l
QwnS+Y5ewuzDy8vovGJ918X8qvGZiupHKD47WgAUIJjZK3cyM8koCsc5u1GPDsi2rI80lTmfyM9j
FiGVr87D/JMI8E540QNatrVMZ7kn3qqhmY4K8XQIaxoFLBdZtjtvd/4j5J4gghQ3fdWgIc0Cl+01
t7uTTUzt1RqUNcdM1QNdwIVHcWoKto8CwdXalwvVujiCJIHMVK2IBhypWOWwMTTU+a1/tCJhhURD
fd98GHzBISrT2wGhAa13B8iu8FOFHIW5vGEDDttVtyFM3nsTcxHtid0hCDVj9ejmId/sHQwYR3Gw
xJuQ1pUIBhDCr9POycB15O8Rao5N56/M3qexY5BY1ByW2iJjJ25b69d16Lx6izoSy6k/ulqAEhDz
fuYqdF8GtFjrDHxie5C6FF4ZmerS5oNG7CvkzdWKDNwvumYVUcTWnxzK6DLDsM4ge8f6NAbSfspg
5WHvqmSQ3xVXbVYKXHGKMXhQM0Ywhz5Jp8krqajEx9uwqVG+Lx66Wi7s3evvBEM1pW9WUP3a8OI9
kO6duZbizWaRYVRV5ViIRDezkN60X1sVMyBWLupT/RQF+r47kr4SF0qyQTqJmwuUIj0+iCoMTdfa
LNF8ZW4GjlfEzg8MhAzn/e/uen06N2r6Jx23vlt2oODrlLkUN7LYWlhjoRyIxkR/cA8zW6g3uz9M
WpJOwrPpXs+UXKMu/i7d7tNx9Qi1aPvK1yx3ty1MteMG9Ex+CyYG5un7SO7YIh+88upc+ylfWNLP
nH16XazFOezG42jHXNMVvNMXQGHt7o2DgqAr1Z6oz2gipZlwOGLGRylq4NyK8CqD1BP58b0/5sDX
CEgyWzFZMe2D0X3UJIruyV5cwvCeYQje+X2N9H3nYkxfg2lONYWEwxsMBSHSbsR3lAGw6QIXGtbm
QeKHgWxPzU7h3Wn5SQQ3FespQlqaZsr+fx7cTxUHvtub7Fr9f9hWDaWIDWZvT38Cs84gvyw21voe
gI248Fk2M/ggOsKorlEqtBactrb16dsrmWJNUfhmSx8QPRybuy/6PjYd/v5CHmZqs1dt7PfVDuEG
rZAz924yBd7VeyjrEMl8rn90fllGb45xuf7Lok/Cqlhv6sOfjbdVhfwLofdHlRxCdC198whA4d5k
K89cadA6ab4Tz53R2LHHIdOwfaeKSG0QwXUn+l8vEyrmJoklYq72WSblFDQhg+M76BuBAXZxsZDK
kvTmzF4giNiHlIg3EJYiyxrtxUF8qvY27nXFpNg8q0wpEl/L457xMkNPF2Io7ZcVx5xGQGBpKTjb
pvDr4YQvdyu27SeNwsT9jx2++yJo4QR1p8sh4+oQWOeytX3A4BH0esIpfLpUYYT7xN3du6hxGRJ+
l+/0p+sVHkWFAosA01GwYrsFgUSBHW47OwSZWQnt70VjBPPbVZC2R3IJnnbP0RaNGrQd8hUMuNHp
l0z6NEpm6gMpeH4Xxo6W4h/sZq2pgaaNz4KV+ljJPmxazYZ6GukrcEombTK4d+myRBDYYZ93JxYr
ELC4mIw6AHbi/4GSuhwxMrJSybZAae/3Fh1FVEaj3DQt6yYX3Q9AknSqgyx6b/XEDb0E4Hb/IwNm
oAj6C88ZBVY5+W1Hge83uG/eE9Z42cqQFcZ1G0zZELfF2hQFUoyb9Un7tsy4lYFybeYnypQFbzYw
hX9S4fqMvAxl6jsbH3k44ZEgVlXspArdM9NOWvA8cUvgLmviexCVh2ec5gBhBenNyEf0nR/DR8di
QIiWiXWkccfj8h2l7yTCtAQoqK5pL3NRLSRRzBIQf3DvWpnsn05n4r8kby1fBhDU2GH3E7I/ong1
ipd6SEhIVngHk6So8spXaXxHz4a3uZugS+NbtN002Y7euK/HjKXhYpH8ck8OGMoNGC2EVzRZUIxz
0gLMKo7/QIyi+dlzg2Wq7tYNGabZCOsIzZuGOIyLcqNDZHeRjttDBmX2utgz+PbwAf95JUHQITMD
mLqatSTptX5YZ3hLA5Bfa6v2mQQhp8cDt2Pze/WPDId6IuoPQPFBDtTGcNUMkHAOIUN1fdJOov80
0vLsxVUpcAQpHh/qC+g//+YFDnqOyw1kMBKhNFm8bLpoFzSRhi75U8+5yJnC7+PbaPGHYM2oXkB+
FkU41zir37/0TUQ+iSIl5PKIb4Te6VEL9Ez1fuW9ZmE+PZVfffYR2Is/2x1r8TXBoSaEJcaz8FH0
pDLHmyNrSgkxkwpB6dMYbB1i6F3UhMacsPP2V/M9Wdxaq9YP7UTWqlytfhhV9kOMz9tt77OvYiLe
+Dl4wts78IVyj7Rh29zRz6NFivURE8vsu1dwxTgHNzVjPYY/iYDJNw0freUgH5jCPEcM+/1cNUF4
z0cXXWVIxCRY8xwRGhbz5x0KPKSA8O8IcRlvEs1s90wZRX40X0TSqOASaY42kC67XOGMn4SLcE5P
NwHruz0LZADN0oTosRswBC6YgdUIjkDHH/HECFQZk7CrsHIYi4pyjKssQzcPEQJ93mpHOaSpjVZA
3XmdYaDqoJnX5ZxvyEY2GldjhRluv9E2HaRmzkDv+J0Yl7WscBE0Wekw+ZOfl0aYL9A6hrMQ5eCj
4hOD2YB6cQtVZLOpxSxGnC2hxS/XNIELO6sx+wZzB+9yfWw+xO+RZVuQMdXx/Tfa0HUbtHaBsmiC
ZOBLQBbqKCnBTw3d7/uzilqcKh4Lw7alRNT8YlW7bCq0VVv39e5QacoFobnJiO5W6WfxDnHWtNg6
DXCwMNBkqPJvVfrlV5Lnz0mP7HAEsiWy7C+tOh7aDifD7XhrVHwkAjhrgJJep/exAPROdnICL9Wk
fSXG3v+KTnWEs4wt2hCYlj49SeGonzxGe4fbZeeJs66FA5tfHMfRh6ZZyQuk3TinFXhExAcvVE9e
SCnzvmjASPIhTCTf7TLSTsQRZHR75NQQGv6FS80m5Zi2IwmSV0YN/1tc0u5GPl282QTtSEsBl7W7
1eXCNNo0gARK8B89uARsXcUojBlCVzKjAdYeuI3xNpylDHgn9y1cslOxTXt6OVHEU3Ktx4Y9yKdj
JfGeKbkGl2iyEhgLU/G20aNO8F0ESBZl7xScMmbCD8u6onIdeAXR0dP0GN2FND3XkGXHYD9K+Uh9
uKdMHaz6YuuADqXFJyavYuPDfMxCN70viGCurXmL/wIYN7krP1LGBykKrKAE0OI06NWfMvTMJFzp
o/5b0x8UTpk9ixlOoiW7dkK1BnyZ+Y45X9ps+vBb7BHo58IzwRhpiQvMIi0muaaic1k8fCQ2V+qs
LunPF73XWvchH9HYfWRLHyt60/a64/ptd3VDNLk3aeTWgFmhmQZ9aj5z2z+/ITnBgPUYQzoacvhE
yhpgHc1zUUEMolwmy3PvvFv0+ui6hKeu2w/ZL2VbSjjn1U6DcTtxVefEC+fKR0NpQW1A788h2Ak4
/1JUMu3Ge6mysWDCFHnokSN/6aTU59Z0JFZ2j8dqMgFV9s60o+gGvlZYz3mga7h0D/oXU7evpm64
IJ2ubAMnbP9pKOFOC1SrihvflwGWCmQY6AVuVu0vxvaDq5nBSmbG6smICQo8pXAiiHIE/d5Caiem
m1zN9C+VpkyZHwK6voaoZGPDM5Otqdvd2ZLABrh/cQ9L16zxDPgnXWJMd7e1n6KC2sOmarEDSvA5
xfjHKriJG7TXuVe+iTW8IeCaqOJ4lfL13GyGn4pPczHExSb+8L+c7JiCxzG1RtEZAAVRpnWWUx0a
7nhBIFX7Hr4DFd+JsaG7hHoKnB1rZg4dAreyXdon4TN/m+ZLci1sD5W9UleUZRcdOKjJ3V8wPIt6
7n8KTye6ztLyuqQcrCGdbd1PBzKDsy6hQdHMlnjNmrxWiJRXw896P/8HLZOaNT0RbHY9R461JWhi
92n87HOafgJ4LmDZR0AOlH4do8MF/VKulmvxtJXw/RzpqxBP0HUOaf1BkVQEV8+q9zJWNKFVaeC+
EnMjmuiQtu4yRnxK80xqTTlroZKLzPQIRtqxumnimXA1RULGZ+h4igBfX9M7VhA0/O38vfIZJfn9
8YETTjL8tkfROb43VTC64TB4IoGWSpF3BiJHzm9oGmoORSkUIS2g6CF3wWXjpJM3nyW7pfVYGGLA
bO3YzGkLFM6tWIFWbVG2gzFB67xl5W3Qd45Q9K/v4AaQ6ekSP/SxBJC59NkszGe3n4qE+Xv9wM/o
5NRK0BuwgjigFTxuZaShul9GezcPF88Y0OOi+bG1lmtOSCu5tr3anOlFVMPZOcZPiYV9DlxHVc38
K19a1pum+dIjZiN0m1or4TZ+mN2QPImuERwf9xRvjcB/dP+Q2H8DDQfmOnLtx8yalccAJ5UBkV8j
l9Ask0NdjqEAH4j1NdEsuOCpHzHZeFlcQiq1FSLWq879dBz/brC2i14hZ+82ikOpjWLejfYGETz2
DSqe1m0CprPhYOTSldIrwFXDn9HNJtlS3Fr0lTNVV1gKvjzq+QUFHgrcjWg4QPpYaOrkvLPYrP8h
+fGqSz0cPZO7WP3ZCEQDR4nogrsqKHrAt/IrAPc8sSAio3d98IcRIA8wDsGQ2VHCmSOO72uQ7mpw
T22hrJjfwt4keC2/z4d9Jjdn/lYp2vKDVBB+NkUE1hM/+9lvH5DuicYGt6fKgeqFMlCRVTjBsWzG
FN4Vtw/3Y93/bTL+S9MOzPDovUuwto4vAPw7uXgIuXKkFvdW3kYW82NOzO/uuQgR/u54B7jxxapX
5gBJkAZv5zvy1QyjnW2K0dXjjxG0R3DVSFDp4q5vR7sjU9W6LjK30n3osBws/l4OM6jvJCffm91Q
xoNDun52xvo3tnjQk9mZF4TsuUz2fCE7JYcvcWyEiINWZA2P+04ime/sQhCTErqy5UhTG4uls4pv
OHgLtYj6gynEmbKYOIZg2MqRAi2RDxKKLB2ggcNATsFnhulN/atWSzOwVsLXqLEm4BJWqzTSFz/v
BqY9qQPqOk2cs+vQWyMp2JNFAaJd2/C2fQk8EkHjOOaaLn38yQayZjQ1uOqbkvZgdssHC4Oy2cpT
kHC5sxZFjRXknronVSdv0sCIOpTidE53LImGxSb2DnHfAsyc25CyZ9uM6U/2LG1HIhrMtiuXlW7l
1sdATB2jPoyQzaez0i+bIdA0hVAT1aayMRl2ai8XDUkgz7vFIw+hQRsdSC1bUZrtmEfzi7nnBpjM
9A4cLJVgrzZtKe/VMPfHNSalB5+VWZYG9Evn5G5iE0/T7yvdE1GV/pYO6nWLRDOFhT92pzFF3zk9
nN50jpPJb6r6ga5ba7vEfxPkGhEJfgS2NBNwuiZeYYaVFbEF7CywksELKoyCpPbS+vXkV5CrXcRj
dnuW/HJgN4vf1SO2mUoTTWEUPgYvEgUIB6no8f0Y3ZDXneV4F8JjjJGw1ik0M5qmhFSM72x2qEBs
13EWhEy+M46vRPZ+XMxmD/AVZXUwmrcxjoPiw3LUZSIYjb2mr2jfH+EPg+RwmWl5uiQH4qBPm778
rkXDJFOBXyDnHfHtMuyPKtZs+R26ApvWBMOmuOoy7a1i+RLsk0MJhyi/Ta5sHu95NPFGu+fIz/6E
ISQVzQl2kkWrZJiJA0EN0URsHmYtrFruLTqh2wXscy74UFBSju7Dq1Zc2zUDeAsWbwLVflSYFJE9
LVtIpIOEaBy4hMx9cSXUziMNyKFnDelQ0wzDn65XLZS+eNFPieRzIFnXUMtkVRKbsa0aUKYv00dp
SBH8DgXLL9aHpai19yjhPRx+yiIfpFPdH0AryIWGehiHRMzCXb852y6I3pNxoL0czZze9UFja8Kh
SVD+xWRQbdIi6yqTrzYziYDGKP1K9GUapb74oGqOLM7ZU6jxAswGoPTr18/mo2CXWOSIdM56JEe1
7MafLu6HQtbmBwFQgGClF3IsBS79GJA7PPS4kpLdLjI/DJ2iSJMmYYsq0Qi81B6i2rjVtvgVjK4Z
bco3wZ5aV3Dj5pTRDXlK9dsHk0Jm8PHwr867yC0TTqO7knF9UswMEsmWwrYrH9XYm1kfYqVpKwHb
Ub6ZduZsfVOr/E4VlyrSQrFqTN/AG5hK6vXjnGOjBEYSQbQePRGEXByHaugE97HJxriZDvEHoJXz
72MB859NyWl/vQ6tX9Le3Eq/Jd/l7nIjXtMLEqxvlp53XnUCs8DvnMlxjw6D8yBzFUFuhOXZnwhv
UyzFPJwKdb4OFS7hyILupXk7xrCPN0zehz3vJEDucYYU70vISHsKRQyR3e+ZBDdvipK2MVQ9uBjD
j7eJnWakwZxbAkoSdwzQO1hjiLWCfPo466PxO53/HiDwQol6941AY89cEuLkfMVzhKDSxOh3w18P
SLaF+F5zwcVS2v72aFHkuj1Dai65u5B0n4GxqXDXXtMqao4/fqY8XIMnVDik3x2G/DywK4T+HjMg
2yxyUzH9/SwBmVODPilUbEn/63MRmY3XjU1oz3yCf1cD7o2Z2TLNMBmqI36WL7VxW2bGOrM+eKgr
LKnGM0YRAUZ3iSlIN4ggkXaVDeDqzLUywAI+TyouErj6A/XCaWB/BxzxxmegLeoFosF1QjvBCTTt
NCdISfFyK+yHZCEawO6IM+DhD7KBV0VuVDP7zLRgpSFFU8imV/Nb0UTEbGQpCyMlVFdtDTdD4cQ+
P93CYKkxaoDI45+mtLCevnGucb2mAuRwl1kCYaxqcqVPDrFTIDM6C11haYoQjvaSmgdcuZoWq8PN
cbPp1GBKANIKSU+KFSNL/NLMXZSbAY+sXTz2H3pOIJ3JBLKlRFkue7s/X1cqZChkoTjTXPC6y9FN
tmlcpapqQsqvqqFKYGEmtS3VxGJt8u2qwFZaCvM4kSYJQC4hTd4ItncDxxDLC4btdm2WjJOBc6R/
HYGfsDh2xjJaXKTzI0lzsArHHGNTGTeDItm3DM7xF1JMXMPW1IzLmjYxGIwFREbAw+35xH/Bzsb6
+5mDVb3VjUpdd4qe/AMVnjdo2yEOjGdoe8ldzkli4/2IRZjvzeo5ZQbDpOsL9jNYoCtJAU+mrDlK
2+4eHuHEdBuQRVon0RC9R/QBoZQEC3IkxnrPE89IuykpAYsh3Rcwv4UWzACqUEl66A5DRgMc3Lnq
GQjjrhOn+IXz1MuaQ4w9Y7GJYQRMZOZp83++vJu/cxqG1bP5N+RMiF7r8ZNmHNSKYgcmd6jqPVUS
fIpO3D/XZn9M7rdpZVnay2RsK4LnKiiTeNu1D1xntmlYHHXETA3UZZsZEwP977Ji72MiTDyWTur3
NyXWeCkO0l/4cdFTu0Ae5Hf7uxhAyXJe35yAcuTWU/RsQ8rPuRnMSngb6CXj9s/FJs96MupO4J1V
XJIglX2Z4khNK0RzdQT977LDPEbnXaL/F/301SYYxEy9kE2X61UpIG5RpGWwC5CRNz4uAY27EL4R
LrPNx1EYAHopH2GUUwbxlnUPf/1pp/udgffrcg999aZEXS40pLv7hn75OL+yW2Mbj9IEIn2iXrSF
eDpbiIb4642im4C7xHgn/BKePzwuyR3wwhpmApmFM8plY71C+Pws1aiLf4RbfmjCoB6NbNJOnEBv
oS5KLPPJcYRkMAOnwhCkjYJrCaMMaebbyrLVZsYXEME38Oi/90yue9HD+1VqwlakwEkJ7a1OVfMV
7gCbE7XKcvHf9F5rw/a99kKfq0jQAwfGy12WH0UPvzcKVzQlz8NwmclER8Uu16MG+vElRBi5XBZY
PsoCqLNyRdhi4LBlvezlL9sCWUq8Ni3U/dND146MD7NlGDr/UAgr1V9vIvzjgBfc9OUsxb752PAm
IAl1QBcvnhq/ndlvwpH84V3Pv8AXdM50qF+p6rKP89xc97UuCrPVoUEiFvo4yvYQQXiwYMaboHX2
aK/7ZLVjt8PIbhz2eWzlRtTegDaHa/4bDKPEyPx66bUi7O39AS0xGVGvkZwbSzg8RZTxr7AjMJHM
pVNxDPRf0bIB1mppNgCyOIwY1gUZXNFkmumT1evfopKkxMuRiHPYVRH8lLwxnfwMmRpK1Ccnf5kZ
zkxjHOP7pyjp27fpgc1QUhZB3J14mR3dY4aNiz3d3PD2cGFetEHVCxOhLf32xSz8cDn02wjbCbfa
ebyA9RU362KJ1QswcUBNDvM88Qnbv4n6hwdlbQQLAUplg4fd2HSvqs49XlbMPuO6QqrqG+arSgGj
fojAT2JqJDbDLyZTq/qbypgPWRF7O4QSBZWOlx/sw7iVm3CoURG3UqW4aUKJ6lV6s9EBT3gojIJl
GL9+3u7dj9v422oiGCRHMXfqswsndUMFK16sgjcfFtsredFKYmxaDvP/ME097UJpXVbd4wu8egqR
mqk2PYaNidLKJsUKo3JPKVbxPe2gdcgdNMoEBc0Z1hQDMU1qlEsdYEIyBMeWnVQqgwvuA8I8LMRS
JM53VJDMNUjlJU6nes5TJiAtK+Qz6nM2niJ5H244kYqMXJ+l9LTDt1DmWtNdaaZehEtL7OmB3a3Z
T2avoIQXko0CeGJ9pnJ4re5elwfz/0F+ci62faombTB/x22pSAlZ/38sBV4vITTSzdwNvL+2i3l1
KlVHQqfkZn2DYRJiytQIl51tvOd3XxJ9O0A544Rx2Wzqnvys75rjOZy/RnY9gyN/MdW/8uJGEL8K
xs7QfbvcKqyozl0MV9VPTyzcX7e/+eEn2vNV6WupiSdwIKOLwYGM/ZeWYE/VyeajdJSxSdh+BW9y
0t4WkInNo0nXGkXgmG+ki2HhD5WFaR8gmKe71Ljy6IZU6KUb1oARxXMECEihxpw8/AAkcvUqjqvH
4pLS+9EzvptvzXpHXVEQr+DYv0V2atygyLBua8qKVJtGksscAs0JFxVcNVasZhlpkVZahKZKm5IG
E/msCTjslt3Zyxw12BsyvpSXOFP4o4oyW1JTDSpncg8Sgy7mcotsrQtNkshseGBuTOKolE9EO/Rc
O6I6LwMera6uwPS2a1gYsKfmdMefTC30HdGZMQMTSm6Dtr37i/TKcyTyuWzIBAO2+viuvaz+fXAk
KoO7RgxZtUhP/oFr3y/bpngKIFFBt8os51GAyGYrOQaEsOVLMNuC4Wvi6ncRpccJOM1XUFxDesVd
noZycgXuMcY15QZ8hzMU23kWFuJ4pb6C9gH4oz+o1qIQJEQMRBrYL1KuKqMd1pWkMHhpLrijrcfx
KXoGX9Ycdf4lT88hOissmAQ5ShB80v/ULuQlqEQKTpsNM7lEUmrF41ifmhx2b7/srDQBmWiW3T/u
gWKMZ8hhi9Qtz+o75NjVyFhd4vnybzjkRB4UgulkgCMVKHHOsmnWcAKW4nSfCUief7UwCAbrKlqd
QFPPPcS1BnbV21QMUSDzWa2fLxyLFVXw2WVsfV012wLfC9O847i2FmSgY0Xh79Nqkj+GJmKQo/mP
q020fUNPTFtPmd23RfTJ5DFNfsrzsbor1RFazqDEcCjW0SnsNaBiYq4AeFGscSOtRtlR0AUKln6p
BF663fhtJXnf20jl3r68fIKXUY5XXhrj/K5A2ByNuElVuQgHSa82nRSHafqN4zpmED5qxviTAxfF
4cwrsZccV5HEyD8m51fVebfaGQfhHjZ4SLkJY66sr7JkNa5rw10sN1CNxsyeVHfJsmUJcs8YR0Hz
wGLGFxJ8/fICHtRnfqAysu+6vWvWehuPDx8KYv2SLQwpV5s6ipvjc6hLJGInMrk4u4sSvZgjDnG6
Jj68yHqtcoFF2RcsUwHXt7MjS+IuD7OmQrfoYsS5NdK4vSyk2dNAQw5akTdT3s6iUnvdAtbNrOjZ
cajtOnRjmZz2PuAeCGvQExxJtJwUYODwu2uauZfXucgZhZ1Me/Pnfulj2LoqCDkCbl9uzd+65OaQ
T/xAdJFvuF2QHT00E9LuRUupske4HGB13jaVFSIPm4hfzyq8UEeImDgVgmvQibB5PJSl2g7QH312
kPg1/faTZxWcvcCRhKtB5ir8i2xzj40/ePwfFPuRS7kx0EdaDnVzysTam7EY/qvCiUyiaY9eVIjU
D24yG9+S2nu+DEyUOFgqJ12Lw77lzuYP6WBO+JbKbxlcALc1e762m5xbNcnH08S3opvuldOsR9Ad
HC7iaZn5EHnf7yfnZIES/h6vHvA6sd6/46NbY+5cvChWnVQZxMXDku6q3zVTomeVEMOI1LCgyAtU
gWVRywceLNuwNWtIMg08qvtQcaEFEQE4BO/bN0QNSyNGcP2YQca084GjDYxv674We/VMzA8SBHq/
SDvokvVbuxpOVUGLKOrliA+r3nXAu856yUh5qdg2OUltNQrFaBdYZoGHHH7l3bYM+pJM9yJiZy2H
IAfCzd586NnMLVthasn1bNwts3YM5Nkn2z/6FhRtZX/uQ+wsWuLNt5fegAU2OuSgn8TVMjJn+F/w
nIR0l1yq7sCURiS++ndYMaXBrHF1c4l1mC0v+RxcLPgrCNnKI6bBe1z32E2Un6VsBkZXa9F0q9LV
VKSEuP/Aw8UE6xy9QNTK1pxZYvLlqFXaKNiQa3DVAap512mSLAbu3O26Nf1gJPichlujQW9vJwgb
RcogoAxk8Q2OUj6d3aJialjfI2h3qP8JKOKGTj0e4oZrru5cAuyRfAB0u4GfJ4MDLtLNL/Llcq/7
ppMrpzjNukwdjttT7ZpVml2gCPD+0XaFGP9Ya9kOCGj4m79ioGnsDGaPnXmOm97YXcurK5jBj/fM
yAb51XsHOdtZ8wSChgSBlfNUmg7ex3KM7tMfIrbgREMKNK0IX+Tq/+QgLtVMxdbbVIb5cz02S5Ng
ayw6OXtlIfPEaG8z4QNHFsIyG0cU/PsWODf2TJ6CpS0AlX0PVWpxFQkknaWS33vcob7YlutTJowq
36ZX0LOwoisTrgFO92EOHYlReehADUxbYyZLvzcLQ4BNlPI4x/mxu70UDLeDWLpClf1hHebqx2JL
Ru3jvsgJB8c79C/2ShPReLUrs4GWxs0+qIg+G7OJDwCYIcxqf3BmMrPvA7Kx2mBPPnwi6mRHGr8c
xMmWlEiP5PaT3PX8IBPHGL1otZW8FqX2hqdzCCAjqmsWu8xlWQPYPqItY/mF7cUEr23n4X+kvVew
XfPvRHgcBB1sohyhZ3fGe8QcnrA6VorFRRddrKsfkXM115jWEZhG17hIJ5WU0SGG/FxaIyhL7af/
duow1cMQHWhDs1oDYFTh8waiv27pv+aF2JLFFOKfUMXBJpVDD8Y5OO+bfw2MwKxC9Vp9MF0j72dp
+UenjqljuPTrhkByf5xMaDUxUk5vo/cXWxBlgKd3BcdGrvkmBbc68503jq+y7o4xrAZafm6fwa1n
DNm/sof12MSUh3+wd5U3xncmbHmZnQvNYKrlXzBDejybnjLfNNHK8lgEleX5pnr4Py/t03fmC/zm
//sVNe07Mig8WbrzfhoJJYO2xDVHC/B5jisq4YCF/OqYR8dqyO7H9TfKPdu3KscRP84/M43YAU3S
RbuoTyrep3uaCCQ+UMqfvGPomwGQAuOoYe/0N+KwIglWBSqXk6lo+BEWgEu0yzH3Ss2JQhl9Rs6f
+LSl1mO7lzCQudahFtpuLowUXTy3gi9H7C+oJyFmvDFBsL058pU0ZGWQfMc+ktKHPw7MkhKJSCkf
GvBHh55LZgJxHKsstZTb0LJxvP9/lZSyXdShJOsDtJJWZ+9duoqN+lh3T3a63XGTJSiiTSk+56YZ
++wQ5udkXA5boB0I4cydkZyQdJ+agx8+EyYxZC/5Aw7cnKsq6ePSHpNfRLgAYhfoEuxBMQnj7tm3
R4fP155gb6rpqM4um+XUMWvAfgVkf9uFr8O1q039GERz9NEzzJLFLEkqfy6zZxRyZ2F6b6FvFfo+
5EvcrLETXyNT9rn8F56zAwkKq4W+bDNcQ4SuYodyISfuc2/s3qUzmpbtunQxwwqJwKLwY7QElskD
knPZ5j+/uF0K/Bx/gjShLBW+YLyd6KdC4KJE6sT+7HYakEFs6uyrxhgquJtN9HW26lTNrBPdu466
joi5kt/fQY96uia/hNWIBNJQLttwhqcHRnbdeIWxxj31fYpHHaJzSXtmnabvjMm4W080EiwU3EKT
3qfHVsJ9Fqvnj8BwMg4SCqu9eYA5YA4z20PtzmOz+QOgQFToGhJnHyrZTGY9yMLobHAvdjWwUu2F
Qk8CX3Zj6993uJQMkHFM4hvO4v9VdWtX6fA6fiLtPIUJHlOAWlReIdzRpY51F088YJx4noJ8fLfo
Dljits/6tihxpf/n4IpEnyuUPkwQEX31IRlyCITE6ClC6BXfqzOc+epkG3/yFkPiFEb0+631ZMC/
3T6DOmn20dNO2VfAfSXv6Vz5VISBt9IGXcA8GAw+w5vromGkXhbeaRv60WNgqfcnhzib3LsMcorh
CcCS+BjT2zS2lf1wtnCluL++epFcPuIwe2Ks8qRhCmmlCMqICTcClb+wBEpoYFdOdjI7cgtTzDGF
J6z9bnKrsKUr1PvSG9MBlIKzsFjsEdfGiyQTwNYE7InmLNom+DB5FBQJrzqBcuVkZ051VmGDZLw7
ldXtZyjwV6zPVR0q4/GMIO0UhjN1fybyTMwLl8XDkIHjQak11NK7puITYqfwc3//oAkUNc4YFXq8
DkTT9vLPtN/7qdnEMEKIC0UxdYMsq5IzW/jjQc7VeBJHo4WxZv+tYQdrbSgffs49uajaZnnqyGJa
Pyxyz7b7s+ZANUCCZZYYvv0yBX90c1VhqmH8oDxIy25V+IOpBZLVE8X/0xaRfkF2U915bpE6R631
Fr806OwSV3gcZj6N26eXkQ9aKln6sidG4/9j0oQLjTNf9RC332uFPcOAH4PfhInj3B55QEEvoJEV
P5UBmy39a21S0JOz0LwoHPe336woh3TTrzsvV4qQu3HBOY82oNsXvytvs/F/AKLMH2fUiP452Xk3
6huRPLUnWRvP4tok/PvRaZAyixLIi4G5knlKOjOpW3T+Mb/g9ZalFV8uV/JFvvcQcr4SZvFFqBsg
CeUcnxj6gJXa2BP/pZjZI0hGilxxmmCEwCuQ5wdB+P0EDIflHmf3MSK5jWzXHeCJykEt5f0CWJLj
vemUWWXo4XwceYDj8fyJHGS9+T8j9i9SEv8tulaRkfZNO3QUu8LkgqwdDCcbDgazT9Hj78SqMa/O
MKpn5Wip+IodPAMeKipJjpuZ8BmhUbB71GJv//EVehFKHaJaM+jra/pWFnZZ0SQAFL8KXSi5moC+
t/tzNMPe9sIo0kjstzjfIJCyaU8csdr9WGxKhGlZIqLk5SuCFgjLFQTPSByZpWG9922L8zSK5ZVt
Eaiy2KjW7jho7Dsiaoa9Y5PBksTYPM/rbNijLIDhZbmqwl0k9QJA9L5RLCg+HQO5m0vMYqggBtgh
3UooUq6dSLqZ1E9pK+X6GWWPfqx142onnAHRoT94ayRdkUExsrU+Pt7tL4UzIYmaL7JXujRhtqdg
QzZz5RFyb3Ud0AAy+0htQWszCec0yABPQtQC4w8wR3SJbzJAKGNsMwaVkF3qWM2WAYJJ1QAqquhr
BKvSfDSB8Zuqb2jAkccOlEigUB0/jFT+NXIUz/6DPmwIamPZ/RBNQMhfExUvp48tuEdeLgmycwnZ
M7f1XBSTOc7l/FhtX62Edc+bK2OhumuS41lUb90tVe3V8KEbelSjaCo9VOzzs1T0F+pPh2f1/NFX
NgZhv/jgxrRVcZPQKkmXl/4MjjlRyvpWt0MAV5yprMRGVnWHfrB52qVZDj4jprF9IZzcb2U3g1Ai
PsW+Bxqnvm0RhzhNlH9ameWzT2Qv49vsyu3Quz/rTkUio6K8sau3ojGaexIRk9qxeEg+leFkee45
uXSMzQr9LqkFLaQOtvrkMoynkxafOBlNR0vCnvk+vjJfgkmBtlZ4AeGvL+2XAJOnCj75XcW++O3C
f1ei9Swtca3gq4nOoGMGBr2KLzRd4I2yZF5G7pd9Ffksc8KkCi0o88MiC9yUzdImkAhoEeogRUkf
Gxoch48ttbv99m8q8uwsN/OS3iQGfKuIJZt8M+s3DXK/6pNflI7RTZc/gFuid2v3tE63xFrJtv46
WHkLhJrFt5ouWO4Om5nUPzGP7OE+8zeAa4nD9kiavvZZxYQW7hQcqQzscAKLWgk1lDeeHlqVtMSW
SVMCU3mSQsz8B9Cjoqo/Z3VoiQrUEZSY1P5XUwTYB7IPqQge2Q5Le3E6xCpKozTRPwZXCjoTCnqb
hFXNjclR4PbhKgq82fdGkT0I2hFtHvD+EEswaFdcMD79uBv5xKgPFBdTFPZevZ5bgKcVY6aA9y9m
wEoAJ14fD1EN59spBZ282K9ozsgEMxqPMoDYsFBA32O46sidM9raO45JG52c5/FdbYrtWVaJxYUb
SSGmnpMuZfc94MOgYlSz8tu48GfSP1V/GlAIm7xfD48wFUAv+p27UtT+3fWH1AqPptnx93f6nmdI
u1Y5081ZdJhBT+emQHC1TL95bgADtPLnkshzvecpGm3tUmuypALPPOT0Ty24UghON/SnhGGkieTE
+vf1kVXYDqASHUlwj03SFZtFfLKckwfriRQPd3XTJxRMatAdmC9dRlfacdS2h5JnwgHy6cpuGUBI
E0o+X/T/CPr59RY7Ghpgsj2wG1yXBIbG0y4eqNOi7swxSrztmj/O88rK7Pmh9h/kigV1tNlrBtq9
fEw1FPDPuU0XM5PM8ibDtrwiILCU7lpv2y+gqGd+XpgqFYGaZDc3RUZXj+KkTfMKOKNFgKr5PB5i
1iTZ6ZA90piREIJHrQSZrER48TkvHjbR1KcaRa1ZtmOjJHhwVKr/ioD98xeRkV/VTtsxPki5th7q
mOjmytcDecWtIm/xuxDwsLq9SYTGYn8Onyq/7w5EV4iHqagARtgAlYEwV44HodZHIZ8i7ytXrt2y
5i5ke1Qx/G19iDfcwTaejAmeUHmTB5LFsKbPFIZ7Hz3K6esHv/v7JQpHr2cIWNMWvHzsByrWDCjS
GSlV2eICyB7lwMq7dHBnQRyDbsMYkFQPOqRc2kTsvl07EEFQQMMeiNU8+tYV0brNkk7UxE6lcqSm
Kn0MCaR7he8bnRnFN9Rreg3XLx9dJd56/bTZVuJMZLto3AXGYpg2KMJAGkrMJa+MGD4SOez2UtX0
IirDBU13DtbsusVJwpEBgOZh2V9ScMmBdnAjToiDpHWrphI2yWqRMAaZ6LHMTHhKDiooaip5V7gA
qU7hAr6vTb9WZjDqUuW9PMIIR35oN5oR0M3cIGZTTMAwv4P3X63IqgkIZYhThdS1y8nZYycBParD
Znk46+6R9S3ImxWSpaJjNGjb16SFCvPG5Z/NZ3rssh7uDU4IJYd2EvsVsMDmBj4ZFsRG7bP3vaN/
s+tBNDz7U/6LwPIZYhkyYW5p1iPyjQ1f8wWtVh0zaMk1zmp7kH7R+mnJt7CFytS1lTr68ozS8F4U
eEz+gAak4lFMyWVQEl0zP1oo7VndMr2RCFKkvtetvHX0AvEIai7yqo10QyrcFtzIKZmZvlES9teV
L1kxGcECbon2clFCERfBItMYvQ9a3YuM/R6gP0dbMNzFhuZKNeHGyZ+5FGHZIyDXyRR6T1CJ5lO1
TXwNZOaOiM8ly3rdYh/0jqxGPUBG5YSGw0VELvblKafGD3YOmzvS6lyYRpYz2H1lfd5qSH3oj8+V
ytkmqT8ZEXMdMBc1+X01CuqLDGpzrQv2zerjF4w1oRajpr0FuEr19+atytSB9mgkQs2FoLkoe63D
B4KWEbPm8XMgY0DR1orgM3ZosnXx4uEnVKi3ViqUsRJRzYlO1FzpqQ66G3AHkOnSLsBgGPc3q5QV
SJtw4S8DceCrlK+HVKHtU1BR1T0zMMtBm3hDIfi3BJpVoXto/qCGg0P+6IsZwFQH9pFiPkf82vBI
ONEF7eO/PvT9OnItY6/NLVFadn1d0DF9GeLgq76I0poTOcHR1+Bsun9deYsTsjS/s/iDbjxgfnfV
8kXbE/emxKDZqI49ejmah9s4VPqWe6dr23h/wDZuINzByaZ6W96FBM6cjBxdFHdzwEGzVxhgjD6a
5xj5pzS+qfw2a0G6hvCeNHzbXxRycOh9noXOrNH96j1tNXOnxxXodi47mn7wUEFll2P8mYWbHUzU
uhruA8KqHtg/z4MbuT30Zw6NnbE/EaC35RpVh+zXZX1qVPe1VkXXrAsF/1Qgay/ROSIg/vohKQuT
VTBpTwqayK3HkkPBi4RCEPnSVCkSpq15XTlhXeqMFD3NqhJ/jtODTDApKA/CY1JjZh/ajsu/7dbN
Vjm4ygWukZ/Ff6UbjEvY/PpeVd0ZqI1I7WadTx5u4ZAS3pbWsk9K2C3qBQoqBz48UxKR+CJw5vAE
QDJjxylaRx7ipJFMYnozHcrZsiIPBZb0hYeC43APLQpw8LY77CYBkQK1tk76PA3utx4ph03dRwFR
sGiKKSiIhd5/YJCiHBriSP1GKSlTgP1t+y30EANlFo1u+cMeqAByJMiCVG3/jD0AZyiA5FPeq2VT
TNWYBNthluIwROAFdFP3xmNLjrc/LC5dnWs9ixg1XNIfqUl5nRmRPpH3GzSF8daItVAiVgsNME4d
wlAG8qCmOqtJLqowff3JKRYifUuKHmefiXt3cE4VgCtefbcPTZ1hYy3QHdkmeekpmfIB+4iqKT+6
BLE/y+eFhUZurzu4Mnl1B6Y9Hiu8hi3aTmNjPTuN5e0k0H7NA33TpzR/X/FNW+YsW/GFzEsiNJ3v
i/kTinFRNDgJTEuPH/iiB9SwvtCvSzXfjPmUzHxXeY9b6el50b1su6D4+FS8tP/iS1i8h8SLksa/
k1PBYMbuH7cklI139FetrAwF+Ak9Xo0NazKIWWOfocul8xrtv/LlDPhFZF5a/Mfo45BGnY5W6B/Y
1DPxkMc0fx+UgjoNXvpXXL35Mw1md+G7+gQ7K4aoqslMdWovQaA/VYJwV9WxSyx8INJpf1vo/pah
Fj3lxmH8WA/tVymmWu8SlyYKNjGV9iwt7sXEtpiBbmzaSSJg7mht0ahf1zH0EFbw2oR+eFEyCIWA
YhHf2tNtGAyXoi6rheGBhJ6uCAE1fYWC+1SVT/oycvmvKgZAw8ocm4vTSOeN2OvvlW0DlWouOGOb
yg//PWzIavd8ZtK4+NcAdn65pkok3BRf04AuO2zljMA1waE8X10S4Ooszq5zUFT5gf8oJTG+V8OB
5jbhxZEfuV7S0Bu1MG4Jg18w3f1vvT1G+x2XnhZj/TtCUWDsKYs8wiimqnXCAE9h2VvlscnZ01fx
xsXLwnZN/iov44IM3XUZPLW1PiuTeSBaISyDwwIShjwkGvagQ55yzb92LSMkqhbj/2v/b1VE7ZWX
vYpv1V8Eh9La4hJSyjyrpdHQtbhDs+1xcw76KLv2vhw+fId2Vsi57CmLN8huUv+l2TvdGXDL09es
b2lhTknDDcDSKXqVJJz1URrOAXOqZs54+wGffx4CqUpQawkhZCRqkYfCO2KfhzRdV4McIblgIIqN
xfWBsjarMU0RkwsPeRBRlDir4Cthw1rnJurUDueEB2j9+gMqubitUAIlpUztwi4KiGRIEu4PK/Yr
QUCddV/SV6Xg63AP+WfyxJS6eAXrmR+lj32yrZZJUxaQYQs0y2+Db0r6ocRZzwKm1oUncUHodqDH
DOv7hNvakJr4xqk0zfaFjmZ6Arkdc7OHyS46JuFeXtgCl9L/u9RPGpWB67Cv916568PLRnRF8El9
IOm9fYg0nrB5JuuLaKgFFuRie/NqPVe00XeMJcTX/Scskv4ibaMHMJ8OATrXdvOeiLQUCoikGMrW
S0/ap1/5JN767Z7cz5PzEkK22RN2CAbLvbLh/zFFHUVlzAS59+5/j38qyniVLk1LqeFMSdZ4bxoH
LyDOadB1ZnVwnhXFqDzCxWEbF8+DHJHRZrWre0PaU1l8JXacZg6M+2hXFvL1drNOZeRCI+9Olmmt
GAd/wUxqjf6PTE7GVIFM6Tdm5207QpzuwCaLkg6ahdr7iPLsr0QRRicPew8Sw55tcUdXN0deeNiR
5dkp++tWNCsF6lAS35Z6I5kh/DivWzyCoeUSar1jFXmJ/pZaq/CoFNS0Dn3v+xRsyBYqbUxFdt8u
ECZJaGv7e9QcYPoepknjx4GrJF6cEGHoG5YH4clP6JYL+zZtOKqZnD/2MiBkbdaxxBrW5QIs1FlD
oeUnoHheGMxPldXthc6hb6jSm7Tr9rlxI7yIhR7xeH+Jb64nO8hz/rsKKRmoU8iNAGFR08smdjAw
TZ5lnQGCMKoiMnHIoui8pgTj3CYkRkNqiYU8FZU4Qh8DR1v7+Xde6naMg3rWEy2Oi5PZ15iv02C3
NO5nVSbybFXmov0OxF+AJFDNHy+8aF/7KArsB+o8tww34tgUrYNdgV/XihF0Ua//UZIL027B0B12
9RMYR6KpD8/S2Llw6SktaEQBNz+gBdAiQn72+eWL2dtkTmeOaIfrfE/8dgHS+Ow2nXzh21o40syT
TMnMjwtNFSy1ZKz/F8sYiTwDKqmmqAiwPvhTOyu+P3VX6OtcEsAZXymZ1wpJ7lnDNx1cnWaASwdP
zNLuqvUOY2xbkgy5TBQ3AAhJXSWzJlnzWmy8TVbTcePpXiJg43vNQvJ4bJ23jGXHY+10MFQj5tV6
1RoLGoeFJBfJEtJCNCN/CjHn8jwgxu7te8bi8TxviID1ky+fPtghk99YPwkgnDnVCgxiK+3AhfGX
kuvrMrugm2w9vlVirbKIcPjdzxT9XSRTQWjXnSfZ2l+y2nYAipHi7ZmgaDOACnpV7qtKjL0C5b/1
ZcH3pdyRsIi6oFEen3zTazb3VXFhSaGexkFd3lr7K+KedpjDJz3CTkkAdCmm1kw5gVHytbJYXnob
CZx0XmKwAS9oEgZcT7tQXJKLXqNJyPf2iwN44ZpOy0lnHTtGqv+3iPud0M08Ba1SfZ5M6v1/tma0
iBIbxdoIh9TeYK6Zf4mwLWygpz7eYfujShTPq5W2rKec6kgJRgdM2dHpXdQF579sGOEFMD73xSRZ
u4Wj+caXZUUFFEbXzm8RFTYmqI8QCOZv88mUG/a6T121Lf4Og0K4BHR2Nx9+BZ0Uyy3sCX9IGAmo
vbFxulHqotIRxheDkR65GkRO403UE1ek8o/52ZQdIpFxY9phv3F7SEQVqI1fz7IJO4FLMHQwA8h7
ItddHsJAbVln9ysKtUFwtQZAohBNx1wvEUU2vVwcfabDDc+r1TgKzXI2we4WnfmcrsWWN+pr83vl
SPt/uAVu5JpBr2uQgkJnOCLJJBmjxUqHdu2nDnfuzh7pPP/C47nWHuKRonyNCs7GD+/avrEahzUt
TRYhH8Lm4Xsoc11xnbyyQon/1YBlIYeXPPmvtadedfh9ro1JU3GHtSX6HscfHbsrOVfDPhklNJEg
bnspejO79pThJNWaAEH24UjinJ9VnEkL/tY8SLyHrJCmgUoekR7V0hDXVPO0k9sPzvPoduLSSm6f
HX3i0UGUBX8ozhN8lY9nDPvZ8yxNNZeQP1pIaO+RASl9m6BlCQlp5D5r3whxRFxf+Fcd/QRiWa9n
DNgx+y0BjMvxEb540J16GwhnaPunkPBaOwXswpW8Gl+Weo7qSjh6CxzPwlAbNhaFK9rit/m3WSYS
e59/7g+lJ7gdaOVvcrdmAI8Kt+hIuW3T6QSL/uSsq564sO+hLXyHJzd/LABPqAh75uGIDIglFDuT
oieMYAicS2V8YRgeiGvhibqLOOv0YYg2YR1q5WTX33GwzGL56lAk9xCc9J1aFLlEL8q1oFDLyZGm
9L+sDWeMYkLTcoRvA5UV7Ed49vDvqtcuKP+V/gsHqQV425qhllDFn8J5R3Pf5khBRV6i6wqtM0vJ
QYhNBv4XgSdHJJVkIOwLAXdTdL35ZsecLDjcC8J9mbR3t6Xjh0ZNrWCuyayW4Uvev55qKYJRDz0N
ZIdZZvvu9vNeb12CBDwjF7SlT81V0p8r07zT82f/iQ3rTqxhMZARhZocLWfQl3XOpTCyS6rO47io
tqbjUO8VlBmkh8r+/bolwIHOCPWu1Vt2DEJ6xRCltFehB57KGSbNjp5i29beBoAj2jX2AqhdaRLd
QrBIjTOVq+qQvkSfeIzWUDaScYOjFeEz4WElfHIChRA+aDQIS1RJLZ+SZ3BW35nVBr0xagdX+5xh
iwkEB9kUWAL8581Wc8i2UyZiCxfK/3ENpglr7QKwtQizzARR+vG6A15r11OPBgYSC1hudEop1X3T
9m7a/rV2Tn74G7nzRpFHTMKGwwv0juEx0qxLxoORLnShkqDIOD0b26jDLSOHGO2EfcBYYiSJwLsM
ABGxpT6SRZRoBG0Y2csgJWDybeAoL0F0uWPlhzX+ZSW0XvkGGyIgkPOrPSVmHsajkSP5ms2Bs5c4
cWGaKkqezmtXoyVvXEHOMp36e2Mhz9nfIE1Lo6cCIrPRlp/asfUaxCOJmH4Su8hVXA11bINgZHx9
aaofwwQt4b5d1bf4mqj3IPCTJtj3gRF4EzcNck1fmXloPwAKq20tb5fCg7UxFv+Jb/dWwo7ijaEi
X9Yh1G5dohIejoeg7z3ciNSAISppxR4qFPY87CYVQGTCjdbtTOP+Ch5AzTfS2+jKSZT0+gaODx+v
hM53hwqP82712iJAFUjijYEZy7ZE42A8L1w9pPcCb+8aDub4VQaLARFF63omJaFY5oim/JMiqOMM
LnGMsxP2DFmLqrndSsqMYK02F3wUTdN43Mr77Pwi/exGpE8LahlIBLB7U3tVZEsJJvHVJunX0EnO
vuFDnrPXmGaXwe2up7PTZOiOiJ2bzfvmeilyaw9S6catfyvNnW1ciBtHKTohnflxC+PCnK+hJqll
wFFR+vcCgqAZ3omQ9VpZLhWlgM73fvfRin5xxsG/ESnXHOROWvUQP+uKVLi730q67rt6Gn5kf/9q
vOLuXMzAHnIIMJv8OLIUtx7NC0qIRS0jr51z9GIjRTQhexaZlfKvbe/X204rrZ7/QKFkiToc5fbZ
DWmMwvrrHoq1u9SyUkHRdV8LljuWHAM79T60N8ya7ddZx58my3CIyPwhrM6EkA3ctd600JDB2IOU
qbKMuNdflOs15/WAvTpyrVkbV/myQl0bwA1MWIuMNHOIT3ZTTcWBQJXporuZF9J5CbHUTWTxelmx
0RyGwOpjUuydA3TlSsbqRXiV5j1ZIq4fkMm+vt8CDNY/w3TdhZ+u1C/aMfqy0FSwrzIhBvOeyBZg
IvkKbWoJWCYndiSihdobQjAq7qiJF0WQq0D42xHh4YdmYa6N48nWaxrLxBOmyn07IAYDb+ZWblrS
YWwuyaC58OFP56WbXxpbuMZdVo3R14gd2jgTRoCtmIAmHnrl0X2kjsSCeE2lgvia7s1caNZPFKFf
IBJ5ANNFK0ZrEc28G0j9GUrKrsxc5WRNdFIYaqPz20lQDZFKqMmpuuupjTEII2k3sewrGGkb6YI+
sGRlRNXOCR6GIHPOwR+xS9kz8ZQUpd+A++k4tuO2OQlySj30tyQPPnlRYF2tYpfzUJ/8CkixkrEo
CTNjIeqqtgxc8lUdt9Aj1nXeIJseoRr3mo6eLDQfB6KLgIAvGG/ItJaFTI9Ru0MEM5HqvtBrLsmD
pUly9kr7a83Gp+d4bHG3pVppvlad4Mud6zFw/zx8oFZnkae0KZZo2XfrNawb6pOrA5qXMWF8rw1Y
XAc+thBfapR2WPAzjbIlSvSqIcv4j6KP7KbR+TKBr8wJWyEskX1+4yUX+X/qrN6boPkBGpYGH9Qh
xrHSwQbUGigpUzqZRKnr0a3OwyWNmWtnc6V283Q4pEJfzHaw8jc+ivbahpwK3uIFqWHoZF8JmgKO
GEQlZ1gwEYMPWT25tE6lvF5s+eyXsGjhUXK7IkUPxPEvlY+44R7bhxka60GFNE57hhYgNL/1yCvC
qsbD12vGBdfmdsmu09n3If+x1pdRMejUIJAKHRBUvW5/XO4Vkb9jSKUK7F4pO1sq5L9R6Id6onHP
KqhYlXo8awqCS7rxO0sBYcxRxRE0d1PfmMjmg/MN00SjDBDGfz1ncpjVVPCSzwy+EMgL1iQPrtdf
U4z+y5eM8GNkkURtLNiwap4wi8YlG0Ps6sh3eMC9/snTIDiII3tWuiEUU2N1jqr/b9ltPONlgGo5
YUgRATPDzfyMgGcmo7wOxi/55W8e/1vqmIxW1u+ZhNNZ+EAdCeL8VTT8I2RmdKhtQwgn61Hgnt+D
YjOUve8UO5FQvQW/XlxrPe2+gxO40K67qeB1td2P/p/ktBTNGpPD/Gd7cRpqYvfWz+nChRiI+BCE
E/g6p53m4L9ZUBIvb0n/c1hjg1fJAeKtFxujpTNPOL/wamxnwSiQooVAWgvnIqMbwK5a8WWfVBN+
qsUdPYvc83sLJlh9oS6fTES7jYtoosOS0wjilO+tsPMOHSVOLqknEw0zGVDiXGGJrKSL5ywM6G1G
GZBY7PRaZoMQLZIhaohKGYsDubVYI9SP1+MRIPRQmTB/QKre82m7HXFHP3kLwl4b6ezCcYln6Ks/
Bpv5RScjItF/Sgo0xnP5BWCvbBS/r/IjSbWSmFhlFt7SE1Q6KnNWspBe/xkj+y1AsRrg3vyzDnUB
Nwc48U8PrCCBfNVUONbOPqnDQfmv1rwVSqJUh+CxdFh64qJWm+6tjajp/ekYiqAOu+ZnjDIe4oAP
h4PQSuUaO7Tbx24JPPAoDKLzQE/nvV5zvl8ucQmZ0KPwyrtjxXYXhL1icw5ke8TvnKL3NNHYra7y
Pk69891ydzubtXIJ/jLmVBm0seEHYGsDpvVXLoZ8vJYTaBerBxXYWB5Pcc4oR4bVscozQiTvmhXc
/s2Hmrf6gbH7A8UcH4TiFSMAI28n2w+DxxEq1SohnfTQZgPWySl6Ux7xn7nFkyaQf33T9Hp+0Da9
GjJ6wfVsuDe6OIU2RVi6z6fR56mipoDpqE2A35UDFy6CJBwp7TaCdzjgP7lVIKP+HdC2hmQSwxaE
vQAWJFTse6QAvmy7sLFAv45vYcveDA8yZyX2pYRmQR8plwJmw6RvXVkWWglT3lE+M+sS9n4E88Si
/jx7UGLVI0wiIf2rkp3xMPKr1a2Qo1dkVN6yyEuJ5PNDe4Aj5AXhfpjtAnrHyjVMC+GvdHUvMwrt
2MBHZ+ILzNkvX/WTlfiaxiH5ge1UNkAjNjQDYW5RW55peElm5OWlF6RVT7t5s+DF60XjGiwQiDDw
ArcrLBpUBi5RfQL5YrOPETCaifTJ7mb1UX7m2Ye284RFQaVHAgLAikLvj0kqx8E0rq/uhvoIIr5j
ILNja7I1w9/QzeaQjCpJQtAyc/4OhhUC5tDePjOxpbVIKbPBMBirc8pZ6mGyDWuNZEE4N5HwcPjh
kk0PSs4avngxQsaI/gXF015d7BqKl9QfFGWseiCvA2O0AR5vevY7WWClderxN8KUjmQWZENfEbex
OZBwb3WBZoJFk5drHLqrW3LhvKunjtBLgjk1wOmTM3GEy+4DbCCuFZribo1DwFMSIzja/IM5rfox
MDdyejkgdyBi9Zg3g4M6G7pC6MQGDs7Ku39PvoS6xE2yf4P1wKjcrval6fAsvfOup8sSVhiGzsDD
BKcBeZ4yI8yUubLH2bn5wL7x3wZsBF8+HFXQYABumITL9A1yeen0CmVa+WizX1T/uNUlA9HusD+o
IdJzS7lPvw1VDo5NBSZnaXkaIG8AdsNGdx7DCc+/kXVxGzUNbz5Nz7RoPRPmENTi0zosMON2t9P3
OiRnmX/aMOPMkwNf1fyW3MLmwSwDKTtjBHD9efaLdORSuQj6Orag4cVwRyXm8Kyt3sHaud2tYN6D
2nANXtOMaEdCmFwxK6Dc5QI/PCn4g4j3issHEh9aDQcwv2c2jVOr59/HcQA40i1OQ2I2bR+D2/kc
J5iwByaqzt1CqfPsMfeo9n3MDyqQFUeqH0pjIa/NA4l23HOz6uPB7gITINHnh6XW3vM69ZLZ4b9H
fKEhNd2PWaMW1XytEBi/akEq08iMEeeELULfgoZTmmJMVMBxyYje7t2BVOG0TfZZ8sSHB1W9opCv
6UTucHncOB/M+KglBaa608dG9/ZQWQY9MJgHTOXabe9TOLlhOClidQyU45D5dR+t4LJ70Yzi/C20
5FsB/+BTKVWqYAGYG/0J1dx6acJkKazExPEB0L661AgyOYGe5X7RPpItTJFzRl8CBvUV6y5ylxRT
o771PemVWMr+7LnT28U3WwC3KhlpEU1HG/IIkPMZS1IrgQSVOz377dqSugUbes33JUwJLxmvAeE2
PVM+mJSfy84hYi2nxf/gBC97yiwVYInWBA7uHcg6Kda6xBKBezj16Zitb7oVfejhd/mN/1bqdTq7
b0UvtkbwXjpYxyzYA0/B1ynsrSC4z3w8XnTt4RojDvUf3g5hGACBA8kVNgK6+rQ9ywKvlrEl+X/4
MDCbRa9S8PeWbj3kvLuZRLiqSIplhEO2xDXJmMhyfnrRTqP4oWqrgLnPCDF3FYAvc+DI/MTncczP
MFKHZ80Eh3yjsF9QJmpUunmRYV/1jPv9f/0CcoLQ80LpFnOTgaucHtpKcHm7Eoe6sR8qDpKoGz0c
KaTyjVa2LaXGboflVR6yLDk1cZTWqy0ArJQ/mrkjGVwlmvHlJj5F4X85/oXzVem+9ZgpoCL4SYrv
Swc5ARGkaiaQicyJ7fylYEsYXtU+ezpifC3gvi/HhMpcAzAwxko5mp42Kg+Db5Aqs3xBO9TGvYuy
SzmiID7sp8x4jIrBpyrdKTsC1T5JT2akONP7UL+yf0EzJ7ElDZiVgoOEgCscY6m/zQ/LvvvsPxLy
y4VNcMfZJ0cze6mGf7brn0vixSualkwUdcwAthTqkh31MoXvOpM0njY5b5iPBz6dDkZnRn7ix3N0
fQNZu2QD3+wcLsQBSFeQtGmiNVHEsStthfRDty+QzvJr6LnvYzu42Eval6LM4IURcXUHdG3uhbr0
PliQBXVTfoZ4yDjGf5CQoCHH//CEt8gI2pJMsxfMgIyUKxeuunT8yx16MXNOkJNp9Ci9BnYdW93S
JA6iQmrmFNVZZiUzbiO1imNIQ2E6wbRL+lWOtui91mLe0pxV5wwVqH91u8uPV5o3pFKNW/N3ThmI
093r7sy2MS05XWUMs7PmhZ7OPUGQEmbUhvwCjBRgiPJhzQkBivhsB8K/Rpj6Cn+Bg1jFKTPDxnWS
HHIqZYwUWY/tsokWSx6YD3etL5qpJzaclC1KLCo4YpCOkZ+YZyKQfeMYDMcjkfCiIWmcGONiRNUU
l2klZfSZZE2+Ba35Dbt9b08Ec60XHAg0215VBE+NFSfLwVEqKpliCvB7YuYrO99WJHd8pEvgr8L4
AHvZqqKXocel0qxaJ66qJkvnGhd3oghAqU9vU+MDCFzb6eAuv/etqYfOLFdj/ptykBEdSGzgXZxX
PH7p+NgPkhJBRzlmdAMU50rBDM/EBn/PJanbehkQb+tZURACdB5okd92rwq65QnXqYjz+t0/+4EE
vOJWCzghex5Xpahg2v4+EryqXfW7iH1cBIQR7IcHaWmTRnoMsAeDVHN4GPAqqEbNsBqqqxspGFE/
p0ppZamh+woJQN2ddeZwE4F5aomfP+WUJeM158icfZUX0UJqsx9TSxKEeDuVnwc/zB8PDsb1QAXt
3dGCiRgNWFARvS6t7hoZ4UEUv60yZc0mCDGCg8S4wH3iDNbEWMisdSHxNKj2VFy/PuvysDqYJQo0
9N06EpJTKTyvUn9TOueHqjtLmzmFc5k16rxTmhNjLcyiHyQNazY7+pi9mPkvW3B9cIkpmssiZM4I
U20q46pFGassCGd9cN7/P2LjB+3wzm1UXWNI20jBQrOYF+yrYeaRpqg6Q9oB5N/2eWFz+O0bLV46
2b9aRsIfVPJ5rDKggxKLfcbXmNw1B9kSbZBsJFhvYNGOxzDhZ0S0OFhgPkAqLZkzmuZlf6R2fZVL
2FAnuq6m6Lt2yhg+4uSjZvOmj9swUypnSDhiTq9xQptN5njUGybL0qHMq3GLR03osPPOYdffzgXr
YdCYPx+BYI/0+lhl148OfvD4HtPTyskzL3N0UNdhH+0QmCCwsAYvpmOikD0dM0gWdaHezUj8Jzcf
FSCJWBIrmtYYjsUFCvcFd8xFwetyYxrEDwzRuhaZsF5hEZ7QV1e+FK+Wmo078rrWnmQC02DMAncQ
qQK62x++adT4bxe3Xp6n2eiXrs8U6SlTwZ2yqVCyATe3Lcjroi8DbIyGCWZhtAxfuud3YgYBpaDQ
GBJNYvjaI1tVgO7k3k9pnABg7MKyrpjXPJRfGXrayuGvaZ5YBS7VyN440UBRUe3Qd0ISLyCNOe5P
L7OSCiP8yHVi64h9grn8YY9ekMFVw71Ybuf7KS3KcJuKziJMN9Pr17GIJ6wQfn9AW74VImBuMFgL
GXPtBtkAsCGsK7cTtiSk+XXG1HfyDJBeneX7KkyK6vm+En4lyRgGVkOw0Egd01jACydQbKli//Q/
tSFemn1yQ7dSCzBDv9j/YP27WJ2RDPuiJ0y9XXmzuVis+S6La0/xgFsHcBf7jl5xS0ULUSxc84QK
qhEhnIZXFXuHrCYF/utXeiAF9xkvSt9o84W2i8gUX/pVjaWFWX5CHN8StXXMBHgAFys0oIVSiCo6
esQetwtkFaDZsZp2HXb530OpMV1f3Gr0p2gv+gteDlhpCic69IfhrBwrGpEHgfBa6+Jn4wPh2sm/
HH9khNekurdemViGYenz/EFB7dughH7eZWmmE6V0EOw1/4e7F1JynQ0mqTkxubsghGElB+zA/2TQ
xO+mXQ29dXJk1GghrdNX1CnZ6kr0Yz2ETOgwdR1p27kf23W+ca5QBV92nuT0YWrjWQuXzBZ3RAh3
cGJKliwBHjxI/RDOLg+XdpuiFS4F0fJJntxW41Mzr+lvI5lyJBn7XPSrNIybAkgs8RZmRtjLBc0X
CRJXXbwa2kLd6RK6+EKImmEleRE2n25SBw8vFwiCa/00f+1Vb9E1xel1boD4R1DypKeLWELuu4vZ
v9kuJVcuET77eu5caCrQD09rNntEA/L3Wf0GaNeaf62OefvGLFWmXlyLd9eqoj/BIqwXLDHKp1xQ
NAdTJknBU6X4HjzE2y3+s9SEoAExJ3DJpHSmbwJuI1MOVwV4yn26dLME2NY3e6LEhEV0tLOCGdbv
d/5cYcuttlgcMgCzRN8b9dHQjLjvBU/elB1VVuP3laCTEhCq+HN/5Nj1jRPEXkRoOAJvvfN857c1
5wEcRUY5MNFRxB8JN97x6t6IyDlo4hGMtiLiBGaUxBswbu5rZLt8EJmN3ezIuCpGtvuHKjtrfHGT
Y9TwrhSWaVUaDI4sJFJuIzUCKcJv0cg2xjEQy5KnNwHW2Eop0ksBOpX0hX8U5Q3pkJBNKDH3xyfc
lj0heGzSSR0WcTDbiIN8Krm49MfLKRahkwyBaTrVfBTI3ewvRq2KM65rr0YbjU2vw/hszo67Veja
pi7EqxiDeUNh/1m+o+c9+tDsUiVC5cpJ2wj+oxYl5BdGcikeNLjaS/pc4XJX1AU0Oag1LJo6Hbk4
Sb+0bJNTLpRFdaArXMBKHOJ8JdtbqsxD3xzBV0tQAmIO3emTyZJvf8j+Bm+9akEFdsqQBjJrPVdY
VEA0S/fQLfZri179acpxCEzMQ/PvhFjmk7/t4u7tdiJ5qlLMTdb+2LduTd/CXUgp/owtmsTxyA3+
UVCCgNNMUw9L5d0vu/8vQNG+NWGcaaWsqsZJZVDlAQXjd+dngr/E9H9vjtVJH4rbhAETJrRS03uG
IrNa7BCccT+tJS9tVyBzsFRC1he5+MBRLUAlIWoIjOdQZkqms/kMoJ9pKSv6y72WjiTSzMMwalK7
Gy9ZFrDFabCKXrovfepdRvHbJC9L0Ptz9DJ2r11kqQfXg4gQ6SYCZ5GA5IsL2gIpDP2j55fbTNvE
XHrf8Wsu8FNEOzamJaIEzEooKdOwwVpsMFNIaC1GsuBBnHDnynP7ZPC6rA88FkdUX7H89Z2P0MDk
HNdb2qtrM/6122QWAg1G+5PRKZr0jcZmRstWeh9YqWd7EBxut9VWlldDs/ZnzNrZdRntF051ABGC
+fKWKhViEPiZ6Qrzr7fTGLyJtjxYpULC81s916wu8gDLlsAOX75RYeK5185kihPU6OibG6XPbkOx
Z6vzBKGAX5mFilFX23E/Fz1ydESA3QXr3rHIvPbeyTFYNYncZkq1Ml3/03sBJEFFJy53oeY3RtRF
y851YkmMg/e+oXjOrOWjP4oDV0Yp5mriT4ixLrLXQExdgyrVZdT3H/KX9TC0Ga6jAu9fZSPjmdOx
ThRB6dWbz4DpESYXhsPKO6/SOx1wa41bD7X/v3IEykjDtM/qKs7tHqiBSI5+RDUWzjs9ZsxYsZTy
fWSNcS6m3fZgc1OSLv5poDeiuSrccmOp7f2ncX7in+wWBpydyew88QCO1UdMrR+ixGEqk9HMPkw1
C9tJeGYLm9r3Ki32i5+PBVLGMjwTSlYurZDUNzmkcTzslGWAqqFksWuUdbPWQFHvJWDBOqQch7cZ
v9ERTpRIZEeTfcby3vGNxfeVKs8BLO63wsj69aDGqPOB7ovk/6XX8vxnOVAwRfvH6v1qeD1Una9q
YBMRD6X/e94DQGQ93k8SPi47JImsg8j/Ulmf3MCdwO4jECisPlcvgBLTJaETMY+aqPtEJrMGbGRf
dAd4f+fNoWZA4hoq+JlLUuPohoriwujgYqwgRQgwk/RHlD3BfUpACW1VNE39AKzZm3MtQzAuXmgl
PaFR/3iGF4l/UsDWnfTY7Mhs1Gfj/7JpAPuL9lOg+5Rt+tMoRCzFJXc7Mj42eI/rfshNMUYtUnX4
yYkRZdUHjBiwyn64mMRUPVDTQm7E49Bo+cH6tUvRgHaLcZYgqNkJ6GXDXMZrS5hycB60YKfCHaNx
WEWLYMmSELWVs/RjSb5KHCGouhyT9HS0x/Oz1gyU8g8tEsM8Qck+qRSly+erolGuzUTs62qyGIJV
aKSyXO400yejTkjSypRPa+FGL8EOXmZ7d3hV61c3GX01Y2PR7PBW5pEPJQf3t3bMfruK0xYMtBd/
98qCCfLpJd7FIayCmk5kj2nGeODs1in4bOB0HRKyy04Fj/n3/gGFFcNxiwymLlbti1L+3OOErJmi
iDUPe1dKcxJSI/pOQx8vGL2nez3qfvxO1rlNKewPmUbTENoMnO2rl5WOGgYgmAus7Jkg7hVzvRoa
ziaLO8m33Mq44TBxXsBfLJFZRh3qAH0ekMvn3AFIrMbEHw8nWMbLHqY1bUebryWPUfwxfvLV+WR9
0xl8NEVps8Kvct+tLL15iMibyrsey+hoJ+WbbLPWHShssg6LGZiubiRDfXLXnwlyiDiHPbS5iya1
p8g9LhVbb4XCNqXuhop834QVoiIoyWW+Yn49m32qFGj+/8gI5V6TQNPE6oT5aGWCpgu0KSW2Q911
fVxsT7azv7xD7o17JBiARQzlD67JWAWkA8TkSPTDzYrewjmUJy2C6wnwVvAdln62WBxxpnpBwxum
3/lsMkO1RQ0fgubxeVQLeyXowv8eXvuRyg34vnZpcMRIae2St/GuF7BinNPpfaMbSUZQvsm3530t
ipIPfeNTP4kZ2aKZcjRIntXeRE42VDmX5tgPTiTwfNxibfbPU4P7naNnkVYPjPfCNwV7+ss8XIcX
g589xncpclxoK+zensaeyvFlFrMIGWkmKWvK4m1Aqpio9vzCWXlx+0HtLUyDFMJvSNlpk4GdJRiG
WH//Q4xiw0SZ2URoFxmVnEkd+ZcWMbiI3zxZhif2gj0vqM5e6/7bg1Q6fTkozsFI8Qrl4HFnKMEZ
6aOLXQHaUBudfSQSqkhh7cIBL0KUNCSNou69t9bBEG1WX3rBOdNP4K8ixorY3atdnD8t4ESgFVca
yBf2y2eLXUWHgCja/UYpvbvfNdLWwWLvC3xu79aO5bXF+sq/bnc3n92+HqH0rl93SgfQRqJD7uWd
TMiqPfth5HYrtQem5TtWVXO5qQFAxVXiN/tZYYK2Y1Om84eWDgCk/zct1JszaQfpnZCle5tuShK3
uy/LA6gEcwD0l31oMS1+18z7HQCZ7qBIa0hoMStbfPB/WIrxgiSbqu9rYTCC1Tiokrfpf69bTs4A
0tYyXTifQyqf6NDQGQjZGvDkHYQykaIL1fgICHnvhHW5aGftjycwtrh+RLEgUJ3cLbcyvRfLQa3/
RhdW4o85vZV28tjvji3tBIuGJhvN2jFpzvPWlTrl2yQImVouRHT19oP+w+aEjgmx0SLzLxCDl2S2
F6I0bhWKwAZyqRdNm4yFSzLJGMP6raXver26apB55US1oPq0d/YTWjGxpU/NCP2XtAij/Px/MhLU
7KPNF96t9YBDo3lQkmfK3k3oMhUGyGIszmcw+4Qk5bhdYeMiSdy8o55hXoUyTIFhfHvKN9Pc5r1D
QPSsGGWTGSOGcXK4kIa1EvkHyd3KB2evt2mToAbdSj8pbtXt4CqcNkcHALDW0pwyw8ZYfx93SlzQ
Atq7p++2mAUlTvH4WeHGmCRgUPK6Vd3KYf3QL0Gra+4ts20FCY3YhFoalOUegVJ1cl2wOFX5SPEd
IzTYNbHw3f4REZlkG7AF6Cpkjy/+e0Ju875zb7CnTdNzTnsr918FvxZLnuXyNWb9VHWiz/CFy9tA
UnD7g5scmNEXjo5IOo9abqk6b/NLbD88Vj1wqgT49RBuuY9oj727U30GbxfYr3nB8xMBCAKgrnq7
vHHwO7wdLllpTtKqPG+1UHsCJ2bV3wSXIrzQ0XaYFHhzjH1xm5lRnkwp7BoJhiuEX9apvMHF2+Ng
Id4cjrHbGI/cUV+G8lkOxaXgIF3IXZh3jW8yVM3L8jFT5LQoLxcrQyWm/rWUkKQRkbUdNn3GWMkD
TegDL1Q5wypJQT2G+Op2f1OBxCSoiZSrLV1vfNiwyxQRTczMyPNDv8zGtyJ+OKKMY1dFa5737Pks
13ltQH78qhF6RCsVUVwtt0qi2PsQ83Dvvd7cCLO4epEQuEgCtSiCroscKCtN2J19UJwss5/L2IQN
5yVM8TJEIejRX6M1G+Ni3I+3rcS4v1aOCHuB9RHlVzf7vzKDW+HjpTp9Y7mAOn9OMhICaaPH7B/6
Or29QCrzWaKOfSbWHCmoPSHuR5cgEXf0lFDQVJ+UwLoW1CoZ7nX7GI/RvKdoxMwDJL4zXPLiqNL3
TF7GBg1IpEfIA09Sy5wdW3unO0hBg9icrbABkMVQDv828W3JQqAuBD8QcKCdk94P5/zUHSDUo1+b
W+c+7ReibIYvi5DOdC7DsrOlojcaTtxAeDwp1NlMWONkmNqqE0yzvgon4Q6gZbbIm4zFTuZeKG1g
Iq2JfxS0MfdqqryFspFSoSck6CsqhxDnSslKSBi+D5XqeWTC5pOeuPONKMlC2sGPe/a7LnxhlWKv
uWR2DTsUriuDLpeCMbW3s2TjXXoOTRSqJ7GG2aEjEfrX7rIExHLaul9791otx1XWvi31dEgomlcf
HsotwEHsKINohczIfw+nbuVmMPOnO4Vaq8VHKrmIArt6kpdBS07vYdxyqRdGz+x1QJDLg3evYwHf
CpcArCqVGo5UXgi4EGuwy1cOkWhagFo8CLMxpoxGf6WblUVKUwwdN/29iMHvgjp7AAhDpDEYkuHq
Bg1yYDnI2Fmai4cGLLEpaL3aIj7tmAsBZeZtTiMk8UOLWUd+EPsIpUEUcs5PwJ4WyNdGMKIelJ/O
SVMxonEmX+y60B/jEKgJnSHokX84VQwHqNDUkSclOLzeNxP+iIhGBAS29O/oEJp7QPynRzyK9Bfl
ge2oxooYCX4Y7FdQ2gTIDtQ4SUz6JaEr3ghdD0DbogtNEYaYppb4gfULvXawPZVRaRAEsn/dQlsr
hgmSSSPDFxhGUePwb1sXDF+nE7VTk4xb0JhcqiBN8FSRPwTymnFjEq5g2/3Y4AQRRTCKJ/jP+WJy
SIsFmUqpoiz3m1MCIS+13/xvQ+9nA9TInhxbnlyhN1GKt7njRA3QT1MR8D7PCwS/6BS7k90kgQhb
9SHqyNIlSdw6rmI9uutWJtSw2JcloWdvp81DZbl52czWMEoQvYcBwJGska4vIgkpcDrO/lDt5UdO
ccEvzHRsmOTkATJ80jzUBzLzndzn05bcT3/7jAAsnEhZm+XPZxGY08drvRpVh/dKC+e9is/NBoAb
du23hEEf5IAVNfE26Kx6Jn4KPOa3WmqJkhRum3Q+OvPFUeC8p+XJ8M3r3/nkyQoi5NQQwKzWs++I
MH6d1A2MEMI5P7osyafTXJVJ+0MUSoyy73MJof+fF1N6mpVoIakfOqWy7mjwu9Uuz5cdbTQo0IKB
+auzxaxszHjSs935VKBEjZaSHRwDh5DYjqdQThO26hsBtTbhzERcPoxPHAPKcPKxV1lgUUGDvgsP
Cz98JkNV89SL6JUv3iWKWPd2YfX+7477fsBJ8dWGQFXhccI0jSbBjFs4z7o1Lty5lzV+RT3yzk2T
ltBvERDQdidrTs1SLHPmsCrBBAFOxt5o1EbZiVRx39qTXGz8ehoYdQWt1PorEy+d9wNqZLoipCAX
o90xqtN5lDCTgIzH9EBme4aWo7bfIBkhqBfH/zdZfPn5M1tsl7Y6F+19LhaBZxyK+kFAa09FT2Yr
Rwfc78EBO5rtbxGWpFEF3uLT5TZ03r/U1OZQA3U7tz/vfKsHPtxp1ktnFEZOp68Hi0U17PNeEuoj
9IieFRIxLSULnpTT+Lx78WKTSMaVDjjRL2loSr0hQW8xFl5BmIS9psKMEPRZE8L1PywTbu49Pfcr
QZz7ydN1SIiQw875tU+piST2bMTZfHPMMGc5eH13PhmPfklxQW3VFVa55fvTqI+UXQR2CAGUyuT3
IEmK6JEd1Q4LfKgeRsRSwI4p0EIQw3zYBDv2HCRcrOz2BLCVQLJU4dVGzTNpThyS8WQQ882DUG7h
blQ/z8CJnb5nJ7ZApqZripUtezagfs6o1COyQyQk0M/07wPgJuBNtfTH6wV/1STlsK4b0rzGwGzj
VvxWIh4yyzYgjBCNUJYN7IsSQ6NTnKRyBfGn+4IgraVX8d0t5faUUnHKXDtp9xjJLilyYvgq5tcQ
S9ayHj27L3QIhBnvQLE7rRiZE3Duf8ZkcB/n+vvlQUO6OKzOQuppq+wFuWTV0J/dYDmUhAMWM87v
xclfppm15nW9gkU2crgK346tZDOkRNB1xGKaR0fJJRU7at7TGZU+8UxntGDZxldGTPn43fhqgwaE
tbSO28K8HJ+bsi8J5E6ilFWmx+9Rw0/cdhr5qdq0CFA6mxDViKgH1nLzXRKOYTRB/d79CuXybm8G
OJ1UwVvrCaV+qKgpJOXQBNei4HQd1oaZ19qqaMMKA7Bn3Q1Mw7+r9N5TUmJJmsbWAeNF/3hQU26Q
c0ApOHddsfyrzY1O1ItH8DdDEEQdA/5rRZYChdlHGDE7bssVGMVYw/4Q8qe1IBc4xZ/me93rqlJ1
AQ0f44hlHwSLM28NZO1+cLhs+2D/6IaWdstZ5Ro7OSn96MpBayTW1x85XJ3iraqESkvA61Ymr765
7y5PPSF353MGKmBFfJMZDkjoMyl+n1C5UgSbnkvMZBuhM+C6pYUyGsfbpCByB1AkVnw9avp7CD6P
HrY3n0g2Z2UJI390XVeJ+hmx0Vt51l792TxmM5nhed7yBjIx0+TBWEpRn+B2Ky1y+ylOlf/pr3fs
R68uPMWsS+SPwJU4Id9fDuHtoiCSIxZj1TTiigAYwBWnf9LMvFtiz9cXHpOzAhms568kbDcK9bea
45BY7lFrKI2qJ4R15sqDaOV+FKAEE8zEUnPD0evemT2KNE8rya/dslHszjCNgtfRLEmNWfF7bR0D
wVAzHFIbLrQ01RuqfuBCz0QmE2vz+Sk5PKWJc3uqQ63WC2EfFmcTIt6BDx5mktogl2czI/jSe0BH
BmssTBIgsAskDmCldWz0hr4NgCovDoPdpEwS9VIzBSQ8M3uYnnKh4pKFHVicU2eehOdWO+GFxOBI
0hLoJ/0eqaw5vyytH/Dzrnd5qE5b8r7/U+TJyo4Kgbe2I46bpah6QXp7hX7LIlJIr8ihzGSyQt28
FzINzWo1DtlGMt1uxM0jr2t8+CwHR0zAoGVdrozGAjJTKhfX1+kYxqr82j8JPpe2yMyB8vuqqCzn
7ChNcto59SfDb3x67oaFGw6vSXC43QC2ZJhZffXmhOtHFnBV1COpTHT1cjJFsLmGKFt/SMzKQr2g
GegxUcBChPlsBc5T064I4ulNQBmjCUr7lycAfVt9Wl+WMgcJa2AiUZXBhy+Z20khwEzKibqUPjoQ
+1LVZR0prbhnqlT7seTdFrigGa47cLp+hOquhk3hPqC0/6WsXB0CkGcf16RIPc8LAkwvDqBX1IsE
RmHY+xyIWcgxID4AAp7T5fQ/zJlRxkdXPzhHS2F8O0MsluTt002AWgNtlk1QHuxNV0LTvGUbr0Ac
8Qgx/mHsbsAzk7bMC1WC78EqljwMijaDDaJj5O2ULIm5FD1ved9h30hjYjQrOfXyrdtsn3RMd99V
dsq+UFzPFakJ/qJOBs2veJ00gju6+gq0M4AhzothO6BRY1KPUB1rxcPgjzR8v3aztMUffED6fmJs
1cyUC+AbPZXAoAGGqNZBmLZHpNTR8PtfooJwnWzhKd4Xc9Nwky6jiaMwjX5vDWVq0RxyUfMMjYlb
ngLLttuTMvGT5MhfL8muhVsNwlBEqjCEmtBQTIG9royEj3TIsf1viCD4HFTbTT18yMPR8qag4Vn6
r17eSeVWIFtT9SELOwD81q7hCLo+nju/AP04GhMtTAk/RHJ6hnF+XJkqKKJ7DtMAsdzZkBB3Ba5f
AzcJxblcfZhKaQHenp3kyiHiRWhXn8r8SveLZqqhO30JLDr4GHIXzvSbiVIJo4TF7S35LNp2LT+M
sO6ZyGG302GVXOaMVfsATYH7GylF5u1ah1476j+Fm6l58UnSoLmuXFowGM1IQcHjn/djZ/WxCQCB
+13A2dvFLYtotCrZEjToC0OJCvjFfdaSlWwg7aWoG8ekmKP9wW8ycGqkP6YF9vZ9YTplS4NQEhzP
oDEequCp8n/AXaLk43/2QSYBIi+UJu77m1QXBgMPFKDj9qVtQAnLOjhehH566G+c9xOULEGaQcYT
fc17e1fYjUmnHtrzNk/MzB7x0o1SwBeauowPlu/6tSkf6KvlNb9ug/TmKa4alyJMfVn0nbjpgxzZ
OiIh7PtiNWs9xqSPHUbWoHlUy0Qqut75+mR4BDn3H3iye1X8ktAa3u16GlQiZqTvPuuvWpOywPHO
A+C7TUXO3IU1YmSOT7R/vb0Tvka7b9TDGT4h4+hxqvSmk0XvHzKIYjx9MxVgaP3CzDFljxWgMOqT
n44gwQRUQjYAK15nJNDbr+giUgkmLTTmBumsh6LRkfQYFgbcnmvsVf58GisqFr5mw7w0Vr87Ibvd
WOgHmkHzpNzxzf/sFR1JyxOWONCP00J2yJhqk5v3HqfJbrPP7XfzrTguu8zqeGvs1iB/5wiSYyEI
LAOxeCBcm4BXlmTfZ/AbnUfRvT23tElmsMOlNuGjhhSAXgdpuFcfOaa8eKKX3uxpSdEPvXIshWoH
ziJ9TtFjdQbTjqhBuVQK0WzrZOaVc4glN70GWe0i469048f7e86zrwfdMlFvdfApMls8XOvT19lT
snKrgQiqJvZLvMCJDctqEk62rEHJKjrG+Anl1sL8ukkMS0cc/R/uAXMziiFWxdVfcyR2V4ZexLBE
1kmVn30sbXvgUaQg5+gljDNrU81ZRQIWUe2C7+W72AcL+/DUc0mM2Bh/xSX6t4UUzxoAOY+08kzv
NIB+JrwXnF89E1EFOOJsu0T+mhmnmEWsGgysmnwXMHzPRaD5J9nM4lAMEgI41qVZFu6ttgpu9HNR
JA2bJ1B0AuldVlYg6htOv1pbNawVw4sTwFfFuQIpH/cAENx85gMyG+beYkM+r4GoqdDFqmkBh4Hs
Whdb1/K5E7vkHiqq798rlmY55kxNWeMa48Z7w47IK/hVx7qCiCRBYO/NCAozjoKCf25TKKCjxlAg
ZrwQGKHenOGztts2d71JsiaghhJnn4yHgD9ycOLPdrmkZfsHXiyh+VIy8Mr82HdF9gcv01tMGiLl
RArr6cVxaErpBoy6Xs8einDdRtDbcQXlR+oMvpy3T0teM0QQSJ6ULvbRo6JH45pw0l5zWMn5hRi0
c/2qUo/3bVCEGrzYIn2wd2yOdtB01HQdlZF71NxgMDPEVw7LH5g5vy8j/4A66MrMSGA0btI82rHc
zPATZxtNB9h5E2X4BjFcDb/Tf+0tBDedcp/TtalU7bhC9mbErftNSd23FBk29iXw8ROKNYVi87NH
7swO9Felk19LcNIClHTTKNIDg8USh+rR0YUngqNdJj8jSW+ph2HW4AlyWWrs/DMvvJ8VNOj+SbK0
aQTgilMhPxCSgkAfti30UfzTMZBknPo/UeiQh6zvSQFynCD92UZ+n8QRZluAmPOOEW8amQ93inEf
6umj9FYzpBTGkvawUkgxai68+DedDe5Z+RKPsP3NbVdKN9FD2e71HpScBLLdBvP64RrNQRcLg91s
TVZITcmMJji7SI88Q9MagWevFN2u6Oo+PkPOufl5wWvIgMQeB5w/eJ2SHlnO31PZn6CTjSQY491j
gUIFUg/gVZ10TV4WGib2Pn8AcSfvfDecu1+zYXRhUkFeYg0F6xIRUF80U/NJy11q5UMfySaaFJQz
XgUTwLx5zppFTnfg+noCn6zJSCteBKcHNGjRT6mJQjey05Q/97vmqNelykvwAyMXq536eYPG0EgT
r3ma/wUdTJ8HiQQRzF6F/9DZ0Mr4rMmj3tSOS0R4kalpBH1Mf98JpB3pSdokPj6y7fLaBwrWdQDR
RF64tITW7cGaUoizfGcQ4NAWNCYA/QFpF9ZzAd6zjigxHRrpetV98BW5sTYIS5FuBryk24Zd33DY
PM/IdkDf2ngWzKmJiKTwT3wfvYLDDUxxTPSlq4Sfe8jiP0qkL/AaNxicq/bKqFK7Qi5Me9KBZ4zP
2Dhu3hxNGZpkjx2xgZ87yOJ3eUQy5FsLOjFPtyP4WmKe+Z9MCTMsIwDz5IzgSN8TKeNbQE/EBQJI
+gut5cxw8SPBUGGAZ73Rs8htluv7EcAOrng/HJDhTEiJYNnQPPxOxOG16GVu2bbxfQBtI6V4sqey
utbeRrzwaDX1B+brAL0e5MbXoEWsOdr1Xqml+BweovrGxi9V9gKHXM6OBPYQEqVKsYztS3utfzyO
YynMkzlKVoCB4l+YhvljCAalEMK98k+PXIp99gKWguhGIOCJ0fmdKHKLTWZsf93/EitA7rkOsnX4
HkbfoLGjSndePYvMNYjGAGG8Z3NT5yN0A2HJ+64gUh2iyxJewpaBFL+zDEc8GM+U8muu/NaCqga9
5V7/IxEc1u0+YKb3Ruzr8qvVc8MqQtJRgMrL3lXZpzF7flwJOcI4Cqo49Hr9q+LjFA9MeLDXAbXN
M8RZRLylrEsPX5xtNtkkoQYVehBv3juI/LulXQrzbV/jTmAFU0cogrj5pHceORviQ8N9Wv1bjubB
LRRFwDR9LDsG7fIH1Xa8WvBHeZM8FXGIwOcWzrzttf/qnpkkDgG7geAtaet2pmjodwyrJ8GTdaHD
N2A9FAT7dQVPXSrcTy3WEVqo/CltTjUUNv3IVnPRP2+ItCrMv96y0qe4Smnmc/7y0wSgyBMv10GD
niHdqO+uNWB/dovbprIcLAEBoYCJKUIR0bz5XFRKCEwnOzoz4/H11iQYRAOYKFkso4mCcZYyTCfc
90EjVR9id25Qs2ablORPe/hRm4dzTCnCwRmBX2PxvbG1UKthTVOO4DCBPlcUvcndHsKTXAmahFYf
JxGKdhkIKtkkN9nqqy9cUfX2esld54Mk0fg/zuh3PCoBR0DzszmwCAAwmdICDjCfVKpKu9LJzfGe
QtOkLCyfAjodHCQOhqgP7/lMtuf25/1WGunk2SLG6lcgFg5jYRSNKrz2CDJSlc2ncMDBjb4R9nDc
n03mppSwA/lv45eiW9CVqyIY3A3dFE6SW1Pa2aty1+9kMGECZ5GgZ3VrX1agcsqCRK5Rh9daYC08
PhfZIQCZnGTqJf2/CFv0h9ndAhB5z9xnqxsD277YshL0qEjQ18O+RMW78HxfUENEofhWo42G30xK
FE94tyLZHTQwnPQzKciqqfIuEFHqM8Lxf+gzbJeHhIgZvtQ+qD9oJ3x8wx1g8qYW2KIukrwFQUgi
5LninQdLfnFeKvpWjv/eO7z1eoR/py3k+2tbnYuuYvkqhcS3wbzGZCnls/BNvKwxX6lcydZ7nWba
ZqRiIF0uDaKZ9773g7WJ+VwqoJGaUgKLodYWsLbnMxkIagFfJ3DwVSRCJFoL8HE3lQ55FTGuwO5i
jyGIp0+iN0ZNkKzyPWJc3PFQ4HQ45MHGwS29uh5N3GaV8Ruvn9r39ElKGVYzp/RkYIKzX0iLP8k4
VcdVtNvfokm609TP4busZ/NUtSrBvxnI2ySzgP6QUChXvXp8XeIbxq2xGfZ3UF3gF8tTsMHZMHvr
vvIDBiS6zo84nnaRbnVxmq9x5EvXjQmtuLBL7a52rgYH4n6zsRCa16D8G6eUGUjTFXFfMCHT4hUq
LLHBc3a4X1G/XW+21fH+B4hR+yA6WsIFq1FfqDL5kkW7BvVL9fFN52NEeTpRXSZooKra8EqcilAs
o483tvYV30fhoaOqPs/JQ9NKRdxp3Qg07YylEVQ5+dK360zRyqaoFJlfTU/vkZkeEzfPUGo9zlPz
g2MWMkVQ5mej/tyXRJ+lIWxbdPkXyMX54xZ+dFjpNDz3m4PdkNsCeEJTDyZzxq6yAintY92EDUxA
6ug2eVQh14umkmdEsXWWRGe+XC+A8xQDXV4vQGZ0uhlMFbSP7ommci1uqYTD8a1EYTZuMvB6ulRk
VTuOFCCT5Zrk8qTnj1BNIewGMZyn+52XfIe4BOKyX7AMzvpjVYI/Cmh7fXEAQXOqL5dTNkONkny3
QdANLdRUvdHPJ5qAQ5sasD5jJ9xs/ZEShTieKlNa69/QYdDHiz/N2ZJZyO7QNDz9W3pAh6ykEPAx
aPqEJnHTRf5710fqDbNmngshQUp0epMsZQQIexNO0ZZ8xiEvxzE7k3ydxAQK903eUEt99dcG6SPQ
Qm2ISavwD6y10/X1HuUvHSYltvgp9xIJKJ1S2nNmIYPopaVPI7Hmc8IRUwvWHOoj+p6RVCrEsJSc
WU90SeM4UtW/eQePOM1zkDkq3sNj4eGKNyAeJPYU/WtbyYXYMQ3+EkdTA8Pz+A+JXoLp1Fht45t6
+CZdX16hQUethDY8Nb5rS4LjC1fpWxZwp7qftMPtRUePnJKVBrf1Cb/+INFYcf7pLm2Cqhgfr+0s
58+gEXo1OiLE/Y7t5sXR7Tcu5HIQGxVjuA62Q33yz+hD3Ufq1W32WxOzlQ6cyIqEd3fT3FMc8kYg
RABjwMhCePejoVYPp2uz6vME1/dngSORgGKvjTAQjEAbJ8/i0deN8qINE9Pi2c/rOXc80tijm8QP
dXp8ULF4vYWB47dHWoFoUSbRUKPI6NATvcfQb/k25+kUH22a+ZOi3IfSWUlkMJ6WkPOFAeRtVBQv
c4MUnGNxWUS5W9O+YapEaBp0Mwy7iTLlB/qj+FbfCfJcR0LBqi98D9IuXUZiZFSOeBZm9z/uyzEH
nB+MgFXZcKDxMb2vVWTo2PWCMlFpc9OriBU/GBEeu/Ls9nd7o1COGEwwMpW+f11E8KyYnioRZs3U
gjV1yMl5sQXJTklOAx//aLrYd07XTH7XO3lNobRJgIMKNrKiUiNcN8Xd6YwHJNqoUuaqX0q9i1gZ
daobo6Hk2z0K83XRi1KsoVA8pa0VznZI+62Un2vL+xrbEDOWTXPg3d+40cScYMsVEyqy2n3tlAxR
FQu7J8bQ0BzGK2ArcEmI0MdiGPzA1LukY8LxB6QhnKb7YRoIkrhrEjZjQyrAYqYcNGGhcDMMA/9E
KLrBOW1mvS4wDobdp4qSMIVIXHpmtMuPd4Os+Ia6aVkInICgvjtLhwm0skkdhIL1+tRQbWISyjal
TI8kPzYUBBViRMySFI7UYEgv5UdOL+fDANBvivGdjEZ1NQ5WLDrYfaRxPV+lM/1fPdGstjLnaAQK
gisdrhzwj5tUttqQyaU9YeWzN+ScYWsi1t3AMhBqxov/vicg960Zmbk2a7+wdJRlBW+f3VBV8mMt
dRuBf6xGKx9n7MgcJ2ZwruoJBBDkvxCNO/+7f/P+8mTwjD1VXW3WjemkArHtaNd5/4OSvkstPMDR
pN+VggxCi6KrYZjSCiIqGeaQGEi9hQfTSR6aKdKJxadZMp43cUdMZWW2xOhe3WUoiezZZMNe4VN8
L5zJIgVqEw1owgKEkZefU13yVPzfXHMTXfFrKoJ5iVL3+QnhzZTBH5n8URIXRtXCiE3VwqhiOzav
eflQUMsN16zO5PgUsV0B5M3ouyrBzQC/L3s4HOU62m1g71Y+JmKkcqk5qnJdH4VK72cj733uoCd4
7/YPDfDs8Gc3zd69ZFlBUrlcTQUzS9/J8TmqLSgKkGmmxB6M/6rVmwmwNWZoWUXtuCmU4ek4HxgF
kChwwORqFijFWPQK6C0iJnA2O14pre5SKPBCjrWs/fzK5sOyU2RRpwNbJu25nz8HCz6X9+DoLved
T9TWL2CMbXtrkUIxbo783r1JIfYGmhsSP25wfvGgPKe/PSoMI48I67YjkZWvf+R+MtHGqAxNGJ/i
zF1GZuwjuSuwA5kUyuCn7ViPFLS0BY68evZo6b+bfBDUz0kbkf5PbVslAx6jwRvGDjkfrdwLAG7G
I4NgXh5nyRlPwiGGuPpD1HpUNM4QuV+ag2cDjOo1/UhY0g8Qw65pquKvVGlA7tfgIJZczgtyJRw1
ADU5WzgX2GD/kNfXbgJ41RwdB1uxgB1icgyIx0eV13LE1flMdPAl/n/MZfONyeVSpX3Qv89CUK4R
fD0kOLXCl5/NUGfBfkW44RM5G3+FxeEiXvTW8G43IaN81eLoxEk7tfchpCIPcGz2DfoXHEgBnKNc
f6domEI3m2Aczvg+zF7D6lVEib7gcUrAiwytMkbUGDGqBWdXYBretWzEcc8t/3tu2P2Iv0dfaS7v
8Br06xdBulXYc1htR2JPhrMB8ox0GQuejikU711ev5/mf6HqyCnIKn5bbSlUPwMhCY90p28ssBrV
w50RVMQxXyD+nD6Qy5VrtFgv8iUgLxnjEe8MTZWW62nKhPiro2EkexjDhHgukIGXzKHSaz5lZw0q
Iu1zkBXfSsR0mWJjvhP7VkguBf70rmg0JmjpcuYz4b2Q7bfba5N336DQ1qUcg/BDkXOaXrViE/YN
fnen67A6jGn9Sz9jobF+gnR5zg/4ooXqd84FehyZ3jN1hnwrVs4wtHhGA6FTbD5Ao8FqGREtNdHS
A2IrAZbYTMFy/Ojl7Q6KTtzGgRjWz8KnBbp3apr8hTKtwdNQFo0/TmeCXOJvNLaCrk7afexiFKAQ
1cYziPqAK/opu+/TrdQiDgw7eci50gdeXZdUMkmbnd8sZX9zxugVanwJzWrjPR3QFWKDOxeyn9j7
QgTA4uFd6ATBB2Xahs1vmXGEEBcFWeNA6iRAAjaHa68GD47HUc67grGGV0/w8d6CQuFOSFAr+g44
p5mZBi4MKF5MNJA5lmP0vLXvjIrbrN4H4nhJoJvDBK+t24oPxKTqFTFaa1ThMypY96KuEqqHIHQ1
kN9UNzKR9h+BYqee2DrBP3AcAtP0PEPaP7jAFD7lzgMiWtJDFuTOMZ4j+4qI1CR4st/0/VMkwDNQ
vPhz4IM6+HheyPTadSDag1IUtPAmxv9ZXvql6sUD1qMguaSRj0uJmtOjUw0cOgWlEFhf+14xLm3S
5OeHS5YFP3r2nF0KjRh/tISrllEYqh8Q+LcM2jBoG494+sFeEUZIiiNXMinsBM2oXP/rQpwE/pKu
Z/+jVsOqICwHAVucdQ7iuv7R7/1nLr4FDl6198cu5bp6HnPif0aaB3+DWGEcGphVWoMWpB77yux6
ri6ShvzDDMRnRsRsm0SPUgb+ye7hYi4119TgwaNnXkXnDubsfQHDo1+1C0wXOUXE9lA1E+PFw25r
3eQ1UcaqYA2QC/p1slqU6nf5jy6U+nOlzrKxY8Pb+oYlpRIvIjTBJPHzHBEuI1eeRMETm7QTzV6n
IphC7LF2hcqJQaIL6dG1TvHfYPwtlAfO5kc3nzsbXNbZiAKTVNYBqcB7pE0PhDXx8LoZJQgceoBd
r6Q50lKCX5Pktiu7xtTMsItnnnvjwNcokEwgTNw6wSwWKeYIrRkzuccGLJyD9BYcZT1wC6yhRN7X
Ppi//jRE4PBvb8Xp5vay4idZygqOEpOAYHCuzUsMHqGcG0xeqxTHpRXvQkb5lURPG19lAH3icF0l
6og4EX6kxDbeWZvXq5aEKV/+u5RpQyjNydYdqgDa/ONb5wSX+55RyVzMRTfWow6L97EdKufg6JsR
ht/VG85UcvtRwUowxeabw0UPM06IufGdPE8CfVnV7vmjqgNIYyKhCjw159kX5YSi7DpEFZ/dPEUm
vejoJyiHAp1mIkw99yK4+CXohT9ZaZVSv2WWxhRHVlfRhbE6dY7KyzPjk7vuJTmOZq2uLHs5XSCh
TG4KNEcPkD9KwM0xeXSzxCA8E5BT8pdMbaluHg8PZ4Z1pFkpToSyzg4Y2DvFSkHj3JMDEG3KCWZU
3/EX19gl5yyPq/LBIIiITXUJUdk6GSQFjq3JHO5wfWV1uy2i2MlajG5dI+bHAvOsBq6+SuNw+Beq
gsD7lBYn69cJy6yv3+y4eJO0sJASc52vJSr1XMmKg0zZfpC+aYh82TljR4luQ8EqSbuoi2RlF7/L
rwFPZgZMiYNT9IaYtBO1V/qV9ACDoC74wCPFA1YGGc7AzQlVn6dHBckGz2pwpfxa0ilvkSFkBd/W
VjqKkrXjcb6f6hLp2GwimxJrWoE2ylzk2LtbGT69pe/XbWT+TSl7DKmbHiYeAzJAZtyKIIthzLPB
bdpghl3WyV9+P8LM92/u+GuTWceb8BWMlPZs6qtPRmHnlfnhwxszxAeReDBpzp7DDWknn+UHHS1y
AUSk763DRQjlU9o/K+KoL5Aqu4vR25zV0rdYUl5FcFTZtMq5SUFc79pXWnwCRttwBw9x8UOrqYpB
VIvlsfF1DBy0o22pbRR329K+E47+nzmSJQeCSbLeBChGnlEcUl60R/yt1PR3jYefSk5k2aScRs9p
7i5OyYJLx10rMleD+EIwfsDjxXQEX/J6YoJpyJu6Nny/Z7tc8ob/1+sNmadEsjHTYQelILcw9Cfp
35r6JtF+rACiWsUexbBWLy3Ecdd9fdDfTDPlQ9mM9qgJm0wE5XrB1bnd7152pD1L+SZeFrwgCB9J
JD2T4kiNVuwaM0UF+931BQPoPL17nYYrxSXrVn7tkCHylT7UadRhkYljBqNeaooWyYAbhxXCknkI
prhxqcwNKeMx9LrLzfseynajhjFDVXUd1sshPYZsotRSoxr1JtcMpDWZ6Mcvs4pczZb9Mheuu+0S
JLdtKCMSMAunbbMMWNFGyXSc22+pQVsMg4P87nzx1CxPDCbmFzLyfIllqCDpmjRhEcxe5pGBKRGE
zOtpHp4xZdQdCNJApwohAbrcdt5UNdeFZyypJ75BGDiD8ZqMoWxglfpXpKeDj1VXkTkDvlTRPfXS
d2dUYFYhV4DulGJwxWpZT+Eb1BX5aVDZRLTrtUv8sHHm7+I1x9ad4gQEIqBI0Hz9eB8BpPJKJtVc
dfMaNi5JH9IfvGwx00unIukAJ8iGfg6EUIpAPfXMYlOoJPJwUftO5NEWJZb9uUo1KLuJcTAtkXWI
sLX/ivxDlVOp3CwOnx8ziFIdSE1BbxyAgiaEAWhYN72xPqZQRDMrjINzdozaxu/6TKJ2MgduRx0P
2QqASs1VhxMFnU2V6u5HoXyZQN8NgYC2W8GeZ/ExzOghpdt7jORpgn5Dw0sGLhyBkQ0YnYjDA7Ai
BOStsg4q1TrBQlSbcgeJfIBBtUAW4MIdfAYqHlCQgGoXWSpKD/WDV2E1Wm7KNI7ckBEaTMKAzaSv
k1CbfOaNXrtMgrdhedfOP3S4WCVK/D6WXiwevceJelmGgDzul56Er3NXDMIG4PFBbC7CmIIR1OvB
JZMm+n59sPZvKv6dDl0ZhzjZrLSJNGX5vM3e1AU8j8UVvvseZcEx4+PFXha1mdaCQKsVcMPF1mus
VlIafM8IWZATwc8Iorb7nBtEJfFu7B88UvrJUOUDHJPNciIuVvdg9ojPVEQw4IzR40oA/g6GVKVy
kMoLua9XLPAQjDjcm4hy1pyU+xa5uyJWymEHeQ+0WMTSoi8ikFz01IC5bFejjLThBUPJF2I174UG
ZL4AEtXJuURgBUsRkHTki/4kaQmnGDC8XB0rCg4f0PcT2qDcQe8Ud0CMBExmvT3NMfYqtwMTzOF6
CeOrJ8vB7ZJgp4Dh8YQL9odWGZv0KVENkQHcJ7gTNPcgRzNNB5g1UIMnCa5Cf43nEYEBgaqSK9HJ
BZg77eAaKzwwvzKPZ9I1zvEg4moCx25hqdA3VKkOaD+bzLAHsfqH0dEgWNmpqzGDcmL8KUu3sA+c
etnv3PwG3Exoq49FORvbvo6h1mucuXOot743jIM/EeVmMgit8qsLf4+7RmTtO6ygv2dr4xHruLpe
uQXzJRTPc1nj6vZzyh0bk+OAMiA2FbpycRH/cXmeX6t49UdxJIR+2nS3DUAq1mx1DoKUg5I5ST42
61ZZe9i/65oND328vz/FEViSAKEF0cdGVISxPRISklWT7+ApSw68OS6sbstgzcBSHfLDxq3ntFsy
b57wrEosYpQ45Emd7f6sy2ZdcPOYpXjZG5nTEq0lF6XiHfP6LJ2GYkcazcUv2ugiJXEhGrAPUJ0t
gep5v12m272robmpiLP/YkgKemA7Fccv11jjaHE3BNl69JzRD31/acSvUPbWHTdfb2cMViypfP4I
rSVZESY18hj/axpa2Jw2XYEcCvTmEpDVlNpil9lwTv1KZpe/GkMfYSNc1cDmm0dZnG3ReO1tcf5o
zFFehg3I15J9uU05opuKep7MPyF/+DbDnisRtWPoVoZRGvKFStOVrfIImj8NglBSsfKy4RMikkFk
ehPvBmC1Kwer4XeJdsos6TIH2uDREhZ08apNjjGNwReJqrGAUBr36t/OExrKVTs/bjQfYkBc2kHo
KgMilMKtO3cEDVPwofnY6RQ/blA8Z+fRQuO+NRHMIPu9EFGsRT3kVGEeew5dWp28euhl7We8eiNI
8/RShDE65u4xl/4TRjDfQtZ2DFAZFBaBUSkYAeiqpacYHlKf/fPIR7zKs2OQpz3f72nV4//Pz5qC
IRHxgWOKqgOi+oJtqNwIecXVD1B1X7UbBTNwx3NGzE5zaTYF1lDwPgSqBvAt8v77K3RBxpfzdxuQ
qOPPziPDUvIXG7V+B1iZGBeyMFUp887km11qBjmefYUlqhyl8rOFfMQksFKW8CX8BLw55gD2wwpA
Cx9NakH9DDl2C7u9Fc907lTgUtVfkmBiM3stFjCAs7Wx7cI9xHFYeKKp0AP0CpxdS1r6/F/gv+Rf
ngTCpdGaiGhU/rmjKWJrtIGL5GNjQ4b+mXmsuA2m0RXP5sDRU15u4jHTxJgo2Fvvl0zKmv2dbUNK
bDk0BR6KovJWfPTGJCmmdjpM5+Ld0vMAGJmOOba9yQ3s3AcGv5aqpSX6aMtJ/+GsCPXnTHIyTgTG
GgzCT1JwwOqlLOCP8fOfqXgVc6WRzLiZIrmkIYuhWYKDvmcoCR4RrxB+IgMecFiSr/leePtZDMgH
CbHmpKeYx5Zo+wFdyUHHeB742oUSBZOgVoJhT2fMcSd8jzYN2SMgTCLZ2gqtt45TzXjWQt8AriYF
HIeTXoGwqd4VM69199ydKEqiE8m7h0UI1DLXRnBx3NFrNmswyrUppniZ7GHTiaBBrLWS2aprKuKY
+A58R6zDUubrn/utyn2fkNJoNeO8YKyztBEIcaZKaYBghQbQBvZoLtpIqoSDBooKE1gIhVoi9DMI
usYfaABM5JOuuk9rRb1OMN/8gfohcFzIsd83vlkrMzDXVExJga0l0l7+dob5jCYwn1+Loz2T6Wul
QfDxGJZ/Iq0wMRWLNLVEOEFw4Eh6ZUs4tMkSjLcgqzJLLi/Vsvbdh0jNITPCOH2+cel/sffmnoog
1PFXKzyf1MuOdLwfpEG1iWfjWAa0emlMntsgx56UPy+enXdaFKazJgUqAOecE/iNAWIGY3gU3sex
WourlHKdEczk2cvZI3eD/snbHEkN6slWMJIiAft5v3YHY3qMLQYppMWVMx/Ia7uFQBCGoZUJR3H4
hMpCG4trcCL0n9R5S0wUwHr/Sm/17y7WOwnDHtgL9d2fHn9P5iIDZTXFlRakAt5pldqexmmuIOMR
gcXcfVwr04W2bd1dDCtK+aRp2mvlEwAbYo9t0JS0zKY4sbW5539BG2CCfsCSXwi5Q8EKXUOnsLfv
D8WxcyfFMWyou3ZB8EY16kplsl+wW5wdLPAyFZVtnAHhtBdyaZdxchzbhnLBngMbHGZhdofAcA7J
Mh9i9Nv8HtdnfKHVDPJGAc5Rn4db0TJ7L4uhw3FzXhpQNrzSEi436VYyUo8em0za8nzuo7KQHCI0
cSdq9Sd42m5eiMMacjo5p/PNWGtjom32F73m5lUSbUNzp9ExS6shmutz7/amjtZExPF0OphiPeNO
eMhRMLcridzH/Tf/yEqZMiIbfbwlBK4JldY9VfF9m1OFy0NQFK6+JAe14bBa6/OlT+mEW5mTvppI
HJqox9h95l3Qz3eaff3XWPHRzJHsnaIf/xtSHeaxPJvm5GG1pd+yVOA5QTc0Q97DK41bvbEDmam/
v8r7Bzvq7erFz+sjB8QJhG0L5G8WKA4MBGkZEuzHmcxq4lxBqQgy/fhtPexfq7EZwbMZAGkczgqx
eWL1MiPz2pdLUwVaklOVBGTOvLP2b37DbU7Y5psqeSkyP/VrTqNySPpYhle9XSxsiNfI0ocjyF4H
BS/BKTbZ+FIP3Lo2nrRreYGLR90hm/KAHtvcpfg1BH+8dWEH9gkJsEcvVhaHRW8e0jzIezxgMi0A
eaLUsHaRBwqo/MIq7W8TwPsZBcNNbDM4TOvly1NY33U4PJbusGCVHpCagGCMeCJhBVzucnBoN5vz
VSB8UbmhIVkw38QHmm23M4xVMJ0fOUDs9sv2aXVxLUq0dn6zXR0fIgZVhnUeTtFFyneaH+bmav9Q
Zs7RRyWnKD+RPlpIfhMIzEtLxsmnJNdj6W2MJ+m1Um+cb9Ha+FexDzWS2uwuBtkMFl7+BbCfoyVu
nD2QqcFMXSOcARFEvIqXLLJyQKUphjwyN/UVaa7E4TjWDrivZ0uJkQF2PR4wsROgXepODNt/4FVK
6u1jKs88pzMtRKQ6cQUfFbbI2tWvmCCZvQtB0URM+yofQ+e2nTAkXRw6HvYx2FHx6OaSW25CrL97
EfFlAMNG1PUDgXxGlvgpib1ISownRKVKxy/Bk/iTZ/2KvCdTVLXBsQCPElnlztgJDf7aE7wc0Uuj
G0ctt/j3jjXTqYxGSZz55cNLbLZkw3cMINK7a86nFb5jTD7qQxCcZL43t2j+/oGLgq1r6oFYbMnb
o03//dOeJPcIWota+OzrY7hXsm4/oDDaHnzSfNtccDGaSi3UwvxkgyFpSfsDGXTjHx0bqyzWMneb
Q0jr8gukKgb2hf9WWOb0dC/0JQE4t8m3IN5CaH+yzrS9iaaYhxn2xWYHegyhyrkFowTeTm/Jn4QF
Np8D0c3vZ/v4wZHHkSw1q8oOW0cHCNZdkAANl2MaL95hTWruBN+9LyprEhiqL8+FWX4fLrdysoiI
vEf7HL/NVqItw8KoJL5+uYgBtV/9o6S+j/CX2PU1MWpX4JsmsewrhwnuhDcSWMGlbbfbgcVd+LXV
o6LMFwp4VoLSmgZ8j95hrICQn4R9mLSyKid9oN/TxN0QYNuMgXKsx8/Jjk8hdawJYU1UgBER4WBV
t7YFUgzVvsNrpy1iAzhfNOeCN0bI2wi4odG6xIbPGYt/uKp2wnY5PJLKFypGQ2o3AICcMW/IkMhR
kIxNT6dSt+gwdEBBwBLYT3nQVjyU+v+5SZ2KDHp1KqXto+ybImaVO6gbMt6z+GBt6cUZd1rzdzNf
jUvxPJLQhlFPg4IMUG6EJfxrxFY+hLj1LD9hY0D1LctPV1UyFmbRC251KhwphZOxKS7PQCBHFEmX
at4wMKbTbkBy43/iHI2i5Lq0b/3ki5F31z6NwhbHPNEdTvj9pHgeyhy/vKj6eaCYL4CFrvgNl4MF
aI31+pQvtq1RuSxQIJbU2Y1IkNG2tdVIj+R6fw0EIv1dDhostwvp8Ikw/gRNoHOG1hN07smNbv2t
FVlTTYooSd7f//KElrYL4kpV9g+58Un3SDyS8D27Kj36Smn1R0Q7AzKeKD+YMFmVyCszIY703MA5
9T2aR/DN1W5q2TcY6LHKJhCf+xeFSBN0xuzw9HU9C2nfAewyDsT3id0kGhjZokhgyKxp0vRHgoMA
nDeOs3YEeNDrb9G+Jy2emtV4332XPaH4P53ft6PT/QYFh++GFSYWMQ20bjlRbjXFFAXp4mrBSu8B
ia/n7gwx/pMVDXgQbmlTvxCMmEBbCFEiSiFk6OCLEYC56m81f7aIY2r8RfVTtr+ToLu4oPWcg0Ha
PBPEF+o1iaC9gbhg07y+bxmuv21ltArzdHQ4XfXdzsAAB4HfbtEXROsy7wN4jmqsmbQgpqGerNGw
6nARmxnpqcfPBWCWDR1ker274c5nWbbC1f7RRdGyBGqlMJ5h3VIps46EtykQx0PlDCnjDt7jdZsx
RwJh7JKmPD6WSasvhSoWQ4Aky0vlE4yNAi9L2Bhkw5f2HC8LB+5FBbSYckUO61T/xUCR/Dn1XXDS
zDTEjYGwcF9PaleTNBdelcKgjFl1bqS5LV/shxsu1BEt7vux2bVwvdzqICwzvxp/jtSnl5bHziV6
uUj0QZSdv81SLXeSz2UeUw05adGpoAQIXXyn6z3N070/VLBVz2MSJsGDvv1sdlFee86KiZOrohWe
rzgZCIKaXWscKah92GvbBXsaBJk47EgIFBqJcRcXMonlqciyl7PygG/dLE8RYpQnDm4N2J8JPKTw
PdtdwvljEVFipvB+cLdiRha3r+S5PgrTVCRw0aQijaZsyzgCV9oiieLizFPUtIfdnxp14ZVruhQt
QcyMHJoaeOspX0h5V8xpFsoDfo/RwralNQC3Eo9stCpKN0+MUcmTuxtucw6DlBExdREz+weT8rvY
GL2LfY5axPK6uGO92bRad31Bt1zi2is+LF5OfGOWqyjLiPF2TZu5oy+y+5HW9ELMXQ4YC75RYsMy
NxLPi+8/lx1Nir3ZmSjbvfD0mMzqmjsIwr0/VkjN1MUHIA146TB5rC4orWDAykYOwEca1PmlVUWW
GepFScJ1JvsTUL1X7kfbfI5HykJ00VPSUWURMs5LPvPdjB5vSBZmm+1tT6Fuim1qYL784sIyHHED
SEyR81MTDul2ZjCBy3g9/s3vNdUsuwTmnSWB8FlJiLc294a1aVG70UHMe/XMAShNKNYFQuXVgfUa
qeaqqTSft6+6uyKhO9R5OfiFrYHwoJp8PGnUJ/rjY4qhinj96qucntN8hMqbvGd27rzFtjbWJmPg
PS2ep9nghhlACMfPnNkVYMPQj4DzoJJvbsmcoH8MocXKj0KD4h3ev42C5zwOo7E2QXTP2ke0wJPB
e0G27KqJLzoWbIedac5pGET4B2m45psf7AwwcsgwtuVfNeNibW9aH49ViAGGLz9lLvfyjlXH2Y+l
yxzFx85Udz1F0zwsf+1lVq8f3fCtFMNZ5QxtVHUwA3yg5Z6N3voE6vgYoz5HtyYCJ9PkptDSqBcb
3hEUMEU9YH1WKa9zfoUx1QCpPvHQq5N5wkbSe0kVlgkDWf0IPASa2BoABBsAeFPaxOKaONOSkgfJ
sTFhOFaf+OwTNmmvEjTTMCWNp8yu8rJt+4l9UOoMpOL5xuJaxuo9eA2qI6NWS/umQqDKPES8voey
PPgPGnyDYTFw1+T4lHsoi5W641GjpCfXH0jmK7b6VDiWmvctal66Bi4VM1S3iJVRWT4Q6oPYjUk9
2l7VFjcZSuq24WNlVPQ5aqEstq9qsM24ZVSGxYCQTa4APhTFhtz2wZ9mGll+CfJSFHrRQhXgyOmQ
us/2Ycm2OvxaZkqGysgOZ8znNg5oD29Pj8BHLMl2vdIOyKbOAQdodd4J/dW9hkEewRhY4iKefjio
5arv2Ye5UWxfHzcXyRcQd9d1XE5mkRW+UO3h3gPfRK5ZM6GPLd608uHVdfWfWpw1Wobx1Zd6zpbK
vRvOZDClvBiRmOD+Qa9DmUnpzx0SXibnalh1UJ+FqvECvNhtw71WymwC8PibjBLHJaJ8Zbi9G1do
49UflLlLDQV6m7kOZQHDCuba4rxfR7+mXSmXEqD0dDMHTJucDb6yCcK7rnHLXUOW8jCcK9kILCmT
LG27RuikZXAdhUzxxrLwXb13HdhiQoT6sV/y8AGfMD7tLeKnM49Fy45ZnZkQtpmkTBsGeVexMtLD
AqAFn1S0Wn03lcB15ly+NlzITfDz1KDD9X9uq1ZW4S4KEF8c1Dt2EXMC13rmsDmZFx9K24a1GDzK
smZPYT5r854y1XZdE0nhe3AQAlD+V9gL1yyeC/5NtRZZ+CWcHKDasQlTmCo7tfMiDPtJseODMvBi
2QQl65zqBKT+k8ewV6+QYgyPt8zy6fQjzNm6kahvP84sYPeq6l+f7tt0DcpM7xemM03az0tumPpE
lw+BO6yTvN/9b5oJl4EvpL1FATwax7zfgffjhSUmYoVBXKoi/FNgWRBe1R+e9YM1eYCjPPu6evH7
uiRTFGi9KW3cdMmOmMzmV+Ys98iLy+J9KDCZGFYXvU7uc90kYqKwvdzTXH1BOjVPMdcfUVBco0cf
6CITxMAFut9sj4Pj7t0ud9xMXzUoJZ1578uQdUbfgxgFh0f79Y7nCEY0qDf8C4Li3aHWhjnkVizA
RWJEthYQ4P53OdcxF1pzGOVK4mnIxzTSzHWG5sLr7CuJE8b86x/h6vvXgEVDuYMeNidl1ZpYZNYr
lCPqgJWiMYQsAxFFI5mrc2ImeAe33mDG9so1oQtmCCh493STlpMHwza8W0mWhHtKrPVLkitMsl59
zcLxaBEbc3hH8EUDZ9Lg4AaJSz28EITzIAICurosMqracpDkd24GHezn5V639L5k/ZjtQssDIm6L
1SZqAsuqVqOpF+GFSsCfm4kQe9vK88PsBoQX34TuVpuB0QxrQIPbSuvMcdh9MfOlVibKUC12DNko
NBXjZSv3lfpwohqFIXq1ZVlgMqpxFOjl5eBWtvlKgT260bYjhaVAyuHTAB7nJFQYNDrFGHxx1A11
onvh1yQYooq0jAd/vJq3iFgjmYWRxXT+5vKYb5Ph1YXw8MiofBb95qviKMqCiK67mg3Qrp8THWby
vU09WZNZ0oHQvfyxn5IB+QNLnCaGOO8dCZQVQcY/IuL8dnPz6bZCEP2RxfZDnM4N9gO3laQBUqqY
vyzZuPp8UN7YMklSRjnQCDGDvlRiYV9BL1+Dst1gV3acFuNDWYHYqRNJnLYANsR6l6LstGQxgZsx
he6VTHG16NA8mordvlFvtlGFbpuOgYLrezIg0HlBcAbX4ljItEcTOdRKgaEYG9Q9qunbueN6vkwx
HlzppKDm0kPc2bkTewqQwnYKLMLzzfFIwdG4NAwBIO3W6pEDBvs8CtlTWiEhmiUUIPNlpdqN8lAX
zO3VzZykXy6Qx1bBxsos4bUKc2zqiT1pBXfansYOJHdm37VHPNw1tr61lXTrrmgwnwzfIpchTRPG
9BrgYSz/tnZ/4dJkaeD99SVEuLFbWF7MWjKqho1BJYaxzfEE/v9h3kFO2MDPuomlw4ROxQLm6qzE
ublDgAOXy0ILw0YWOyvcKCPBzYn9mx5LfUBE9xMNmxUz4tdChYpN65W4PeKIb8ciMMxcGvuo6kHV
v/wrbRsBvy2CGTC4CkjtK9QviUR0yvfBlH1alwB4GhGM32wdvuENf0Za5GbpWtvT1GdoBBiXixDZ
WdR71LCcFLofYFSr4Sp41INjXWqIBZubLOqqz6hFq8g7pZ3uA2jHo9aVSzYVWDzrNYlDul4h6y2N
3ljaJes1dEUp+J/nzAVi3JqIdJfSrHua6GQcxkQiOEwoDira0mCo+VioGdYCPnkXdPoEieDO8zbK
RXTsorvEWRK7Q1tLhPsIttmSHRlJtgj35TgFnEm2OsZPcgrrE8OFhaz0FCNor61WjxnTQVVk/OrN
vupcqCIa3IkEvQAkMuGF/zhnytb0XQCdVORpVb256uuVJHe0HmjeeEQ09RTkTaW6O2eQ1BIHbyR1
yoPErL3lSbBm3rjhwRjDj619WTBTn+qo+OqlXb1wG8q+0ZGm2EEuijpkIJZZIXFNKHGvIVWK0lt8
q7yqfK46A14CbCqapCGy4Cs25U5+YNBudkcjZe9rrzIoe7TcSQwBDLjnkShA20+ClSlf02HcR5WD
U24j3fs4FAuBph0wprVlKLRnPY8EnVxINi7/n4z3HgZ3ULSphK9VrJnnOJZD1lT2WdCR6raHj3yw
zZQ1Degbf7OXUrzjwN5DZu1Wfn3O+bJ9r6fM4MPlBRJZjMlvfhGu88rQzCWgVI4J0TTFrHWrLNrS
onJ6suIIJJz/kkcw3uThXhHTHiQu+u6l4mPEB+V/fDnRH5ZIOYjmmCna7MPTMyxfyXFaAgRAGNpj
y9SXvi2jQ1QboJIghL7JcYsNVPZ8v7fcTPU7heitsSeQb+Wm/l24ijH3FxELUCEmi7RuJEtvnKN3
nXb0uCUJ1IjDdPcD3Kr0L9A+2C7mycHJgxcfUcY3zPOoRjXid9/LsGbwdpj5akw+VGiEOqctZbN0
atR0KnSLHZybwt1jEi+SAVa8pKLJqp1ze+HEDoB31au4WqlpRfAb64vUwZE3jUdYbJQsGjfYcDxM
MDQ+7MiLPkQQRmKwgRvHxnW6z5UQPXo39fk7zqOsyl1HWSxkg6lbNHUcuQ3PgiOyVYs0K4nxLjAt
AMZWG1nfycnhsVdm/ZGdbXS8rTZQooWP91P5LNnEnfBEVRK9TJ3C0hoCfxbups5oAtWxkCg4VUcf
8x5VLdIOhxHYV/TQwr+AvMfF9G1ZotCbwyzVJSu74rOgjBbb8i3gHNc1+1Ut2vD4C1/kdHv7SDWc
qmA9ZEE9GQ9pK5T0iSJHhh3zoOfApc3NznqL8W/OokyDTgOnCiP+R1xg+BQxxoLGFGYq2cXTQd+5
9RmFdBIJ045goBm6sFlwxYbjjxcjB/He1pcB4EjP0yuKvnSeBspNlHiyVyAmrsowtsE2BAFbl73n
XFI3PslA21uYTCCLQsLg+ouZjGaiBjhqSAcjemM3/np5LHkZhdXugHHfzBOlnhUKDuQpdtz0J5IW
GT94dspg4H1/651cogxtv3UfpwrYGOsLq6tgDAcUVBNlwW5IoUAiEdTvZrRZORe9kMkKO7N/yYf3
xX/tDgqQRAhnDqRbrKyiZzlPjnYKBejw07kK+AXyiqwhD05I4x6NBKg5uz/LLoxG83jI5WY7i0jl
ZST//INve5SuUJbW7Pu2jMa7m4PDkV92zVOF5+9pfnOxt+CbWEZOP0FZAq7o9quuldpkOB8Qs5ly
5OR9O65De6pDS1Cg9YKfviIgjKmJlO6lgNqe5O2xh7chvBnSrG6yaYtHNJlQrI5QK070eGd9POQX
vvMH0dHs+3EW/XwgYgSrlxYH5V+1HUSD3UARpy+VtqRuPsXAzeaU5EEEdzVjHEVKoIOh7pRX/Dk+
4u/uql5SbwOKy6usa8Lv9YDKuelCikxKp8EECTN0DiOCw/H4kNSZvARuLcAcQtgULJUDr2oCmjqo
SH5UuVpNfwHPzuo7uz2NulGaG5qDjjZSZZ+oG8RPJ4iQxdYp372FgaTLDV/BmS3uDEkMiJz2Zw/u
N8GQ9HWLpuEBrvLsuT/Jr8+CBPu4goZi4ff0G3A6R3PWvCy8CZrGzfwiPX7qB0CbNKPKhENlVAYa
L9PN+BcMJeACfg4gYvk9z5KM4XLORGcNePotPpsa0o1dEv/7bMjin61sgWmgQMKLQQQZhZAQRSrn
GAh6ntApATwdtCHAwF5S+9xTwrCmY3Y/QlRETr9doS+IN+VT1MTRgJv/FgpJhXEGRAZmmREYgzlv
pQizE66zLfMFD80jCqe8xpxoBjLwa8uCjK4a0nYRxJYZfttJkpvqvCjxaooyT2o615BsnMIC7rRB
R9uxBPkHz6ChM9sDNKE0xdFjy60qsjfhIsprS2ZZEjoTs2no558yookydlm6iFCCQS8jdaoeUkpD
yzhF5qWsZdxOuUkHKVT7aYLf48y5jgVYKkeHOJ+nC621YPdnR0YmcAVZZs09qAT+iUKPAP2neJqb
+DffBG7IC4E0pKARjfXTS3UE0pB3w//EK9DH+Aw4sd04L7bXgYSPGBZQm3VQ0r4KeOQw0xSowA16
JD7IsuZpbl+Q48g96+cYCc3i0+HoqljIKJcdX6+SVc5yJ+RwbOMqwbPPilhypHZ0D6kLxtelsjZX
Q1afnvh9rL4tksG+4DZFM002FhFnohmYse89E/mCK9OFi3S2IZYWyEGa5D+b9pkdkRIBc8XYTA6C
tkNTorPl4UuBZZZKzt+rgZzHMP25rJem6m7qYuMI800fyLRPVW5r0jEbKcs26/IyJdTIr2rjbjOP
/nnDhypaqVjSX7QQtnAoJFzga4iUzgOn09Pysq+SpEttDoCluPktNeqyDjTuJOiv6eCCScjxl8J+
tSJbueTu+NDGKDjikRe9QGONpgL3r4PNX5mNjB10HHN+AP0PRlhrOVOgch0b+PRWOnEvVd471DEB
QtEo/b/3zrIauRb90ZbH18qUhiR/UMZWujMD+fc/Na+PGXpgpsMUt8K+YqRxj1ofuxNQi7tt6nvF
fdPbpoEi7B5RJLc3qNh2VOUE975v56pbGFOvafLC/4fW0931w+loU5pSelR6EWL7pGKIXlG1z2/l
HAkf4RQAo+LPiRLAm8MOxJrXnCzA6hBozRGOioSEQr8deZwWeNBpyNpI3rYsAuerXo5ueUedDOIR
FXCG5PxfqnsMk3KrgaJk67ApsOtGII6n7GTJjNyST0reLdV2np7PtDfWkT9razlWQ2Ch3oVoHwIn
DNHIpdOSYpcfXIupEL8TKJOyTHr+0U8grULdcaFY3vWxBlxR229wYht6uRD33/FGbGCY31zK8XlO
lzRS4Gy4vqmlmPkL81RWXmvMA6ABZp8bhn3XqqexA9iYXeE25UlOBBd/z/Fi6+Do8d/nPTTmtVep
e78oM+KawngBNFKxBU6OPZ+bPHQMX8Sg8qoBcOLxljH23FY7k5Hqp5sgVw9vMHUaXspR3skat4yy
wsrcIb6XueH1I3DTu143/mcbIudDG8LfS7YUifRKGfCnTahIo9L5kp0+qk8ty0NSInQVeb3jWXJT
jWqr4Ym/QJbsEkPA6iWZCA8udaqrHdiNc0Z9Q3lRJrikj/fq8ha75U+F4HPKZQcMlIr6yKKfctDa
44vllCGSEUCqaSXQmmR/b/DMfaxMoKzjK2GwifbWKXzfskXpZrpM86FMjDyEp2AeC68HKZrDT+p1
WeQCtIj8a4oZ4cjgMKEynyOw+XzdiWyErUW8wGXW2wbqM4p5EkTBSyRQYtqYPM5bDMPFXsjFx+br
Cr3plokk6RTEc6OF6/7eBuEvZF4v1h0SgP5Xj6oELFxvNAWWBCSGlqB9GI3eKLi7sY7vnhfobZ2b
Yy1jm5mJM9O9tmQlcbd40+D7HxDbbLrjhwOhNA0zMe6WlKRE1I6m7J0eQarOBvu3A+rqFq5Rb9do
LnOHTnyAbWClZe3v9BiUbEv2AX4w1ysxFhYW1y9TzII3m0MOsupxbeSMysDm3E6gHcb189BAsbfH
T+4lS+LeffYaW6d5JdmdBnzc4CdlCARTSz/PeNiymAQsTeDqHu9TjY8oRukUii7EWt4Y7Ol1vu2c
AXgexH1olSuyO4fD+CHp6ktmgMWwQXJLirLM4U1GRIdMFn6UeN+Y1v8XfyJTxVH1EejWsf/LuEhL
VeqyI+SkEMXyVGbCoK4Gw+bsAd334Us8mp8n2QpuK2yZPA6ovXmLU2o5cCC45LgSIAteY3DNiqhx
v4ejwBdAv9TUEdN+ASK2F/JIFlmjHxaYF7sXjngK2cMKnjUMQasgIs/7012mrWLjAmeBxSokEi9L
Zf/deWB5VifORmboSY7u7qqCnUWkadjNmfbxnTcv/MiDeeuQuFXYQdn+NX0KG+4f2INy0/YLVrbw
dlNZAiWvJRuKDlHq0y0SGuOAs/pBSKo4fCE89NuXj98iXDidOPPTVUheEMqzK4qHXJSaVpSUPayR
uF3PAD9POSpD0Bd8NpRi1Tzz4rCZas1xZHc9AK/RpprriOB0CJNJg272AHW2nPEHoYCgH9mLdS9K
apdXq+UrB3H6dPhrLquITOGHIWL6qxF0eWAbT0oh8x+p7C5YGkufkE3eqvBbrH70HEblZpcR00DC
eECfOq27XRV0dDI+xzBVLX0cqAQXdwJmrl4S/6UR8FEx6BaeDkGfxhtGBUoVajHXTeufkJCOzx6p
LNZRymRjqOXVqGxv8lYS8dtMyH8cEzEUD3Inwp7XrV6W88Vrmir4VwGi9mao5vkmBT4NbTWDKovO
SKtLRLC/Mf6zVtetckH4UD3mvW5mtw4T0oRLUAtIBYIIoNTRmO9wBuXoGnArzvlohAQ2kerljTki
EOPd4+mfxtNrbH0flfamYLNG4j1ZOpM5NkwIAWOYYOI/lVnl8Bzj+KTQxrFynOu2TjPrz6iG8NyO
/8VrJN73TWHi+wHUevfxLy3VBrp4tVJyu7qQbBYJaDBLDcuZxZvcqfQ92g75OSJQhAzw2rxI1CqS
o7YaLDcqGGkTUYxFALuZJdv7gi3riv3HTj8/CDHOgY6NKu8UJNiLYb8QvonjE1SrzIiu4h8mlYSV
pw2DzRkQfBMZ7F5G+g0jha8sBbdlcccN9tScrpLTqU5oQYrjIeTKc9S+9T7s5Fg9U4nwmCM/p8jP
+KtWgky3ha9A3jKyFgH++HJMoyolW1YhOw6sATykJYuA/q6kNtrkOK/hlGPimPNuJXjI7jb/qZ+n
/1SFBkGm1UzGszrU+uRm23lsBhSmwlqYywnVfsbT7kkq1k9YwXUOT4pnGnusmiRNajXak3QKpr+x
S4aarexTu4i0Ps0WzrlXCW9LmdYeunqO/mv2+edqurgmlE1MO0MXTlU81hvTLS/WurEr7lwbDwrD
cFnWKisUEBdnuG39hK8XunWYZpu+rszXKoccJngiZQ3czydHJSCFQxXVSlEM/uOXmyVOPq2xNQfT
my9A7UNSn5AbTfb1/VxXiTOO50558RR5z38et/YempfFk0qpH6EQe9poz4K9pshkJhPeBwtrcF3X
hlVgZhZ78tqboaxmp3ScbSv4t/jgDrIW3ZRPLYok27NbJR18YBju9+rEZSOasx2l7eSF9MbK7szy
q5PCMrfAObcYi+s925S2xX0NqSDnIDEHO0GzQD4IIBBGsxayFjmkZ27EuoOTmC8p9FSdNAhqb+q8
Noth1LgvXn2VSQNTDo2iKJJoNHZ7jnWaFDQDodslFuFJWYg9ueYWcY43p9rCaEBx7kS9blgvOo8l
S7akTP9x5JNSDqxlAJeiHbzgMafD70AdPB3VF3mFeC2b/llqn6Sncdk/si5IE6nbxmY2hTs9ULEC
aDp5cRQvdKK9QZzCwICIwPd50wTsLq1cmgdEhhWkiMfP6NEhtBouAd4tbK0vxTIRfLUk4cwEBjGj
NmCOTgCW++pBDa1ya/ENUCwDLbF+/nPuImiakEIKVPa95Vy0EJrM06XAQHaNXOX+5dX3uniyDgoa
nrOXft9FTiAWeI0amsZYsKW/6TkCb39EIVb76FsQHVvsusVrfsYHr7E80F4jwZK/7LBOPbp8ZQcf
bkGUhfBVbYPLIuClzp6s0nl0ugZ7QFxIJz6rpU7vGiffFcml+RiC+Nw+gbz0GX8CjP8bZld0dC3x
KApPCer1u3xqMFl6QHLAPa1Vs95I224krOach/Ynn/d/Lg3dkcApHz5aWbmogCWAukZrXzjiIhHa
yayhyvXUPs2I+OL/URT3Z5bEJWn4I8Cdgpg4b5QWVsdLiUca6BrXKZI6KpCKmHkt1FSGgI8mcA1o
L0m5jRB7oKfxaO7s0BHEbLQ1IUvU7LBBObhXb+3h/+TpNqFXRyG+QrhxY+6ptyFduzOvJ0xl1QHc
YKtxFe+wNd2KFBqQ3hkm21pJq/rRi79TRk7imnGPMp/jWllOBiFPQ3F+smH6RJgT3Fx4CCsOM5Zw
9M9GYwqYxKq432pflGeLlOKf/FQ+zhRL+j3mc7s/VA2qghgIVfgQ79mOoA0flFQHHRyYUMRQ3wx2
dmU4jamKhFr2q4p8MA8R58KRwk58LXCknJX5U06k/33YjUfaFTvBtoNH7HfGZtA8OeE7p3zNxu59
4LIJHav+tgg1FC9J6HUjOf0/S7kbcyfcS4KOGztOyX7GRS75+0aDi+3xcbGKiN26EfsoFN51a+js
VFLcWhmr7TgMToLKeIPqRaHadsKRTPp8nCrXdJomnFla4yFv0gxawpXtEIbRr34tzRk5jRhlZPDr
omJDxqHr+oPK3Wrs0bgP1B3trq3JG0SKAx8XHK4VJP9j7GQFI+rwxUNYGsYLwV9h3AVdQy9dqbji
DqBF8v5O/XfTT3zeQQcwfLqeHcPVChnQf2pdQE0qc43xOGGS7ql7Z1IZ1MC5R52JUD7O0DBvBmcV
rRkhbs2UD4wrDarSSb7lKWUzdpLSQew57i4xe3DCr+n9mTOKkAH895YZSQrp8gHfYeCBzuBh1eOj
hAr1PpnUq0H3gjxG3EbDyTKPafTzet09XghcjumsWPMMdw18mjU0TyxVzpeue9hZLeVEv/5+T40o
9MxjwoFUY0/us91zCBJvOnc+H6qwCsIsGrfkpQFmCvwdW0Pp8s5WaMUT1OprRKfwxNYnM27DuuW+
pBjZrBGmv2KyWj377UX3bgu+IMH1MEjR805tiztoraahvYM7N7tWB4iuLup0Bb/FjV7oNhHPVTRf
bukx4X1K4S+XMiMPtXHhn7x0XPHeWextNrepOxw8ip1flZa+3Y5+cXU31RVaPYper9SwvUdroUFL
ZYIK4M0AIeQbsUrxD9ixwXkmOcjXL6IYdFM0gmDI2CcvOC0Ym4AlZL64GpSVT495MWSugKEtOtIy
+kYjwxdV4Tk+tYQ+BJSQ6AuUePP1XsuNwRXBMqXh4olOmmjLry81wUmewL1xYe+Z2znNajSHkEhu
55SVDBbNO1O6meFxo31HtMD11e0iyfKlUe8bffrWGIthrIKsWobJXJH1+CXslKIqSgKjoD8srr3/
HPP7wr7v1k1M35RjF33pQwbCebiZTqgw+cwabrY9ZPLqupMYkUkzUfqg4MKjgUdkNHPlkRt2LMvc
HnPj+I4+FczH0UFSdeVy6Cazd5OGYyqLQFnJIqG8hxiIkEA4nu/ZW/SYANYP69K90lKLh097LeP1
+YIZ32Ni8KUttBhH/TiiXxQpA0ZhbKwqJedUWah44h25WxcL9z6S2NXqtuv0C1NqrrR8yHCXDrXl
6vLu4PvM7/EAXuqBpGoGUNAwy5IpHM8Qu771F1mER8ZIHLvysFCTGdNIkkN0UFaW6qygfKPN8+Dq
xMyMcUOJsWn4K+zlhYljW/HVugbq6Z4nBEYAZChY/6a4Ppt+1nQZHewB0Cv+CrNG9FRO6T/f5tIg
6dOxyNuadbsjyqAlV34FQa97ku9C/iDQLEyCt5uHL7OhxzOsTeRfK6VnMgMNsXvrdcoJRLukeJif
p4VecEWNDtYAAkB2vgFnyoPH5Kl7F0wPUoKsn7qHY8QGtGklX2bi6pq0xf+j7/XAe/2/0kEqDSqd
IGEJUFDRIidlzapxl68MBzsdAma7bg+isgz1DgSSpY+69Fxx5sdynI5nZ87gadZC0mEQqZh1nUH9
cr0Eu9OOG+n45Rr3MQCrPT0uIAk61QSGtQP9e9wCjNCBKdcUm7PNUfhjCgKHYVLkXjSwNElBxmxw
KBMj1RNUI8Vi/b7+qdL0iKOv2QEq3eoxwkTRoog6p2P6P0SQSFsuH0kE27i5XTmU02Q+jSUu0dNj
ZSYIj5KTKuFbQsx8HGCSctcanr9JR0pVMkrH6tovZoGf2KNhGM+Go7itABX1fXMT6ltw7hHvjbaN
+cq15JsweHkL0YW1zige6ny/R+5Ct8PoklddJFZ3sh4sMDE8Xq4s4thooRQQv4HNzvPk8ntfI2DO
teb9BTF8IFVmbhOfP3dVkx7qcQ9bMpwfXiO0uCc3xRSEUgm5KZXR6rtxLOhvjDoddqKUBeCGCt3o
pWXL2bZVyYpAHBVyNmYvNYC4XcsbmIV1T61lJ3K7ZyO2/LJVW4EoNPMV+uMrsNOa0s6kpvH/UaXm
bTsyROdccoOgQIX58kaVNZ7annrAMAjiJ7DZqqQIF0/AbmJQb4uznr1M3IzFRfiuNBLaxUlVuHZX
AsWlvKrxXNZ8CvaNo4TkvLO1ih+BzgxsvRK6B72lQFD6okC/rM5H7DTp5Yg+QEZ8txjUCraXQvZg
DEoR5t/6CBoJuFqTm9x8UOYfY+V4XGuJXsjqnyFqgUNspaJ0kPoUqyJ9ompOBwGC6TOCww5UdCv1
/hD/zVU5d9zHaZP2a8024HKNGMMcYRCHskPpAZuHWDMcr0c88dLjkji1LTASbRScKqK5JkxmTmWZ
Yudu1umhPOBahrwAjnQIlTQWPGmqit+5vvaJwRMoSriUMImoLn/mezsoqo0ST9fIRvkibVxHCPNW
2JefLCkEP4yuhcE5msMqNKCSojfE9Oq3LvzkUEH4Gh8dTT43f1tMgoWEnqU/oaLNsK6WJBkKHOQ7
rOvd+pUz3bCxnFSQ6+D9aY3AcyB9HerRRVDZPoL2H6o5ajaI2beJ01rX/CCNBR0nGE/XeJBeZIUf
8M+mOldNIwyu1GQN4h1nuAvaOl8QJiRKe8nHXDv0auMODUVsC9wjNxpM+mksGbHOfeGig+Yo1pRG
7tAxn7UggmQO8RqCK0Pb91f5DYKTvNzr3KaTEw9Db0vFDY78rmrYBBLhoe0eXcIT9PY8BUpZFbZv
8V2TIpHa9ykzxfjOQ43QQJRo2/AcMmNBRfCzX15IUaahjKiVdXYMrJ6Xzmy8pfEbfqq3Kv0FksNP
mPB3e9lhzv4i4dCkXmXXcCuTjIgEW/YL7Dr2OPrjMgPPyNSF+ovpESF6uwoqe+SKPOCBGQpBogt3
Xeotop5TWyeKn/WjK2PaMuqrnN2sH5eI2RpB4gwWNmH/TjUvjO+kxA1Y4UwIu50DTFJ+qDJpWVeO
SgZDevuKAFfcBaQr2t69k7oS+3z/yJI+Yj/KlIct+js2dvz2Vv7df+Uy5obOo9LEqPbY6LyYLoy8
t6/h8NA80Sg0w0tlZyb95WcA7HBm/OYpUuXvznoKm2sS/7eXEo8W7/kFweQxbkbwecsPsa6dSzHc
Xo4wMjXJDfM2zdXQbar+8+LcICCi2v/+sZR11JcvKzLuyXyZjp+jl7RRn8OSNJqH4Cb+XtZdpMa/
Xz3MeHlUN/QC1qy+upkkBxh3Sjje8n8VVjf6pMFMxo7e42f1gSwS8Rg307TNrurBmFe88QsvAjDJ
6FfCI0QU30If8oX5yoyHm3FNkSEC8yhjy8LY6msUXZwoHO20N/FE9UHsjGS+cObsjAApRlU3VcZq
ma1UMd8fVEe3HWoAZo2C7Rwm1+s5tNi7ZPciQgftN8OcQ5eoO3NoxAuHFon4Vc+bTwdQINnmBk+/
foUkO+dDdTghmTc7Ej46bMerKGCp136uev5Oup96sYMox2oOtx9MF71VQLQpsW8k+D+Fp0f6BoGf
rsN34j2enx4xxoSZsX42kIzG2dZq/TtOaQr2VqXXsGYhNzCFAmX6Y8oOBqNR6A4YPcGOZ1AQpz6T
ZKGvGKVDjPm4n3bpe9v+sxWYjD5Gp1rBpIZcYCvkjM4T208wVWQf0YZYSI00OsqXxgwg+oLAPdbT
i0Hfnsxl8fRqGRbiWoMTJ4jrNFDVzU610YkUFQh+tzDkuxf4D/3BcL1CBnADejBvvjjZTPragKjy
FEqdcsuiMKAVzBpnwOayIcdHtr/gdVK+NdwKxtl9+umiOgWqLlSqzlHSKScgBvetMrtqQFiA7XPi
JPXoZXotCP2NQ95n6Z9sIIaozRvxZkUhPdEb21aFoy5jutQGhkGa1/BhgJl+wAz6RsHzNgohIH3v
uqWTatZS50sA6lwyr3LdJ4GblLvmvuJqgpBkI4UKJ/KcILpUJA2edJwbSHUyXztKRayvz9o+dKHn
sbtZktJN9hgQypCjUuZ+0W4NSzvA1J8PC6QblsJJ0pUWjnFCwR3/6+Fh4cQ8jZG/lWX6PofRFk5Q
l81sif8GjioHviMRg6ctB0OhG8Pli4PDxtk6y5eBba8IV9c7oFqEBRgC2tdU5AuDbbkazbxRRqhp
hjB5mi/DcbZbkV9Rfj5PSgykACOFohtL/C/9xNNQStYY30PrQnR72sDEdl08nRjfCKshuzXMkyvM
gdakzKWM5TssGdrhWZ3blOV7xRqYtjhCzt8pcrOT3PwyudA2pKWiuNbeDPOlYfPn5TrW1WsV0JsY
SCNyu9ph+MCu90SjDPtx9OLpGgn2rX++kmDRhoaQBhckutYzBOZ2YeBXgDauQ3iucYn8zuLVtqGi
35tE/ML21ruYGqaarqwuKNwjlmP6zsLep7AtmusDMdubcvLjFa6OgEovWJaSCvdEIW2SwV+kQylE
YFTtIhDuWaRjPo1WFw6ODULZoUXJ1lIZd/W91SRe8jG6pRsbBWhDparMVmRpYWziGqjxwRGIqeO0
jK5Eq6TBH4Ezvk55N8FsyFZofVg6uSO31zYTAr5fvhE/cQLeXkS0AsKlTAuZ+XpRFnjZFwyhhmV3
N7QsJWPaSVEX7P/AwfCDJxBEz+TBkztCa95WoJJlPc83SHhECNZ8Py50NwO2Rc+kQCclFLHJDthu
dBhGkwfLplNYSQlV2rFEiDpL3HzQs63XIMjJEsuxgbpoMCkVFckpfEzNBIvW+nLIef1wNt7G1I51
mieFbc7JWqZLhQp8C/zJgGP4v30CPfPKBOyIvGyfGzTMhKzemMLU/s97yQZDZP/KYsOMpwNj6E8H
WJKi2LtvVbe5NeMt4SfwW5f3Bbfue/V8PmGjWtL6M2zTovCKYwbW0LRbCcCxu3xGkhpKNoPSllSB
bw1kTSWOKIlIjpfouRTA+eaVp9FQ5m1WyTWSuXH/aLsty0qzD8XUrfjeQ7efEfak85TdPSYUzGgX
LskMrZon9YbFE7DUWbrlLs2T8BQ0FEjndGNCvFPcubhtWF7PXbWo0Abl15y3wGclnrl5QPDyQ413
Pwr1DfOVQvL6TMjY4MnFm62Btl2W5WNmN6/z4jwupL8OMuisrYvvIb93aDiEbuz8wrdaB3G+7LfA
xXeOimLMRCVDCrYUekXztLSC5NZVb+Gw8Ss6LyxiIG17rCFvy0oGaciy9p7Yh4mYOT90DT+HxqE2
f1lnjxLWIiyFUE875WO5Q4kyr4kBCp6xN4fi2Giw6qfcEU+ILYRyl4Ij7QNuHXp7KQ4spmBOcDCC
6l3WoShe7VEZIMcHgrDBVD4fl9zR/0BVRjV3rIZjG+oSZwnkygSGCMU495gzGi6HnTMQGRJzIeBt
O0Yl+U9QRU8YiBbZwXGxdYHoskbIgJkoILl/l6et85B6lj+Q/UKyVxijdk99BqImN5NJvq9z9yDk
GXjqAYArdswHNPFYxPWyy8Zt9Rv1uT8VBMFHgGVLgkMGkPaD+bVaHNR4GIkbw78XV3VrGdhPCNkl
8tHrEatgy44+S0KML6eIkBGRmmgynVeda+iYj4jY+drRyY/zifLu4vAK852cN/c0UKlkrb0/VwB9
6uasuUKIx9ki74YJtA08Tsf5w75D4BEV/5hy5SeCW5qky+9xFwMtt7bLjD9hqCblWAoQEP64DiYm
n2Eih1kLq/V5ZwWndgyaxL53aVF8GedzLmRArFx3HbXK5W9dLpBpgO73vevXvquCFtCeXn3agqg/
sDsZEg2y7aXW/BcJwTpj5+rsdPvKynHytTKrY973uQu+jV2/EuX17osxRi8Flzic83CmGwtKbk1R
OoiemJYcKD5GvMFKyUTudaoYxAo3F82TBL5A6vdFR3E4p/d836QAWszvLQPKlrYoBwyKSVgKcpOP
Hh3lv65usPaeNqF0jg9VhXt9GtYFfnime/jdYceYhjDTU2bcmnN85iQwd2rv2P6pa6dRwKd0Iyqu
nGJvIhOYx2ASFAX3ngt5Zjz+HcVtiU2lAAb3/QfeBoIJwB+Esl+fI+fbiRBQ5oLJ7Iz2rwuqetBO
m/AVfvuaECQgMiFqyUHMMWXFGzgTXnp79rd2OaIH0gW+Qto6wfoPycCAvBvtxlRjLELtNXM4jbaE
2IU73pkcBI+uh1RJPvI3LRhWtWdoyBNDjfNRIYNb+k3V0PHuM1yyyobsrMy/znzx/cIVt2fvLUVN
QxH+91rLBUWPvQXUi60H+VX+Us/51bR0Zw5LhEXHfP3UCBNuZMfcIQKrNQU+mUGoNrJxneRHVemd
q53xLzQf79QfZdu6zOSS/Wp5/l/BThkDL5+9/2R+y7cgBMIoHUflwjbm5HenCpamvN70gtwVue0b
Hde2Er1afxfWhDb75jW7Ewzx1nxc89OktzQpqHQJ5qSaIydVpmlnwVB00xSWj1nQLhRWrBryF+V2
WRJqSEEFVsBHNBmL4XhTi/1EYqturjq2Nuv2Kc+YAG2Ot+zaaI1cCtS8mW+H97vZg7GE/wgVWDq6
gP0eKOBtvipeZNSeAGD5aTNGT46WNDjbL30jNmpFg43ZY/waqGKA1KTx5hYtj1kT3Rd2lb7TSOng
gEHGbHfYoSgrdC3pV1cRuSDIJlN9D8Eu5dBgdMFeGmyy7lOxU6eZgzeQ1ZGOPNyKMKLl5+6lCzrw
stbWd9hG8oV5H+oIqI99d3fYEUUqvoWlnPFZ38/xxY7/iD5AIl7M6D0GdbQoGQGfDe/QaLoRy+I9
DtQ9UanwlDrTF6iB8iFqb4IAfJ5+DjKgSYo7h5Yb0F5XycXtMAyoAD3pP2tSjE5cNeIkxfESdAlH
jo586/Q84zxJAnPC4GEbc66ymFOMV0Qz4wJZVFAIGkHDbZZyF7XdJymmw8yMRowOW6RhZ2+U+QAB
/QrLySGA9EtwoBceMiEev1+hqC4/yx0Vfj2umGQOSw3qG9++C3R7HqK6e8CiZ0hXGK0Y0pu/EBPf
ClGNGdlKr7bV1O4Qta2Wzjcsblh8jN54RudCTYPqCrbK14WlO2GU6Wbuf+F//+aKjRtMps/QvgQ3
WoH+C3lKE8Pf2Ha0Vc/Ql9345pfUHtjTmrRlB+LrKp+wf9sqreuGADKLFDH8pV35LQ5J0Bu1eUnq
MUiGYeOOqeO7eynOVC0TezrD/riXYAyK6iPd47odv/Yc91ZZUC+GKYCEOKNkZ2YNwKksnQsRsxNr
ydFsCjekroiN4d8n4f95Zng814/NtVaG3BnBww1I7MZG73JkFuZixbK+P08n99/u8eSbL2bjpikR
GfEJezgJVQK9nb7V/TtTPZIfc6CUXYj3/fLQVTRBE3Agn/+L31DwxKkhPaoXb6DQ12rMgtaEfbAk
YhcAB8xuB4/q9FGmmFMzBbEZTAizEV6UjnBNmZ2M/Pie6+sikVxCXFqMQrleXYHmm4SmPa7eYzHQ
sm160BtKNK84+ujp4pFI6K5neVEgGda1EaDKwtBaFqmyEVcHQ7X9lV3KTQ8VwB7Tw1TpnHAa2qru
Rcvvay2+jXiTffhArp2aqgt15Tg5FU+VZdV+/Et+No6fdXPa9biVdcVdLc3pcvXu4l7eW2xfEyJm
Pv3WvIOdjLcsx/yioQWmF/92j8ce1tugljcQHU3z2ZiR+xMxsMp/3kuZEHpNfr/SAZ/yShqkFgHa
StXLcmR2pmRazDUXvOS478W7aNRJ+0rxXRVwL1GQIBjKkjdz3x0tfKuvQ62i4VlMuab8XyYRmkbp
RH4eyMbduaRV0EMb0x09/dMnECHA4Y1rjsbQ9bSafzfm12JPxfg5BIQHaIwFKanqsosq/R/kMZaU
cmquTlmgtq96D3/Gea4na3BvE28BAPzfVz5YwYtvPALm1cEtBfTmVouRUNZ5VaewHkbi/ip/qRYl
n4/mv4b7wkO4leRjxCRUJX0BlAkvLLWeFaaZixPuzP9LvTFmbbuTTGnB2rOWja7V3Z+XWQe3Qs+h
EA2ebXfyT/vPETaCy7pShKT6K16m7IA4ei8YU2ammMS8Ae+CX6TnjaJmKysdTIGzsRK1AqOlL8ya
cWFJD4FlUyLLA4xjRJo39Aaj43VozCaOXVpDNFNK3WtBX9IKadl+Ka8oSur3j8yKQsCY+iee2/I2
FQwjVhKY23id5iKci0muTcdDZbsfM0e5aKTs5ehykqWmnAG26qw6cGuLEd2MQ2LnzrtsNxkwpYp/
+IE37PWgsNXZD2fzGkRP/CGq3RB+Yv/Nb/VDfO6ppj83eYaKiR2gIy4bl+XBTzI1Rbyb5ndn3XUX
9KgpK/PqOwb5Y18h/9ydklLF+DO/MFRYaynZCQWeoBhRsLePcM9GuQdcZ7csLmU7m1RNetRswNNS
HMduIHZlXCTQI3oohd3XPyYAx6yaz6wn3M1b/XOv4ZyJ5IqW5EgO42wJ/rIXxlKyAve3P1/8Dyle
g7UoadH8df0OP1sDfZIihS1NCfTrLpTW64NLKdc10bBKz32bkfidpMUJZD3PkoOn6yMtn7Ouygn6
86N/6T0yEOo+67Jf5f0aYmBDnnUM0XxuWfVLDqqHeZyuE2ZQwD2euMX2jmnXh/0sM1+t4RCT9pvc
VOctEoZxKNDexpqH3FVcBGBlf0aLtiOrM8qc2YmQp2TqO0eK1MjU9YZwiPgfTXd8Ajd1INF/Lj7e
tnfy4bxFkH5S+zrjRHaE1BdwLNA4vL03faptL0FEBrHUTO2UY7g8HQ2LCV9MY850KnqaGL+Rxh9m
5TRadKrAkRaQFKtSgV4gmbkjk2rwbvbsVKxz14ldGapRbT9yuEfBREFq37B4eiA34aFWL1jn6KsQ
NfxX/tupVwogagkyw+2GW3HjREMDiYH+K4AXDhEcSpP8PLhjURzyu5zSv1q5hmjOj3OvDZuV/Wg+
IvzkdZQoMAgvXSCGAaSR+uR5wo0U4ZLDm2wED5XrmFTg7wxkMAjViFKDsQ62cKkMl2pnWBV6MLFz
BjALiFJ5qg2D888NTSYvI86DgpWwAKZ3sGQWJYLsi8Bq8bNvOalsTvsitPwu1cqFsLhrAMne8utA
Cf7DQ2A9K3za4Sa3+AY6+gu4XOEE8YyjNtVpVMSMTJsgO/p+KLd4vqDNcgoKRM2/QxFmlqbqBK2y
0bKc+68mb7XqkqiHM0oBvGBULIHl+kcDxvDKNL+MNMI9x0RtXZSz/SToACOvCMn9yZyu2xkbFd7E
7SNgQCbHhSNTslkKaaToYZrAn33LSg6PavqA2Bk7dQcEBhCFlj40Ntk+YYlfBfGhXbRUuNqBWdhw
MC66917zhhXVEfUxpa/seWojfP2Ygwb1W/7jRTjO1SXXsm+Y06lZIO6qhfNI/g4DbcqG94k5jHcG
iBHusABh7p9YosHuQ5fKDOT3CO6UXkJGGgVxGqRXKW42Bd3FbB4NZ/Z7ZUWTP3ZpXSiAM2n5/sJH
2eyvkr9ZG72RtKl+ntxDcJdDcycKQgWQOmWCETCUStZBDJXvOSqUEj1KS7OhEAe8PHavr2/W3PGf
ZRtLfBQd0YCDJho9SPW8RGV769UWGoPWqyqcuTgH5JkhLORLFJI9yrvNkUEm9IUSQKH9okBQOwIO
cuxzuKfuHqrF2rxjLYluMCZIEcafaUh9DrhpaH0q7la+NWEy8Z1BcTVKHFn0TmUEC/vbb/gK7D1G
LSBN2+KqfLc7/jLc7NOtB97IpPZfD19qYAnT3P3TMNmukgiO713s9BjPIywywT4TqSWr3RAqJ0K7
WjlMZzvTnN8Anuocga8AOkFa0AA/pOalJCCCsy9pYiq3bO5ykgcA8EEt1RBY1HNhNQMRvbhnNeDC
Xgb9R/jEkRL/qLgDGuAz2jgQTU56Ftprrp+xv0+cfrUW+/nDxM6f6xnJ5JLCeV7+2Y8y+r/JEmPU
508ZppwAJXRT3JWkXnMVM2XJHl0qb3xxNYu6Vk1NC/og4mYxtsz3mmT7JY4/BWi7gyaguJimetLp
jE7MGDitT3GggcPa23ClN/FBqUjxm/SEGLqiGTQivujQ65gm19h5jSyHyuNBVQG2TgzE9aUXLraR
mIEbgnUvrgChXwKWW2rBd9sLDu3elpvcaTaBhQinZx9HcvKw1SsWqkiJEVxvfMkj1Z5v/ZNCfyrN
5Sx7yRvESHR/tp+yCscE0IfeBKod9k78Z/myYfmSYE+dreXIF+bwFFqYeZLywV3WPfBMSUQrOMO/
X/ZSCmaDOlEBZZzoTJIqM00Y3tpH94rVxyWif4diKhLsDrEo1TW3idjQdabzumCLHb/UQjBTrJtc
G1mQoeW1EhLXhSlKgningE2NaucmtNDZ6DMhXegiwuFZUboLMXpRpsAw/tt4hPSUfiCOjTl9uuTH
0ognSQyBTf2TIdAxdjohBzrUvl9G2rEdDkiQlFBntKEe1KyB8oVkXHyaCXtLZaTmN2A3s48b5vrV
Sbna6mzrHkQn/w8PRUd1MK6By912ErzoY6qYWPCniKQ6z2Lz3higADk69fKiwyZbqnOMaNmizdQq
DGp7OjyW0qPpATUU6ErbasO8owRTWv8RjylEjrk5y7xHerQb3ukNob8fEeL0fJrYv0y53mEwdDxE
kVsdzUUYE/SajXMpG8QsJHxNkbKSDslgFEDIw1oYmlGqA6uFCVnhjR7aur7bpYFGKt35iT/LENeR
rSlQHa8EZ+lCnnFa8fH8WPmgqNqC0uLjoys3MDQbr5Lf14vvq8oyCMWcNw6b9oUd5eQgNC5iSki0
Un7jsEnQ/9RyOVSi6AgjSCHRMEzmKvkdiwSJxOqUG2cwJLiZnuiI00UZWurg0dqP/BPkn6zTcSe5
X8yxV5gv1f9HFgzs6eEWqldBpKJV657aGigLV4Xeid1sao+TDauKw9RqiBHzNLJZOzktHjpybLUi
hEjJq7P8Ty7M6N7oXhf2uDqxFrM6KvGO7cJGUjBeNJC64OSlEt9qm7UIn+sOVp4GGHmGy0b0Ygea
4gh1J0CCkOPulBk+hDGhEqiBOz5/v/D7GqiLRN/ajDp5TEbEbU72fF9h0VfQwgCr5uXS1zjApZpB
RfyXKri5sIsig03qGfk33rQ+Lioo+1/0vP9ZML48ck2LbHrJ+/YB9yV4V1HOfAyKORPy/3BqcCmi
uvcuHU7rDjj62eZ0SHLxmhLxDpLc3DUPv0k0CSPhs/IYULXpOwtG6Ug6g7dtHDTnowd9luNKnIHV
DadxJwPMIe9eJrSNHniCMAOTX1Ft6BJEws24z9zikx+sXL+RQfBWUYZUwbrBiENEo6JXJWQIZHlp
GoDrcW5l5Votkz8z91mrpIQYY9pVxD2bkDgHocGH687o75w8nqH9IQB7C1Bre9ukJICRvpeOunEO
wEY2T8TKxR0yJS5WWwVUpq6/2AwLf6As6gJI11eV6geaeEqKH7qza4mRN+1XeuAZGMaVWdVfoj30
08I9g92AieWK+YCO5vaoXH0alizaT1zT1YPJQXnNK9iNq5naTzkIJT1O7O4rcFaPgN9jWB1r7eC3
TaUahwdiEMOvvfKrljqk1p7SD3hCsxP5Ur+DwCIj+coLI0FE1DHz1DLxNfpW8ibRqcv7KyWT6hKS
RcTfg8v6rd5nocV1j6jq3Ai9uWIavpu1LTRgmqm1hkT+J7ovmIQTl2E/MeYqu3Xdwro60zcCk8yW
wI6N8980zViRBmLFjahCwXphHeg7RBBQXz/b/IZ4vc4Ejp3oC3AipjwNdRqmbQwhDFEQJsvM4yne
J3fQw5CDfdN3EqWaubFDCZx7y8Z06LzGeOhTeT3U61D5DUBM28X1xhZdpQs8vNfiwvdp8ZMwOiDn
vVJu+i2CRugfC6Fn+gUtB8rcVzZI0z1HX9FBKSIKaiXbQbn5A0/PU7owLQDdZdxxt4nGSx28FiML
q++jBNnuMz8LBTUPQ0NHInvgjr2CRBUAncphr5favxLEF/S60Q6XsvdOAZxzlgWMiwMRxMeBEW53
yZlV7JPi3M/zD+OTQX2IS8O+HhTBfKzaY28PoLdcGqe+MUDepAmaGo7o8o6LP+XWvD2I+qHtdEVe
IBja+oQXXSTlhr8AZ22HYgg9YxOQevZ9199yL369Ue8lpuNCUsmjbwNXW6z64iacdvxYG/wetyDi
zswai45gVPARlRlb2tj0QyoKeNXGpywS3lUtcbSiED7f/+Ldr6y8H3vWnNWx15lSE8TU8CiZ1dH9
TfvgrYwGpkSCcsZ09QVifSoHXxKQX1qh2ACRE67qC6TA5LPMjSNtq3Q+UwIghKaVFcuhorCGpV9x
75nzfmjxP5CtFHGuZuDn9OEaAhpTv6uD2XXhM8cA6PvtzQM5du3c7QIDfC18XzUNJ62Lb4KFL8az
rv1qAakZ2Fxr1tG0cFOxtsqIe+r/MyVmk0RNW8d9NvwEO6K5dK/eOMX9P9zGGG38/p6hTGlcYMq0
cS/N0tPYfqH4W5PLy67l0MxfvgqZoyb5JaH3+5rpJGlhcgL3Ssv/+2tibqcgY1alFIvXQ9Sa8BgK
Gf8JKu9VoK8+qgyNVCqmogpqjA3lIQaqiRz1vWOOT36tHmcj9hpNndlptwByHkjXfCFqBCd0YzKS
hKopIISSPHY8STBNvmVp5NcCsgsBKpQrkSDcQVRcFSaPdjSLQIETHIt+2mQ7TXEO0VX4SyakY8r0
TUQnaZXyaDZk59lqeFNEteE59MvV5UPBiiXKfTkcfH764cH1dPPw95g/vWzvHtTGTeF4EbwKqyLB
lK3smLn31pyxBu0EDmc2daAOLAn6zUU5lKnR9C/H6f4WdWxnX8poGbyab+1eUcfq+YQ1GS4cTjZ/
EmqwXb6RwRA/LQbChY4j35CJ4HMtOJmRoCkCrSlrdaV7x2+3HsUroQLE1AYlNvOe9tputBHLX1ec
rmKPVr4BBnJppXddVq0hMddckNBsNIWUgLcfVeg4zNbx1Je4ZqWBHzAPjWTRf3ZWwn9zTxo4Cx+O
d/qzV1o0H82s9Yf1TvGzQgpVMnqzZtrBx5zRDERWKJLJKLsS9/qliD8H1ivfU+OjtbYrasN8gZj5
36/MgnFww3cqeImvztgrgzwbIyxS5curl/qVnExim5LejNHjFL57QBBR7X6gxlHfZdx3E2T4Sc2w
PQlu696nqgABMTSaIMNg9Pfp6FTEQIBel08Mi2rEihE8M0gVIQIVc3+ao0iMmAVSamwHos7KsXW7
tDll6xaV57rGHUiNuaUD2AzNiH4oVWCX4Pqxlf6SzYTvgoPcQs/0S/56qMYSJ7QbJh56c7DuqvE/
3nIKuknWa9N1xtd/r2/eP30jfWf5d98a9WASJJIIpXuYpYph9pHxVubsYPsKp0P0X79Ct3xnskcm
OmjxTD9ZawoU8PoWQ3L4kov6EWZqOo7WOOxzZaK2u3OB+7cbA2klqHFPBsCvevCoQJTA22FhqKiY
R+yJ2TMsO/tRGTm42Lar+5AkV7KzJHiCur2Mrz9d0OWVVjVyfA8i+l+xUDkMxDII05gsJRgXrczD
qJcmsPBc/jv03AMkKY8Vh7XXqEjqy296lefPp4nfub5Fu7sZFEe1yThbIMbtu/KEzBJADrfwNsmk
bH61jjgGmjLb3L2vJRPYtBEeoORKP0YnJO+kAdsySigDi6nxxq5xnAPrJDp79q4g5ayRhuHhwiiG
azwLqH5iTeRkjKvz6n9bPFPI4KfsM5MPvhhAZtzDemu+/nkM3GiuvOTttDWdh6TG0usKoxtW0tFI
Ab7VO46gVItamccNlDq34DqsyWrKcIismt7MQW0obB9whgsUbxQjBm8U9vX1qXjnW6SFWtDdi0km
V6CEoSvS4DIqxHCbL263kfivp5QlPUmtu3PmGaFlmty6bLCdXa8kq6yfm8AarCsinGp69oJx/BFz
3ulszR6op33b4ENOVbq+zKPNXoTqs+l5sXSqcHjFaWPjqbetLvfLADvRAHkzRdcgCHw5VsVf9LIx
ukzAQunzXZGfX6lWrKyQg/1mssv4GElw8eylgU8sdXMS82y2hOlCXV69Uaud5AYZrFBoawzs8ud4
dcKc3XFkbu1uvT2T663ClpE7geJZG0O87eztbByEUx35E9U003iKBLNgzPRH2hyFD1iBN/Ddfawl
cCqEiqFirZWQ4gW3ytCRbHpGjmOd1TdJ9Y2DSlDVcOQCHDXGpF3khOryssgaz/xhKBz6a9TBLM9B
AxXANclQF2+ubtBeN+4NMnsxbrtViuEbshra71Iz0W7u28XkmcLm2uos8SAw7GW2yUUA7RNj6ETL
3Tj2VhzTMmWtLCtNzjfSmhPInvlqOaPVEjmDu0/ejTiiVzZ7mZ/nir/2WMAhw1f3Yw78iE0GTFzw
i3g02NMxPNiU8b64YeJj+0Eyyf62Yw85LLIHfYwX3loF8M6/HJuJToEycNlLalAItnXZqgTgZiPL
8rPeyLLeClj4O8ybBs28q+AaGOQIDx+ZLKDC9fDaWogUK7JkP+bzEe2JzF3E3Z+BzM1oRe17E2TG
3ytVhd0Xp9Q1TbhBCC3YroPqRspMmYpb5fTvytrRF2IJ2/sKKIhBNiId/NFDHJd27mxlV31oDxSZ
tosQ/ZXxO8J4UlyhVxgz/ieS9VOENFw6nIvw1fIabYtkDHgbHVfy7J4MD8CRJWTwvGx3dixw2GJK
xvnsi50OpCHm4mwrVuwQWtW5dErh/jiGd/k/pclRMXfpLDjHL/cGnHWltON8fzF4d1hIN5m2/53/
YUqqXB6TVC6mybKadt1O3Wl7UQRaD4L0Hk4MtVn4kZDMK4nDwnktiqYWt6YZxGjIJXXDOymA1QoS
R9P3D45vrK1d655DRyOuqZaVkG+Pf0xUzvo5fqt/wjSHSD+MJKOKAR2fKusdHlrS6fRaD6a8Icme
2IuHLIexdC8A5oOFq1gh0Xk7JMPYwEOIDO8QJ3axuqmlf55r/ndlD06xnmef0TUCq3StLtU28R9K
4Y3LBGYBccSON4n/I8nLt6c84HCY9MBjhmUVj1PazgoxnFDPCcLCFA2YIv9VPsbwL4txT/hJgquL
q/9Nd6dO9mpGsaDoyrnrlyV6h6rGYenFMVUWx1oaNaoFxfel5RnJFNwMsiw7QMAvbo1EjeJkTKzS
XDxjP8i5FsMmGREmp4wz3WEy/1Ex0ufVrN6ud7UYYgcv2OFs8lrvtShHv5SzyPYYAZpGOhqVYMbX
Xjyk5iIDrGG3AsHV1/70OP3FWC7B/JISBQXtR6K/A5zQoD9rlL/R4Fo/TrPGEj5CntpJBqG1Akck
IfYKbJNbgStAPOzPAdaJ+CWMrTtFjKV7AKDyXQWpdaRYubN/mdUOyb7+Vg0xgKP8W1hbXpyrZisw
QRBkxqCqTxzLFoddcetIs/4jq8p+nmx11Ca/05IrCVfpXIVlZ/42Osi6A88hGRPRjheV7NxXQgGX
V4tTrrSiEEJpBc8B1yYNaWL+Kk1EVcAbpmLvyMpbLpj1I7UwsYVLqULaYbhJFTOu5Y0gjuFoTT8X
W5zZtI5qm6/DkUSnvf9A/KiUzhnHOsIS/g05UgJwUd4mzRu7IyT7K8iW99fk3ozK6gjBqFKyNc23
58EdAO2HmSy4W/Fit2XEB256nEe0WH2IRdQbHAHlJfMm2PT2I4cksY9PBo9ILHF7uiptvR3F6jiS
Eqg0ntgj3+0tJ03bT9+EDO7YjgRLqdcSxKnOozA0o810FvWdSPQYBaJVkLXBabyzgCc9gsHuB37Y
axB1Ub2Y/OFb8AY8y9xqYnMkmpLQqG0TcnlRekjuoqZEqnaqBpx+EAdAsmEC8ds/22ot2J1STSDJ
HV1qvf5CNO6BOS8i/7qaIWHCqnyhuhOQtgEwThN9hOq0DeTImiAk+1LfO79NEaaJxpg6DdSAOcz5
6u+I2RkQgaSzj7r/AK4bV7sLJg2ZrhoKbNT/vztDWOUxYqOnWWWoFWjTgUMxatjtkLAVJH6F769I
MS7wwWz5s8gExUMUpA9H5WJ4JrmANNsaE00viRA7ZhcaDqMJYK+kSufKHI9oovVcAc2S6SrsuD7r
d273tjN3Du/76wfu4erZhf0NQx595Z0NehFgGkJq7Kf5374t0N+d5cNMe2Gf2lrXSExifs0FLPcU
frCdA77TLq69qQqqXOGTztGjv+xW2BgPhWKQMFZzFaKQgCsRSFC+0229tt+1WfgmFgM/1mCQaVP/
BcFPjvQDKl+0Gr2YVADsj/bdayzJ7be+DltGc0WFUbgXshBya+Y/XZuh09rj93DUrxPlFHPUMFFl
7E2gASO/duElK7iKVaAbFAo8yTX8oT+g1wydxI1c9Q4uweVH3n7AiKTm2vW09lNAv8SaE+eViR1b
6M0j3D8Z+07pm3fuCEO7+jtNg4ExXeug76qyvfarFBR47dFw5DTEGsepQ75x9VeDr2McCNo6tEAK
9EsBrGMjo3dqR7JrOfWP61Q9sZXFSRWaoDsZoCLefWM83JeLbinQVdfYNxfuIHtgQ65DNP9LLWsv
qAOJldLouUITpuFdrv0+TkmujNmubaX5Fj1B7Osnq4FeqADX1TkbEkCKHd7c5w+SmpAyuxDmcNmu
v84p9pn3QF2GXuVM0Bz7dq29breZf56YV4CSMq5LZnDpCdtzh9Cggqm4PXBfJBaOfuY7c3KicejX
/rWVpuXQ15KQOq2aWq2klF19BCPrAu+L9lJDBuWlHWKodPAP1KqtgTgNlZ3ygRxKSS8PXeWkfl6C
pDQ6UgYFEimg7QzO5CH4g6ksp332d48YG/pkzvNBnmRl/B46+HgR6/Ilyqllz67sKtl0L51+NqYV
FpBidYdBuLhsknzJ7psF/V4P+70X5MEJrLti9c9omKpQYJzZsmIHAi16mJF/HxHaE9wXqn9s7FTZ
dMl3MjFv5FWgVgOAjjaNkGP3KPB92CUnGftHFnI4SUaikvn1aDNsUxZQR8QTll/4oTqE82uxobF4
gVJ7Ep2skBtKpMvGiXpL6FBgdGusC3tg7G98MjoFQI7QV739t1m94s3ZcPFCV6zjTAVwm71h+v9N
YQxllGOJ9mXGz7VjEZRUvYwQIU839LY783L1lO6V41gbOGQKnHz2vbMX6l/WR+0/s5HdkqDqQIrw
0a9iLeOmqMUqhv1qPa14x1plkBxrgrXwHA3JbX8vxhVCopOIv1LY2+T80nUrvBJa6mC9CzsNX/rJ
D14fj/x7zLcwb5qUlfT6WO2Tb53MYmxK2NAinhLDGn1Gl4LTYLGW/CKkBGLwpF0L0veM8lRdWhky
v009FDaOUbVopSeYkt72QWj7Xo+OBKb6xm6bJc9a+A8svdL8vLNuLO8x+iqmu/4mR4sj+ebW/cL5
R5xumgpbKTq8SZ7qTDX29f3LDbNuWz2NutBk8RUuCfheeCwaI3En4BfAQ5IFyRunAc0iobtMaeD7
0DSUkaQ10bHJnpyeJ24pvqaxKp8XeK5kDewi7376FyLBv+WLvY3v8BqZX1SbrHKgShPR/AYoWLPE
hVQ9Tordz48nVAuiXf9LSAu319d4fkv5sFD6dOtvdFtAKSma8ErKO0zOPlmfgHw9TawGUUocnb9s
zZf42enLmvwqRgdAxdduIbHsoA44++c3UrQLr5TlrsIL107IQfyI94bn40E+BdP6US0uV1dlfPco
52fYq4R3Kc3c0SOW8vJ6sw+WY5XVDkWY9Dgzut+bzzgvusO4x+Wl2YiPmD5noQEvIFuPVhpP+z16
ppXqeG0V25GngmrlRTw1a7A2pwiPMkrSKxQBDng/U4gIRz154xs8Vw2pH+aUaF7sLhtRvH4AXSRd
8hI3VtmDatO5hgWo3XaYii7p+KRL8amCW8S5KQrnHYRNMmrKlUaVkPqZT8o6rl/QfYzNfBlRpfrS
YO43wj1xeRD3BzOD4qqS8N/AHCR+LLPv3eA8pe+wewyLu58xMnfyZxzGV0Y3y2zQGjaxNCx8o8iJ
MwdFFFMkcty07AzE139WfC1KzSUfBwak40ZClR8mpzlcF+w0d8RXwLLPYkxfHtVesk0JgGJgo+ze
tEZF6M1MdweVZX9AX2R/Oodv9O8xQ1mal8jjnXs+IzVvWPWz0qd0EI4qThk7USLOHKA7E/CaaXj8
9gQdF/7avEps2AzblVxUv+pyeEVdiemoRP/McEXeg0zqR8l1NyrJu2728rT+e5KfN0JxeHBcCxvN
rLfbnYcjhD961FH676sAWO0/9HRNr7gc+f8lkMnOMnIs/yS6ADXqBJGvRmJW9IimlL6CZbyw1g+L
ThQnnxaZcTkGwT3hPRVTMIqqRc8BRCH6oA6bIsEewrEZnYyyxKogzDEXZhATdxSoSuANyaIgUCSy
Ec+EpPYYINIa9EfKe8ajFQZ5wZC+cW5VWr45HE8kkEFTw7pgCUpq38v7csPXmqwa65R4+Rl3m5Vt
hr8MChz9B2wUYfbMq0zn4+ivJ0h+BS65JOCQneZlV2xSkFd38660dk7ZYCxTQKBO8X5o6LQ2X1wd
rxH3VKd5OFD5CV+TTlBMz9d+nGNy/n+nQjWAeQBpvbEXsyqHgZ1ykeXx0WEQqdEYuW4t86SpxrBJ
us/Z1RMnueCqw2HnDP4VdMGhswr+2w7XFnRW5tQzTpc4s+3XO+X2z9R2UOXVIAyhTIz56RbugMs7
WuRHBfYCxHdqNfqBed161EljzUK5oRKVDGBMQvpGDX6At+A0aVtfLh/Tns/1ZVSQZo77Amv5TrR/
vU8vZTV6M0sm1Mcr/YFm1QPXYfuZwc4VtivXCNbN3xFLQb0fOjwDIWAyh6aNCR6N29aA+wo8m71+
2DKV/R4e0LgB1ifTlk/LpVogIhpDBZGxCcFIh9yrDCAQtiyIN5Yze7mDV/1lKmJg7CN4U6lAB1MU
LmeXb0Y9AReQgy8mMOBu4hUsVnTdANVnDQpPjaNDwuRsul/5g7MKJqe6M+p9S61de3WvRTlZ4PRd
99y8SR8Tkx+ZsriVW+ROwOYboKvzhh4qiVIvXSJbeTFF1N9idCbBPpQ8RPU6l4zU+H/9mSjWRUd1
AagewQsEDUP6+IMJ+u2wDUIeeXGg3hTdBX/2lMZhPEMQbwkQCW06TJ5yCRlKt6ZWaYqftrMlj98f
NfsvWUKi4dKsyCnDC52Ii2KSVx3Qfv6c+q4HeJFfXE/dQ2hcJsbOoLW6Cgcu9rQafFtaVU6aZyrU
LuPFCowavrIJ7Utt+PYMi48KBHhtsKlgWFuxFHo6/KhI94klq+y/Vp2sGGMeQ3CCeGehv4FUKZ8n
p6/rSMgPuWf79qm9C4YPP35l86hJdJgGCyeLuZzA+dXIRzvvsGj2fBuzvXi9rYb1FvDSHolzFzFD
i8U4BlnHc+9K7pvymNf7BaRt2VC0Ei/BM0sDhuKO3bE+d7BvvjE1gbIhzxnbVlYGAoc/ZXilN20f
LoF2JztfyyP2VruAnXtJiv6xcmXJZDl8OahY9u3xYkISRQvXXcFjFgmZVtfMKcBmxX3I1cUehq/s
BBW7k8rTVqTngXGhZ6eIrcsPvT/9Um45j3dlK7l7gQb4Mj4d8bG0mx9uw76EECZoPTicOOahEIPf
hZxHK13O7t5Ql8nE4Y6Wi1GUSIs1s2eE42ZMHVsQS4hi0G5V7GEjPJQ470XPvHmAmLBGbN2U3C0F
KK/G9scQkht+X798Qro6/D2tDn9Ffk3VFhsf7FERiNjHnbyUZWFlXOEF5dfTgcfLShEOCooNm6eo
fMqRbgAA4o2PteQkRYd2tlDYJapOVQmoLOunu2vmvUJWvK8PjsKX7QTd6u9ailv8Lw/WXYcwEmDi
yRi1l4Ma7S5Kzwx7/QdV408rFi9zHVlQlqmvOpln9oOw2YK0aKjyCdVeM4TbIDMwRjoOKS9Dtl5v
qh6uAfNg0rbRijhO0FApbMIpEIg1iaEP3Xx419mzCy/N5HAwCvYqGxWi2e/vYPY5MZV8NFXNoeIU
I1OWD0AoemzhoMtVzTMJYM8Lg5wJNvEh/mLRcQRAVtKabi5kpdFtbm5RmSQPttMIl3c0iM/J6GN8
RmpLc3tlNtzG+O10J3uT3BkNRY3f1dU1IFuij45KsBOaX6Wkf8inI6yvw1zAl845gorgpNzKc0VU
p7Z0vXKc6dTypRO3fYSCxVe7ACApre1WSP3EqmtISHnawJz9RizNw9ggf4e5HezxigMUv5DTsz/h
aTwZNG2rOJLAQDbz9DQMpc22keJIeLiIy4AZg01TglW4um3DUKkFesNrAfHn6o9yyO+o61NldJPF
Soc2+FwCJGHRkjNxiEcgNDhWZxLTYYbXoA1K0gRHJioBrD1iijoOecCKcO7tWqgeKpBxYMT5871L
RKHqq830V/tE2vxTwvRBOoafsOzjEhBW6yJtQhk2TyZnN5kMub9sGJ+1WW/IrXojnNjJNH7r0d+e
E5PdHl1pFVYN1L7qzTkqgCgn31m0YLWIQioFfw4vE7TQRI8Oab2Cnv43VeloS0aCiEXuUZdxf619
8+i5RZDI+pWyyaeSP6milXI0vmrLqJpiR+Nga0KbvP1KnG07SNmffeGqHfJQJ4Vu4fq0bRkYQMhl
oLjM8lajEPlnHyF25xPLoDg/+R6ZYNgNmaYRsJeQ5ySlbXoLaaA1xoLFNJpZXu0bxraUz2jTQlna
VyUkChvfSoNCSvvJZssD/vjtkdB5hrPeQE6bz5PK/bPtIVVYHqHO/RXG7eLAkJeciE6YerpuLD/1
Ck3VvM4sggGhwoHuMtv6M/JfYuZG40+r/OC4wBtAP+dFkIDEnHqREit9VnNcU3Qopo4FenYkxc6U
EV3TsTEoX//7EkOx+YUhTnnLhClMWHLMdO3EfmIcwWoYCIAWbOdMzl1sv0WgRO2c//9YuYy5Bn8E
/VSlhVGx++gy9My1okgmYebch1Ye5HFmQJKtDpVNdGfX0LURhuxnEPOfCr5D0B77SZGncZ+Gt1ZU
hT4milxXRnsBEt8zcsG7O5yINNTSheSQAPkQVO4U8lXtXG1WqzpcZGV8Fd54K2eIy0GB33kjGt0P
+iv7Y3Yp0xAzzI4f2nvkHuehqDu4aq1vtd0grJI4n7XK7z9xiuUGi2I4dROSXGXGw+5ulLiLkr6p
Ojjw0Qe8UEwWgWUE4VmF8ODaAXeDVdiV4I3MyDZKtO4m29gyKw0HPw4KFQk0CAW3fJhlYC5U2rfs
+O9IME1yyA/oCmE5GbZWtF1WSLILnSgJ5B/5zLDHZYeR8HbN+PX5MRX+3Kv46SrMKG+msZyHxyl2
K/WQMxrT5OFZleR2VwFpngy+H2ayS/JJy4ogh3vLfQpbAe9WyIHeh0uTz/WTWz7vqa0/0fZr2Ghq
6r8v13y+kuqa42Kez0NyEcsBFjVhmAI7zHQcgkHTtpVwfOY+Jn6is5W14VTMQtvV6irAqeTngte7
fIWaT0M0PXowHNyY+EoIM7At/8vYnq3ioFCk0J5N3jaJYqPT/apmePEn21RyHLVymH3TLoU7c0Q4
yCv7t0t+/7YsrtjGHYIKDugpkJKDObbwxQSbrTgbg06D/Hsdy4I3um2OCA5Hoo1P6KZLTp/V+g/I
0x3HP16FVZbfj51/ViH4nCO1DX7E5X+dGQMGI/wXgd4eOfFBXDwY+5v7hMKHpsP/PjBjYC8r9AnD
AHfrYhsph67GZcfIUR4+VAn0e9jG3xz2/+dfN7BgYttVvRrGfGtZq3k8DWpBOhXhl8L2eoJnjhQZ
duf5/s4bb1WPzW4jZCtE64HIT94DskyUpS/wdOt053z5OsEcSE+S1vBo6YCsuWpW72DuuZz3/3dZ
tUxjEXCaE0FfhJpxKETf9FIEyWEvesezGLD/uDPG8vaHxsQIZB+wrFtVN/bmDXpIjdDCir4eg88B
Loot4Vff0aQfJ/3GRZzxynURO2YGe0KX7DVsAzGrz3ALAZ9IGegcFgbWqIhK+7oMfu4qwG7BBWU5
ClWeSSvl57eQkcGbWYkyb3LN27uq31mmQ/j9uQkJmp7g/4DeMx7K0mCWzv+Joj+zkqVgtLVZ2IgW
yl86YR+5BoDGBpQUM1JvtDGBuFAcJqzrKS8S0VkGfqCzMtdZWKl+zAV7MwcpgRI74e4HO5y6sTie
9R5azQsJ47E73YCrVhNSK/8mAOEl7PjjzEK4wVSw3/ehDjORQNY4COOH7qCj2cdDMR3BhUGkgWCD
edRb3CyQyp2mEbP4CiMjDoXyPipbK7qE+GZxc5ez+Omye8vbpsMd36mliqdmXXTrkYpsLCRoohVa
l+OkDfuZrXo0wGy2an4u+gjwW0cPDo+LPcZmAR6ae9Budifn3dsvziOicucTilIIHXXhRcmF7Aq+
7ieEwt3CVzXhorabA0jOtUaDg0WdutHJmFiHarxZeVdgROR0JasvDmlYLpkx1EHnnnIOzyJP7dkL
cXm04It1f9FBri4kyJsh3A4feYAnTyt25jnKArJQ72T2QC4WIeT2BV8BFbp4+d90m0lpfRcYZZVl
zBn9vT5EKloCGxS1yQH9RzrtZV836+BHTfV85Qzo9uGSyi6YSoSRD7ec/G5ablIbNaP3yCvQw7sm
RqLts4NDPztW7kdO4bxtJOAyHtAM65C8CjrFwZA8nAzeqBe4M0Iaon9bdwbcQtkv2C1vFILmgoA8
nfEaawBDb9Q/c/CQTnPxUZ9iqmY3W8qw1ARPaGuWUNzvE+bSzSUxt4L5I5aOheq+U1bKTNKTkJQz
6cFu3O9Ua2KVQiDqpRlzbW++Lzcdzhl7/luIueX0dv+xMqsQW5KnK323J0OoGAkH9d8GICiTFz0g
8W5HDkTuLdWs+Q3JuWkfknczkQaIh1OzMe13PTYwjGHOlnG/LAm9iEPZ0TI/9pGZ9ggtF2/o/F+X
l5cRRM3ZgT+3HO1s34ZCdYJHSlVpIjSRaZMnEPv42s2jB/u6EtOHm0PopgnBER1uJ0jvWb/LJxhy
jnEEzGf0bUtPfDm05ZipmaUe7XhTOBs1R0J0Vcgd0byq7jUnAjg7NchwPQ8lvex+PQ4W3MhkMnjq
p8MgTask09pfB8IknFJyTsKGPA50kKnOlzEKb+wWkONJzhPnEoFBU69NdTgtwltJQ0DLO8uIkC/i
fLjYk1aH5tHc6SL2JO5lyOjjlRhZQWtP+pEUX3yJdNEcY8v/FAOyB2+A9UnsVw7uXn0V6All3IUC
Gig9+xOFUY98u6IBTWiAusnFVCROBy1ilr+Z2qKMZnfV0pVrD+JBDxS4w7qxajwU/JxvOBu92Y9e
fyyZgDDC+ot/7sHtB84DfthyXGV0SSLO++LQihJ8oEN+nxFT3N+Z5EfidRRSfGNajhZ6XqpjuXCA
6P9IaoRwU/gm2nCnmqz4AnBOmPq6oXAn8YucVU0SAZfbZEuNQD1XB/ECDzpv/QxsjRwNEAo5kh/P
ErKRLAzrPfBwe4zRwueSLZ/zubhirH3YPdox4S8+WPXV6DtvwHAPHs4b00M/XuvFbJwtg10oI3G/
W2g+E9gzLeQT7JR78b7F05mGGkpAGekBe+VQBJ6ZUPsylrR3IpcqadldmD7EdeXZxFVbzzwx7nzn
MbDbztJ7ko5uwqZBxpfiM/z+r/tDhME3drT63Iqbt2HDv2E2UwsvrFzSmiqK/l1KoGXc8bg7krzl
WRd4gStAEi1PsSFED8FCfFtTY6MwY0yk177DObpuw2bowqqiW4ePM0N+mSOckwTW2sDcYlQidM2F
2CytqrpeU3RSYdj3SRGJlVUje7r96JGKrcmRz+elebQLP5S1VveRTtICQrTLdw1S5yGfUGvlC65/
Jf/G47EdRKtBv8hNRkOWLC7IrYCoKIXS/+4j/7IhQFYuPl5CHjXztBDeGrZM4yvzHPSGBTe4f7Cc
InF/qkZDFM9IMMf+er+ucQduCBKTamGYotKz4st92Iwze0hnqfsvFhDY0r93OfhrYSZxh9Zzaki3
HzgoVlKg7Dh6vG0rWftLCPZg2NTsNA2zVXhGK/iKRNjkDdtaqA9ajayCEpOVKcTOmkhqRGkI32mu
JROGeWzKW91C6mC5ZSjqgdAZWMoOG3Rq9PuLQKabuLq4C82SuMh/cjtOawBr04VH2iXG7ob5AW1O
gHBN+zBL6zu2if0iWTRItz8jNSrn7pBZxoA19c11OKsnrp+Xd4pa3pnyzMd3hga08Vk4iegl6i7F
8Jj5PGIUmDpQleOVSIE8I8U9KfFa6h6SCxJgtmLX0k5ALgzwCJ8WerBFlZgP33UhVaseGQxFVE/R
+3dkFQeP+4Y4q8dhpcL9t6M7lfwNu6Pb2vgMooklEkSioyiSaUFihIrtP++s+R5K5k/Nkqde3tGZ
BexJxuZFFzLXpUvEeQlLCavYR19wmnbRf+fixmZybkOZNYY86RGh6c5xv2TDWxJ63J9b9J9d3A1e
rzoesKFekl+ll22FxSR0cOIsRhV/i26hr0YbZaIc/43qXJvtdzAphJj4YE/5di1Buz23L1t0PZNL
/iA9eYCb2NBvwwLdrgLANJQd5mblAJ14hXVQpMmlEt89QUmaaijksGmBMtwK/EX+nXq1ehs6dIFp
hmbYL+F+jjAseXTBdNxQ9qBpV8143RgrnSROui9/xSD8Y39TKzAVZsgs8ZEcujizMLAITTMZwPtF
stblpkv9Ayme0qlpyPjtcy3HsBNbKKO+hQ2CVy1RtCllg6CmU9pla5McM2A2jzQiU0vRmB2A9ZcE
qWic0+Zew1581DtNwbS4tUT/RfDBxdHoCWzharmPsHSyK94mzq/aoZn4iiUTaAF5XUD7KQZIfue/
8KcCTZrOBkN/UtsI5eTddwtDnyvc4jgw5HGXb3JSDkwttPu+kH/ov8ZEMJw2WatweEjOB1kSrg6Y
hrr3Wj+KYrkgGjN0r8cLlmweSftkpE1JZTUTaeizFxsR9LAoH92FW5HdkTf1P1691GPVqlmJKYUQ
jVcjQLDlZ7g6v3XXnvN9O8bXpRnWg/S4JB3eggZY0btY9NMuV6pInMN6ka3nztZgI5dqfx6CGzXr
docXpH6Dfo1RgTfw7QbcPhoCzqm88joZwWg74FnPwU6SAsJx9zS01u/5XqoaWzhHP8/y/L7bKRcI
nj6gnw3ypRfcjoMZChrLMymWkUTZ9KGP8FiKFxI3om2i2bE0Wgr5ob/sZDvyvTFnUT61UEH08tWR
QX7gLjmqvDuRP/lXbw66cUI8xVGjs2AyPELPyyRSVmFcFbhUzK3GmG6JpcREjW+D3+NsEzJv6BRx
bFqXvQnJtLxfSkXE3CWJEGxAeMyqDcVyXf9CkH3tVTAHB7SDJiCTDLKG4cTtOjhf0YaQckEZPSSI
8klWrEMieg5Bw/5966OjIGMhUTUEDB5KE1ay1GzvI0GuK4qP8FKRH7iXC14lmabIezA10foJJbXp
gwJ+VzLBm84FplWgBhTNkUi6c4zmXtEUwM77YRHJDBiQ9AVcz3wmyZM8buBHVkeivZt95BD67DCs
/gmmX3lZ8lxSSfhgOtL2HB8mWteJCJJNJ/7ASdp/nvVBwsNhfuCoeTZC31itXoiMMNmQk7FKFO/f
ns5/sbFomNh9/jVtT+dqupYD6gElZ7MFT3t26pzYMw+7o+ObuuGMj9mWAJXUK1uekYbaSY3Xxt2p
0uCv7Ic55npR2rxqWN8vD+/+pvR1H06NQ21jB4UKLHIioRX44xP1RO7pzy4Rpvk5zVblfZ+Wjs6J
09KBWh2HKRiJOBHm3m/qJXFXFeawlhXHyGBDBBhIlCEHL+sZId3KW7qrH0obHF6cv2A3l9A7kL3Q
oQr4Eupx3p543vwjkeu1S2TRwc4P/QpgA6qGF+H0ZnqZ+6vOdnIWgu54vbEbuL3Z5uRS2bH1GOkY
SGjbHkB4QAHLPgA57mnaiIBNnzERPxABebjYB+Av+9bIQxqHNOyS188t/Xru3k2CToyegaNtWC/u
0Jh4lWw2d9n1tkYb+Sw77MxXqo3EqSeJOOt0DYZpm2j45pwBvRYxb2MTuKrL4ltsqPDAzgd1x2M6
nLcVMFusO2YKOIZ+UlAh79uTfMoa4/6guT+TD/5Dfeq5XHXVtsTy3SCZoetQ53YNvk2CZfDqgIhn
uD5pwu3AvIHJEygW7VE/QAb/pmjy6TTqMO9RURQ4/YAm/Gh29yGgOXe9daoarNUdTaZ3aVUC856/
f4GVLiE3YJyfBu6Jl43q03XLUh3VCAeBy8VWP7kr9kgt4r3FMGbOCzR23zlAyxTD1n40R/2CnU/U
HpawmjezCEplvc77oEmEj4EhE5AFksAM83KUUzflUbJl9xSRQTQz8n7DYU3Lxf0KXOszvUyOyHH5
GM/RBcjbqgzDJejkhnUMPMVWYfKhADQrG0xmq6gaqo47/qlH9L0K/vT2SvVSvtqBKWFV7O34h0w0
vOqErTsqaAd6B4TXvvinqUX5RK1yp8YcCVVYbXNWA8Irs99idJ8gJ0JRBXCJqw0uxGa7dK+Eqr6a
3Zb6dT6UraNdRU3WcyCzWumSBit+JzATCGZUhqY6c02M+tCMOZdr79jUvieLKIteNPQDd18=
`protect end_protected

