library ieee;
use ieee.std_logic_1164.all;
package processor_1x1x32_Type_Package is -- 
  -- 
end package;
