

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UTmxs0OkmJURXBOVdUGR7t0vPgcBU0oVnrXWTlGh9ogLy+aZVadnSNImcgn+4jLE3/0AXAxZXQ82
Xbw5u5ikwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NDHq9z13OnSHCjB5ixLI6v+O9siiJNJuJRP5KO7VWFUgsdEdfLm2msHdSHMZWHSOwKZ3fpyDnmNx
BgNrMCYycBeI/rO2pKL2N4HQAMnhKOZtiPFF9n2RUplezsx3A1KtfrZPlHnD/UnZMT1dsl6klarx
WHWoOj2BdFWF78jqP/k=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pd1c/MzUc/ohRsjBZ9c2FYMEVEx0/T+c02CO5nj1hjCkjBTD1iExW4b2fGAqq2hXvApptvjN3kao
diEYImrFYF0oK+4fJDQ0NDCFSHEPkV9IuYgpAy5fNfC1Dx9rVAZAI1tVIUXAIZsy7oaGc/ReA3s3
/Ev1+YSM6X62ouq0EXc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ds2lszdMaBUWm49P9ovDqEJCNyznNiiJV1s10TsqQV85Goa2s6Y0q2oK0nkUurPC2r1U/lFQ6UkY
FyQj83Ie6eOpnawKkK55JF60SUgc/KJzJ7bDwIpaZjrpb+XlrqrzZU73J8jBBHKLoF1/Njgvn5Ad
h9N2MGH8gaas+uT9uDuZCA+ii46LQ3K2yd1YWXKK4uzoENDnOnWVcV9omYQiZt2WoMmuDtnHiiD6
BU9fNvTDJc2E+yqoRZLq/i7Vp6O2raEB1EabQzrK+1rVqoRBidd5D+df98jf+SVXW4uK81yOCvMA
LOV3/ZU0qCRQoJbwjKLC39h49ly0sWjEpfW/gQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
df0vCAvcFSWs5BffbtXlfaFIBd83+wey54D1uX3YAx267SlsUp8LU636/ulbSzkGShRGyHAsajTQ
lak4/g7ql/uNS4cPDTprvz1MsadnxOACDABIUOl7lg4w0zjMlnHliJydcn6lPMrRHgqJ6QJh1Ypj
8in4rFzqjprqSxw1d/10YsZZxkQoba/tmtftne+6yGg56W2Fvkku/OTLhJ4+2k81Et3P6Hl8rQs8
H3zDC5jgcWutFMz9ATChQpuoW1Bt6ol0u96wp5xiZl1ORv7DkneMNq66FiXR7uQAikRnfSIiT6/5
QAjuFDJ9beaONJ/7PX0YKv+VUGzRFq0ZFYEUEQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nCZ8D9A90hmHjnYoY13nJu1ipj+rg1ZVc4+qcqLwK/I4sVkFzYXzOHfQZXQ7YKW8qcQwr7Ja8l+y
rmS/aej2Bl+/GBm2e8OPwXjYQfJZAcWrX3bukYUhs960X48k+oy8IM2fpLqIO5UjCHWUKDAmMH8s
veeZjDOkDvXS6zx4x9hZL9OB3MW0oK6L//tk4UtxPcVZEJmBR7mpHfQdetJlD12R2NEAOMEs9GYi
egJoRgy2DcxVo/qhMUxikMoNK8DRbPimHxnf/gi8Ss6Awc1pw8Haokg7dho4WvcGQs5jULvRh435
wbmLZ1FnvnxhHSbLJwY8aBTSiBsD5Jozey23DQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504800)
`protect data_block
yscLJS8Qa5Twf06eCa/udQTyUp11/7Y4Rzi+yMEEPkPYjthSybsKjIAurIWQSujo2Y3CRrPB5xDH
B1iHTz1tj6ivacFivtigI9ro488ar8qyjb7GCd0+jdk0gE65G4ZbeNUEQsKt7L/dH9/0ZXhoApCt
9O/80lK0hq1BtBjPj0EGEEzWFWLlVPdJ6R4GjI7A5oo2AvZUG39MdjqE5Gik1fjk8qaBaYR1JqgH
GA0/qYnU/BVU8xipxESY5IMXfEfwsIhfuc7oh0GVx1Ab/dNeeG5IQZ4AkGG6k6yon0ASniGx+Den
AuU8cPiluXp1z9Q21BhacQ5ju1AAaLb/+XvYxtvH8pVyxzDGG1l1L3rcqQufTz0C98r7il61Ni26
JaIa/EOtGllcrIxyW/B8IByVHb5wI3FCWOiEbm2r9L4c0V7w3mwNmjMwsxr/BED4xvatK10shcbq
hLSQBW5lo1iGn0ZYyWtAeA8HXxUJLq137x+fb8V9KdG/zkaZrJOm++gB03puBo0AO3FhRLcu30LD
kWZiwWs2JdeG9sKZdgRsqyDcram6zt1qTQmObVggkF9K7SbXaCc7Y/+IYEBSQbMIMu+ACR3k3aos
dRH26so0qAqfAp7+MWf221io/As517TKnGGPE6DtL8QPl1U9urZUqBfKSQwgtMjSNRudPcxdQEId
kHCccsYbjmAjNxAfeDR3GXBRiZX6oiokHjEgmsbslQYQbob2WJccRb2WOrVJ5FtKIbXR7cj9sqxL
ymYctQvnfT8amVhh2Ig0rsP6irW2mn3rRC5YNw9rxUGVJJCwwnNlZbKfS1O+D2hp3O1GsYM6SXxC
fsNVW4W++eFU1bwQJhmlCzY2ZPzP1AzqhbnmXEq25wHe74c/+DM9rrhYJJkfcHUkwD44nvZAB0lK
0DKDj2xxwr4GTM7PnDJAxCW4XDRx6FUZBPeaItp1F67nhuA7SxrLYRJR34WK+Wi6ZmYUiZ5aJ7Ew
hvvWmct9h3aA7QjQl/afKmYdBU4zCoPdldAfkKRw+FsBTS80xLvl7chhr9MmdQ3jIqkc8woRM1kC
OKSuZ/m3NqMVCHIb5dE7CtxQ9y/cM1XD14uTdNlKxTLwU+yOVUCynK2KlQPPZRIINiZlEaS+fX1z
QWykJaj0owIM5LjHiO9m8hL589WkimyQqgF6xuBHwo+pNh19GW+XSfhAI/uWclnAgzFYxr26434D
X3x7vllxrp/ZbGL9tvQXxaGtDXoqRdSidtT9x+f8CYw6jlyyJSB/lJeKAbFFYDMgLYAGD4+xVfmQ
zcCdn4PG9SNTFl4ujSLrzGA5FETSCt0vyG6kyKBVtoWvRHXHIF9tDT0dsGzytL9w0AUf/deuuoC/
3Sgw3Pg4x3XEkYZQq7z85o7zrY7ebOLbB2TCcODPoou97BkBW7EGgz2olX2Tht3upMLiXOO1ULWi
OpzBZU3Zpm+iwsByblvWzoTIxX2HagYlI5g8PtNBs//Ptwb4NRZulTbOA5Jjc6PO1pL4JN/RSO30
M3pqe1ojJ9sAUfY6GJzg1DbKEY7rdhFnJHlJpx11UCx2qX6/W1dnl2E6ScKjrRkwrRZ5wToFk5Es
+nLumVwl8lh0ZL8lEkjsRGj5Foo8mlcv6PoJi/jHhhVWDVqhSno3AHnwrd922I9uQrC205VCrj83
rD/BKjGUHXCW+CuK7PtoGyTOJPqDw8lfLYvMB9W14NDi69x8BOAzk34ocMgL4jpJuRGdFjoPPjh3
NuBBPgEGGmiOUR90RYuPmjqz4Q8AVfZ3txW1LK5PxdF5LvJ1aJktVAhsXjHHRj3rmEEL3K0fJt7P
bPaLl2qIhS80ZB20rnHW8n+obyEb96mfaE/i+/tp01zeZ6SPjO1xTnGShNuhspqG6bYw+u8A73Lx
AHHa7n0CfBqQnBuGCViaMMfpB34oAkG2q914bO/Rc35mUqvjJlL3k8hXaGK+4ZRP4fI8Ag3TRkaS
unn+uQj+iZ//foK0YxOFRf80vdUyo1GJfQXRJ0P4X1ug9Y00DLEWhgQnbXdH0lZUaAUmSqCR+7b4
hhIJLfmHffzcLETecHJ/IZjxTEKwHhzSjgwyRmkwC8SLcfELXcrjSwC/LCHi+zhzPfCFQbyquL8/
MdW21vVqOLsYDHJjdXqO4P0cCz3829RE8Ys4frTOcRC2ESY9PY3VAUaRGckMifwOpiVIJXbgEiTv
I04TgPrh99zM30CAEMg5OE9r3/ohRAaKAP1c1fEKkNparOiLgMUBX7Uh3dRo4YfC+QFHkyr5FLiL
tFDBrQMoIvNqeqCsy3AsWavoGekZeVAQlBJlggKhY6xK+cotAsP4qvSXhDv4X2KzDXY1awhhf5f/
Q4PmIu9J8BBqHNwtj/TmmNMDEe9fJjD1jyspVjgzq+efOQYpDE1UplAdZkRFzJVQMbpHV2JtEvi7
qU+r4maMJGdomrrI/N6QChnnJMOm4oyIjg7fp0/4Mo8F7jH6ogGgTpFDzbPtRh5TzvFNyBF2zxWs
c+uDWhgF7znLLxClHKjPiA/WGPUDe7sRtOCQkfzKrNePO4iHDuYw2mGIHnK40GUnDo6Kio6X1+y6
6aFyka6rsxwNAXEP6hVRG7uv2frD+ExdP3LLRBuKh6XDUfGrVQ0W0Qav7VzjdsouzcTQ6XJNQ11K
VS6E5Ej9m3wi1BLcy3tM5+xiVGscSCXfbFp5weFGSUIS6QlV7SqoUfroyqu+mVHFUsyQ458KcUcj
RHod3mR+AFonsxBUYZd7fjZqUhLiI0JzGATz711QP7dHb34a1RJXt1v+WoaGgaPRJDeYFu6PhME/
xAVTa7lWV6muushNibI/BwJ3JjDEbIAOswBKeaZsAZvVBHE6ykStu8FMUfNmck+JONvBFMBmBxFK
/+XISKdNItXRJrWajMgV0AR7B1QYY/NDlPtvoW9bj4hXu/hQKVd/wX2KjtCFhCrjCp3O27oXBAg2
+EXwSxJ5MsA+/9POLRuuh+h8sJY/Sc7apj1oijI6OTFAcSTDtrpfiMsd/edh0xMlkD4AZd+O1py7
SFKL4V8giG5lTmpEm1QPaF/E00bJiPAv3rK6RD3u4MTkQ+Uvc3xUxEiRmZ9V9KK80DjE0LcN2254
o9ednX0007c6XCTCmvMfEpmnw7gMdYyl9tW79bm2t7Fo12NLV294lzpFQkIknD2bERfXKk8YXzlO
ik5ys2Dzemq2dap7BoAyLOF/0mzDo+RHNFe3vSr2dXgyG53xZCLrHPlMFeHheWnA9W4k63fYqLcy
J2I1i1Crl38TUzC9syCjs4QjFemPk9Wl33IkGA27rCGvK1qyhbXCwsLf9wspFAPBKJo897xCURfr
VLPYgK5gmk99zog5+2zM2jJc7IlVQDGAJzTgla3vkTpZOXs0bzqpM2gGnqSpkCGGk1PPwsqXAkFA
DmgN7oONRXF1+gUsjVs+hg8jPZgb6m4l4fFnCMlMQxl21jqXU8rxyr7c2rtMwb5BDGb7Vgar8yzG
BUEtpgK+rdeOYnLOdODNJ3D6esJX6aM5+sthckgmUisTUAv9K0WuSFlUSA4JiWnDrpP8ukESaurJ
G/of12ZI68XOZk/UYe3uzHw1BT758LALkm1g7tttsBP8/ICqIETV5BD45uQSjYWVSZegP0fcb9Dk
9VkqcfNsdNuLcR+PCA8YB+mkDX07mLmOeVOIyTxCxNHkfw/xEi8t//o8klqWAz7ApSEQcT+VaveA
lVrExmHkeZep7w93UwTBkxa4pvA+cjmyDqg8pa6SgRsOodEoX0eGCGIhUEy8yJBQo6pzEHqdnorj
jaJLREQ+h63buuSmyuLFcDTIRemWboRor58zXZQmmLW/AhCp4up9iofvja7e7epqV8h5ECxB2FWm
fPVgfwRyXDRQPjBA3Uip8lSUAknBSitmMQnrCPi76tnaJz60FE7dsLH0TYgoIuKb0JUlB4XHw9+o
ytrz+xKoAy1vTTzbmEDtsiohvmtVIMwaKEJYkQ8oMHYKFQlTVASwiUcVoDaY0yTSBPR2w385UyPp
pclXwwJGmDVjaAJnhKatZ6cGpdobL73OiANpyGDsB8DH2V32qdt0YfCxeU3JsXhY2kEJKFXp5uei
ag+So5u8KZjJ+NS5D6MQN19d3Ej52++a7VCIvTXlvT6Cey45DfxjDFKsmPNZK0VF7Q781xqwslr2
gCaJyf7Q9Qem9ChgGV3R0k4Uxe7byCdt+XeqDRdsT62/sy5fwxYHloyU4ebHLNjVEqnIvxDwzaZc
joJLMt4VSPu5/AGZmYP362D4PNP5tsQrxEEp1mUFmOu4O4U6Ecai3EuphxGxQjiZFrriIulqLKge
NRgCeAkvfGweuTO8vuh2Kni77ALq47ADRyf3ROdmVSkLf2odGBQswcfLtpikh6ekFwXLX6lNNX+Q
DOA/ouZjl1lT9Ktn/P5tOkR7H8Joy3/nrN22yHHC4rwgOeVQBF26jVUJLs3Bc2hzJPZbr8iBSGeH
BYZSOkW0GwR6+NJuWAYdT3ONIyhwqM2+g/YEdkPj1ZUnX9xGK8tZIbtN6EUnocJeJm5vXQNebs/R
jSJEtLpMMgBtsutbews2KJ3c7jsnSf+1QRWhAv9CLZbdT9N95G/MajEiVtw3ycw1tjeE/2b45sfr
kBiZEo6+1woy6NokPbXRtnT7Toc9FMDfKTYao27q10igxFx0sIZCW27UldUAkVZuuSG2orJb4+WZ
mUR6Qy7MNidEWV/K25r0XzpLf6/cU4i0HVW7V8u3drbjsUFTVRvnNNWKkW+TQSbeukddvfl8kmJS
UbRksm9lUILClUz6QIa2W7oUcAwbl2KWLN8PYOoSwffGjKbbB7o2LmahohYUqY6qDKQBqw/P95mm
+d/R1hiLEpeB6G18Kfj9GwmHd9XcxuIcozX5D5RBh2zqtqaOXGWj8WoaLA2RnE+jRtPwAiC0+SyP
HD3Ft05VbYN6ifPZXnJOzO3YwMKwZhHVGXMwaQtkMKEaVS94Z0X6b7anyyxkGa1m0gimmu3v2IGu
SNgHtK8ombQuiUxbbyFHq1OowflpDBjPFQsD3xBQTZWsC/Odeekm0T5dRJoqnD5PRtSZXzocqh/H
OgGp1T/gjPxXlqREinmIB6IbHY88lV5czdSHm1/0Oi+pizVbWgp46ZuSgLiCvfRvjUmoFO05FeD+
YrB18MY9L+7xz0SsEhPd1vPdX+4ld+tOjPfuOdQFXiU2bQEOnSuzSJBS+CdqslxuoJdWlNNpn5lN
icsSVH8pSByHSkBrarHE/oeWGkjtuxaIAJCfU9okS8K6J3SBNJUKBUd58PPyV4aNI47MB3+eMgOx
ujXvEjYXFU4hOQBzcXN9N45pjeMelqQ+bZJ4swiIDMLbHrar1o9at2rMN0MGRF9J45H2weBn+2HM
vcVbsTjqRlj0yUdfuuxr4GWhKi1nUDPlfdGKsGW3PYEWxNVxQcqhVf1zU4FcSXT7+wiqvKNTBDIp
BZ76d2CmC1SjX/qw2nWgpp5aXX2wo+9UTcILDxbSJ0niidg6hDzXKmEmMsyjUHs6Rt8oQgwDYpO1
2a/JCaO31ppftxJgEfBQhNjdrxuZlJp4o3ZAin9IqmUx9DL5Hmi1v2wxEtSxLAAcnRwj7u0/j8pX
c7ZJtH/98MkUmVOKtbabfkhkjvHh1EnDfVk4DbMWSRmDGaPqOAPB/9/PkdvZL64Y1MD/jeMYl5Yg
3blyjg/Q1VHp6YJVHAkGTJthf3VQJXn3qvsKqFvXeocrEq2IuYitO0ve2BQbJEhsWliVIDXTp32I
wYV037QpablVN5owykwQeHNBwb2HKfH5AscPVgJsFRsoP3qPSiDmBiva0U3gyzOgPThyWMr9im+K
g5bJPP1X7HGb9/hgOPWl20U74Z7U3fl7YH0/561vTEq/fN+VFYZxC2uGdMqb794XMnvQ5ubx7bM9
54jo/lBFKKacUBWWSFtRwjiVHZ8xQEgO7QYpsnRqqqQC8luXPDsrGolCNEEraUikFI7oHvneWH9g
ZU7u5cap0ssLvLmJXKpEBsNALUbQZ/pUSTGzHzc0SEV3t9zDoLl3lINIHNHCGaXKoN31Jg31NJkq
4io9DIUZrcgUqADj6sYQYsxNjP8rkoJXRLNpXzkbFzbJMP0JPwRQsACZcsltQn5fzSoV+ZXRDsqM
5wfw5WX3VRCAQLs0unsl/iQHCCY1DX2hiRtMpeEJeSwdHxHP+8+Dx+DVNO8z5Z7qWQrSnpZEdETi
ffqKSWFMWer2vIpGSi+3heu9QHyVVFsD73z2ypS6aflVe6Fls++4aU/W7YQbH5ef5inYnewz9ZIE
LuGxD4dIAl4vGv7NKaafMo0KgyCjMgnh3JkvIM/5JyVXGK5NoZ4bT7iHU5ymJ2OHXfzNj5hDPLEH
Rqth39wrYK31SeRZdSlbapbTz+ELZgEQsg9M/cI5jR+ebpDNkx7lbyKw98glBHRBhyiJbhyM9LVh
sOVfs4bOTKCW4qy5XxCd5zh0q6taOcD/r0XYwMLzeA1IPy8SkciTq4CZ3QlcuccPMXOwpFKunxA+
1Ie5S0hp9I7O/CWRMu+IRkIwN9nmdQVZyRnC3C7oNjbg/W31y9MTjJaRmO25BbN1ruow/pzYGfHd
6EuIa0Voyv2DtTLfntzkvOzYZg3L1+T/MBGly1sm1lpkVWjuB9t7FbaGEOFjyWDGWuvJ/yh6l359
ybrgCYRuQqit+9mC4v6gJCQtZtoNX4+TPlrvQifTqAeg0mi2BEXHTmGPHlMxFE/LRvVr69iaGmS0
rKgV/Cu2o+Vg0LzH8WrGHlB1ixJ95OXwrDH/0XbJp7NHUSEDpE9wK5yK4HcCvtXG1bkqfC/h0inu
x+gcwhKKdi9HVQxlCPe+W4tCDoPa96S1D5TZmhzYSFT7kqsjIjkjERKl0GOh2ILqMmZqVvqaNoKp
VmfZUlPkQnRtktFTTpb4it6D1bvwjDPxDdWqyO1Nb7NycyG1qytwmbz7fVlUh6X/bBv4jK6e593Y
Psjx1TS2z/sY/WWQHtS34MbHRrzQp4fjaUQ3E0QFC/3qLz/9w+OuMynXV/fn5tSev+t5zEQK4yEl
M49mM2bZ3waJiy9kpk7a3V4J8N9NrOKZgPZXXPXrWF6sp7JWjXLvKnQ1nArxIIxsM0czn9r8NZZd
wa5YQDvFp6aNWmXtHs0gP+GZ85QIRYjHSEa8OpHHEQbyBiQ2qpoz8CzTv7/oWeDlLJMUex0E3g+f
8bbmGeR/21HXIReWLd3Azsw8hq8dmUm3dD8vQV6f59ceoqF/bTYgW+w0n1QUSlqGIQCOgvjFu7/K
Uqwpzkh9kDJeLoRhjfopV565LxccGnla5q0gtXF9f7ZbWOc4bx836ceVexHsdFE+GyJYFpsbOxXE
QwdYl04Sp+HOsh2q1oRaq+DwNml8Ef4344xoaOLcZrwbfmCccZ0B8OLofyt1tYKwvVrbH9x9yAd9
Xl4rqU8GZ33tINHeoScdDfifjDTh290fDQ1ghlqfUmLEPUlQg4O/xjMwt9RZ7FpG04W1X+3z3Ht4
HoYI+4hG679b/CQ5m5Gtx2zK2R2Y6BaclTXw2s2SD5VsZfPIpo2/eWeUYShUGKRANLJ7e+jbvV3Z
Or75Nt7tjlbFlCyDPLt0YudFyj4Xa+Evri3f0xIYOwcyJZAht7w6/Ni+GOiFvZEHc3EOOPCya0Mi
Xu739WbB1cIV2v+/dHydKknqIlhBD0u6HkGCdIu2rsQJbKxisOI5tkgeKiAgz7to/k3MZJnUs+0P
ZHG/isdKy5D6rAmXslqZaH+ODCyqYTew9by0PG9bRxALTq86SXXFGG95gzSOJnZt6OIRQRqkFaLa
GWw4SGAtMRxwx9X9Dtxjfqg1Uo8swNuUMUE1h2fakKZt/7VUQtABYtMOxTaWvUObSxk/rtxk/3sR
iQgwcaR7gUhe9PKS3phNdwllNeTfztX5i9onmf/3OPmg/uQ5GpruLWKbTTMUZdeEDQmSs9q+II4S
lg2KEQ/2FYzxiIoPEgjxoEXwOfriGQsalnaEvz1fZ6qxOHqpGDwT1i1nUWFe4/uMVCjFeQbFTgeI
ffKgXl5Fr8Z9bj5LE0ILLzdiqIpe9YEx1w0Xy3jmRssWPV38p4P2cPMnXL4A8aLbK2SfBd6s4wg1
OJDpedY+XY+vNpFkpAokgajdxbV1VcTQXm3xSFI2ar6zD6EUtePIq15fA4WFmFID5cyZQtBxbrKh
4h/NKE+1roVDSMuhp/R8oulBX9x9FrRDB+fxaWSPCjId5UUqTbF9RCfSMAtADLxUcKpEhaaFRLMJ
SdsheQhVV0dWBLxF+hoxhEv0BFEtuSExbVXyNk6iQFF3s+iayUWOzeyzREo1dFz4pDr0j3BV1aV1
Bj8+nR8HANJmNAWaQkUEKgJWP2w/yJO74PtSwxCC3xa7ytxwnbcn7oQ6mCvEPksaom6UhzgnJYW1
ll2YcHuHhVGu4OTsH5e6RW874gJEya4s+yh8Md5b2S3j9IerZCvUEukBGvVw7ezj86LIbEIiv/Mq
uPWggY7Ht8tiTdrZ52j5qDSPWK/DKlmGnDST3+9LBO7M49s6J+nr7rS9aAVwHHIru1yZ1n7USCRX
2oJ+E5cVs1/DnxhMAt5LN4RCQPiss//c0sVbruw7T9BPw/AIse3pL2fviM7PA/tfzlGboxflxbBg
ctg5781D/pZKytriXRwMFczG+P0MSzH+t5pSCZNUR8t6KlHxAIkMMya2oGK2b2o7mYQHo7Qlw/pw
4lee5nBa0aHwlDuVHqJcM20flMiDHK5G6axahCgU877bOWjdVmeV82Bj8OKTQIM6UPNgNauOuTIy
FdzqiGoC2F7jTNdjZ0lYPpLMHILe2+VL8paRianOKxYqsxbHBdU97Jvf83mBVCtkGDIaG5xPV3Fc
lIHl9OLrVMymfaY2CUbabeLP8Atb5DXJ4AxwHMILhhXH+JW3UAXSfEhA9NyIXagitHGy6Px5dkCs
RIWy/dxX91X1YwYErbWPLENHnSdz5Y7mL580O4rUAUe21jQL7WRtQHXHGCIa/PO0A5dSuPv9QOM5
+j4BuG+cdbbTx9EpiAwrLboBkgelx2LR5ujV3GP/bd7ijJoSEZyfVDsfF2LNHHQcOFN1NvD+SruQ
SGIRu/WBmr/N4vpIPfdycN/q6ojt00FZqj1GWt1nLkiEo2iZVxFAgXp9tJ4h3BxwUn+B+Udb4WcW
dkFD36WtgL3KH28hP+hsLyYLnWqvGht9pPf7PJBiuWlnJbokxPg9AuR/WwIKomM65KVnxuu2D1k3
WHhKo1blCzn6020crPESIANbaONfLevcloESd6iBSwTLtQB+4Ogj8lminjOkDn6PLMB6dLfBu2h4
MoyjC2dl9/hHDxvMdJSTFLiULq9ST2m31mf2O7rbu+Nt+uPfI7AhLxAuI159CoWnS8v6aQ3THPPe
8CPuCCCjGQ7wCvPGBKP1a51v5a84EAHhwmkaT3Q5mHCsz0kDEHf08571thbW1NpVRoaTJ46HeWst
j5+OD3K0SLD6PgSYo5LLL14KbYxgLfII/tSqfT4Ch2eGY4GtfNrESzjfU6Ug1xOqG8QM1BTjou78
/nZDD81ohzeHtRR7i2XzgqCEKbxk9xAgDw6pAlMpgu9VU0EBs/i3UNIw/1MmjGrCLrhGstwd0ym+
+oV3vXzeov9CX8Yzg/tYFpj1DVLu4ArtmObdOJMJJRyMpQ1E9cKL5sZSC6wC2igeZyV5DelxW8I3
f0nDPyhhbDhjcsKFf/lwilP++T8Gzrtfo8sr5F7st18ftbHCBeEHSeH7sJcWlM9hFXud5QvHgUia
0a18sQ1IkjzQ3l+R0E9dcE+tU/GPiU3NWWt9pV7LzBZR/vKo/Sus/gV6ILEvO+tgfm6/3C6R43KH
KUdVfw1Agt7fkynXntFilALSbusAlWlyzo9NHLJWUM7Qqant3bZPPza+WMWhBd3mIxiX3yVGCsBN
YuHOzVdxtnkG2/jl6Y2KUqlaG0uDv1uWJ8hs32YkzNOK76nHPXGyjm3LcoUlURY/BDq5bWsieynV
S37f8CE1Pd1FdgSAw73SVagC1C2uWwJ3DY4AgWHpZOqNhLhMwNXzYtnGcO5fKtPRHKBn7Ai/QpDL
Xu2rwH6ZehN9n0rmuWIn46rVbYaoaaltIlTuTQ0S2ECP2p3DKg6L2FmatgWF9g/UDz2DvjS7/VL9
cfmNdt9LL6jT2mFyqzkhjmodJujz8vk3pnPzBFejv0C/1xKWDcE1AQaEtztsCu6+t4yqXVmM17Gc
U+FKdHtzMP1GoqVOM1G2bVbjPdKI4WgDfqybgPlT/XHr8CIzoKXJZ3doLuncWdctemGZzadbERHU
2dnROZe0IApScG5YuSQfkbbHt/2M6GYjldLczfPiWw18xpn+Ro/WIKYjFzrWI3Ya3j4GvReA+YU6
EzueASaJGEisCRKgT/zH8G2wUJfL8f6d7bs6cRvOmFOk/bpYJnRSMBlUlcAUK8MQdm1ee/rsLyKL
kvQAe5Y+xJB+JLQkHnUsFDdnE6ZC5ILRgFoZhfSg20RFGXjV0c+HFIYPj41lpg9+v3kIhPQ+2eOg
sOoAGtXHyViobyJWrKr791cuDd9BoI3BvfkT5wDusqN+2uKZJlIoMTQ+A1+w90FIaDWBFOYCjTP9
+ubD3VcLpES7oq7o04etzHrEQolh7LRuaASlNfGg9D2/QHwJiqwJxwOjfa6pV2YJ1xOVGOk9pBin
nqe948cZQRvppEteULW/FCFpWyGsfWPaXtps5m0rJZBrkxYVP74o3r78Z6w4AmQqGofKGy84FITZ
MnyKY4X1aGJIIMOWkTQ4O3o5oqF3aIT8PfVc4zf4ecBbz32VEEA3hIM5a5AwQRYFa10WmFB2WnmR
9FUaDtWvmHy+YxzVmGjZsf2LDblqrBXmBCrdxhNIp4eFUIgq/Guaxxo5O9DZuIbnlL8P5mLv0t1Q
Tzev5jHaQleC5a3S7H9bv5L6LyQ9QxadZ66KqV2XMjDBeJZtbzHaXUYcYQSybPsTn4yBDSCyw426
GZs11LAG1LEUxGR1le/3bhoUfYqsDZLEKCA2w15BIm/XEJh37++mgzAwo/SXECSFd36xyXmBbVTB
XADFPvjvgVOVuZUeh80bPul1Y80eZdSufPZoOxtCYKKGwUa2BpKBOQZGsoAnhcwhDdCUM8XzUtLp
8WAv/EHwcQ4KhnDtYdAlIIa5+JCR1yGL8RBguF4QXhJazE3rw3ptH5YgMdkmi5qncb5e22eGHerO
wuo8RYoMf2Ey0yDbcBQrD1y3JEEziZWzOqrvoUtGjUGB5ySoG+xAAW/s3lLsq105yCS3isxSP/Fs
C9VM7BIwGWFszLEuaBLCN4JmNBeT6yJtgdDV+VXJyDUgPmRVzuLXdjs5KYDvBOqx2sZQNTFV5PRq
7N8em0utdbGT7fXPOUcChL6T1YVaV/ZN+ejcJXJlMKv/xA/9BFxuJpfDXZexFDLisprHNJaxCqZx
wueVwrIj7iVCjX+NUWar7/Kwu5Deb31R7vL59Iomud0VJyq2avOHMBXofWCvufQc/tw1s69ZCQOe
/k5jHjYu+h3rRs0g8daLCxyjYZjsi/xN/gJvaID0OC3zFuOdgmS9oUSQTpFSjN/xWaJz9UN5IuPy
ISTYHrlrCF5dgMut6dpHp+V5lA+HdcnRkpSYBlNkV8YFCWoNwimk6/X019dbblmPFYmOIZUfWE3v
185hsRWpSSQ2Exp5mxSU9snTfBmnODICKdF+P4aINsWCui/Zc5ObLg4N+XrcZ5BKr8m7vfNOxQ5M
ExG7QLzII0ffs+lFQFSJcvgTrX6iaBkzb8fUhklz87ek1XabHH7/1M3KNMSvl+Kv8dPkza26hpsU
kXefuv4TZNcSsVGf05RyUm5mSoUzn3XSdZDypox8tDh6xCim6Ugf//gtflr9OmxnVnN5GvXfMU03
3d1VeTbh27NvrsQEU7+vWReTlyNAcaW6c4Wloh0aQMlrVfyA03LAiFBvUMcmCm+dsZgfGdPmkJCw
eNFDwHGa8x2sLy0sSCjTCXTySEegiX2ca0txcpYqoZm57XSemL7KbcTxvYRp9wTH8464vo85d50O
Za239tAZJoL6A5XVW9BjTn0oUnHzVHMmriq8rxB0hhPbOGaKinlUAG411avzDxoXQ+lFLcESiMIj
3/FJ53lG1FP0hWMWSUkizb1d1S1wDGUV8bpcYgROfKEMKeHyLDxTOp5TrwBDC4W4HNVHIXNoKlhR
6z7wMR4ywbR1FnbvEbQNuxhXcpNJdV64s4Iz9v5G4eugSfzLPmOYNBAz880CJ311G60PQ0JTwbRq
4KMypP6nJVEVbC1JYhX4GaFoA9LwglggVU6YBOgsJGsMDCBV1SSrjRUZtTkZQPZkj923avJV8cJk
96dylPOXFGWcKXTUrQBzXbmVl+501XzyF4x+rAuD9uKciBVN/HWjcpzbKGmnP47FTYNWFp+wrV+s
YLbNlZCecprVkKdz+aR6U3YVp8AmjOut7aWDqwo0uGqwr7cHP4ig+LNz7NywdiLJDZg9AoUb0O+2
Qqr3WUT6pTG1Dy85x5ZFojj7PEbyjN+Eh7Y5pzj1sWhzW1l7IZ1zYhTj4+vLdz8QqJSBx8w8788K
a2KhCVZEGZEacF4q43eW+NeCSZlLCbgP5o7aolQ6SP3uV668aaPeAnMFHXusxF4QSqJJ3C/piFRn
zlNXA8Lxmbv/IGU/78Z5DyqTNaBfOpd6AvEvfLlyeTrDpUxFdLoAt+jwJt4y2bgexo6ZJn6DAGA6
HGVRklfWPI5yxbT1FYDxVsB56NMnMtPkkIa9maeK3o7XQuEYu/5exkh9LjRxQ/jfueVPSNW1P2qt
4vF0OzrrP1cZ+frjoy3SLNgvzc+DkcJ/zeC7Y2IXNuGFLZMl4Gyi7RMtRQNE4cDqp1oSUNVdSXOC
I9aPvBjnQxSA/Z3oEbntV2Kw3j8mN83WwnVX/p2yFWcg/SiDus6mrKVHN0grrxGmEt+oQ4R5xNBp
knJmw3G1B+naZ0gWGx6m4JXm4STiUeJfJBmZ2yNRIJzbOjQsu8akndlyHfB6iqLG1hzvcobK00sG
K5fOMtVrWScbDfX4o/AXTSbxTLqSunB0+DQLZqY1TFPVnwD+ZaAYCcP1EHpgRC0fgWeIDnIKfWmK
JJze3HQmINbZWLZ71fFNCJ7dgn8TTrTarxI+55QyC68UK3vOkXMk1OK2QBB+G4g8X4aOnIqDfimt
dPXm0E0XrWypfhP6eUPOQSCYimXVguEICRixD5cJwKQWUk3IsMv9UXI3y+k7HDCNsbfnWPwI07VS
WaizJ4MHGWZg34PUY/XoVIjSRdNu2PQhS/gznLFrK2vJd+T1a4gPPtgDvYotg0wBB3uNWl9/tV6m
R6PuNWKgBfbTMZqR41B/yPIRdFaD+tImXQlL84L2ZL8AzJcfqadX7ni9JIZaIhhRA7WIlImG9AuL
2Ncest3dH9VXcpeNWulzm09J5dhwbHzDNd7LgHAZyuDcLsP4zfbDKAy4Ps1mN/8VyB9puGS3C3xF
3RfOpQERBAn8DqAAK8Hz0075hKh1LAKTql9sEBefGgxlPPa9on471Wz2MYCUILR/6z+EwFaGdmcm
Jxaj/vUjH/6RaOtOvCZ4hNidNpQz4DmpPmwDumdMuOQyBg7twI8XHE+WWY/K/o1BxuH+LyFY2nuu
opViAOedSidtU+61OQPzuZHRY0rx9QjqFgNN0X8NqN2lYC27cP/j2eKkfG/RuVNKtk4mpQ96Gs4n
ukhfS9kd/AY5dQHTDolFZdcnlZE8lGNqoRqZT8lJyaFdn6oheunE0RWAZlTSfLjFO1MQUNXYoiLD
tCjtklvEMxhwitrFNTEMHCf/xZ8TKB+NF5Tac0+I8m/WrtBgINafsHy4eUUpYF9OjT6n7sNFKzmw
vU9onfXLtHpqZ4ZtwyVoL1nn82MIhqvv/hdoslk0iu30nk2O5g3DpM+P65cY4j88mLaPgllx1ud/
wp1G+7HqA8l4M5TFsWf8aXJY5UFUyvqIkB/by0vyLA3NovpSQwC/zlNFybCxSHF+nZ/QLYcWGhZ0
y2Bv/dqtrOBwaaVpb+DUoEdlIIGXn8Or40GCfBYTJCOy/t7rOmcLny1mjLlzx1PEOG3/Ye03yout
UO9BsvCDHSTgtHBnwm9h2ypvqwKRsZNct5B5qMnolHVfQXgnFxdtCisxKAMjsnJLxa46Q0QEiFtu
gb0TRvWn25CfccljdjTfSsmycHE1UFZ6wHxYZpE/SM/QG00UzN/EuVaBRCdhMS72k4TWpExI/cr/
83zLc5AlcGRBG6hkZLZMuifo7oPZ76I2cUo4o29zVw+xLrV7qDzT6a5XMZgPskPlDbQjT1KA4IfQ
ew3QZAFDE/OC8v2gLeoSAQcDQcz90u3U/GmSch7kSn0nKnf0raoC30TBtfWJJvJyXAUNvRotjcr+
Bn8mr8iZW9uII0VYIInG4MKob2PDyZWjn+/BJqB1GtmuuFaROQ93MvSHwiwsjkQ0JcCLUQrrlH3P
SETLQFQxDLiqjJYPeXk//LZLEUhZ301+AwdDBm6IYAg5KdmbZpkjTMTEZcaByRP5UrAY4EbIBzoH
zhp7sDcdSgEhem4yK8cT2UKPkHGNIajqovS6SpyZ8K92t8Jg+IlPRnkcjJFwXqyJ4FGiwR3dkcaB
1ZSHQGzXlZTueolSIFB37uRYFhsWzOQP8Z/3oLOCxeZev/FyjGbtqOIBPtOw0Ljc8XYvO/tT+Egc
JEv3BBL/ZtBoXEUw6YftaSniKg0DsDMHNDGWez33f3MepFkpgrfJvl9oXUXpoMWv0i3/vK7ZjJP8
eQ9XgnaRYx0OYaEL7iQ4rLnW7xmWvXQ6wCBY55FTW5qouLEb6GDnIfiJNobvQzmR2dMWDCr0v8QL
Acc8Yo81AqSeJM1AUHYVKtyd1m5yT8my3qnn6s6KFtL9RpYttWL3vp2EyOjz7v339QjnyJBM8MnG
aSgI8JvcbJ9h84LAoSVmakqjaIgRzxEeATtXms4E0QBBnE8MOj1M9Uudwby8svoqMPONSGXRvJw4
8ZUJJvmRrdyri2sdQwg97Q4U6FI8eccUEPLCXOsFJ6mDbEufpjG15Qx2ciR17zlG0nAQsmNkFt9K
dlvaHew7oy4Q+Mc1iCHv0vGqPDNiZKkKxtdNFGauBQk2n2AIKZUXMNsgz10+0BKRZwIwXLtDTR/j
poR1UmBW/PZSSoq6g/pIr35Iq0kZVfTRM3qUirCURDEB+7ODaTKxrhKlya4+Ub26VANf9swE1xZj
j/xCNY891HO7LGWUkokEruFXdS5gorhVEcaqMslC8WSsHQHqZuBmASItuKEZccMjATxZio00AsGm
h3/d6qcWiL5n7+CwMpLfrs66j1SV7i2yECigo1of6mxdyEGvrmtMh9SyXdx2EX5rIE5o+XFv0qsE
CYJQwUtCx81xiZED077DZ2uUqi7JqifGGWgGJkZBuHyRaHmVziiY0T4efU9Yn9IjcIAysXXsMedU
7qYr48WdjYRU8iYx7Q/RsG/5+3x3Ygnbz0II9ojOCIbTpS75fYZHX2rLgbnRts60D1McboM5iCbn
Az/rcf3O2NHla8yWjiKy8l9IWOnHu8srdusFU86Zui4iCs5iYk8kyC9b396yd0+Q4ZH+ZaD9L39c
DdpiV78FTMsxIXx2/ygCtVBvX8CPwkUVzfWLgRFSw63OaycEjaa8QZ86r/JqCxgkx2Z9eyj+gzmh
3fBZ133o1qEQ+S2g7i7sdfNXW+Ekc3oM5DiMYefrAnufE4RHpTCXrD/PUBtfTRVIinjLVFBWccNZ
QBbHwR+YCi0M6sK2i63hjv3eo1ibarevCXNCqHPYmELQ7M3aaIo009M3Vq4IDCtnlSCQmwzuEcIn
Qi1QNWY94hWjDJHCsFX0VkF2/RVgSJ9LOHmHQTvLmuFjFdo7rPFhZSWlqJo89cMjRkTvXVd4aLlX
UQKX0U3xkOnqblu9Krblmb3TqCoX0iwbbNTmh9Ioi3kH6Yi9L8cgj38RGhM2JG+cwlhI9rrEgStP
TJssmyjtdvz3+EzaImT8hLqSU/+6c3LU7xDvUIHlw7m9ve1FbWvdtOwnaQrE8yd/yQfDUs2aGJW/
GsqRLGxvjk0FRONIsgjHsfctEJKEjsXk6i/fZeDgDAyG6UyAalT1+Qr2/u+kSI967VAgeVUKKSpv
zMUqpYe+wiV6P4CexpbfTlS4Nnp2GAf+OzdIP7FaXcWT/R6pzOaaTWHXOiQMUkziPog18K73gri/
dTd3DY7gGdrbxtasla9pxUbQyZXgxY6xZfnbjSfjveUzFZV9NoXZd9AIjdZU3glBik1e9CRwsuO3
CqvnkTiWJ5Pbic2cw0FoJoCcmi7SnZvi+qtECejy5xde9uUjWQG0yfIy62GYj9qwhFicfj06QnOB
vMQ0rR7CgahjKeM7vLqZ8Vx2q7EYzXl3gEI3HKnn42i14YfbDAWY3ZghVWqO6MyQO2uACJQhHvTg
oSdxVCivd8ilHdyRfmTY9GZTS2LI5jSwmmEUM+i+5LTcaBnnuFVkkFvqgE3954l0LfY+ieAg8Gl4
2Isesni6Afnm4r9DdGZxawtIWJ9wtKj7IjRkVj/XfsMF7DShG2w3POTBfdQX2VgdNIgj0W3Kq+/W
WS79mjhsl7S1QeoMgMwtdHr4XWq0ke9ukF5CKM6XnQMylcO9tvGJLwee4IlpmgUrbbyVEXu5FRS7
B6c1BTXM5nEYz00B6CNDqRVQssa1De5apCZQYrPlKYDbdZ++49lb02/JBNDnd8vC1D56BzdexmJz
kFdfJxxR95rKjOEpZ890BezLtxjeQVGt5vhNtbsKehh+gFoqToVaWhzm3aZPK/HFywpfdDQwFjBx
09Rd7Nxt9b6Tb0Kk3dhnwBUxxLRiwYW2x0X5tZf/ITIS8onEgJ+74yp88yI+t/FNSfl80mg7Rwz6
wUw69Il4OskR5WVxqfTgDIiMu0z5QsYhYsjvsih+UOQavZrAhTPrbSi8mSaw8amkKQ6jn+r2RdOU
DHX467UYhcXKZqahcSkmX/RR4GlTCl8o2eveJ3XYm8+Z1KfDwCLEbTGMoYSPSImWazoOP4k6kHEY
w95jiYo5PXQIlj4ruql3rWYClL/0mRiGKKVipBE55WkTF87CHn7CG/RMJVndClLrFF6BaM63g9Rz
Odlt/LdA1xAw1k+/pTucqA8b7ypl3ayDVmYlp1OrK6ng04u+NhBVR2G56mByhnLhCn80Ps/5lYcp
JUb8Owm//Hcne/f7LaM4UVq+47bjzkuV+AHqz4u22Wb0QQ9s0MfNJS/279f2GmJymmpMu10CFh5X
0rcAVhNBGN3MR0yxB5GEY20AXe6WNEXqJ6bC6gbSPb+0Z2typjLjm5xywjFO7rfmwJeRuGbqos2i
J8q++B5rFY4VPr4/tY25PucmQYmADgs90dVeDxTnDZzPmPtLhSW9EiLIcxnIpKvVn61xWOM5p0Wg
qeGpZGErn92y+igiL2JXVnyS88jNsFnYEFHyK6wCWfBCO5QarCxzPlddKiJM0UBmtUfVvPD4jhHk
Lj/81I8B80Hc4ASBQo6TK+gjReH8bka/E1Zx5RjBE1AqQko7T/LlqNg1CqhOnjeTKMJvxnmgvnzX
tQ0BMbyPoge5Ku53pou3zsE9RCSyXCKaowO9Lbt5PyOh+YkXZpwonr/ksYu4eCxaeGzxe7C1xlKu
5RMwxG6SBFefM7V6+T/B9+tqJxfYmCOraEX0dXzUMBQoTNDLkRjGFeaERNKNMN8KPH8/A+fbIhfS
H2kprH4CCpTfi/Ss6Trzhz/pZ6IBmTMJMQh7CX3PXWsjGX7xC0XdLPT+Aea+rMVW5faDQcuhgk3/
e5DWXrW3U0W/tJpI57/R+nrCuY1rPPEGpdCEz6yw2FrI1KZHsZshRYxyhncOifyBFmeae25cdPm3
uvCzk+cJuwhhP5145BVZ8rkWGW3Xm/BVMZw/tDFxQHBja4XReRbf5Vh2oqZAjcdhcjfa3Ot2tf3Z
VfYnXhDYRb4OrAbGArivJN12GFuht1fXEVac3CFFD70LDZLGp0fpXHMjIsnfEV0CDc74aobAxrDh
+cpiyEPmfRkYWBM69uYxzqSWLABAK5Fh2t2kcI9AEO2uLuISP0VPUMsUlw9aqgycurN5bgzPvqud
d2KgZwCSr02ErNLAw6EkTQ2JH9w6/IuI1TbARI8Fp4FWvlACXs6afRBHutg89qD+8rMsqGjQK8hO
Lv2DitFtm2f2OwuAl7zKm936g1TI73/dY5kMozqeVMPAtkimSxb/EEcOw87qdt5Qj/1Xfv25shN5
3ru50s6UD3rQZii30ZzX2DJz6pd/FIAHrjZOOtcYKbywQKCwSSc6uhOvlE8vb2WgnbMnq4eJpxv8
Hf0nijE/0uMOT93mzpPGpZVl7rnOQwV8VdmGpGRoZlqQzRXu661L/7SsBW3G6H1zl+US/8bZwBp7
Olx6CPcKEyIy+ZPmIdz5cQ9i2yAjq2BzM8uaWlQMDwt+3rJt0z20MGpyF5iyMHJP3cFNNmIJC66Q
VCKHyzyfgu00Ce/jQ6YKnwDDi816gDIe23R813K/9CcaWlnHJaMSXTK/b2JaKeq4FvYpv1zfSTkw
1AZ1qMEfkQy7bA2spELw7qG1trXSb1U3DD1d29ERDTCGPdVfSGfDtdSNhUzOvut+M8So+PuzRyLL
dgII8ukRQDG75tfPUavHohD2MlW6N6TkfgX2+xGrr9MfwqKAFUqJP5E2Huqo7o07ZOMIHuV9pFs/
kmDZD02xgYOLoHs9EUEwWngOPLC1EpxvvkLo9gaB/qxRPmGwkfge2T/novf2aLgtXPk4tl3oG7RN
DsvB3tmQcbzR8VuvvwgL9NUrpfj945D6GIR7q6k1xxI3r9q2FjhrJjv/o62p2/TXmas++37rnv16
tEdiEBqrikfHW4WgncKZEVcpvilzLqOSf2DeZcSEgGDtO9rImO2F6ycM0aIlEPrq9aTjbAh+EorM
VqQPZcANMZqsNGSmur3ljy9uaPDT485SHH+VF462C480VuEkUPyxaWzAoMNS8DPsyXLC3QVhU1Q3
wSEyGii6xtCSAHtZuW+m+RPnHIBSRp3W+f9zTycleA7dDGKGdXoQSBqpFEzyWwHmTiJhwx1vWWrr
c9LEKRgjoL11bybJoHk1C0NScxKAZvkH8k2Yu5Hx9lKxQCYsR93vlq1XX1Uek6sGgmKGs1RRLYCq
Jt+y5ii7lVHlglauo9ayx/Ok9CgxO7SXLu6KT1TzhuRT6GxKIZRt0pJRtAEj8cGW32gpxBVlGsxY
kGnyF+ELzNCOonTe8yL5ANT36R8jxPMjOxV7LlPcLmHo1CcaDl3UZcqY0t9FoXcyBv8csE9xVb7R
69YbPxUz/ptSgdGOCNolBavWfzRZPpnaNO7TsUlM1npyXJvTRxlnobk5zhwYaIJqPpodCuRgoa7F
CXLNGnPk2XLxGSzZ+aUpFyeW3pk9NJH4BAp98k8mOU9UUuqKqsO+H1gjfgp5YNSCCrrD7FMcvbpX
FfDwxz9s5b5C+y66w8CzEiH/fJAMDnPPCk/A6woIfIofUCycsG8Hr0fK323OWx6sBu6pMgnkwU2D
jB8VBzzt13R6E2EozyZx+2SYjh47+wGcY4yBsKE/sSHpUjG2lFy2uuRKVrsdlCClPZzJaPwCRLAT
UtL+EuUUIcC8CfA7tVx5rb1sJWKakX3UpweL45pHx14WTohdHNbD2aRpIryU+EInC8isAE8E1kcb
eCzFC4qK2nKxKv52aYqRTgr/T3Et6xNLIKo9oPfox5CKJ8iqYHnzQPo2zUXqmirqF/i5K7c9mx1k
aAdlsGSsoiL2BMe+Y81f1fuzmLM5XqvqMiq68h7CWVLP/yJfp9pB9BRRPxMzI8Vf0Z0TW5OrOors
iIg2EUpOd9IKvs24HKjYuOlrRbG6nqKZngXsxlmIobcmnzIE+RgLpneW8r5hRB2qJbo4Ovc8/viI
gryLEHWYeGBPxZNs0slA8oVAlLz3d8FSfb3VDLuOKmdsyhj1D2qk9amy2pNqoZwXTi2LnrRoTSx2
Py5swifjZ4U114djC7qI4bDbomyZsmRrL8euw62J56tZSWW/eJrAW0ixZ8FcqqLj66NZ1MGHnM1w
gZqW+6eFknuVCSh5cnaXsoyR5N8yXPt/91ZtboAr5M+kxl5qA2o1zQ//+35zZI0WamqzIn341Kks
f73TuWC64HrDEI4rGscae/7ha7pOhRtnpvj3fyFrl0cm40dIpoDMvYH6b2cEb2g/wnpc420wGmB2
EizMUJF6dy7M3B93VVmhqnZDvkYUDMCa+PRPvtOhLoeLHUtKF8fFczyevDI4yEoZ3Y6fr62oc6iM
xkPQ16lFYUyA9GW51KVpiEOwft9mbe3GdCd/HeEIXCET1zCxsBPToCXkWhjMqfziwuPDUjVoYrv4
4CmkU60FZqk6u+yLovL2IVV/iye7SljAD2Myvz5PvvGyMWsWznmoHq29ekR8xQ3Vo15PCOEDnL8y
3H05Rq4tI3fXEF2SC89X77WpKzPtIdGpEbNqhm9mQ+B6G2iYrj3lo08WWAHeLnRWw9WyVY4GAEHG
lAf41mnBJRVYKPmE6ITnxIzmUxJQ6MHhMFf+sonms9OJsZ/f1pCfnGryYnqBqeAoTqpHTADTciyv
itOpYEyZWcxmT0gyNtFDa46U9PgvsuKdGM855Ie95ZX8Wq6Cg0G0FAEVAO6pgxUn2akjRL31M9VX
wIDHwcJEevRmh4fSMdLuWV7j26VDwG3FGLk2P74VU2xxXgraBVBfO9uRxiXEQdHl5VlWaYD/ghfD
fz5cHa7th9tUJ4a57H0h3ch+ADoq8umk4ZS5/4MxyHhFRFnUM4u80I85ETkgi1JIN7dGoW8aywCG
Rh3xE2W3XeuTKxlWqSZJOYwome5QVSWss2UpA0RLqH6YDZiiCGuLFIgY90zEHtvGWFlLT8kk+EEL
sVOPXWDSIxSzMVLr9a8dJDrJKuuFLJzDflUFYLKIPWLZt8MaIKHHxSwSx7nw+j+EJr2dxLI1TOX8
Ia4hOg4gSrEsh3uZXYUvQJ1I/HW/CiOGCs3psP1yUrT0ekJRIVvA6QRk+l31w8LeGq062Za2byz0
unqrZEnfyHAJ1TQipqep4k976rZO17e81ZKnNaVSL/g5N/GfYofl3PAk7PLo6060P3GHa+Uig1gh
ldGzXosu/RETbhPFlsiBuxpxhS9DMT1GvP8A+sty/HBnzNfSeByW/mCxvjqRa2WZG7LuhCm1URnF
lqXBYIPJ0gFQdHFd5PsTDKvhCqcHOrPjbwzxA/JqICFH0/SBq6dpn+mYE2qe3OQ1ePG2ZsnM+KCQ
1zj1KS9viI4DMbmxL8Jf6SizpBFM752MTiQOfjalWGK7bNeb8BSoyKL951rhDjuO71HSKKM9OCgt
XYYNBjFac5Rx8n3PSkXZEakd/1c6uQq9XSg2plnpg533MkONIKw+Zr8nKcl3KkPPBdQJoFxFOljg
p5ji5btWM0kuLEa4t+bT+Y/9MM8LJ8fmRogNALSAN/lFQdiNlM6lm15/a+VSjl2m2SzNCffKUnBm
gFYmFpiaUKWvFFhUmIKkez77fUkaVnoUOuT1UET0f9wy0EmE6fK+Qd1VsSBWc02+SMjbdypSLp8j
Kp/gavd3tDinpVLqbrKA9ZQsgJ+420J8DrSLo/Xs/KBeqv4shlGPhVTGcCfn1j/QFCT7G59P+JdC
A4ylOJFm7AFReTDaF9LGPymRYuqWNi5yF0XspMzla5axTRsuCC5QGWVLDnD7IdKuMQVrRKbYq7mb
vKLOXujB5Jc0hA4HrBB2pJFGDnhKsfwFbwS+ly0DNLaOGG6VyPtJRpWM4JyY1wbj6lvSNAp4VyKt
cNFAtVOeu9hlZZPWSOzzgXa0KyrjWa6gROfg6bwe2S3xk+G82wtdHc2X4g+fAbXgF9yaffvytMlg
teIryJEqYhW9V2xGkY6oZTp0ANY2aa/bG2IqDy43vwBItN+CUbzQWqrTKH1QRAsJ8kVu/aq9shjx
FCmWv0hccq0qjrBMPk5bitO6ccPGWBrQmP4eC3/Qv/u0V31OSlx/ikgSIObjljvW8/hcDcedTDR0
xdRDVr/GAkQ7aIZoySHfWJDl5KOHz7AHRvIGmWz8Xwmmt/WwZq5KhdFSXQQaiKob/GOhYTd4U3t3
RE0nfpOQLs97bzIit+3COKj3LjWY2duOyScCxnGwzBI7vxyqL4loXtDBE3ZZlFILpSIP4+mo1YQD
QgzwEdz25IrQOLajVnv53txNNqzEdnvV8fK521+OlupOkMtmm4lKbF9a4LBZ/CORXJ+AzyX1je3p
NtIUz2tP7DJTBwuNaBbamQ6aA4eDel5A8Rde4Tq+q95pklcuW0KWHWozU+HL5yjHYE2n+4AbRbw6
rVIdKW8bbuECGC0St3owHSwZ4eofnBDk9IBsoZDzx96aTkHkC6lxMdyx4nmfKRmPus0eZ0OgMZzu
4Cue2lnfgffjxwQQsksqkohxLjfMeJugtyF/NyWzPpJGOwBcXYAGo7tILuUaKdgL2cb5V0tZvgCI
dlT56GTM4F54NmoVvC0uKhTQxadbay3ufrUHetHH9GVG6xVg+hl3RUkkrE7JZnmPrZjXoB0HMEV5
EZWuazCwZRgy2f/sPnDRAYDkXjWpH0gRVhurjSFAXG66lc4KlwZUCorxldKMTCyP66PHF/8YnJKO
W6uGNJlpkhgrekFbJyt2PmP6modTkENjwOPjcxCrWfFv/XVCmHkYVgKJAcMl3yJJ2c/9wNSUVN9q
9bUh99Y3GGjoTXaofpsPMdB62fIwbwGX7Kzz8gsIxhY6xJagb5bJDF+2J68ZNcF4FHfM6kGQUjnU
aFkva96OWW/eUSglSb9oySQ1+i7Y90ml6JgSsUR/M3ugr0CqArH2P4Ko2SSYoJ+jFRZn6h3y+1YP
hh37idTstHAbZ+CrAZ5UZZhuNsOeFEG3pB7KYkLC6Z92yjHos9LV9T9IK+T/oT/ERvHlpmB0EaU3
UhAZmxB4De8ptt6KQCf0wm67+qY4c7NYj/bzT8O2HcBD0/yLoVysyQKpJmg1+vUh3grONo/7llbN
DVgMxu68R1CU56uK7F5e6O63EwztDvOP/Kj3nSa+X5+SREwIZG7mN4yH86Oz8xznbX8j2NzlMqXV
gU2a51XWhL1nMpX/17G3XZy0eSU1KpVD0sCq9tjCAVGTvPxoIPqwnGQ/esqGoBoeaCxRliOe15Wr
fytVb1CfQqf7Y3B1ul9LkofqscGM3SVtG+OGHVpP9q1gI+Lk4RCEZKwoCnPJYrjrJAIenDyzAixB
vpzLrYf/lbbjl462Jm1jqaoShfjyRgoKXwejdB27BFFDOd3Iq+zHkqYS5JMXHr+/u3j9I6wjsjPH
7hY7NJDhmMFv9+X3tFROZD3FpmMc8fPtf29aBJmA+aKvGUQtwXZUZSS+nzoF1WUBdtogg1LhMVJu
d8+tbqE2zLOM6ncYyT8XNCuIfuT9unBExF/bc4cGEE7IUIOvjEnEqFQRTdka4kQY4cSHAS8dAKij
vxNZi8my5xUnZa5GtCPGyZ5yhYb4bpCFu3peNWvEhZHevxH3whD60e+nFwof7tCEj+aUeqCbEl7V
aQSng7iFMU1mI3nZohC4aFf/vKcYu2BJxEOZUwhwyf+WQQvzYrhx88w+GLCf/dk3o2YZE563NdGV
4EYvv+YfE807h8OBp/2pBd2Fd9zLTWrWG5G0c9l+61+fczonZORr5y+6oT1EtlWZ6FAJxwwLpTvB
74lAUgZj0L7DFg4kwarX79SLHn/DgqmmanFcE5lO1jTVX3VTzo9ASKDI+fFzIX1bv2lN4EegdeOH
CSUlXSP8uTT0bp/b9qkwpnx+ZyrjvjKE324g20IGZFMQo1dua6tU3yMSNASgIskE/864xD1rZWYJ
YWMmC1jiwruUMjdJJq9tkrnc05xeqy2ufJn4AidoW7m0FtnTcOjfQEYohxJbNoND3g/DSQHTibEi
izWEjrxJQvpgoE4hPhPLWooZ6nXyhM/M9ez8jjBYEgVjHKXZr3VzJUWwnqiV04bNnj5uNxTbPMLe
bZJx1ZwxVY0qVqdp3EGIcHnYNVbbGZAuhU2CsAghs5JQP4FJnipOWobwP2oeN2mtggN+srLgBNJI
qxEZT1yQQNtU2YpgOi2XI1IeTMCIKmSajZ6NV5RlGqNgiWQaLSVHb38E43yE2JjhLn7iQ0O7WSNe
r58ESCanXsHAa93nnkO7sDPDCW2K+pgZ0pIlSL8sdyblFZoTYO8UxnrhoDANHdykqgNIpWyk7Ir+
OLEWwZXVMjTg6BawBMJU0NNQiTqw9HaPgaodIsJ0fK9lUD3aiDmoIQoNr3tgIcOw+llifw3Pe0yn
SXmvUu6JVjWdLJHCVC3FmjiOatvS0itv1z3woGDPl6Yo8w4I6gh756v/mzoRr16JjOkeEUTsIcAy
/qV6dRmhMdLV/3gbEvunQ/7sSQJZdrhNRTbdopt9Vfx4h6BGLcmrQA+L8f62R6L0qldLXqd/LUMx
PhCGMZ2HuX5U6j4icgeXr5Wuzzbt8ldW8TNrmoVaodBG6VDAWnfdPrN6dmvuzY27sJjxunZMOsYi
QMm9BpP1hH+Kj8b3xwAWydmCuPoX65AoDU70GDFDLdRoWc2iWcGFfbOjwlKWDf4BXrak+oL5HU4I
EiEUyZtzx/mpvTAXTM5sq/OMMxVKJFTjHJIXAblG59j0FjYqy701q3HpT95v3PxRlhWbW/QXPh4M
ib3p7pM6DR4ZkzRYcHwZEZQOli7+ItPm9oOXUavVaqRS91yTv0+vGm0mFm6msQX/38Dni71PvSNU
K9FYU7jdyiSGCULkrdfwthBojKfQ/OQQikQ1ls7f7p08Ue7BUVg3O7ibjzrugmdt27VICjXY7l/M
4Ge+sXcllin95RAYmQndbwMk/LlIWEn43C9vI1jUwUfxgPeU+Qr6Q0B2jl6WeKFxslGE/u/PTj9j
Yf4iErVWFwKBWqy2fa2IpzlJr7HR+/wiZFk9fVKCLu/4BrFYfpclyjnlJCyVV6a3E+c8VIEtERCl
mcWLAaTqKvKqHRQrVJcbfG0WIwrrFuT0z00bRSvIqPYXY4dfNEVqLhdYgN9svhZJehf27iLvb/qv
mp5lwuVa/fDqueIvPCd5wEJ5cpTZ+18Sthlps559uz9qQwXwxOXEz770L2Jd32kAf9fi6/6IgM7J
ZhFPQRCd/z9sjy6hUBITDrdfxW/Z2dJaxdQcUtoGY68pUobszAugqcAJxHokiLEzvah5Tdi3FFcn
muNN8GPpGDGGS5rVge2yMdMIPr7i23URK/KUSwj9c8F6a2sgp1yabAyyYVICpIpyRWXYzbDpnmND
yu0dl2j17MiMBMvc0WHGc1w8CuA7WoR0SbhJ+H8ukeMzGevnC5IpWwFI9CjieM9RDR5B2SFOkzJm
+LJWOOYGtSCtoRgxnwgK63gRaa4wWzp+ghX2OhEofkY1HRNVMqxQJ3jdBSAilg1l8Aej9AL85dra
LMyZCdvW74E4Llb3JICzRQwnlnmqXkPV5Zk8GvrA1u03tOmO8+p3HrevuyzbhQQLWDKyXsMkzMVL
i2Px28zyRIRgLpYcZSYz7rcYBNmUj0DZtZ8aLvLG8GXw5rTwru4xdidmiZ+5J/x87rF8IDyzmVpU
WchenE+7wmcBQTGxgaS7OZ+ttMeGp/UcwvB/Xb3ElJ9Yl77AzPahFv5vPoLiMb3jZjuqH32vt/DG
pc9ZQkqqIzr4Mu45ZpbzC3dlUNeOWGf6+VS4Iy5mupx1uYcDYE+pRVF/ph790xd5y01D5OHdCYUC
BMGuaGt+pu28bCOQvNTH7sHw8dbudvEhDTBRXeV/Mf7wl1uynDkTKyo6x7d1lkZtwLnxi5pVfZ5H
xT7U3U+qNbn1NT73f2tJgFzCvQLB5uE6Ow5rCVGEvi3+EMhvvVTq5NlXvipPjwk/zQ/8rjQoxCRn
U6VEWVx2bjC+imywaBaRlHYRpe/+9B8lbWHpyyfkFCIoO5jQ4/A6A7E49LSGKfjpe0JwkcNLXbUP
6VKycv+aHF3AIcZS3gMsEsuZYHkuiTww51dJhJSAIDnbrGrHc2Qwpk3ZDwUL/cpbOCFDWW/9jmvm
ccIWO/jpQY7Wouq1LLrT412FJa8Df9h8XVDEtSYk64F3gl8J4JngdYhkX/uwcQ+Lx8RK9KOJJtXe
m4n/JjXF0j3cuXGZ46MBFER2PzHGMyu0/CUcL9ND+wL9HeIg3Avo1BMqOw6zZ5OHgiQIKIkG16SV
4nuu8fZ99t9DGF8s4dy3yNruBaheX1c3QHQhPavN/ghbF5keJcxj5tDwBM2SSm1qPZJ4mJIj/YoC
PifKhN4Iu1gZUst6hsbNAF/GbGjPsga/qVLZY7lIkne3WOmF5OezlmOQzA67XePIz6j3vIC6r9fa
/vE1RfQ16hqwHSgBIWVPqG3pNBfEk/c85+nD7HZ8q0r9ztjxA5WpleJLBhJOD4Gw4uvLBA+3rw81
aIAKAfyDV4NhTbVWYHYFIipEcZfnifaWB4LxWbsBUED5jo1MZwPrF8jl0wUISBXeegnHC7vFeteM
OOAZ1vlHlXheQfPuJ1ltoea5eLqe1zrPnxAhn4h7skSjI7MtcGLshi1SV5EbUCIDqSwabAieb8Kw
tni0rD3eopm0p/O3nKFlg58cTjA+xYjf5mpMY8DbUeQvjMYRSvcKD1m5wAHHQbZR3WkfuPYrNLdQ
rh8OxRWGWC1cEj85tgPH9ZrwzShlNiRW3L4zVoQrMjD82amQ8giOgBBajtIzFStOHjd9+v51NUTR
yLhqTz73Q3YMOH8okyJm5b1iqIHBQ1YvoI82B5owC+ZnsZap+dwsOk/w0kLGTnt1Zd/CKwdSrCxA
Dl7Ucbhk1LpkwN+7+EyAYZWxV90yMfiB3LYGoic/4A4rR8SCRotyZDPcWhCPTZq5BEGXyRDM2o3I
hJBaDaieWPIfkFS+n9ttOzgFzWR7m09uVZ5meEFEck1HfpKII5+Zw5WCpTf1crRgjWT9Wv0GE6dR
wj0duIOpEVSS9l+XZGlSRE8n9ufRW+lvf2TCeFLwYy+egzKku93Q7rozL1GoSaC6KfU6f5ITIGu5
6nRYF6ZJUTWBO5W4A3Vy48gtVq5o1xZCtWUC0COQcmi3k8s3+949H9YpIYaufM1EXBoH8vZUpKea
gbzLW8Yiwk8lYojrt+xJ8pobMcQmrDHuaT/3L7rNXDZd8e0MV0zOoSL4sHXfe2QHnFEcH1uqrcuX
G00dH++OJQm+WHswoChyRmqnFI5s4ZVH8OtKbS5iv3/JazR7Zf7aOK4LIKe00NiKYQ3fSjscwOtf
9VBRgs3mwAAWIZrLz8Chfd+4XzEEgec1FJPnYQF9jow6NJ+Sjq9lIT+E0GyOp0EZuYohDWD6jEfi
mCmxOuQHRQwYPmmTGw/nID6WXWyQ280d/sx2+n2Q7/DGW7eFSpyNht45vUEjBMRuc31Endhh/U+t
q8LH1swlP781MSKeB8yogbPcEfknEI2FmeKZ4lKqp32FZCjSJJ0dtuLn1ZFR4oMoZvCFi9JjCfQ4
YNWVTG0DOynFC3NfGsp4njsVpeG3rbjg11sSLr0YgrVyOxyjsrUZTtDJ250vFWr2mCuv/wgqDqdJ
DpaEQ4W44T8XJbQ4d45IBvNMlEx67Ybsx+Z3PiNKYmUO1kJCiD/OUw9Yq256F+DvdmnYkHtdA6Jr
gy2lp22s6hIncs8fIso243UWGu5+Ntzn27TqnMyt6QDpDpKniVCC+uNMikQMHvnTDLpq3fk5qj9p
ebivh55LYNNPA0ju+mG2Vz8FrXxoXPaJKc+lgI0qsh8awIkeqa9DSZM51EiWiMJyQbW1pA8OQzw5
pQSPO9eURAQx3l7lJZPHacMIHThjB6mj+U+bsLhpvQX4/1S7AvJAqgeTzEB6vG0Sa8adE0ub/C9D
oeG8zIMP9nG/EcECFUegiAfRimoSLiRWYTaL/qNJv+Q5HaiJWsDDhSmyTrcrmFTjUO/b2VKN/SCn
YBECOHbywMY4oyNMlCrEzKVxhyS80lpe88UHFBDn6iimusWLS5gWqysX5/6jJvmasos/Q95O6Gzd
pNtCm5WBOR0D9Df76Cfh7I5fkEzEGXZipT8tYKNQrtyVZNFxiVqAtZbN2KpEZYQYcs0uX2Ldh2Su
8X/HTGEV0oAI+zh4Tdi7GKP1Nb97ISLq3J6CEVHJtBaoaZEjghDK5aKFN8kYqqYbKpjv3fQoQWhs
HeHjRIsCo6M2PnqTKRiSK7EVNcPAxbrU3vQmBD4XlaLO77SSMtvViQltOnrHy2i0ahzIJJoJuOt8
/oyhqYWlHLANJ57RiI1dqPC9Mc5d2VHHiNsy4YMCefjqXmS+0JcWrnYRTJ8bK4lEfI507fryP1ZW
qx1QICqeF4XvuKXBp3djG45OOGNXTGTov9KUe7IZ68gZgfdFSR6+fLLhCu3mP9kB5nNiepzCXice
7iYahPDstabznvnKFxMfuuf+aBjeVJuhIwlc+em1440ChSeY1o7WhMbDYUqqL9911DRteUIIIZD3
ho32EV9D9GxvEND6U+J4QClDHu2jvUOTdqUrBAHd8VNlxe780WNG6Q1q6aoo9+p8Du8xlfOWjfQM
jy44PsoHLPlRYUltYOKnED/YNb3snPh0IP6TfIt9F/RoylbrXYpwFX1fLswCHCJrLNqiLrwTlycc
t9T4PZfLuz+RD5HHgzdd6fxbP3o1o7E/WkZdEAhBTZNtdGXFRPaM6w066RxCzbTvt2dpwsx5lIr2
iBMqyUbyt5XqoEZ3c43aeWjvIPVyzOUEYfR5O2utdsGfuvszxrzDHyCCsPILCudbh4YxoSCQ0D/H
HKODrBl4T7tWSZTL7i/OFE9oOyLBNCBWk4dmfPlodJT4OI4ssGg3uAmnUV6nqd77f7n0L68bn1bQ
ASQk61+r7GWBAi+C1pbJgs9N/rmlem/bwWBqoR1/SrvnlbnFQipJxEMDAcnIkpznIDde206Mlf7a
H/TJqVIApJdxoC+zJ0+aG8aiWj0e7lCwVF6b4gEv2Y6+nCUfislycq+Fh5/KJOD+OsE1ElR5CPC+
7glZrXKRDckST2L0iTSfDvkeSeNRETCN+WD0BOm57vYv46XPjEbNl+3IHaACzoKHLhxtnN0uqyms
Ct7w1WR3uyYKtrl+Wa70+XCGcxtErL0K9/QNPh0NEpeRcrgOXBDJhhsDTRgOQa1UIsPxmKdVeuC6
P6Fdmmkb4dmZ857/9pVlJ19NXVhkeHwpjlrGBYAFdh/mOQQIe7VSbxXy9bJ8DdwxjveobIvnoLrB
52qghvEkenrLytFXx3ymN1zKrGBJMsZh+7WYz/J8yyTh+OrfxFxIEsCEFLvqA3pR99y9aXfGuvKi
09zNcwLSWJEmrWb9gSc/3dnyvqA38j2n/SpjCpBudzUIjs2YgN4qbnOxL707IxudKc5/1GixJqqJ
rrlhsoXXgfwmb+7olIt413UXN3nyytRola9cOUrwHAfd38mZgPK06xwg+KHwbYfg1bStmSndwq/j
uPt26zW0Hx5xRpy809FXXQO0W9J5BsIGTvT+I0EZlYbw6FqIHnIGSFJ326+n5/HOLDQinxJ+meFY
96+SGupiUCjzx082+cmAOh1y2ROmP0e6ntCLIK1wXXlO7+8uSIMjdZKq7f1KIhr5pHQCGe4mWjT1
oEIeRpgGn8y+IjAj68w1oZ54UjxYcF5xWACJWLodvpQkEVgZzolK72jk2GdsWY/sgDotU/d81Fl2
7LnvoPf/LkxxzaCZcPY6Wbkcgg307epkjubfGuzp1EklMcVDUitMFGbSGpxd35gZSXed8on9z20Z
WgpeGMVg5WPB/1t4ElGpV6U7Zhki61b+cv14Fs0/GYPnmHXRPf8N4bZvwXcKY80tVX/SKEEM8r9/
AbwlBjULyVLN/7Se9pstgjODCdEjYmWBG7QUMA0/LO8lRT9OD0ehCt3H/v3DW2DWfs0TnUkEDo0f
fenxvYpVlo2OHsnQY9nlqA2H+6QQWEkTPVxwPtIlAQ0AZkd38j/vJDlFHTcHIwp+p67g6aEiLBZj
buTYene5GkKR1JC/fng4/bD3zU5p17GjX6MxsWdX2ZF1SQZWtzDP4m1fQWapQ+lrIpvwX1zU78fN
z2SF9FdKlzgM35zqIBdF2hX+lmDlhekjmZ5DkrjFTDkC0qcktmiu6ond5XjYvHzhmz4+Aq3OeKS6
JbyYa0lUe5Rl64gCNPNMSsIDuYFZ4H9eDvpIfN0kFKjJO+xoCKmhpzYgSxZLp+cXE8I3wp0T8yb+
5vovtGk38oBBeGE6lUOuG2gRvmanDMxzqz8tZqh8SPsEiF7OVpKZOr+C4risPA/TULR6+yvXJcZr
j2pve8prY6yekqhci3Msh3zaybnG9+RSUu4lGdxR7rqnh9UAlORaVC30uddgKMdQf8C0iqR/1YIV
8rxJkyq2zY6GRzcSt8op6BXetKHqAb5OhZSvKHfTq83PifDcbtObXAMB33WI6ORR9B5idKt2KkzT
7xPSJZ+c+JkvXya7Mq9TlqznX3uLPVY9ykn752qhYlRABzQWaOT3ynpZfhE+QDC5sPyg0soobP6I
ngMaGqkIiAgqRmgqoXE5//iHafjOOAIOX1OiQn/TPlVUU3t+kKVAkMc8V3VtVKoeClxfIsLC1FGI
YlCUgduA5RTSizqScufQcr/ixi/s2qFduZRDabOX7cc7piLMvhMJGKTWDKNoErMTIJWJLVs4lg25
hKFdRCGpEzU8pKF3lvZEPeZ4lO+UCNjv9ZUYmB/ipcLVGuuRPsLLS5MAMkmKDuO4Z1iG3dt+CABt
gmz7ItPWcq/DUOPEMNYs9OGu6rPWeau9A7cxHvpC3tLvrFmV7bpHla6uXZtuNKdY4bv+WFL0Q3I3
SLk7XHS+YQnJCUCYsioqxVIlxPReTHGGFeubhACxwvK1xZht9Gjgn56kKM/wIBTq3Zj4dNs5OMUJ
3Qp/gEv64ocBaTMPck2YlNyqVKEbKROsjjE15oXqT6ThERrMf3oJAyxglbSBLBaE5NhSD7tQM71v
P2OrPK4LLMVv39Ym9g/5kCchgOPk3pxA1jpTJE7O0D+zl5SPYLOel4CvfyfThvwg0BUWsBKfHgf5
9nbwjWOMAeTSNJOj9Rz+UTjTtIdFSRsbE/xOPStEsGk4cmf4oguHaL5NmFtpDtdQAlP8xcbPTZy6
C6tMo7LSgyrvA7QEkuUR+bi8Rcn/DyWOau9wmURmN9eAeT6NUP5O+paDXdsQQaUE6MCk66ha8XlZ
PWa9MKp8h4zIUfWIlZXRjIqx6FMtcNN/uV0lvl6gkxND5PAEd3sWHFfntYquYgJnnhN+f5rVVCQk
ci9BW3D5zepRvZfLDKLRnPDNmOb9iLbbeZk62XwXcAJXFTqaG98h14hI3WOuoJuxMy7Q9VPA+NHA
0RKt4Tri+gnxrRMeGOAufbnpQIztP/sV2XvZRWv6aTeA93gr5/awECKhNyAcpd6uBCCScBLGFHbl
WPP/WLG0aJfGbooR1cl2Pm1KVmhVLf2Knnxh6WdJfMINHTE9ianSuOx+FpjlA76brVrkCpf6+tmm
Xzxpkq1rhgiBM3C1kbXM91u3CsqWQT0dPMEq2ZIQmqmnYZuNvJCHYadAT4dHK+wsjEGlSwGoYV/G
5m4ELDc6VNQlHIfRIu1Dfe6HArYPAzkFQCIcXdAOdBprrl/4aH8XO0Ay2qg7MS2eoZgSY4KiWma0
dQH3C59PiP5T9ogW/ScPtvHOqUuWuAvQdEkJ9Znah0N5cq/jD4F3pFbok5ArWHM+qJZaKifrkL+3
lWVM3aSyBOdlET1nbXTKix5rnCSkwf3o9JWH1jLeCE97MiWUGdy8uub+UyyGh+PZoQFz7fvRIhb4
97arm12aC+DjjRVkQO2OtGnW08l3ErPEa+SzJsVztAs3DXXdQU9jnC7aMbmFr0Jh7nuysHGemgIG
u/y8UOqGM6RnaOXWYgZH+1ob/+ANzKStfk3GlwOiZl129JhA7fhKQQmleny/PvXIPOcFIP0hfU5t
VcXmfzJQclGnjFv34EOO6qd0w+6k2OE1pBAH/LXGtdMnW1gfoaWq/WvlUs9oFMdRMMG9WfJz1GYX
b2iJeeFJ5LZ6EK6Wt4nE4MnS06g27opARvDqhHTcN8+hluGBii1vHDkTs9J9JyzHtL0QTyPkBaQB
aMjdmhhGkZEk4MiINEBo183ESLjikdCYjA9hWX8RPw8vo9ygVet+OiCcWGxh+XNV4h8wbfl2HICX
FE2wrYL7NRuR/5HY7ApxEIIL9VbpeNm69rmwAINrlLovUjt0dUWsL6QLiWks1r0NANEYLuqZN7OG
RZ2y2jWN8tXbmSxKqKjdnk1Ae9E8+00pU/Meuxi+gxJz7CUJUDUZQqTox8kFIOnNyoLHsuV2cbg5
lCPSAIkzubhy3oDDeQtLXlYDqBO8uQv6Ow7QJk75KNcv2V+jL+H1EFKJhL3gU3xamOzlBGxykYNm
JOpTr5v+kxzPz2cotJW6MOKwc68o5JE8U2C7So8S1CTdW5XdMBhigpbYR1SvrIK0k3igZ2zwCumx
WyddH/ba+66Y7Ew46m4Ij6CHdVECat1Ola8Y/euyyITT9q1oJs9b91ejFAcRceyXMgJscZ5zb0GZ
OqJOtyIR7QuGrtc5GxzhUvPzH7SNib0jrfShmKoMRs+bkq0O0lxfyDGSuVKvyS3+IBGao75NneDO
/+6hadOqX3vo8hLIMztrpbJPRJVi5vhHzH7hwwbm84MDVVWKzOHs6LImaSripNmQHo5jow8HHId0
EMmRm7ZoaD0oOwq540uhX7SildtQKamSXPp7GildwL5VbNlyEuO2wOHAYeLk3ut3LEuCFWSoErm/
R5pY+FOj7DuqclJCIsQAxGPUe0ChaDtHdS+tpAhVHIKiGOqrFcF1X0mAJlBSB6sM3TmUWZ+VBcOr
JK/d1gg90Rfi/t6d3iq9ep7KoqgAKFxbCdiakWrzWCexsejZhjGu4eUVTMAS1m7KnmAqmEgh93Nt
rj+6o7YLIB1iirP0hSa9bPQrn5KdvX7eRVfhB+SsNMkl5HnbZMq5YALpAvmYngvp/Xfmb9aeH8W1
OtfCrogdJHTLA/93EWA5BIDtruax5qWYDAx1a0GGSj+1RNwskeOnBiGMYHEQ9VYqQ4ZTTTrhD86M
8ygUajSFOMkmKD9b9TVtw3tNuFp3PiMy1WZgezKna36SfsBxBHpvSYQy8vKCiaYoZ2YhktuvWfqQ
OND8nAHz0WC+gNYil2vaJcXdcBjmkFsgeAXTZ6OF7hXp60uZdBnOChCUihKyaBGgfzwcTnHhe4qW
C3uZCTxo3bT/fOPkAPPh3aBR1Uhu+a0VtHeaBRsR49/6Q3Hc80/JRYoPXaV2oU4Sm1eT3rN5302i
UgoPMzSMWl4cgBT7C015ewaJ5HouUdhM8M3n1uzgdeiv5eOS8l6vLkgiYKcG4q9HbbcWsyhtbMS8
Fwc/kukfeuF9bdIb5QEiuuwmnM9gk2D/mf/8SsqatiML61kkZ2uNQ8AGSIxahNYB3b5Zw8xIsSvQ
KQDtQlRpRMPzE3TMDekPWjgoMHvRkZeRFZTS5bxnULH0PJF96Mm56wQ2UDAe0IclDTLrWGvN6zms
nwzoI6QeRcaBEqSJv4Fld8MuSs/AoXVCoYbKdG8Hxk+5cYj2GGam7AhZnOtzIElVxSqP5lEpNlCa
S0KrNm2ws5ljjq7LQzZncIg7XMfZ6YfBT2ifG8D+CETU6T1OHs9uuEj9pAoq9NEDx6bjbxpT9Ep3
ERnbaJeKrbc1mEb0a8vZiDbMEPDIj3GHZ/dH92EyjIo/ZkzO6wEn1bWGx77E13W25yIHvyk7Lpy/
sbACYx1e6ZOuwLIz9bJAHozyJ0ufV5/LKC7tAOnxaWTVtHTSLXLV487cfPo3IGzRnEiOxZ34Q83U
EkmaCay7Lta/i0u5MG4zkaOfudh5IP+SVRvfzMs8lfOtCX5rmLkU9U+UDXRUxcTTOuP2/LHhZhnm
4O8CtAg8XDCWb/FPQSQpxyqemYJirDnKlkmP2DN6IGedgZ2AaclxZ0pMHnZ+GES7aUe5EkQ/huIp
zIb2slDTO7XWokvf6gKZc6Wl9nusaKCyVVedFP2YVoZmXRsmU7WwqMGOgqXtl6et9DeMr3Y8HUz8
op4uryihFIW2kIfjXv5l1ytJOFU3QEUz+4vNalVdxUS1dae9EVF+1Fs8VIjBIo0Vfyn69IDPt2+J
zqvFf/hnpit/09xcnLaIDhSBrvZoeK/ey+tEEPGVzRnuUhtN9PERARMG6/VehiJWRyIdz2rHvNVy
9LMSRBVBKOPNz8pFJugWZVmyuNDzotbgqjRo4z3AL3A5xJwYG72mk+L3qvC4NY4DUXXeMAXNvQLi
7RDRP0kKC5tKpWW1tulWqxMPj/i3cM+vzdRU7r66+M15gq2LgqDauQmoWOOGJnT6VOPmlxJ/dVOS
pIH9nfl4be8OIjZrYH6N5M8dkW6eHGfXosHOLjZVJVT782QGa7pVLFi0GSZYNXPVLDV5R+SDIWPM
Ed64mTSyraRbpw1/ysy8sqprBhTREhmCCiVRIIP9HUeQ+aIns/q9Y+mcFlGogGzOn8XylJ6AV9pu
0Qw3dXfThfovK0Q0MYhXQKtVfnJSoYNNmoGya/oaNrRz31jq/6zHWji/87sbzOBLwXkFOYaVbvBt
q0In5zQN3Pzw+LqGeGPHbuD61r2j8O/aMXS0eBFfjAQa7WnWaeVKaKbof27kdLxlawzBhYBP6XV5
1uapIN4Z6pEojxm3y+imVVH9cFs82+uTQ2lHw9wIC8UzoSIqVdbunYfYCPQXhjATL0XJ1F5jTme8
HPcZ0gvLFdTrLQzM8INgeIC4W5QSQkkhOpnAVq6PxaDixgDo0bhpDdH+LwxXlgzexZ8Q3PIs7Pg3
5ZJOjMw66Bqe1kvcQAVsf46Qms6P+RnEL64U1L6vQaJFF8+I2YoYEGRxm5Wf0OPDJxF7SvMMDwxI
+hYwt1Ww2H4a+v9rM7sqm7o8z9BuTH9Y92J312yaC8z3g8RsW1J+zWAcsUoTfrRQc+AJPObpkZ8l
qnzHN53pgtF2ydgpzfPanecKeXmh212Jlri0wOvIOzMEbOubBuBcBgsa8QLhkmWLEFMZ1KCmjTlM
9h+g1rLNTFfciaOcuuqhLamvQ+EQ3+yeloyJkLM1ArB0nn4wNusHZkHL/5bm91GJER2xMqX7/tL6
8VaNFUK6QbS8rCn/LG+6ezJ3avlxL68Pw1onOl+ZnkDHopzozBFbJCWQ7h4F6aH4k7ttqRRnmKVx
o9Yyok/vc8OiKXcTMPM9AGeyyiASmo7T5LDC3yp+l4Pc900Sk9WU0A6A89dYZTbY2beFPTO/LvMK
wjRDgGvqF/CSByAU5G8J8a2xTe0kE5ueo7eokJBqK9Tn7YMoGpiB7khhxl3TUZ9c5xadHDt7Iuqm
v/+jJuldMG4G2Cyoyt7nxs3ZU8CBuG2f6d/sJqA7zakylgj/cylsJ1uvAlhcqjs5A2vptGCVf3x3
dds9tIuKA1rUlmAoJZdouSAUT2Pqe3c0l//LzQE6wz1YoDN+ZJ9SVx3ZwlnltZz6nG4cnpbAnmz6
5c5XmRQe3LaaAp6A15ybhYPG+0GW2FEAFrkkzbB2+aUITxtPBtVyizcD7WOH24evmJV4LaOZ0ZTm
42QEB5iULnH1XE+kS1lpo+NitC2MWaC91FvFR/gd2GkhbYPEKcVLEoQqKSsrWu8JQcQGkCQT8LEf
LbdEf09MSQUKfvyEmWczE1f+xwo+1ybUxdeJCnCBOj2ocz/M78H5BzigJHIi1Mz8GLk6qKyBnHBQ
C9EbeEaICm5vDXHyiSymK7D4bDyaLBOrSuaTX/NvdHlyRU7nMxjEO5/dNk1qeTY3TC1fEkIfqMyt
OpE5OKYLaKQhEEbaMHXhAFRkcEjqrddACRL/hwVgDn+gUb99Wwst4kbj8A2gtuE3g2kZ4aRSWDct
Q805VmhR/75GZz3qh8/KO9/vQ4Idz2SKd9hLKUjszyTNqEj24a1z+PdMYxfw5dFtPL1SgUTIQwYe
ijf6vO07aB/+oi9dIJPsqsN8OuYaCC/fMQKhKPECMBVHQozjv3JdHCM+XlSVacTtfeZTUY9wx076
ijEEwZwBAn1z+sNPVgmkXDyq55rgATu9LBuHvbhyBi/ZSHz1FgRuYW1NAq3SLZgyPP2szDlvOV5J
Eh7jxhbhG6nbI5c1UVKqkuVsuSKgCdhUPKXjKd2CjHN6/IjHNgVlCkJeZ+R5a99f5SUP6beBEscD
IPDSqY3KtQf812KMv5BiF74izsZEH0lJW0L9S8zHJ4hQ3dFq9nhbUWnZCZarNHdBPNUnYjwEYdgA
YTs9f7skDGvhQf15yrtRObbcUUMyLApSRvGEYvxEnysL5RxzUqE8BJKjHkUPJVuzKgFfjTsB+o9E
SaXlHpyLFQHqG6iWIQZLDjFvN9lMhM7sUANE4SbUESAj2NGJt6LIOZnsly0eLGrnWQ2dYo5ibVJk
n4fZ/4IbclDMp3f46tAY+O3AyN4/8/B0IIwJZzI/pRNuhnDGGuXUKQVrSTRQyK+47GqVxB8O/j91
3zjvIycHhzfZW9dnNge8nbPdfIa+KPd6VC17x2xPf2L/OXTPRUcwG/FsZoERMT5iVZmrGLlhrPw9
4O0Tg9+7XpvRiiNqHBw8G5CP/krFEw3Fc9NOxzaTbMyNxAJKxo9BVFirkN6/wANxbyvLcXzqPGqj
A0efsGUvhYAuuqY+727H7N+/Hcd6SCoNXq145DoGTjyGwdrKAcX+7+78EpZGed2aWTNdvy+G55kV
7ykL+u0Nqk3EvyhC/Dm283ydNKuABbHyh/uFzq27KZ6UBhYPCT3fzNlout831SzK/KXW6hWgzJj7
zdgS6Id6KGt4WvtsTzQ4YAIY8r+IihOJ/bJRI+RVB1YP792pCzHdZSvu2HHUshFFjTDrOosgq/+5
qFLNbxWdnkKtWuh4aO9NvKoHn7hTYY7Dn609CV/lp2D+IbyH8s/3aSg4C5CbwpHeh4SiQX/an82i
ipY607+t6W5swTbtcXBQ8vQjiJEEe7sujGLbnMSoHePC7p9P5pjXAtIGXxUsONxHagVusBcLS6v6
xzqiFz7YYGFCui7DwW0J7u2/RKIemRCcBwggh/YmgclAKVfpIvOhrtW5m8+Q2B1icU28rxhUqEuT
06mvGf0JQVKoo5kVh/or0VN7ASootD4739f8/KgOTaoYVkRAayNELm04yBXondmoI8vPX07AGI27
FqcTGZFZ/eHI8WiKvwpYuNPd2t8pHp8KZjQPPJTtmRDWHiPU5T1G8vxV0aLvJcBZ8sZ60H/Ux43j
HX/cIuj9Ue4RPd3YplHtnflMZyxzS0SKhW3qO6jpVT12OARCRuuUbE53cjTPnkrlWRa84LRaCugZ
fW6njCPtbaXmwRXUuQtyvbdKva7eWT40Tz4fRm1VSHECniglMv5WVWsvbvRKXv9me0XQjSIL6i5x
0WKGQGznbPK0Eq6OOV5mQN6JHS/USYjeVpF/BaF3+P5PQ5LnXROEIoebN9tanA+w2B2HDfM3ktyo
ZMuNiml1Apj/cfaI527q0bq1KkyA0HhgbMdLnXjN84vB5fAw2tWH6SdHPUvDvZyhfGL9rN2gaBBo
+fK3p1GLwrrZTQHLaIKhP6QWpskEZpqsxiGOCjm4rsCR8WtPpVhqJbrTC88stz/kobbojG4dZGH1
2ZzDRGr9dXZW2KYYE1qIC+7KsvoZKMCmGFXUWCJDZIgIzjwyCzzKCNWRqeIWlkLRVSsjzMtjfaGV
W7S6yKx3660Qjcw7EB60fDcmgrJE34S4z6M0H4Yf7/TYs/2mm7ckXLTKmz4XLCxDq/ziqCv8+5vK
aH160PCSl2UtLifBFyejOWdanEbVH+bPQ/nYi35+qoau+B41F2llEtwWPv886fOFwoxIkmr4BXJ1
b5vV7u+dnG3zyXIucPh4Ag6gOT1fOhaO87gg8+KPEd+czNkxT7FV0fVV15UPHUocFeXLQOLox14D
nWfbgPWcIe0U0s/LTSoUNGkarj93gzwrbxnESmkFtkbh1xcvYUdEWPlmm4eJ6tCvu84K+1NV14/g
m1u1H1l3aYmYoUxZy8olDZyCV4fJvz65mdBziIDujjpcSRQhexwt9azJqik32EUxLGKAh0Kage/3
DdeTaZgl95ERQNiDAJkAv/lH9Kr8ZPt6KMBHVG/DeaqqzdUHEifvtVJbJw492fD7WgjZQ1vFFX//
vJ7GHsMG+El2HIIigfba6ZgoJ+ZactrYNrLcloj55qe0tRfGa961FYv56j91MwRG2dQR+gLQR1BM
lYPIuLg0slyVGJWsp4z3+D7XSirOKQFdjLqeP5myQr1BzasgmfLmG6wow4vLbefX5enhdjG0cC3h
rP9k4Mdmyp/5wWkyynVV6NshV9s06vdDTGySAKOspcuhjcXiRXTgZTUWMPbMAcXxDTKaz1TYRM3T
XjXL1WEqSdgfFrYsO8Ps+ZBazVQnMEaCGjLgpGhoCdP7WsoOPUSXWrEs1ox8IreYa4kLK8QNmZHL
nT1HTCqW5V1XocWGsSTc27csgz9kGnDTQj4EO8Qutp+vJjJecAoBvutIIvCbzqeqWV9a5h2BuVNz
OHTADgLVwFmhk+laLSHwfLZQuveUACidLyXSD9huUKCsuyrfcN4cj4Uur7qxTKEXJ/v3PntnoOXg
w0Ymimee8xgLCk9YixfjzVO9hWIVLzjTvyrJkx9ndtywk2k3y26RvKHQksUFusNAD+gMstE35aSv
Ew1bxUC2o+EgXJ+k+PmG+7skFHZ4uij5jMbp0KBc0yf1Eg3H6W3HqySDW9tPFVOQ24cZl2suF//0
uwUazzafyBwZvsf4XHerwXv6I+UcBMIt4GPfhHSO2OPCigcs7d3glaCzs2cD/7XO9QUmjIBGlOX2
THr7sHCIpDp6Jn+jVWIaenSCDCuddB+WL8ZHDQCeGPrxC8pFX/Ghcoe6gk11jyxHDDtqcxSI9z9p
Bn//2bgXwybFastzkNsbzTEJcCwF2shz/pyy61uJQjgVeCotNSq+DS7TvQyXiTW5YvROv7Sf1PIi
64Oys5C9bJgXaGCZuTR4x4d98RBDkieNDJl5uNwZ+pEkySpquV+q3c1EwVBCc7UNI/t4Y0qEl5tz
g2hORBDgaxJ4VjoFIXpvcwfr+ekjiD4vmWnP1K52vryO2fYK5sU/b/4tiuDpLAO7LVUEghPmSbUR
WYcw3/Me0XkAbb099VohZK68oHRp1pKHRtymq3ZgCAWdiJSf6lW/NSkaQb9Ko0OI0ML2BYkN9Xqj
aFbK8fjoveQkVjgUuaUTImArBwPUTuq/KYxcP9TP1oqkv0w2IW4tqRiLOdS4pRaJ2/C8WEPQXWHq
bJWRKt1eq0KMrlJnb/PW/lDzciqOoqv//112OZwE3V0L1SVdmXct1AWlBz59OFRtE/g1t2VfaOMT
MAPin3mAZzq434YISY7LnUdQWoPvgnY4B3sGvWODX3vIUd8mTsedxEmpTy9M1+aphrYb1BdKwVi9
VxpRV+/u34qgnfIqi5Nxgf6m36bRU5LOULdhI+CDkHDWtmv43z7q7yOd4MWoHeZR8Y5cMCAI0aoJ
jUM1CcSNnFmAwbrnjzdhqQzya/tqKKi97e2MQcbMRGDvgSIx9wRKcCiBCW2El0rpCy7VflEjB0hA
2G0wD8yIdiTFvPYottgX1s1lwkMtkppHEAAK9dUELufzlnXB3Cf+lFtcQxAQC3xDfEfjSfW2gGDn
m1rcAx908BFZ4B7DDzHkzeWrf7jIhZSLtaWW+xhEAHn8hULONoLPzg5IaxGtq0ajicSf0VUshald
TVcKCboFtLbFVsZ6rmml7fA3JCFF2pUQtsDshPhmiK4V4/h5oyZjog8VN91XIFIZIfLdai9tht+l
C/a056j8caZLrl1RncItRAtaSUsIePGA/45z6l3CxaOB2q2bu2iMt1J0obrZhbqz+e5uDfoSXo9C
oPIyM4ZHP9TN0RGVoIIMspT03+NiacmFYNuwGmmhTpo4PpcVZwWPczmSX0J06Gn+EicOJCt2pzY6
co4/VXrROwkNgZEce/cPURB+s21Ql4S+aO6R/5GZCD8KixoXLXWdNxkf0vnVdW2K/4WxnTepGAKT
nDKLRSic91R4qo+x1wOnKei+JI77d5jPN7F7fgn4WCqSxVZxzouOdTNzONvXxnbB7j5+jfd+ggVW
qZ8kAviiR75pP8t2ko9V7k4e1ZzthcQ/GXBwTxLDzUNOU7UjheI+T2FZbz/tdpXafA9sQQQymsJA
fwBkntqxmAXmazFNayf4LSvajUVHlKa/fBsohvBPS6U1qKt4Rm13NtEhkUrM2BpqEaK7WdCjIMqp
NsBaHiTt1iLuBgK8/E9AV7tOYYLiNNy5Sq1EWIizrHX87l8ljfclDvUhjBNVjWszYZ31GXVm3r0B
rjUOe577pQatqbj8NsK2KxlagTHWvTM9TbxQ6/StoE3nUZsPqViwrvMb/Ut5i4OFb5P5O6yJrHXd
wydmN2EHw2bkA8X2Wuvl+Pozg/CtUhDbXVUcQMBntd16DMtz7y1bpQpPeeBrsLqWSpAdMMqInRuN
zQL1QPxwAqwCv2la7+DbkuTMT4GLq/fdPWTqEurjSckpf38KH0d8t0acubkVNYXZmG/67ngdOWyF
RLCJQymnc+P7qlvCirTJx1BmZpqcS+80ag6FwVl4yF0K1A4Qr6Wa5eqv3b81UCicl+gAUSKoJadz
dlS5ivrJp+AUqe9RZbBR/Z2OepkO+cSLsTtGw5rH9/NGtgT2c22W3ztF3z9v7uXXOA4/eBubyDjN
UvKEjJyodLfBsQqxKwPbwCsRWFZb7PDfxGkV3b5g+uXVHffGScnUU2XZcv+su30RWzGmVA9k6sn6
k5uApuGzyL/tP5Ldk8lDeMywKt3A/s98DQTe8+CyXvKLwhkYalgVTFxPLycXvaqlE9vb/Z3pa+sa
HH5g/e8C9RZWG5PJOMvoe9I2zAnS6+Ml4ZZze6DK4JrpktCLIRy9aF/FF7JpfUi8r0V6ef7j/aT4
/4OAqB4eQ+kmKZQkGFcS2+HmccpA1G+U02tIlDfpoUrnyeJano431G5V3KQV4QgVYNawLMGSRTXY
I52EwVxlYgoc+71LRkPwRoh47OqHRGQKtcWu/AeCS5gt7CbMkM/QpHFuYsySe9r5QNzuUqe4Q6ie
dqQS6I4SFyEVk+zFnW0v00svVPBkeqA/22wKPRCynWKjktino5M/WZK5Ft3Qc62Njr5Yq3n17Ph8
5PnidV0KlPHl3J7Z2uZdObRFionQh2+Gnq+F2IQA52hRHilV8zt/JTcZrdM4a1uxaX/50kre3BrR
Q52m2zVWMvIPRfyKxbzqCnu1qMcj2mLc3/cW/YNDvur3yMAEOpdVtCCyCH18RpUTOCwleHTcZ8lf
9oqZf2oap+x57ttas4o/CGNQMVtAMAMHC1FzNJMeF76hoDJVGQKfjW2P/q6QZNJPUevzUSz1P3VJ
uBldlUvMWKBj7ySwwOrnsp8dBxXDpdLvas16NuDnDHpDS6qmIJ59qxV42+U1M+XRp3dDByo+7pY3
mYzRPx/jTRx+E5fj2TSaaEYnXVlc5GbIF93NaFvEv4mp1HcoUtdsFV9b5gtLgYTELdb5J3K/7hr7
oD+DzygYXPIp0zZgvXTR+bXniqklyyBeWsxn7TFDN3LouxN8Ww3fdhV0MV/XwGBt9kcbfesCfcHr
rleiVjFctL+474Lwa6CbmPFm42HXNz4Sw8ioG6nOxyNpV1v6asPSvxWz3bLbENOfY6Dhd4j+sGXC
LIv7V0qrCRMg2sGmzU9NKe93Stj7mGqrZRCTpnCLiuXaAHsgxwPtSbl4qk/IogedYyCUIs6SA2Qo
HgkATKGw8BjeiOPVmNp8mG8AaAwTEkXrJmFa/vuUlv4A5ICmCxXDqRA5IVYzWQlXGXjdCh4r3Dmk
a4sMKriwcsjjdgMWmXigSkBYD9EtbU/rif+TLXuFT6n3/49/OQtsH3Gum724Ga2cYLKN6cMUC0Kf
jBYa0/ek0hlAIWH+fHOXPAcqeqawZltY9rJFnkCLog8jL2nw4jjsPOUicGe7xy/GVyjROkiphoNK
zdgC9rFceHopgWG9KrCx9fEKwq8P5+p7hOm+cJA4UvXLYrBVsAGT69p6mOVSGS9vvlDg8cMJTSnC
nqmA0WslYvQPqcy7rCKPGgkTK22zowKFxzXG4bU87bdHc3Zk+DCIjw0eTz4kvHqY14AvilJureji
h68THlF77AGXM3fhMwTA2gidPxEuRgtSe6uibwqykjZGNp2J4B6krW6VxMEud2cKexbaAczS4/2W
JMRT+jEoJtNny88ZYYgWuWca3YS6Fb7smOuLLq30i38mcZOs99OBoyKNnqMBfTTsMdCH7lCtIb4h
A3OVfz+/wM1PoZK8Np9xo0lIZ5b4girnLPZXlu1H8ehGxufn7O3q0xKCE9lGlnH6YXErH5qg3K+k
j7gGqxtsGcF1fYS3dfJl3nbxISG8h2coCKARUwYHo+sC4HdAnEepluRQh+x9ye5yUVbaIA8xLk2m
U+LWCePvValqq2U8WXQbzlgmq/Yw5+jipDir3GujzQGWC9KJ2Mtb07CexmmOZ481jNx0u2j9wiC9
q9McozaSgHGOGT/xZ1lkfMK/ZPEImwrOxNwp/jkcczUCdjoYfBLODlRIYmkXtJlFZ6YBlEq5dKrC
pY5NeVjnopnndrdwCfwGde6AVePbZ/gThhyxmObyGK8NcmNe3cTwwPPBgfXwGKzi9BbCy0C7S1Pi
UqYcK1+x1KYhbZ7hUv3RPhq2lKv13wL2kMJi6mI67ZzMKyDFNFNogzfzR1Ge5Dap7h9xgSDxVFoK
Rp6w5fWWOpAh22hCc/ZZwMLizgIA7RklkJ4Kn0BvluT0CTNMatWMZwvXrY+8Hw6l5d2NN/QVSaFq
8xEMNSUiHvFkG1ufsiykPfRqnWknzxWzvG78HdPB+AZI0O/E3kYm3jlDlqiHikKPJ1qF0gxcfaqQ
WoYSPLHeD+qBjnbv1ABQvzld3a5yEcOSzN54wNsPOTYjMo4JdRbL+Ml2KnDBpXzi8oDz0w8ZmsE9
0/OxhwGUV2/HIDds6L9NbrDfDxtkqOHSqVE/BGJ67wwcXZMtaXN8wSAO2yjn+dDNlU95CaNPF9Bg
ND6jeNzRPF9mOsxAS+nsHlD9RLik1NX3pUdOCs82VihjaI/HEHPb+jEny+IZtT1NPaG+dxdmrtu3
GrKARHo7oYRzStENugEohymTAhBYP0gy+MaGE6GYZ47TqTxxbuJu6RGvrPGS1romxU6rpfBfAOWT
pPyK9dRNj79M8t4FWKxb6DiTHiQdAIiuj0r2OlE7uyVHoj4RSCZxLxDld9vhrt/2HpckrN3+BhHO
PChCxkIdUnk0S4fLy+llkDLwKUil8cTY8iHpQYoy13PJ3mxPRVzkLPebd9+DPFfWJqt7jXu1KluK
MdNecG/9k9XCcBjG3L1DFAGlZXrzPm9S7/k9sh4msTH811OvJhJa4XMFCdrnpw//HWNwlACpOYAe
+adi/XREiyM9sfJtqzrnheOId73FDjmMDyazNfahBBC1qEEcUSIWZpTuIvczixlSs51eOn/XhJQf
2P6nrieROY3BK1kZd+bqCZd+3sBuJfIO/brv9zHCxOYCOOh8aKzAyYyW4IOvWA3Bj1tusmFXS65e
a1cjhriZMsoxwRQeH4P0rW+c95PYfv1sMA6MLozMQgn2vLOxRvsFf8wcRXYOUsULzop6aRb3fn3q
f3+4z6K0/AueuiUtvczzAvmQHv07DXU2gxFhHW3x8oq9bxQj2y7scQk0i5DRFmjG7aVZPZwicEUA
9CqbSOBXtGtOOEjDZ0JlBkMt2spPCVnssfMmCvg0IyqpZdlfSP1zEhuseK/LJAND9yVPBF6+IfNz
zUbnJ+6abNCVmUF8Op8OU5Rf658qL77i61qQvpYD6EP0rIh78gZefS2sJT/dMUdB9Um3b+1a532O
N4Ib0G1iSb+f6TJsNy8+w0Leyn/VReZbl0nkSruwHU1LVCfkg90K440xj9nRFqAe44OsyK0im6Z1
PS6mv9xzBpeBRzWhqxo6TBwmypKZ/CEX1eDkxFe2wjPfJDlTGwOqLh/CNOaeld9QFKdt8Ey1b4f5
u8tIuRmLv0RXmkiNwj6CZZtDXTD/EZYZAa73IaAbxLCR2hqI7xVUq83M07kWZ8WhHiUYof1uNFHl
UfU8fVU34wniB0btjATr/HmMsTtAvJxiU+8I1osk3lDUTP6+GQm8TWjVCx4YYwtGq2ipdO8cly3U
7oQC8ZwbqaVNq+aClBOm47Ut6PjmjbrJqd3NyTI4tj5P1A0Z2FpV1xKhH6vu/HF2Qhsv0kBeSKpS
kmFF2993Bk4UF2a3oLp085KvNpPb4wC9Z1G42pc30IhRlbsVqHPJal4ioBTO4uLTEoVIMyVSQ0aA
S60se+Gcx1cnrogeeVYUzuqbcFPsqoTPcr0026MzSOKHVHcZXJGDkrj8I/UiHSqtgTiVO1pSHKGX
abMGDfE+XeC0TJzkbE1mywtCMy+BvXUdKbSQkhdZeuJ8xmBzKSGIjbIF/eeB2iuSUBIcXydz3ZIZ
okZSwN9/AF556CWjOKZ3ekNj2XFwLoNy1G7CxZUCg8z+OF2gPEvAAZ85sEsC3O0X9M/pNGIpmPh3
TuX9O8JO0UzriwVBNj6U2wYYHBix7cbvCypZXQY1f9qSKPPPXGxHfa1HVp3Z0wbDNpfyibTGSROW
okswU3zadm+GwbB4jJ/+fnOQ5lKjJNHQVs+PGb13JKl85CKU2/M3aOsRR3NOclyHwCQv844EyWDr
r5HZPL913VGxl1EyH5rr3Xumw1XSu6m7F2ybXTxMqZtPRTb9vGcF4bJxlPj2G3D8/jxBVYSqkMrx
PD+VFHWgr3+sorAJoHIgM7MIYGeclJVK+6ERgzg5hwSIxxsHFMDA3PIMRGh0lNblONwpeKnDDvyi
7bdDGk5DzqZCagkf1s+4eoYAz1Kx7SeCJC+hC8XSPgK3COy5P/d+EQeXW6dS0kd2kILmo7oijDV8
nNBTKfWXgyYW4s4pWwvsLSvgiN+Q92H7mLfFcaisVsgrX/Q3ImPQ+TtP41AkpjiM3GPT9697oFp5
jgtk6sfVSl6I22nkRU54QhTeP7Yu7qWfe4cpwxo1BuFs08HTT9nGfqXr8gDW1zZA+pZWG2m/qp4q
I7u2vcc6UDgPPW+6UDxYidX/ywqzS4uZzAaG0fayyGZ7qvszwqdEcE7KTCmkYKRhc1yj068OFPuc
+mvygnnK2ukLAu6pQw49Zwsanht/5bkwJ/CMmiPoHysS0npoVyTI+9ACHHdkZMiIRCVzh0m0MtRh
VaLuIuuXqEA1LPt2MdVGulv2LUz11c/+1A8Czjg8ndOQ41DK6uiRYpWAhl25g79kQWdwrQS8WapP
LgGWU8FvwYIVOvaUDovCfgCO5qY7bLsHZk1PZ2cdkKhlURK5LPVK4rEoEBBSnakwqp17Dt4AI2aA
x114Qi/KCyizLxJUOjHz+v4QK6cpxTZhEr/bI+gd+Kgv5h82higK0lpoxVByNBTtsMySPtAjvRnV
vx7BckDWzJbPI82HeDCVLkEtRNXnYZlBQfnsC8k/9izLe85oYLv2aIL4c3eVVAIofjUZkJ/JaXqI
t3z4eQLGyx5BHAvNVAm2AkLT4iTCbjC9hhOffSCUhjLIsXgSGKacDJ2fFtUOFO3Y9X5UK5mAJSkQ
7aN7bWGIZ3y6bCEawOBX/S+PVlLr+9xS/qVfZ52HOOnsP4FX0bbFvNK3hqC6nGfUp7BTIE2fg8Ic
T0TAgc494EDkwi1YVou3H07RQd8+EF5uA8AVfSywIBN0Vg0jNF11pGv2oTPJluV+9w32dP6VcKCf
gLx18W499fyg/In8Qq1JsVk/GWsBhaEOcabFpL7lWANJaNOO9Q0OiWHgEV46pauRLSWlArKoRj3x
Zhy9udWpKgSbJL5nd5WPI7X+5LuVchq0Y0ZwJmI1F4EwrfOSrSVyegL3wyr+9MLDmrJR06jTQ4ar
DqSu+12zH/7Ndhn7sdU0gOxKC5ivsrOG9IdVO/mNY9n1Ndp6iYDngvH8BW5M0ofhtjC9OjE87sMu
JFOiW4oHliCtSzN/FW2meh0aeiPHjmiT8Gi0uSvFl5EFa3gVYUduKwwmpr2etwYKPfuSy5CMZ0Cp
LHLXsx9ROyMrNR402B6ZbSEpYeYOsoJcanJUWnMfZLIgXNLd6NwxQjhPn5quSCZzTupEoKfszllp
RfgSCq5zxi5YHLvyT8wUG5BM16CniGLvm27hFRNBEAI3Ni3K7VAVMW9JV8yPM+or7tuYXNz4eOyj
EV+eN5aIp57FbJF4u8RhNi8DRMVeDzcHu53xAbcNfcieU7pzr7rzl4CG6T0O8+gCC8fPQbA79UHT
zecXR6aaVx1yaqaUeTVCGvoSpY+zvIjy+3K+/JMePgmVHHWK2L21kIzQaLS4+jFgOCdLSh6sU1Zw
Quc5m6u8Ml2C/b8F++Kb7sn9/GocsdWutA1sOEIe6XTXg1vDuCUawZCqBWa51H5yiUTkx+g/bmSk
e7DywtCTFSec7Dox0Vn0JRX/1nCMaHeigB9M4eQ8bM0gzELsZ2hvaFwmHOJwBuk/SwXFcyo+bR++
yjqxkcksqf8jhVOE0ydua9PI99nXOH409Xb+MvgQu4CJXilMnrlJHKItbopAQoylq9x+xZUP05EY
nA+l/4g2luVqQ4D+QT7MjfodyNM/2VRpKGhjWMNOEqt/HQSayXiE2DmpCEZMeEkDsKMnI4bhTVAj
2AMod3Q1VRJExAcBQQ+ag2qs5vK2oAOZvRY+O4ytAuNDzY9Ej284P7BfQ5avPosFBGRmebAMihkA
Wozpk1c0eJpcCS9QAubOuAacU+MKN1I41QiUKDECiJJtgbmmaag38qsPOOycFx9NWlmQ7z+bsvjh
jdBloZj5BzNkjQ6feVIlPBraooSey/0Y+x2pFkfftvTPWDDDBcWtO5NUg9K/ysHwDywNcCS5VYa5
z239K1mjGtyB1lLItjlQ3KBy8MFFQHIfS59mXVtZXBCo0vn1x4dJq2An3bb6A/52orZ5Ct4RmjJe
bL/q5knDr8EyoCTOcEDoYXShm02XGhEo547zHxj36G9ZRRmZvvPgUE93wBCGyu7/UU2ZHUXp6E2P
vHmKvYQy34FKazNJYs+sMFbU7qY4A76IhfU8oFipWJLPmn41KvrjIlmpiv7RRVnH5RliQ5/vbHNa
7qXVauC7QcxrCwvQm2rlHfCBjIYle0Zl502zUmOhX3/udrJsA5twSb8VWRDg4RpWm/Rb64vru74C
8jck/3ZXp8ukW6wMumqcXHLdknDPs4W5xkudvk8goNEM3g6urj10VhZC6eWHvWryoq+DpwtyBp0t
NFTSfAGH1bPI3QmtTQ/iDsB5xYq7qMGVhisXUCc5qdg0Ph4KWXp2C5VkeDe0NQMrpz5JoKs144OH
BHYIhlOLs9as0W9imr0Ip1hC2Mf7MR6F0D48nYpMJEiytCoh0hIkBN5V2nUwPIuLPkiqFR+qLzIe
QUr9PjPDGqegtFmXTWHcb01fq+EUz01SXP1sVYMpUR/XoXNTCokgiEDNQZjdza/5rXpFADlNsrZB
BJE703qyjMvpaAhln35nZxBmslebxlk1/F54wTzkNE/uTNKidOHBJ0wfoZs5eX59uaao1hYMgch0
FRHjWZBH9TtsHgq7K87SyqU6U4cb7n3LCTclt3OStKMrrvF84CnXs4C9UICsvGwXleZh4c/ZX/8R
LjE4v3Vr4qaAekROIkFYGFgJb/fmXFL9BTGJeMRoJukgvE3NufYDR+1AGvW6bmExYZZXE266QoXO
yn5+L9WIDoY5JPYrpjOvbSZ4g2SNVJOsd3FguCIjz2dmF/HjznqnLv56Mds9tI14COfbnu6cJK2G
nMf2UhBQrpzzYi8ypWXgH8ZnHQqj5TDhP7gmOV6gHU4QqRlDE4R15kpYvXUKT3TpXbL3hjgHGSOi
+n81bVDDfcmSCC44dLsdu/w/fVyp3nnS/Eh6vBfSNPlwMtTjvMdYQST7ftysrhZHC0Kj3bNgMFuZ
Spir+VwWADSEAFtDhKGs27cy7025rse70W6lkY5B3wj7UHJU4b5J5eZS8Wnr0D2LEpUIQuc+9RTV
JZjDur2K+c9Ge/MjV8h+XdDmOqmq/mYcF4lfF5nvowsdfR3sp4bV6idWCuesgi5vW77bpEWNwKHQ
yqhNSIKe2xMgZWeZ2GZ+U5l6xiwErcSRtGenH3cG9XsZ/v8bfgPzwVx0taA081nhPbxhXNrB6RIi
zurma9+V67lJ+XpD18UQkWipsxQIJgnA7fIn8B232IMO9hLZR3B+3NIBdzQSxxx4epiE8L4ORe4N
EeMKxCegAQ6l94w9DgH3Gil7eBfBhF6wvWpmkHaparbb7hXqvzpvyE+rq6K0PfePO20881B2kG5n
Yz7oxjwIq0Dc1g6y0Kv7XZaeltK6nR8WJcMzx4hP3GKKLY7q9F0xFp9Xo43HunOetHLzhhyKjBIK
nc3jAdh7JmcbWoZrfGQdxJTZyhAGbG76H8TWyYOZTWQmbmV/hhDbzaDGNe92wU/mE0q6GxQ1Jk87
GwwlORXoYOBMxi3QA7XmM25oribiopl97GSBsM7WVyzNMEvlpcI8Z7EFO+LRm3w3Zf9qxFPuDaXT
1FyTsimIc6Oo8FxzNIB3Z1BIrFbXm0pS3eVXRKHl8JVpfQg3w2dt2CQbVs4RHN8YEv27JUMVAtor
rFQo9vHpTarV1b6VVH5U/8OjmzBVky9tCHeuzJhklqBBnTYVs4kLaKeEKY+/BJN53f01ttqtvT++
uFDFsJf8LFom/RaWSMpqlPVVrPotTF6wpQThLC6H2V039dEaT+GPQ6yKHiLAwbDpHtIS1rRj0AV+
HtdN+XnOss+yBayeyYvKPrIPubsnNM3aDug08mFreZaTEq7GOwEVor9wZHJSJVzwz+faxaRKUvZe
R4XDTHgBav5c9jYIPXWuJrOArpjEmc6ol9FCUDkhQIPERDJ8AuQlfOtlwQuEJ/qoyf6h21DTyzo+
NX+5ZLZNp3NDcT1Ddtq8awe3S41XWH3+AgXxFAoDFuC4dRZuvd2WEy4PYoGuRNi6B2Jx5Af2FsmY
SfXU5aSnF5L4P2cAyvhGvFafxPFUzD9d6j8FqIXvTHhcuNGONT4FU3J6cqojPQo/QtLZF3sbnbz1
+hTCsxg0v4Xb4hVOYgvds7VIkxxrowynad1R/B6xtmydTX2pvEfczWW7o6o6Tb6eHlWkgoiHj3zi
+Yeh+J8OcvmoS0p4+WEbe79Qpj+twkg+w1jrBpCKrtdixvN3EAU+e3sHeCmOhp9aQ5muowkmJwL3
+jdFpVgtR0JULsZFBk3QqWROuLo61Blg7rNGFSoraHwznTjqLNavBFzFov/aKCciRd2x2WygOe5K
Jl1LFv0/hwT2Pb5/wgJBbQNf5AO1CGyQ3b/odtoIt4Ur7qzbSXqof5diwrCeUzRZHAwBE4ROvizp
8Sw3UZhpCz5YvoY/vhfSQkCpq7Lh0OhCi/xV8J3agieRht6cm4IZPtLeqFghSGrr3E81gCsS2UTU
FChUly/wS0pwfAmlPZylZPtrbOLL+hD/rnW5zbhMmE4rfsti+VbfgbsI0SW6VcdoIR8SF0tz3O3c
Vp8dUihxbAY6fpfPlZMdDgtRQ/dqon026egQum+Eq2fX20iGSeMdVvI9CVzLJJ0bldgl1ighfvly
uOPbvoonvnXKKZCsDWjIHujLoSsdmqqoc/lyGnkpU1QIUx9SNcEwwQLJIN58LCZWZq+XwxGPidnA
oLfanKGOTVR2PxEYXZDGVnRjRgPsc716G0yKXspnrXY9qxd+1wjHYLMMbVKyADWKBFe9YpbCWJWm
Z5aV1E8rr68grHO/pbQ1R5LE39wD7f6QtNdv0K96+4yyFUzQAWyqJJRtugg3qE5Rw/70ZT//SmbJ
Qxc3AYHMGXWqUUocgC25QNezRY6gfKSDUSmr9fwlr3VXAkUGtIiE2K0NACEXUaI55pX5TwUVmGL1
QQMWJn4pZ53x8DKh3blNq3UX3mE2R40quvmzjU0/UNjpu7pfmr6GCRLmoSaCsw/IxmtiTawoDiFk
NoMXQa9USHn/OtLh5ZwSDrLiB9g3RsyPgR8XHCY9AjsYMGt/atoJD5/npOP+jwLssaEDZC/DCFTb
KbY/PaK04cRMkkg6rCEQ7f2whvDhWcdUKsjUjdhdu/7WqliJP4kunmo1/v9qc/ylmxfK3s38E93r
rEKC+wkQLQ73Y44/1+KPF2pW+PsOsqPS8d3KT9Th0Eo4Jbtorz5O25dFxoZ86T79TuoFE2NQShAT
z+aLRo3oGM03QwUSxaD0HnfSMBGhKrFZ0FxPV4trQpQovRYlDctfBCtFIUzbvA3ZBN0AM/pXK+Vz
6K6Eq3C6vcjjfpz9SwAsryZ+Jz8HK2psOgxiwLDpCGQdKpFOSPkeT6H72/kjGPpUytkyKTQl8VOc
fLuXjvPPe6AS+bZLgmMOrkKrkwWvTu+s1AL4kqKKFchVsZbDBAqLzCBakl8bLke4MghEVlNnUKye
rt+Z6d2Lb2FSVuMsutPOZHQAMPBQqANA0XMs/t8/+NxUwdOhkgYX0SK6X2t4ds8OqbwP+MGYssJC
VoNxWnBB0FqK99YZGuzp4nMcm3dqpOsU8F0U4KGiQEngsb21IhYheJV77FuV8XC+uDe1ZWr7msYy
mSdpOnr/zD1lbGMPq7mixkAbBc/oVSdAVlDQBcUo75HeY/a7FJmvjNlsQ3RbkT/h/e0Ur2+3H7QT
49c+mrVFW/XXe4wEaDGJTP7WqaI+GaSyImfeWwlLy1e/o1r3lRCQEd1ToRnRcoee4xdwYkNmUHrK
hq6FR1EOS1HKsPqflhb0wpYFwxS9GR93oNG6o4RqamNsV4uT2d94elTEiBEZhOk5MYpX+kb035cW
80ANFlRVvgzXTZiyxA0huH1wlsyKATdkH3tpM5Y6OPW93xIZ7FEczm/fE70gOEN25DtMHQFyAzYP
MaIBhVEUeC8eznanrN+J4Lc8uwNx2yAP/aJXxs2v0P+MJvzGESpTdXZF+UIjti7R+h7H/PkwHGld
mORlqdsI6DY3mElbzeHQfjIFObwFjP8hcNBTZKKwZ1DXlrOohI7j0CHYFs0UE85UMxURILrHM5l4
EBDoWlOZ26j1QGVQD6Z9P+B/QlS6oT2ely4W+7H56d/7z+GmWOJaQzbwAyJT7V7Qscg8QdfN6tdJ
kvUNRChU5UDBCfMf0S6G7LcLHgN/p6oZv3tJ+K7o8a97F1cA6kc3ilrybB3uWLXrsgevVdNsOVt9
71Sb2ysKrtXG7no+y1Kkx2q5emGyyXFsqD6FkSI9IW1JzvrMLIXjLhkOO/xrXKFfV7MdqDQpIbCo
YSY6B+TpkUpf6/oQNE6IKEVpv2qZIyMy7y58QfLXmdvdRdGZcgSYs2C5IjUUbfweoW86mG8uw/jK
uc4jpp8t+TXn1n+y3a7O1wxsN314X0YWWHILWQzdvJLVl0v/omlugr5Um2UXzDfHElllI+C8wgIF
4d5s/gFEASqr97sWSx+llCOZ4kAXKqc5jWuEzy+ejUiYzZjSWAKSROQJO994L6MZjMvoXQUBWAvB
HAojGYH7W3xCKCZrfo2sQtqhTGc0SF/QTRvHjt1DVFc4b456J+rOyXR1vSMbYZX/xiVQlOqQeYLt
2NuhKweHJkRTlo1crvy3YaRfA1IP1UpHpipQFslB2cqog4rS3lFhcrtP/AVMijPIkCXPhXee1XJV
Zk24+3WZ4IML02/PlgD3uRdQ/4Xk/hzrpmzuf0k164dmQIKVhh5rHh5XEUa4Mlcti3SON/JIB17h
siEu8W/VMwOR9P5JP1p9QRTVsnzG9UZyFKcweAErMhmF2ay5PDUB07iLQyjbSof93k4WH7kk+Iuw
sEPAyD2hyjnNS4CaPEGav1EFbStIOqFaUXEXxSIQnxdUKBzbFSELtTGHXgtcUNqgKKbslDRWW32L
7FGOdNIxxamXWMHHFPiQq9eFvfpdx0AuNxmsptEnN9Y3gWnQ6jEY+NDh/Ru1TB8rfOPtS5PeuV8X
szpoUw1YFf/cwLo05aZEuYModr82ZntlsUyY2r/y4KFlgJ36wmfEcN304+f17XHIKosTryFJUU6Y
DQ7q/tBAXQILEiIzxT1x2Gh6mQE3+lfohiXWBZzls3w9sbqzHKC2SgCIU0fV3isVs1CuXN9mA+C1
S24A1NMdqjHNj+iMOIMx3Ysvg9wuM0nG3/OgfGFKjLsDZYUn7qELm5hZhjliANliDJvb5S18mWs5
8TTHMl1h4K9RwhirPa8b/hvTLaqRPdq2SyUuNPfQE/o4Qa2M6yYWIGMWnVl0yNmopSLE9XJ7Ysff
66RQODvEjiCmlqSCYHpwjlr4U9MAU3NzlUEoTFPbPnv0B1AOBl3Jl5Kg73nlJk2IoO17mcEV8JPQ
0butHudOK5YmvgZQgsrwgp5Z7yfEQZKwZO+5w64hwRFykWggWeE3HuoWYsxQmOdtZEIzrCu4oJjN
EjAEN/MHAel+yGFF8h3OOi5aTS02SoRYlSeBrVaQzGyPZwytrC3/XUyo9AzqRZv9QdeqKOzANBkH
8zgY6FOUBrCEobLphOUJdBT94SfR+uGLKc2QoqvmnqtF0JG89kYJhlJI4yOo5G2s5AByqGGp+Wrb
52mhL9styCe2MC13tCRivHwsPm9c8QBKQ+Gvbgpc6FlVIffSwQgZin+LiJL/smT5t8wuuzydGWYQ
tgdUXvgTwCDovYlUmiwV1S0DEWOSuxn5ipeNDTbPLVFxUhvBNHG4iUJtMu+nL/LF3T6/dNs0CGbX
/6CM2pT+ji6t0uhkVEA2ZQZtdplr1fLZt0V5+fNuL2QB40uz3NctZQD4XGfzu/ew+PKiHlZluFMu
n/PxVhDS7mJX3AXBYmtXkzAcgew0RYPMEprDBClQoCwbeO1ZTZ7OMB/9O4j21Zp/yQZk5JKfmFnO
G1YEZZkHbkkxqEruwhrFK3x2sub6wSnubspOyK0NSOoQl4flaLMx/mfoXoTWGVV2TqtfZfLi8Jiq
AELQ4iT3ZRqHt46DD7kioGNTaAqhlDfcPqc/aD4HTh/JfSWU01b2tozExEqECYM8B/ShorecCjke
u4tZWu7/nbuhJ/LY/sTfFuiyrQcrmypRG4WMVIiILGOEemLCkoImFEd9XfM5CyJ9xsKU/Rv1G5kc
o/T35TB8IexhlK7l/Htnh18BKii8puRDaUYCCE6RjiH4kbGIxHtn7hqapN7s3S+mAnX9yjey9cFV
rBNumhksm4DsfnTD53UGOam+r88Rt1a0HaHyARDw7xsY3xpqCXnhDAhCUPWlRtaRYuUpSvPq6q9z
N/CA6TqN/vuds4jNrrXiKSny6TIYjsdMRYP980nvnWTXdZMH5y378yScxiliD4l5qiIZ24y1gy2b
eNSFBjV0imiHuAqRl5bDYBxqCs3Ez02xJhwjwXtYE9OJL3JeAq+yalDAWu2bA0mJ0nxmm4kQJGs1
L0aBAVCC1aCnaeOsqOKbnZ/QPDYsJbqa8g5nrqvMbnii3NXhNoH+9yqdsO8/1bXAs6Lk/J1PK2eS
XZMdk044LIPr4mTrgPjC3kpgjfmAUHKSyN8HTru6CUtTqB8yWnLI05g72BRcJKHZzua8LjA5M68l
Q0P7Y491nDGfYrurQdgYfUYgwbFWNHLUwlsSYIqWsHx7jXZkyXpu689/vTEmPN4uGBkm+4UUwg5+
yvS2PK1iFetPrABbIPWIrhzaHNRxQQrICA899YdVxbDa/Kvu1XJWaW3KPXryix10NcPXD1JxArjL
nfr7bVWAU1PtEEwyzlE41i+yXEeOhTyhJePmMKpr422mw+m9nmraw33G/8bd90qlVD2VTCPdAwyg
bNMLs9Xtadp4RbNhZkCCsvu0eABQui2HD5oMNdT3vwhFTV6eFPuEzpJh1Ixd44pp93iZWXg8RWwz
1mx2n4C7Qzrc9TBPxqfFbvi/9/HjNVaLNp96wa57Phht0OufJze1wAuxv3fN1NbeJrksEAiplJV/
Ck1z1o1ThWbuLfx0a79lpIdrAR4GA0a8ev8oveq/ZGfHotqa7wywgcaBXdflSW97brAkjRRoMSfR
1LczbQyVWFIo7OshkQVMtKCWNEzwOQbC8mn2n90U2XnNv6aZCRiZCmS1GJ9OiFd22OYYbqmZ+UnI
hjWuUkATDfqy1/fU6Mz5a308y5rNdvP1n1AUd1L517fShBX3ppDNqNlI6jyowERWJe3/+lbCR0/P
yXmTVkA6i1ghNhGcdv24hKfiQf7Nnl3iZsJ0+btNmvqbIaOQGK/XH6KXtMZMiBBAGrJgaOSm1GOM
a70VbIIbX+eg/r7jkhmALGWGnLgkCK3exQhHzjW/E6wHB9qQZzftef3JjVORoPEFscHluMn8HEH0
lVSTxooBg3bvYogX2uj4dVvgSjVMh5tfdeA+fXjPDTLgLigY+KlHYmpy8VE2vgihm6kUkDVBTrK1
1YEswVpVuYckqGIWK9o7GbfzDCK6P83IDOr0qh9iYObqMqqEMxUHtjnz6bG7a0JSsoOAlUFaWtSF
YQcxfLYKXaXqaRK0TV8vm74lLxAgnNrQ+yGTbRFb0HsGorqxxXeodlCOsOCNX32XLou5+DZ8WB/S
x6jXolJGvqg3L65y6tUwrXykSzxO1jUAmkZQa/kY8o/y0nfQ/cnae/VVF59cpfAVqoJVjhLRBXYz
e8NAEJ3kNP0D+mKhnbyVi5jXXm2q00NmO6ptYqD1AAQwcQOdyYgnf6oAz++PtZFPPVt6Xg1pdZqN
BC9eZ9SieD9dikOm0V5eqinSNCSqoCy358nU35fBj717cG9mWPH2hxu8UYdhhIKOiWVv4w4lVHuq
OqyPnj8xmC4iT1PgXRIVj5H9chMkxs/ZGZrmjLsxni2cgnfkEPvddgVCVljvzuOSSO0px0gARVCw
DPmdEA1rz86wCPdZOuBQeWQkrbB7LnN3ma1xSdW4wYbVSkwJXBOmBP5w/r5cNKqZGy+E6gGVV4ov
xtz0t3mR8gd5JbE3doHi8UwLKBpz5UzhNGf7k8kfVDsN7u2Xr7ti2bbs1oV5ErTVSWVr2Z32VU2r
cgtCL7VZGCCG9vAD8icYAVVNJiCjwsZ6zoso5Rp9tg+sIcvqqtk+Zl5QcEFclPM14waSaW9hxVrT
YxeBc/M0HhSc4H1L/xgejDI157d5dIwbRbuSGIPFbxMajkfZ1ePmQekDXEEne9XhZCdgtB2TCWfw
RryVeRqg2Mh6iJfrL4r1lRc+juwAg3KYnXM9lFGLaRGdBEtP/Q9IO3xJaBR9GZubOHqFQGloSTL0
VSKUR+v8ylhWlWMoWChOMBSpyU74A0jSFHn5C/wShJ+FncaT2PF7YacFGTnsWe/BCLijSltRnNb4
sCfd7gLfZ1uqxUewGl82mus+NY8UHjINUBSEykdQB4mBxt9L6/7CBIIx+QggzuJWClVh5VtYvHhP
87F/+318PnfZj4kMJaylSd7GVm5wL2kElzcikTueyU4s/50Q15QfclsnzjsMB1+mojZS/rX0HMty
8oxmGGeZ0/M1/v/CXPiUFGFik2nkyrYnwCofLyBcXKIXW2BRU00OaU1LT7fNuIL3WTXC1aJwM/2i
5d7mrHHDE7fXK9heqkCZ1aErcPY3irYGo+DAQTGAa4k/yUqWD5fuf62YuiJNa79o4pBipunqJyyE
M8bEzZwWDyJlEsZUBwEexleeoTLGwvb8QuK4T19FKUtWA8nZyO5/nlDndn28TIz3qI80IfE6Smem
jsAKKjFQ5VGACbo1F5kBmbHjrak906u+tQB1MVRNi8N9PwpS657IB60wLFx279Pl5wOoobRuruVk
7D1VNUszrLHb+Q7paZFR9BE9qSPRomGAoCpxa4Vs7nfH1qvVSaTR6+VhUjdnZkFt3GGpOK8Lh+9Q
LgmJgRw+G5832XYRdyir9c9SwfhmWPbeBVRkIIDgNPFh/1MYpVjM8SvcK5qVc9DNOItZWuHmoJzN
0G26vn/zyzloarlqOrAOgwcLSL6Cyorzke/HKTpFVWc2z5FTlDBGcnegxaKOCuuEEtiGehmI/QTd
7VIAJZh46qRrbCvGY1n5vfep8A3debkzXq6PVtm/uqIIov8G/Q7g+Kj6OZihi4gt4ttDUsaOE1tI
SZflOcXoBoa9VTrP1HM12luFAy11i+vfbd0jP7/BJlJbgrRhociBawXllS8aa/oZm4V7yUen+kyj
i+Nl/59kVjpJts36WqcgyL6szkVPutbz87diorrrLi5PygHh6EnlOcmo7wrTz7qrNR1lsvw/oC+D
MfFb1uYQM+lQtnAT+xPVkf24c/gOhGc4oATpmKMaAffteWRVA/6qIgMjMr5W8QokL7f3n3gSGt+l
9uRRJygFRXXm+M70KkklJHHY3lszoyzzQ+4eiEkiy1XzYloSvElwp0BYkhVeJkRazBCfYESxHDam
DmMSuLQrGubM9/OdzpYQD9WlQenPFzApyEzcuvL3hOcyG5vTXzeMmqZhquijErRO3buIbww4dhzc
Flr3T4S2R4JLKbZdzBF6CfVkotqpC74e9zwzyOtyTcpQWHeWYsZgonILi+eOS3dGOuAyUPuG9arI
0Hpl+R1e6m3HQ3o1Z8MgrWUUPa/jgDlWr+RHd0ALZQcIiJjvm7VWCEJBN1dhaa7mS019RchjSZLx
o0SU7kKtbZgCel8gpHLZrsXLu3C7Ahhz4eOzDfGj/o1u1I8Hbvc4bP9glM5X/gZHJdTXTpmpECzk
uHKtysvsHXuOV0vE8yMb6J0y+KxtjxUXGDiafQiFS5ArCn1AVpcHGl007nXfHtiSFmn7ntOGBg8e
xIVtflBPo5umbDvRIf8TmD7CFuieoLIGACEMUcK93ekw/p/HQm/pzEa6z8S2HMXGfauB7ODHqIjN
g5FsmpDKIbofMl7s0b9tBQfoEo6UeSunulSkWQBXH8Y6UYUYbSgVSsFxpGMy7z8lzEaY4npKxrS2
kX76MSm6CGnWwUceWLFZqZ9b/FmbJoAiJ36lIAUw7vAq2Sxk6FtkiXLiFBWNW8YA0qQrr+y1PxcR
T+FwQVtU+YxRA7Qjo8L35DRRhRKn29UCW4ePb6j2HndDOGydcIJXO/iPLZymzhV11Eq3snTPc2U3
uzcURVfAA6eaUowG2SpXY4ph0y40HSw00aD7Of3GwFhsaJorITn75xWt1I4px6tx6ukXc+26Jpxr
ixAuSxLBSqY92KDpsvjZJ86BxAbGPbp3sxoEzXPQ3169b/FqNR6pGFup00j/KiV8AYsJFg75oG8s
jz+GZriPFcwxH36E3PRoK+6B56l5CSNNz4VRp8hX5YcA1XMSqEJCnEWIak96KgwR3asQa4DPLU7A
MjFh7TLH3qnlVran29BV5ijxMrN9o2T3BdTjvf+ja1F7XBkDgmyxe8QXsyp12lve+mS3J2hIGe+2
sjL2s4dFAsplUC1nzJTcOW1Ty5sUkFlX3XBuXl8OovtAE8grnaWM1qA8a+uXruCdAez1rN0YmOl/
wdmymr+VrMEXdxB3OWjz871ZcA1Lv/rE6LWZdHW/nbXXYuy8Pdl7IGpXmkFv94k5lSrl0nOTDr5p
o+WJWCIkaUI83sLTqUqUhfZ72a+HRhJPFRgm1MgmirhNZHDWMcAYT9q6InjwuZilfkV0M5xHDRmI
hC5h8SDdCxlXUi/xmq/N2oe/cLUu1/IM3SsvVFzK2d5Gghl8h1ondfrwKZnbxA7x2938+NpOW284
IPNfEi0uNmSZ0GDYiGbkJWmINP7oxujpSwcOk3+JcYBRsLNOEiTv/2Wve38Tmi5y3/hKj8bcZbF5
zJD5P/y2bHwfBB2RGr1uMSkOdqh/HkhWZh3l2Y30XPwlRG0BJ9Z1Lle3Wr6zv0/9v1VjZfR9J2sh
LSVn0RvAfrKqrgz4R0Eb2h7pVE65kKgvfprlP+Lblbu7hG2hyZGv5S9Hx/9r0TIb19PvSNh/LqbU
EMU8w2Plv99aIWCv5MlafotsDprg1yUVtLWnAtoUPtF5G0pcAprmhXmCN3DLbKrSCaHJlTWHJQNW
VRrKSLW+lFu4aylvBr/qxxDoqD57VMBbzB+I+3KXafjO0wW/5qjVpoM6+XnU+Sfx9RM29vtix3wb
/mu/qz7hlJyjMDyuix8Dks7g23ieUVam+u9DaaiiVt76gMIGZy+mCkMqsz4wo62qTeANEiRTQQpo
GSxHJfmsmJhLej9CzcqT9b7bPMnIBQhp3IfncrqNAcE7fVsR+LxfljyOa4VQNHYSzb2ee/SwFAnW
DFBsX/KO1Bh4+bsJMOWe3jaYle/npvU/gWfFewnSi5ocMnZ3HW0y/qVwObw8BeG49srW2AeYkQaO
Z0noe+KLCTkKUsy7HQTXVoMvZUWXysP7AwKQAk8guGqhXhQKxsUEOpcU02c+++glGHdHiokiviaU
t97Ea/GOvqCgdEs7iT6EbHR+cPdEv/6U7Mmy7R+Jc6b6ZhxUQRP78NSAKO+e9G7f/WatuM38EAmh
fWysXoAv7Bg9hCEQFUxfLdr98NxgUpQ/CPK1/WvZeeLoJP0LYiuMmPABGc36S1XgL+miIYkLLYXF
ywhBR9BrSB55SmP8ptXrmE3KlfUstf50uhD/9EroGsuRX5Mfq0Hu54/mEScyPjxpskZQONL2hnOI
QBsrfJjFQvd2g/QBkSrfUFtAs5dQBtktW6c/i2t7lsVQWN8T/ACuKmKh1KXT3jDeiav+1hz/qvlm
tW5aljeLUHy6mz3fSffCQzMA+8ult6zta+4llOQRqrAay9sdqiOOOV7Pvh7dlt2seTlSzCkZe0FK
DzT0NXMHGT8fzVR0Jmr7iEBhDdAPycl45TGOUEK8VfpkUeVDSK8rrtjeqtBEW5IPWsVhnsU8ITDa
JbDsvAcsd9ajDH1sh0IuG1kZ6kvrii9+3iW4aAc3+UOMpNgAfbz3v8EtD2gTvVaFnvV8aKXRhRrW
6k3YdlAw6pXUfGFM+zgq1mSe0ghrFynennUehIQ4UJFaYnqL6GXOX9GgW2jzQFH2IT7unp7wdwsW
YJ/OXwFkcR85gyia39lUwbXWSEk5tu6ctrryBf7Hb0G/bCLyyaBtOfY3qYrx0oeoDejo+g/CRD7T
IvEu3cBJX3zQ7At0fVjqwcxMp8HaMDV8e/3mToWyyUByokCEaBDFbQQuR+VwMMUb7Rz+TH62rXiv
MC3HGt6zx4/ZJL1jCZaLwPAdKD+PFQjDvEbJcxMzmZcINFGaPWqc6oIP/1JXJkqgci5/qGTn0/Pn
DqzS/Ge/fAkZHtBSRFf9vcy5aB3wIqZQSwj1zeLO49YJgfWr6eSJ9g3rZZByQXDANKIYgtFTbKxO
9uwWjJXqrR1yJkLyptFlUuQMLgIRGWinPmarAaPE0mEJsHt4Hbu6KN+xfidPhnQ753kZby27EaVt
nGTPkXGBIeFojzJnXDtXNUObeveavhiTXwLZyTH38boWYEC2q3GaTWhhPlZm2HnpPIzxhZTPdj5e
PkX0q2L8JPkZ4Kio35VcieXOyAoqqfXnVIReevAv7qOqzD72oQFo/rSkS5QgxuVbk0eiWlAjoiZT
wYTqJsCB6Ugi4tpZeLPn6235ywtxOEM/sDiVmcceUIDzKGNhCcZt+5S+FFlZbfStp8pHMHm/B4ZV
QegMryvzlKIR3aNhGtkCrY0WYMVXvkQfbMY+epw2nmtvgHrx9s9aJ9t/K8FWEwqKbVrzk0mhyDEQ
cYj4AWYffSDapPUdeXiPfC2kkoVRsLSbxjqzrowkGKB5NChMFgTJ3ypQN9aotHzn6IX8h73adlAJ
QwqX06ilb7MbEpS+7zqEn5HqXhuYcz2MNR1us7dyw9+2CkhdHEfOIAxY2+b0jEgUZiDsFfbGy+3K
FbEAoCDP+WTFyAMPw9FGRdElsvy61VfpAJztWwaL7LrCMV5xAJ1HJMBI569NIEBMR4pcxlTwY4O6
tUPE+nye4aTyps4oC1q/mKzrGGU9d9v3hNGp+nw+wv8CFCONptN975CQoMhJQQh2e4tQ6tsrt/ot
sfCRcv+D6kOFt7FI6ETJ39ho//RXu8yc3vCsEpmNjlnnvZw95xv/Zf3F6uwlRA5vfmNViNizsjRJ
uW72u+gP/bKG37EUcMwsYOQ5Fmid4AKM/tNIix68Wcbtf2S4lcviRZeKwjlK4jiLi2erg76H0z/4
+VzBvmevLtSN+x9y69u3ccFo987yO+XSNJoXArIBS007d4NG+aQedN9DLh+q9HKF/X0+d3wr6pSg
tSGzAJYphwD1OiLwz7fnmIlyH3LGphgrotqFsxqx+q5dJXMOD55SGsPOdbxP77QBPn0YQCvgqfO0
xDu2VQicNkhmY8T+ZNVTNBac1i5lZBN9F5nq1ulIyJqfy28ulhQzp8m0MDYrWuaDhlqB2pTFh+9+
OLopHNl9TT8Bivjza8TXAF6WlKkLaTcUYV9nVi1MVhTzkRSLXhsjEGIeA6TsiCN44rs1uV73FLHu
BWb2jj3GRYgdxsBvMiPRuhDqSKdgT19m7H3f2baMrlOPXON9A+9wcHXRNcMWyafiAm54YyuKQ+mW
AvB0wqsQO9nVIsagBI0E6UbNvFkBwGZ38CyCfqdn2DGpbus7PdLz5jXppU2I03n8+xrKbw4YTKJv
GwP+nRIdB66MXa8oIwXQFXbLwd81FLq56VwCGolnl1yRJM0tXBnJgI9a06PXewcuAlNKrh+hKkSW
N3pN82plmRVtnb3TGZYxiPqu+sWxc4Lm7Zfgdx4yaz78GwNCzWm3aGkF68nrvePG3N35K0iOAKWs
psQq479lidMKnqCt+RElDNIcX8vNR4ge+wjpY6RsbnknxKS44hUGG0mhbKwf279UYFXsotkP68sB
6ZkQe/DjBv7NqPi75+e6BTckLxzvL3sxLNN+71M42w1T52eHxpoX35+xDEDxc4wBZ0dMlUfmYVpw
3pgsddVVpcjjmqjYsgI7Or8WEv4aYQuaZ4jMPctTrvuEpiTqcDtBgrDpBTyaS1f/pBdcofiihJ0M
aWGhPqZHJfS5Kx9f2sxu2m7h4H9/87A+ch5xUb5geW3hQFi6ugTRp8HTqCY1mOUWbe/abuq3IwtG
4Q6/zIdQVcGBvrc+DPyO7bR//Lw+OtaAso86CJja3c/yFoZNzyHNR/dXhwqBtsi0OmBrfYdfAjDm
E/MzWR1aaduWHKwsv8aHz7ozJip95aAvqK9hFy3qglKZOKUZP4PCkJxZzL3iulfz1uJoWBWmelDi
Cj0lQAIUI3DUxx1r1JE+jB9kgKS5izT320BLwNy7I3y9ymzHXw+g5o5vf3Mu4wzfvaIQ+JQ4PrHg
M+w4dYtCOVfANRo6CQ4FVIiTiBa2ZIAYBQEoAHCcLsdHR09XDxJGlykyfueKsoL02czrzRVWr4eS
ZoyF7E0yqp0UmF8VC9yD9eurFuAVunlVc4fvsL/0hePDVzmu7ECRQyE8LN2riVcsuTPtGZPK4MAW
RQ49LpC7FGGK9L+Th28rPuJX+sjhFOzBNb/eiyiyexqQJk3QsUSzl0zE4ssCpyOzqQidL/lFV+Iy
GSgoMGlvAoynJ6yonVyvWLeQQoyHqVVSCs0LnBr4tm0/3X05A/+cSBaF8V3aLZP0ADgHe9GtyYgi
YrTcut6gwEYjstjnYR8mdr0yxoYhf92gw2qlmTHS/JljTWvd2eYRIcsVVPNXX/KSrGd29WYWBlYm
LrqbKt5+o3G+4+YXBXkEQmEqWG2nsXoLbsOK8+OrF9BvRwDK5lljdrDqwBmUK8ysLopmQYPLhzO/
1CMWEpVOYl9VX5ej9qpioy+hxCjkd3xxwmEBJjM0ZqZ3y3DTAN1n2TFlj9Qu+Xca8kCKK0EYn8zS
QzgKZ3U15fBbzdUct5pzbUiOmRnEKdbK0Bc9Ax2xfyw7t2GOsxlt2Zw/qrmf635Psmb/cUbNSL6c
pm0npetWu+qkuqkWqcS5DxryZAqImE0h6v5/+h4/oOaTKWrfrx14gHPgYNmrGqkzRrYoMObiEmTY
zi01AjHgI08rBKs7HrmvpLs1C4nHU0MF/zpttGutDQSPedQ1eUU3ZH43L9CjNGZhAaI9K+hmywLv
8DkjQlV7i3zG5Bd4M/j57d0OiS/z8f5397cxUh7zjiCvMZkcwjIiqflv50iDy6b1CPi3HHalL9Zi
zzZYU6uUJG9lWfi9++K1dYRtbX2Ll6pMVsxX00v993CARqWtN3O4QV6n8G7Oa6z2annNztcgtLOI
+IIOgZkiFdVb5erCCuj3Ev6hD1l6TlV0WKX1+gfdlJ0Xp6bw8io4Lzr2Y+pvddLsHtH8wn7Sdgc9
UpGNRBx61oN2Ss/TfQQuZLQ5fR9q+0jYnD7dbrukYeSgQy8yc/hlxExKR7yn9/f3gn+QukZCuCWN
voGbhrXtNBhLxJAc88AwjsS5wgiB8hEPb5+v201wkK+GqV5OvW8BIYaQQxwDQlj7nrf8TOcWAt5H
PKic0vY9arObC5uH1L//q2Zvv1q3Cvz6ECqlyGuSXwAD2gyuF4Wxhsuyk/TP1j0xy5/EpSGBXSnQ
zzaa/Bu+RnOOxEQTu6Ag4kQ9K88UFMQRN+uQHVuvDBsZdMM9Lo6RI+/K1dxOmZpX2MxDzqa4KCHL
gy5mpPTpQgMUsaoeX/HqqCX9hwfExGbge3pUG7FBW2DqxhiQqnHf/PEQ9HzD8tHatBogLbYhPl50
dMKm/lHumRJjrvCiE/TcjHMQpxOti/TwoCCFdiKVu3kfBQ3OyW6+TG+/AM/7sgPYnctrfroZtC0h
6KgeRVDnxzCkuET+7ScvtLeTmhBWXJlfUh6pmisAnuSuOKL+mm5GWkC8TBzyUlOPDo0YpNPY92QW
vAv8O4+avAh4sFbMEUVjOnpIsxAtch21CdKSS8vibLd+EcPBUyCI8J/P4QONM4nY5o2WysXEyKdY
+TsaZ6NuTGCuYzpLSAC0I65uAwy1C3yYLi8q9vR6sDX2E4KACQUiLc4laesyElaTGk3ZykObEvxB
gyqw5jeQ0Xxf0m1xR33SIQ73n5zqin1F+ZBJXshu+/P7eTmxVmP8x9U2yfx/H4J+nIQqFkwGUkFW
lT8FThiyctx8aBi3xwamPhsQ/ix0FqASbKEfzTaC8M/klyOH5vhYuRZXLLX+DRhS6gCbg1msRp6h
884U0cQkfLFWDJNDkWEXL4g5vywZxJnwj1ZoY7FAsoDI8mKwwLGjHGtl3JJkcwPE1bmf/cHC7e2g
Sb/PoKovumyeFTNs7Ac+xxIcNRLH96E+Au+VSN9ziOE0EIZMN9mdsPuOrE5S2emD8WIgYXJT5MDu
vaqibzm9jvfovo98G37XZ7hQWp9JxY19zQtB4Ovm8sk1xFaV7kIwXfJruoKN47RJJ4DlnRBKe2ym
XeIQU6zpSnLfJbFryqKNDkpKvmqd89AV0508KgPvMA4bgXnV7R5ghJYxoeEvKZpAhujG5KBVKzFC
83dR8ZLft0YQIiVoHgXZXqeoIkdQsWNuCMOMhD4eh5y8ioCcbo8IoxhgavmKVJnFpfA1c6yPCqOQ
a+Kln5ZCEG0GHFflkAH6Fc1Aoib6Ou35nZvUA9wJ0T/d0gZpTdoZ8SQvs0E5MldK3z9EhPUicecI
RqIos+pH0xfXKUFE1qW3vSsLeT8jEwuQKN8Hxmfer/Alo334r1D/8hIHcQ27p68BeEH+QLStyKXf
8Vdb5Ye25XdsEjWqI2bTwwiJoCoP5aI2XQJ9Kjj6YcjjnptnhIwDX7KCzsdyaUR3qOvinaB4prVL
2mkq985kKtpxliwA8mafalM4wP1lxndRM4RZdbDXgwl2ysiMtqzN9+aGVK6uAYGbV7HXJNngjXas
A6bRn+SfiRpsYLDk9oYYBvqg37RNcpcZLOz0qK2QqZhKqO09ZCmYfJzClOHfesieQ5NA6fL5CXBC
YikxwEpi7K6mBL9TGZqKoDOhguEXHr49Omar5T7Squ2tv33DJ41/mXlRGCxnriPLcd7Z97tjFncy
GHPurcpFAgznYAsn6yyPfMJ7vEyhcV8y0hml/2jIjYIU9fCLmzLXMFwR7hdhy46DVpEKSqDXKMXR
NSiq30ek81LramSa8Uw+1xhk0Zps5QDrmn/U8NcHPq/6BCmUge8jPOW4PvgMm7cqjjE66WEpR+eT
914jI2vZtSQ0Sqm3MY+gijX/H0AAntfMVMVS0SQH704y2LK+SQ6HMh2/iNe5Z9YpJv/BiIGEGXKm
9Rx9N0QbNV76uz7GtDtLvf5Sw6TdE2WdGwLj1tfzqyIJ9DmRCezYurrjq+Tw1AaaBoYiCaPCEyg8
HdtuKB7IqG6Am8UBQYMGAKJJ3AylCiCb+wd6mV42NzWZzEknE9NCyopA9+lrvIceYKz2VB04FWbz
HzhQiQdtie/K2drv/om5AtDpLk+gdsUknPsAAd0zAprNVdlIfk64kZizfoh4036gjZNE80w/k096
y+/7ZcDdLUZBTlFsGeC566EAZCWefp4jJLZNSO00Yr/xTnpnd94mVhz4yG9W/HMwRjo/TUm1zUMj
rqWNgyCaml+MbFyP/EpEv1WOB2StraR0uNCaXKD0OoHrpnRaiaZBlKdNTvWDr0X1TrhOa1aYbmWk
61YMvlijsESDaUfcYM7Eti0Jg6UFq582CrrR2UcbAeO1m7XJABAEMbgxiC7fet7BWWOJeZXQb54B
65bqBN4lABXLLaTPyDY825drm8xqItLYc2rz3bYZ6IH1RxZb3jMP3kZUbFr2t0w1mGVavY+38DPl
nu5jDNhba0QmNy4KJFvOViyjo6zYeMDxs6kVzjPIK/QxHYtVl7pzUqZ2HLJ9rfyBGvkoNthwAezb
SFnp+n+B+kog+xIfdT3RDwlqhDlYutx1kDrjH4HU7FyjUiPjkbUeP5ytiIff53s7ThzRtX4iQVsm
CAUO/HazjwAO6IWct0Keeo0NfSyECkl7tjmCfHLHWGqmdAQWhlPgoyVhfXRLsIrP+6CW2QvM9NLy
jht7whTDfY7K+kIhXNP9ECs1enC5vFsr3epIjaqFlbiEnN+o1UGNJTmBvXR1pAYBKBjuzMs852x6
DqZg7rlcCtcA1bFZhuOfhB1jjoc3sI5nnu0DNJeQisYG6gbncneSQT7SO2QDU9vYKx6A8dFWTn14
QLHIO3MVQMIk5uMwNmEKxUy+pUNQ8Z/9HC7kokxL86ZXZa1GCucipGyDZNDIFpqcpyJOkcbIN/Te
sVzGsNxABfUtEmj1S95uLI4/uZwl6DQyd/CdMpCPT3iwuI6/2sydB3aAXseouKLgfJu4Nl/k+RqR
ib7lB5Pdj09BQyUqXV49PbxCQI10hqfjnfSDO1zTE/u/twa79EzdgP/RBVUaCkNqiZmRygCnE4s/
FXUOVSW44On0s+ZTXZ7TpAP3/gzVfdaqdsULdkKrSpe+Rpn5n+tE/zKqfBiIEyJ9hN0rmppZkh87
kQauc8z5nWBuaZtRFoJMU0f23HNbfq6acnQ9GyUhZENuf0PEi62mMM0hZzxJNTxTRWz/XZoxQRD6
cLWKt69HA0B4nzDMkj8htJJjl3EKp2EUtXaykyoE6Igp0xMdkfIJE/AI4yibGtxbkU+er09g75gY
KBC7+HZPQVOxGLrAiTUtzIuSunHZ914svzsnZlTUB8xolg3OZ/vb6jEA7cFODlgJHyBKjE7w604J
g8rk/KJJdKAaWfkhqB5dD6RR10uM/dkjfhVzY7lJqhKSNkgVuf943RaO6N1Y1dGD2qD00bdXIrmy
mYE2aPuTat+6Hi3AnfFEqkGH7TDtbocLQCE1wtAP/kD4yLvMlm4yxeNrSpSUBdHHOVP//SHnUT+D
/+LpctPO/WInil7MwoQzHbOB4RQn9FcH2MQtkHkzcuy7lbD9nBMN5FfvaNkzsoijqI65a38ywXxl
rQa7BFaOqojUIipRAMwLCDgiIDLbul8AsBSCz7PD2DD98TceXKIIm8T27bgeg2QnZFoVHNUFHd0a
VfH/21yLWYz1Nhuhfqw8EX5VWjLAdPfIbyqo1+iJExCZ1ZKrct97/qHEN6NKstTbOBvmd+frWiVq
lDLwE+FIfYmaWwkjQiIeAZ0o0Phis9YiBURVGWAhlT7lUkrznjylPu4gUL+0CH6QmdFBN4EtIu4p
WfMxyp4iRIR29mMG+TLWxtYSM4OR0f38OjYahsuJhtjRo9y/JVMhyGMcvSg5O5sZayK+6UlKar+Q
5l/HnZQpRD5hn6wt1DXqc65Pt8kz3Vhx147r3TU4iDxSBihj/kt8+OPuu16knLtvGrc/moUqbvt2
wXdilDBKCoD33n5cHnaD2t4/KBTNmBpznnDthGzQwZmmvqMpN0IYxuCDOFoKTbaq3CIsPNBUnmAC
fiSAPlmbvez9C4W4RBkZfrNNPsx5bAQzGYN+sMIIgB/F/3GhDprCS4onotA6jS5Eb1EbvqLhjMPr
keeE7rdroMrBh2fgFgTgoos76AhK2KSrqbKbQrD2jlyf5qffGj+U13rLiPI2uIWfuwK1/UCgbD1C
BiAczgs9dLSDg4BztWGJX+Ds95iWEMhQMFhPd2Bez8RkedCUfN46Gn+ucLIbFMKmLmD1M02pSbms
Ax7EC1BC4yXcpmPoJEik8nJyltzIjNBJ3vDlH9EKl/vzqA9DJ9kRewaaD0+5RMk7E71ITPgIHuzz
emnz7SjaYGUUZn2RJCApYTC27MWc+hAYevAvyfLE6tFyejX8q4nKI6wi5g+9UCUa78krxl3YmyMF
S19nas6DsgvYB7uDFkZtfMqCUpNFcZr+VL1q3Q/Zx5H2P9KeLrsjHYfc69XjIxUXjrFBY1D2gzR3
aSCIeI3xBbhCo5jwTehR5TQwHlOXaDlHKyqgUGrIri9SQshVgvuHV2Jvm7CUxI5sBFg004C+e7HB
eRLmDlnikekMi/AoR2H3GLcj1u6ucRK0MMpv2rgFWgoPpsujcGz5m/HpYbA95YLgqp58OOQRE8lg
SzN4BB/4n0y7RrDXTPrMWFcrN4u9xHAPvk1FcAXKlHr2k3tamMK/CbBvrCBOAC01DkfFD8KATDvq
xbOZv4o+D6xvtxD9+BJyq4nCQaLYiebLLSgjlyDeyVM9sOle18jaSXcQA0Wjh+mEc1sNElwZ/HwD
Itl1L2iE42TSNHoGfoepdE85ELAhHZZ5/1/idr3XNZrP1GPN919r/KxNA5heVXhcQMDCcCwxL552
5jTlpJHtlGySgz8NSn2SQiAF7PtiCQc1NzhkI8FXfWG8nm3qSnzLmPpcaz6LZsGRjaStHooaReu9
6F2omDKVZ+Y4WzQecaj2Xc7B40FVy8eNGEG8ldt+Y3l3gASCTHdfSbW7LEgQ2Hkq7LQrkMl9/1M1
trjzCoWMyaK7zT78lDO3WK3EQF8AEyTxiOpSuCak2lCPfxYqdULZdvia4Y8zHNLlL4COvddROzK5
ZO6AHwsUn6cR2R3l2L7s5cx4wtFNUmsnz/03wyuxYIQS13a0CjtAF7f/wY8F2lnEHtAr5SmIZrqs
eQcNxDdcCLsadW1paL/ZUupSdSSDhXx9XnBdCcdAH/MaT0/0+G79uLrfdj0GblM0aDsNvDxzaWcK
oCm2Z+vMTkV5OM/ggXPXmhxpbX+P3yUEJahgtapy3Zf86l5aQVJ95m6VNmqo4moDfRbqW1Efpo7y
s9TU2kVP2jLeBVgp9wesuEpqNiF1IC5eMoWGOTYMgznvsQErIYMC3UBY0jDNFLthaFskfhZO9wh+
GARK+kM5/LKXn8dNaRKaV0uXIROFcT1Xy2syW9PK+wEQr1eMMbDqmhNYm25cvxe1ChEJ4RnT4Mth
jSD1X993DFmRzzN5gjM2jlyn0/ra1t3HEE6ETx/1ZinDh1Cn+aEe8iWTysc9pAjYlHrBFysVx6AN
esVxE92XH1+4tH5tEnanq+tlNmtvx0kT2W4ths2cvPNqMu9DD3fUbycZmtyd76Fw4ipADYNJiUqW
FzpzxQ7RY8dZ9c5YGmspeIaicB4FfVYmfPzhhl3sEf5E0eJ0BMh8I4IfAIKEbQZkk3ZIWKHWC+Ca
znSvSgYpYTeiBik5FLJJafc1R4NBPZy5jEXNk6nxCfW8ISuS/oJ/u5az5tC3hp/y5UMXjOkReQbf
OXik7Utd20vOn3ilgp/f/zROmwqSULdAVpyfm6i3l1Hf/WSv0G0FUY4GhYVuzyNkXu2coD4+pApW
AHH+fNJo+cTE4qWWzv49d6xHUiZvV6r4qZiKyaw72T7JYyxRvElmtv5seJVCbaADc/Uzeak6uk7T
0BeRVauO6GTNQVFi8hePtf+9JHLvmmCt5MreeukIvFcyB2KwWKoNVYIEyuQDxrVyR+EefaSZmshx
V6k1mksNPFy2krm/IWmsN3hqrR0OT/DO0vAp9Ai+gT7KKWnTxxBLBbmAc//JBI+xGEHVcgm5+r7l
fCfAmvoy07hpUneChNzLnQVHXSw7dv+7NUWXg4Z7CGDIn1Fj3NJmu9WDGbpaQwTA8BAp3HE54ARo
FjtjB2TxOXc5xxK/+5sIDhIhp5mr6RCcJllQYdK0PteLGuvo++DdJZdVumdNT488IOoLG3S7cN93
wdmbm+n/f/9zUjibq5He9F7RkoA5wb2x20z1Z0+MSVV9REUIVCLY8bgiMhIYUZnUyuf34YNF9K5J
qfpaZO4rBGluHMbh2d0ZfAlwR21m3LUMkKDohE/GWM3hxU0cFatdaL5opNJGHDUIo1wQBPnNv8IO
cwH32NmvmJ0ylRXuRJJWYJ3HkfjEXndAKCzd1drtx0Mpo5xtQNiuS/AHIqywJbUSNjB+NfPUxEdO
xb83ARx7utRquGFkVVKCje9855hcsEDK0wxZgHvi3geg6F04L3D/qu0N0h3GGf0+JoYrugy74iJ1
Bgq4Fqs20HULJ9UbZE2uDX4ISOxI2uEVp4Q3iXzYAVyS4sOM0p5l43NYrARCRxOA91yNYzxWGaUX
iPhYUdiS2C5TL9gM0CFjmb3gG3PIhfjxba6OZ4Kg7iN+2MJ61lBAIV1rEj7u2JIRNd+OxGFDp6xq
Kh1Un8RF1dk1Xc3oCnzLyTmMKIrrBk4mKcFc79XiS+I2UN7HpX1XZLL8EuPL9q+9BM8zBO5Md4Vc
d7dDoiT0ftTYNhrb1vr2JAwzYpoh8pwxiA0LuCWKO15MgpQrwBShDu1jtJJfu0hYm5lnjn1/NhYM
GzUMz2Mad9YGRGuCJz0shAPG2NFcPlr6zLWZACjrcBiJ8kMpWlSEzKvGgUjZRxyokDR2FN00E/bW
itQxBDOw6mDRmoY9q/MV/fKKN8a4TvmCDj8wIKOvLKzuCSicFegc3Qi7b9fX5mXs0lDHuDAYFWmr
881TlOE1c5ZXrhqQGs8sLI+psZvQFI7Wp8G8jN+1UYDYhFYwkYINb277ibt4cjXvuuKJ9Z4TC2I+
NK9ghHeQhE3/xiJSeyhrwbx7CJHqK9TYDciOt3xi9DILwofZdSgqvhpixMghAk1mbrg+ChilUfef
eMsPj5l+l5/4FrC/SM6oUrbcNHhJhtM4go7DF8095fYAMiU/THdSaqMvU4AdAgCd8ObhppYAjJeW
uUMaKSxpo8Tg3WiGhR8mRP9xBz48Lv5oFo4hLe7C8OAyXGpugOboR/lhIOfr0EXlCZicbaCDemGl
sSusGYGPORXHCU+uAZ0Vc4B/HV7W+DlwsFkpAjNpnx/JV0ipCMiN3Pfi1PCkihI887kaHMzMtk9d
PUqBndjXqX1/opTfY1pFyxse/DNLBvfTzNV8F2X+VCxnm0RY2KFukxtUt5lECgb71Q6PoLV1SpOL
ZK4eiYgyW/B1im5mjmpQmopCOat4RqevY8XoT3gO4R/hTCHnkRC7Z1n/t9QEjmdfOasvOy1nJWld
92rpX/Ms/foJBBGkLrwMTk8cdTOJi50pzAdfh8FEHDfcMaq4xEPk+4IyEg2rmBzdBPm9h0TlgGAT
ZTClgFQAKPzCCpbY3Y5t/IAm99U4DKTMD0Qwq8UvQOUWJE2hN5PBk0XIqeBsC/afQQMp6uOVSVH8
zdbFLHSXtZHahFc9X3oHsZTpSKGGPn4mQQwz89XH73pFvxBO0saohCjXJ9DF59gKrxjStpbgq9Vx
259NbX3DfW310+768rQQuDSfyoxn/EtqyvhzsQaixrMsju+mJ3uwaQy5TPrjukmk70EHtyiP1pXG
ZqrAr2S7EzPEaZl2lod/SOogmnG0APTFga1sfIsjg0SU2/RcDb0cYtKrJXxkbZRCkKB6Yc75Ookt
3M2zHL+grMH0X1pHYXX6pM0EItxkTZ+hou5ZLGaG98XNjU9AaUCC827W0BDFu1Ub8kFg6cPddRx/
uVUcONGceIt0rmQjWDmW0nJEtWQJEks7/Pu1vd/Ir/zw8ikTlbs92LEtLDtm6LNde7qPma4FezpX
CgwVSMJScE1AkoUy/JgzUZL0N8d178LVZ9JzVl5em9cLxcV/Rqt1iHQPVYHXxbPc6cPtvPe431Gz
W2gwLlMQlyRlnjlpIUYv7o8IVUahqK0a8s34YvtO8lRdlDTZqLVcozd9kGS1aIHPuRZBk7O7aDmi
AS0xcv7XjiKkw9LiUv0YaVTRZcM0jRGB1d8Q1NMJMYWriaCDpBijpW5h/+myudPzxdCm6Zerr4vm
AWGSlV664cq67yqU0HsANjGVOOWlvOiBAxiXgtDqrTKuHjaHtWyb1OwQPkJixeayrFEMPRgIozQP
rqIvJQRl5o63HGFQQp1/ZTNKaHuG8bNEytaOP3YQvc3Ggmp2gFUWy4FW0gehwnea1Qn6qdL5aXaS
OPDTYhTeg0Mod8kNb6A7n8GnFsIF0i981tTn4uIDZZA5z00B/hzBpW8cSaFOyclRWZwL6hilFl+/
AUkDq30n7XUIZE0c/qruhhdxvjSJhprOroLhLf6RDbizzjupOnhoKZgyeAHHszSzfC0u5v+yby+H
pB8nOfTGDSFuoF1gi3t9eLfi+igtrnW0ubw+iht0JtEhAKQ9EK7zS8gxb/mLKe+dIRLnJgKlKCS2
7MWYGViNrd3pNlMgKtj3y59pfytt28WIAwYuH/OFSs2D6RJoqqHpr2Q5+t8c6uDOh8aNNAg2rePP
xwPcq575Lk3/4EhSDvFYZrnDDQIlWxiHYjSIANEZCupLg4k9eZU+hEAKwooKkFs7DbCMAuPFFn+J
P9jyVj3QEI7Mh59oQ8uX54XzLQdICj92io6nH8oxRnYMfo+wGm9mBJCqPO24Azkb295Mmcb5Ph3L
RUAjcY9EzcJd8AbfJrD9b9ZnM1YbmIvz5T6DL7ruNyqSMn1oP19yG+MownNvszMKd+F7u8L2kYgY
6muU99cNBCOod2Rv/oDqxpV4DJ5qTR1OLIVwc2s0UroLvJcpIJvE8dvQ+Cle6Z9YSYH0zfBA5zLb
C0l2i+YhvPI+sgP/buLI4wv8Vd31Cll95tR3LRT0CNIq3IAoBsZyTBWshSXu/FVMYeRCbSNwD1kH
Sil4KRxqX7/tPRxPwjxCTyZbSTg35B6+/iU9obrmFxzi7dfvwCQpplKO25ouZHg6bhAmOx2r54Ro
gwry0dZGIl9yupu+bPpEBVzpuGB+6931jKbxtBGbM/syn35uGlPd9DLKc9WjHUlH5GhQEF44Oluj
mG228okXji2EApESQK+C89cJ/pCG1i8wV6F2xtjkwwRlHp0W8oqojOC7G2YUCD720Giu9TygvrHs
+vp03q1V6gqEMt/ivOnXZyNVeMpodAvMe3Ryi0lMc3N+9G9Li/X8k5a0t0hvfyNZK0/gxq9jDwE3
A1YCthkrm9r/JIulHV5+FS9A6plaIuEZXta/rfo4ZJI1jis09IWBdTMmWO0koNPogZuPjPWcJ3nj
CtsVBpvDTrIbwXuuniqNCK/4wlCvZtdPo/4FuKiIHwlXZTB6iu/oDaEFsp7o9m6maG1auBQAqLvH
QhWBa4cSaho1ewC0HJRsHdDnnw4sP5/SbsAC16dCE6Zf/cpZp9lGabE2Q8hdxjd663QPpCZ9J+At
zIgy50O0FPJ6bUmlIWXHf1v7WgYQW/XfeVh3juBf5GScttxAvewRrc6HV8o3vkvcP5zNFTPAlFPq
wpFvrJNtXQcbrW7gJfUAXb6Gi4YNd6C0qUdlCBUZbaYPjsQjt1BU3w1gfhyCDZgafbsE4rXpn2Yc
k4qtQGhksscRm0KM1k7rxDlxJaUu3CiwMuHDsk/idvhmcqicSIxp1QyYHNYWZ0njaen+wQ+/3ev4
99rAf11t0yHCfb730XWER9RaPGgkKDZdlbWgrVyiWpNTiRvRyNeOmNlfsDOkVtIxLm1oIWLuP5MY
sEhHYhnM9k91Nd5Oc7Gm9KYUnZCNWv1x6KAWwL77Cvi4q/5Ia6ZQ6OXIOhI7BbAkcJgjf/CASYXA
JoHWVmY6sO5dDA2H3fU3t1Y8kBBhvJsYfPeQavea8i1Sx85BMhVMsJchKGy0tVAqsJf75tD9oWuR
PDOwK5HG1KIlkWJ2uXGpPZrJDaYjBsP4e6qXsHqFPiKVZewrE9OuX+LyFS8V9NDIJbr9TfaD5/er
Z+us+4Xe8d/GbcXlMUEDLeKXYP6jC1xBJwv2o1AuZwwc7OvT/wfNHmRnfYaCoNTkO9+XupgNZfQv
Igp9Cn3k7qrKz7B16NIjd4Ax/5qj3H8GiWhzoAmiHBF6qVsCSzKA++BlwGC5gI6wVwd1EMB2m4kd
8IIRcFPJIy8ASVdgEOWkw/pPgvEeJc8Y4Yw/D95B1rDu16VxI3Wc2W8lFc3q2vdl31hAfHsKMlPC
i3SrQrTHvG5D9auD0aeDcnqjT9P3KLMjop1O11kGwprCdW54XGzPquUf/zPO7+J5HGMHKRK2WYQK
1jQvN71YQITUzJda09y2ihXhhi/2azyzURZz2fabdTfgvukG5Un0U+ejxEOt24eCvTt3mJXSrvkT
8fOaQE0okES5N5Dn/cI1+nTDBYMVIqzxaTPHSY7f8uDHPUjnLa9RrOcri41YgQfZYQRm9dGIaB1L
q06jVxbNFYe9k1VFh5/PldKJqli+HgpS9wjTMYEu71YH6eiXRRLHr/xlzMB33doKkqMnu0tl95ID
8URimD38mG1EQJwxKEcsmSEZ8+kA3eGMBZggwY8FYmlahq3bNLi/FoYFzY0IzDrER7aVQ86KQi9c
AtmickMZYUO/pLwd8v/Zwi0gch/TVWNI4VX1/JkIuhVXujZQOizOv7EcujuQbBAyCw11r6wmZefp
cm6LI7vUDvWLl2Po4b8eRzMV7CXoQxc0NkxzU6ICw+b0NtHh7tWebtAxlLfIMMNA/jJo37lXZ/2c
cLNojDkcF+QNjyIFZ2TzCqVQ7JZLUyv3GAwkDtpXPL2loKGc5H6jjj2mSGWTFD++9DcBVJZItMZn
9l5VFpCa0Jzc0gDd2OIUzJQx1HRmPwOjK3BNJz0ssqmzAzCSphso+1sQEibpQTZCx9itxeNEjnIj
K00pSyrAeVDhYRssZt+gVZoxtMSqTayFWy2qG+VfGqGbP4ACzjepqdrNkSTC5LhYPBmlBPtSD04k
6EeN0CBDe+J1A3zow6wQ7ZRTFGnnv3lN8FHNIiXoz2k99moopESGlBAeNYpiIAL2XPE9pSUHBkl3
0bNBrC1jUeu3GZJyn3oUuzeJA9/NHnwc4NL2l16hmvVPD/uo2QqArR8/4hIiU2ewiWa2IyGlQS9l
rU+JOS5iGF4SiZY970bQM4JrZdgE/oVmKve+AnnPzBiTzXZ8Qk5Mam4jzCCb8vZxRtI8SFugb0oC
7iOtmYAFxmgbac/LLoPHzvzcyitjvb93+OfoW/onw7DMLinOpUAsceFf9ygGFgPpIImnfrjlmWFU
z5HzDueZz5lvCDz1l6DEboX6sY+R6ia/9ynnLdvwyCl5AgFuB1LZybyWk080x72OsWK8T+yS4hiF
+9mYAfYT8B7aL31VUxINpV19UtXW28ibrfKgvOydididwdqoBXPBTj8PkCY95AMxpS1VTG/l16B2
ElLxiFmzLtV4pWWIdEQC0PRVYj0wyfHB2z3s01b/9DvW5U2dZWDZ2AR0mREtJO8yHcd11v3ETnh1
iAHIlNB2pRj4FumqtPnSHcawbUXS9IwJYe2nRQmfWQaNJnh9/ZxIRohFWEgPErekQdAmFsP4SoJO
9wuxdrkyCVCklCwd/CiXvm26tzAutTiJtvLhwcohQeJXxrRGKphT3K+7HFQpUwus7Jkz2ulInzbk
Mw12lGSeyDBFAmCgbrhryoK9wmSL0Ihxp6CTP+PHxbYl9N4QExeMME/KLJrILF8yEl/4D1bow+1I
npaM0ht3PFZ8+nEI+JJvnDCG0xL88XrILquamFzMLQQv/EW6e/O62IgsguZsVZrvF5vOBC7Dvhai
TzzfIlUGjJ1W6SGgvpnIb7B/ESc0GjozYtsIXGxrSB9tsZemCCWsp/Q4id5u5+HYNA0CY8h8pUbm
q+ddcvnRgeKexcA3yI6dTF72Ayogc9DJMEhjx3APTUoiSjhknxv6YPpZMKbZTFpWGsZX81gKvS5D
Yaq8HDu730C9wHrw4kSZx6sGi5doE4bPq5vNbUgIOFnS8MKPF/eLAY8XD6IJsQmccLnjmjemtAbW
Qg17IVs67x57lRouywaaxzwYGVlXCwdCM81qJvj8eWActpBqfVhdWXNXurKWC+CY5+/GwrKd5AQw
Mh0AA72OOX9f7vU2+Ny25YDprAbs0NbqrsFUyYDf+wCHYbnWIhaaf7swMxQsiUIytHYxYVm7ADDe
XfkRwKQBEOQ2oBZ5kIsrl+HscIPMMtdVDSkdSK4aKKa8YYMGcelSN5Br/Jqc0/K9XkJRgUIxQC6c
3NWJvA7qeZ79X8KCPPArEHP/3XlUL38qzzAnd+uW8pOFjvPuv8a+dRxOYQt8pgP/KbLlogmqnsPV
0A9VmkmwJRGuK2d8OunAxcb5kWS/DPu+lShYe5eYgyODvH3qJgVSBm8lt4jWcsaWj/u3i3ZfcuKu
2yv2ekxm+qu1nPJRAIIgQiCcb6FLpq6vleIkh6AENtd2pS+ikthGEHxWU2G0QZdXf5vpjJ0FMNb/
lGaDnC1/UXYId4BBpVDQ8ywS/xmrVWw4HH3thFFY9ed55nvP4xc/YRc95usoPRJFvnCql8n4i1Rv
gYsmAE/BOzcm2cznw5pOYo+jKWrrfGcETzOwFA189J+OeDqDz1BJ/yPXgdorZfgDYSuzCua0bVmC
pAIbdmjOxgJZJ3fHenGlt1nmjpqtcMgBSKU4Z1u6hwfcY4HsTSwxHxUlESXxIx9bdkXtBmnvoc/9
Df0HxpTsr+6lWaWuKI2CUo8QgIiSwA+RoL/xN9C/fMBez71I5MRfi4Vp9L5D0b8ruPHiva4kjBfg
4ICN3wswRIQD4171nmmaXY9vQixyC1T8BcjL2BaNfFXtI26wK8cEHC6XL/pAgvQT4RdWUyQFjlGh
iz8sIWMRcOUcGLmTjlFX6TUgWhVQu5TYqP24lvTVwXHKOmM/3DgZ0BXfjPsDOu+Ctb7ulqBs8+4h
VLMZoE6tVxDZ8vEEIUMwt5Z2AUc5TEAEFPz6eYZGJT8IsOeFU0QRvBCAB9z86J9nli7gutLW4rwE
rPHBx/tpnbgrpPyB2H32y4Sa2Vy5IyKgNR7moIJrWpJVyu9K+qu2/KjcNykAEZ3focgSentdKvhk
kKVXYnpMaGVXV4D2aiZ45EeMBj5XPbz2nguWqTvdMwk6lh2+5zhtuD0JuVENQH16LBrNoiv5atdV
WjZUq5hQpWWFvsjPwdenxnfdAigz2wFiIEvpYyZSbH/zOSr+j4hxkGY58vv1jwvnAeq/v41neQN/
iDgcAs6gEkLhsM4SmpBnl4VxZxTiq6oMZLukEQPWuepYMDpRCSwqyTZWAbf4RPYypyXJnodgmLZE
j+brBG4MjHN+y0/wO2C920lONM8EXN+uFUmbY9Ke4H4/y/M/0/8wNQZizUk05bxfGyanGKJti1rG
8hR7GKuSR5NDUBW3zXwd1tI6zIlQgv9GvGJPxi5JRVMtgBkXj+M9K2nhiLXNWj6Hn3V5N2e/aVZA
0CMhacAkeDlcKKi1mBB6JAeKMPs5BHibwGcelWevpPOH4CKEFe8XO6PjVZSzI0cKOzXvdGp1g03D
PRkZY2h0yzyr+3gWi50pCDHgLGtj/lXNvvZPyKUoX6xa3CRWGHotfWrUIRJmHIg3TMuxkpzMH33L
x6eZ5OujPEWie6v3MtUhOeQtmU7QP2Bl5P+zP4wPzTJWzi4Cud/zhkqYGumjaMBid1OrjANhBGIR
/VDiR4rw5UAHDEqlvVCbypbtkff7Jw3P5z1gVMx6cilD3Sc+H5al2ey3Wh3QsUaEmJBlnFYo4HvQ
ZoXl9Ku1ww+BGG3C5n6Ze9Uq6oqQZ9pEOalvHYihnix29TNnS3DPrB//bhttrnIackcFBc31S6EA
iBk3ypgfvuTyXGU0BDnlHR4b3y2pI/cAzrIPFBu8dGJVQhEKR/mZTC2ee77LrNhaWkKLfP+sCtc5
Ru8caqf6NZuRgkJ4YvpW9qmgGZrAU459/GalwxQ9N8KBLyGvYtjNZfy/x9saICWLuyK1f//wdA2z
Lb6Nb5q1Wt8U9ugrWjHETxp+n6DrF697ADAUlvLkr4NsHnUPqhRSK4nU+QWETbDn0AbySR6yNQIp
JiivPhzuNhCarnvGfBJLBZCB4hTEqc5NLmX+cHeOI7uq2zIer8BunG/uA9ZC8k5QXWEbnylcS1Ia
uVUTnihcjmj09AR2bysy37g8Y0MMFkOWI9hw0wzIOd0187x3NxD+CPIoc4v6jiyyw5Qf6YjBh296
uokHprHCne/Ilx4MiYTQmrPMODad8gIwGzZPMRL1rVFVPaUDml2dPqeTS5Z9OAzCAxjNdXUdF4TO
SzOEplxRz7tk5hF5l/9aKzD4HShCNkSazBB5/8bBpsq3p3TG74iBgpbrhgu1xzYW5WYN7Sns0wb3
mpRYNILWE+fpaek74uBJyj7UmEolx3aiyBttcL5YPOqYSWPF6rS/Dc9wtsTEOhku2GxYnJNi5ZnR
sQXeHCgNY8Hr6HrpvyXr6TadeT6h9J0XCsIaH/MGBSasMmZ26RgLyOXtTlxoiZKVD3HXTP12BIS/
cQUd/wXZD65Dk1WhMQ9G61LUehZ32aYX/kiCiE/X7jYn6Oq9avCMsgZeoMPoEcg0U97CZkTXMsqP
OGnAQ4l1R/J7iuT7pbCmPJPzRDhc9whoMG4XZXJBsi09AB+4DaoSz+XnB5ISfvss48/4S+mFDDS9
OPtjZ21UVCcCj/dW1Qgu4iziRRfCFU/YJzTPjscRKrkr/OfwW/+53kv2NLvHrnk1jdqXR/8bTVVA
4vdyeW8jGJ/xWvNEuIdX2iX7xEF+tiXd5YkJwZC2ldzA0b0bXtq+TOIJKNfcVqzqtwrt0lJldH9s
aMC0SJSFeUR/ftflWhJadjXJ2UmPr5mo2qrMepKLlep0LPw7OjRepz5hfoKwEbiyuRJn2Qdf0ugq
m0DFVvzEzt0nyZe1m635XHDz6Z9aU+D7OQodHpCq9nen2aTRdql1a9hVK1fhRwBFwpugVnsEgRjV
fF7s11RuHk7oVtZt7pOWAQj0Me2p8+TGy7LZ/enHt41Di4qopGH4zjs6aeGck1pbYhLeLgfGR/mm
kmf+SGuD3VR4HrY/Fx8Wq3bEWySAfavTPQpKyI1vgJxrgetbg0ZqwM8yzKsELOP3pOC6UKl6lBhP
RdMbE51OmVZZ2R7Hh9r8GTZauOnwYa3DOxRJDCJEhWUgKFKm5cR07i7X0S3Q3OMx0EqhAJZ7rhRK
Roues/DeVwYRT5+8OpeAwcjD6sOB4LvV+ZDcOxFDhBiJtjjQJqayKx7rfOnNksJhE3J4XysLvkjp
OrfketwsuCb+kq3BXW+C8cmDDrSDEfd98kpp3oboJqbaxgityyogRGKr2iQDgksat4TOHaKsZ2HM
CSXaLasiVUr7vr7uIpnXymWohE9Hnd2wUaqsbIkY+Yv9O/7DBt9uwChX0bY2DtPro4XApq2rpZxM
7r4QNPheUpfRLaP0prbLRlTArz3zAt8MT4nPA0iOLglpnl2YZevFky5AsR2v9kQ0yb2BZ40Tsi6z
Ajam0IIj2Cl2QrfHMq/MCjAIM1jdgQXTxAYljScAnqu6k+5frjb3152lm0if4dUJvo/Wf0HGUrZT
fqjqua62TzxZifvq4/c+Xctc8DMq2Gl9hwdrOJxjz4uACamhkssz9svvw/881i57QqQtKzvEirlP
2s7kQ/zEUnZ/68p6Js/W7xIeJ+Qr9b0VlkiEfGQo4ovkqPlWUtpFzmVtiULQX60IrYSsNj11D48m
uT6LLFqYzKWFeSChcZae71omxXC6c9MITQjelebaEGpGm2DDxaS75dfdapZ6WrSDRV9roSw4CpJn
vf8KDTDYhMMl4tZh99DjohGRi2Tt4SUybSrRyRhO0PnIoDdmQi3oR16CYm0JoBFspOgZ+erezzhl
eKpzoNbkP2Wlq7OSqA6UiRMq7CKSWNYPosD3bUDCr8IDkAVycbQpwZwt9nbzHs7hhoY+wjUhOpQO
ubke2q8g2eBNdrLjtr1jVOpLKJbIcK6Af+i2NRPW+eVCO/3tyt+Z5TNg39bdX6dFY3UK+MIyhiFa
fDiGakhq4xG1HD5fPpe5QKJCuJ9jreU0M/YTWj2JK96qiWrKdx2zbYz69bSxVEMyHvIV8+z6ULpC
U+gnN74OjrJXD7RzIYa509pj0fXwaYbPO4TeUucUn2A6qstFCkvIiknMo3Op9+uOu/vW0gpgi26h
9CgWNFmIOU6ip2bYF2XC2o2cT1+lRAijrOUVtZ6kRY5j52oZHSInxy8Eb6RvPiXf/tfwKVmvw4j4
s5BGjBzEpRXPMplkkRDqliyBm/ElNq88uOhyZixonPRoOK8U53tWETDNWqb1/g3MClNJUhHpEvsy
wONwmrEZj1vgLNMSYY2GdnI8SfwK6RA80gq59C6lDgk4718VWN3rZI1rbqtH6GVsEgTJ2xFokjTG
DmKKnUEdo3wU92kG84N38Z9f2Wqml2O5RaKuwwClGEAmBUT+mFiXKkts8qVa0A6veygPgwUwNGNT
kdqi237mH7sqBPsAl8vCDtvpXJJDyRt4VeafQ6rBWYhJs8GtloL08kDcYBJWDO2xroiI/GLUK0pw
HRIuwQOUqXx/ZBbJmyelNUtrInRu6qfxmwFkYeCwOMhX2LoXIQipiUffjyIpPj4bRT5QdZ1XN2dX
9aNDdG7I7rax24YcMFodRQ2w+VqKV7rz7j/NjHfcKjcGVKwqmV6fW/52ipu95KqyCSKSGL9zSd8m
sHty2E5WD3sm8e1D0QxzGvbDVZC0a+R3jRNyhSgHEL/V0uesutgOwjnetsearLzcfrbuYXchBW/b
H2rbvKZsH11Tp2ZRn5J+ZGxSm9vYIWs2sa+qCwRKyk34IHDLBEy5ppgkkmeKKXX+sUw4Puif+JLS
oigfQu5JQ8CdNt+jF8JAYzsRxiViONFcWmU4Lca0pJofvnw8zNwSZB8PkgRDyNsFJSyADJATz7WI
AUXGpe/6iEmb+ldCIw3TNYrvIrIrWlA8cvi22tyTJsGNb73qh4djbHq2d4R1j5vZO/IxVXTdCZMM
57Zs6uyv9L3+Lftcm1Kw3vmExaA2f9enYX4FsQ3UhvgM6RJUgvV6v/rRl/AIW6tospmHTCaFvhTZ
jAUaFzJHP5tRdG/uLhLBl0oSC+1xc2QVeXbxG+f+ZgL6QSB/0MEAoiLjwwmUbnlwhf/tCQTueo/Z
X4w7ZSLn0q+S4UXraCj32mLT1zxLFoKcsPtCizR7YUp7gF864zzTV3F0SUYDOQmmmWD2RsRl/iAe
H5/yHPu1jSirCuz9NAmMmY1LvDYRgKVfbSLNIrA3NOCvXDfNfhiWqVlKZSdarBU+97Ub2+k4/xzw
sbPYpN7/Vjjayp57JvtkEqy1BXhsdknG5kPNrvll6XcrT7+i1NIvP9obvqL8zXTqux1idbVsnxVW
ICc2LQH4sJFKIH/mhJ7i/WridGlw3yq7Gvme+dv5S984qlKDiHT+/wr/ddJVuw0GjCTTjMferix9
KeWNECGS+XmaMO0KN+IoLwrcmby1UFYVgF6A7VIN5O53HII3WzbF0h5gHKoWKHngZ/GZ1D1vbHjF
WdUOL2S8F9cjxMNBbIrpRUQXITA+1x9Rp2XRRNP3hb6fJ+3Rgv1XhcE4rjq9/O6nIgu3hmFTVyQI
8eFVHrwXlqi+stdFAiX0ronCujeHocyAYZfEvFAnRacSPp2uwSZq6OCbO9mhsfmOMY0Hfu0uLRW+
HuUNNQnkN2JZ2P/KrD5y1fr+WEe9ZTX4n/OVBU2ec6fKZHAT0t2XUcC6AbRCHY4KsiEFwi5lavRx
0Ie8eKRuIgikZSlBILXLa9h8BUpczV0J/OC+Rfn0MBr+YPsrslczPYW8oNUSbHmil0rkC97JLuV0
CWyGJ+lPMOLWF/Rbs5VtH0EhaU/aXn4ysYqkBMEvf6JPZeKPw/9eUyDwjXQb6OIrkr1W92MbaEBP
0FTxwyjIiuExv80TtsGThvJCBZ73TfrcYDIxwY0YJd+2a+YmfuiV/2JqmIHxgsSZ2YFH/FLs/Dt5
YdP+MV4QlMl6sJPLVp5JOwHepwHOE1iwTK9RylWedoRyAYU8qLeRpdVfQJoT0cbLGEM7AtWTJhPx
qJAZ6rG5tVaoOdNf4vk9YUUQ5swAK9KcfzfNpDmKYyW/Dzj/MP89XC2JN0I3tzHDTdOHrcruuABt
VJTvDXgCspS72zsUW4R7wHJpO7cSxuht4VweF/V87XKcAZ3NhpeTPOaGQisalwnJ5mNpVnzzW+vU
VtEGTjylguvZu5Bik1mowIEAMXMPS3kdgWux8yJ/8q9JgoTgQ8rJwwXhd7K1WrbANrLSvP83Afc+
/Bwe2lEqDUL9P4+o1Pwkq8kL/3HEBFLnw+z5y2isxtGzKvcUfX5lF7Gz2q+CRGrcWYMD9ah4l586
sXz2c+nj6XTOMdjTmH9MmPPZGIVndG56Fs/kYYXhgKDbp33wmxaZQeIIODnXo1ObZ0Fni8+TwN5A
py74YqmwQgDjEDpDgFZWLr8SAu4JTE6epQcUvk6lJchzXoX43hEiO5USScJD5laBUNS2+1NT+Svp
D2qKzCOlhZ7fSY+ckowFhHi/bjQDRVI/RJACZkksVgtTJ227yMPDmL3xPkEkGtiJ+L2QO5+I0B2F
/bKwNzqvUX2tJSoRZkIzAcfbijpqoAWCkFjYlpm1ebyURvhz1+sG2CWtkVWhN00M1S69IZBZkz1r
OlenXxEz4oAK7yiSUb8akrs7AY+KzN3QQzRq6PypxjhmDthP9TfPFRTqyydcBdcSsK0cMSFHMzAS
GtaX+mWp0DpEhC14NJYLu3JCH+ZFL2oQ9wqc09YURC3JTErjko3YVLVMwjKdUWBrQPRb8WLFUbT3
i3xnQugaCxrPM/PHUFmd6DnkjYrEMAL9E5T1SHNkA+zENOaNlUdTlr+u4forcCBEgNUx9owtwYVr
CxT8riTSNqIduWfKUK0FeFqrQiwOAE4KkUr/QTLBiRWEzxSWYel20BsVAoPjxrbmYH/tzib5lh+V
hlxuRmg9u3p69gLG0eBh02+5S75F3OdcfaH7DcvDLkewrxn27swFn2nXtzut+czCT5ZiLq6BBrW8
3wMLbcx940dpx5y2zmhk2oVNM8BqVguy4/Wk5zZhMV3GqEb1BEnAh7gmEkw/u7KkS6S2KhwtWjDV
JgRmqk1ZorZqkt0PECIPoZu9cDpD6bzQqHZ4zCZ+RvUoMm6+2baB0tYN58+2bUyT7YABNBLzB2oc
fFzhg2zWaEMQWfkQfZ4FvygLldAnpuNfOazDb7jFcw3MsCTvxWOcNoxdb8+l/lsHWtoNrCEbBbqc
uH8Gfb+qlGfs87tzrChBKTk3Wt4ygbBZE9vGTbcAoYfX3oIZXXcDtgMcYVXjswI28y0+DbP39eyd
/KcFNRRv4/yaKWJUT2qyeObwMurKIAbXca1efXT0wJDNLeoN278VzGwjh2XMZeUFhR1sKWffPm0s
dtDmhbRsV8au6L3qp3f/8XHoHpcED8m03lMCH2F3Ry9GtrUO0N9rad95/YPKMVunPumDuWR+X1wh
F72dfUEs2b6ids+CAaf8tjiLP9kCpZ9GNpsLbXPGitNsn1YZ9O9XGJO5RvFahdzwxvD5U3P+U8ge
l5kggLFtvQ9TgiXMMCnyAVs/vGA9iwxJod4dBkT0bjzvfq2ajvpk0mArj8OcSPhBlQ9fun8TRSPs
3l8AUD8f8hyb+pWEuVeGVcXyKFmMgspKYXWdgf8Nn7yjSf58+of1Fwqz7DFkNluwCl+4zNC99bDO
4UNvHLh7V5UMMQBlAWCG+pAFjGbZH7WbQU5S+WWSx8l57r1Qg/eLZMvcNNPM6ofrCCU+uLdfP7F0
GPPhHqxcCrFQZ5aggNYSNrzYZf/+Z4XCErGCW6xRJEA1mtcFan8TaoCYZAs9kFNwa/rLZ5rAvNQe
SYg5D4MqEzFj9stV3G2KszFsqH3vBYOYnxCMj+lSEVC8D82+oib9BX1nf5oHTnf3EYwymBT1ee7V
ASygxBX2kdZRTLVDiOIdWFOyjPtpky5UYKOdWAd/zGmtpgW4KBzmHiv7kS00yIdyv5sQHl1ByLKa
9yFb2fpdl+qqA2CKlYFhiMBPqdqzZu44sIsvObXZBFLribWqt7W8s3SXXnyzltSg8AVQI3wJMARR
RI8lN2+BCyxosrurdU1USki9cAhLr3LicERgqODCo5RS+TZH6N1VqXpdBW1mqu+Gsg3l4XyuvdCk
NtGLH9wXkIyuB+UwvByMbemdpW2fnTzAH16Ixy6YF1H9aVX6Jaj14mIuIGBT+mfkLQ+aDVz7BbVK
Lv7i5byjT1XJ2VDwUYe+yFrvROEMdVj6ypPsJqg+VtSMMVAVh50srQFuhaVYQATc+Xh/sk9tCKlW
hNkmpgyHiZwiFHvxRF76zsCcPqvz8Ct5FZ8NWh+Apb8fi3MiL6gIbU/KWHnWxmE9fOn5LecPhfCT
mS2F53FdLu5MTOojrE1k/pba1o/nhd5sjumhDzNjaEbT4p6aia+lUWL/FMdQI6rsSqmSNOpBW8V7
BtSUtqo3Z8ZYvLpi4hhduo3ivIv7owd0Ca4DYOcZI1qsPhjf//6dub+eBUkXUWZVKvoz/r7RqZsf
HsOb3bJhhbSqwkwiEeQDTQxE4t7gfB8fb4bH2G8u9AEz8mLh94BHEorkVRuL+yte1MebE50bg37c
4qeT8Cmu60HSVgj43uR4P6dloR9qA1AXJxSZSklBM4ujs/0GpVh0dBZNMDWEpU5oxU417YLOS78U
phlCx0XBh+reINh8ZbgAtcHfMuthMtsa7yiQo3czGTogLGIxL/dYLmbqy2e4900SGY3IOm0LzF00
WgOsgDtHKLwdubw8OteNbydI5ZVrOC44Stlvy2ecVR95YfdCRfMNy12nVFgubjFDoaIB1G08RSNZ
qXoI+5XcRuYDrJZmV1Ywc1ltSN5U2X8vyn8ogUEl7RYLtmxUzAGudOLSvn+j7Tn1Qf27OFoBZF9L
3VTZl9oStahxUELj++F2OXQuGq7dzdDrmQA3Z2Wthdb+0yoQpWwOaNta4Iea+5Ka6iQQ9kBDWAUl
ioNvFPfNSt98UEyoUM2Ea7AjfGZjBl4zYU87IY13iQD5PkDaiLxCRQck7mxY+DKtJ+NRFTWZaV2i
FvGnF9eSS3LI+6wsw6Yxdiqor9WYP8sKzN6p93Pgw5jeyLXFljLRB0TgPhqTavsElbPaKi1gsAy3
rePox4e4I3GCXqFR6qGGTuZ9S4lw6OOS9lU/5s7JkpnhFKd/gLc5ECOPBI8kbGaiL9X5XZSMMPzy
r6T5ZMXSDJ2wnfZ/f45QUUgxnAmbLp+QwTaGrruaUpAaLaUYMKxWzxDdkmMKFG3iqdD/2eHH0beL
sV89scMKM7LORAl30Vtj4jt6QU+jKx0pc82mhC4ssAiugpWPVMBnMwUMpOC1oTmKBG0pVNqJF3O7
y3b0M/INAAjw6CktkqRe8yx/zHTUKtM8OlJctnAxJaU38w3vhwqe9Pnk6aGVGvroyZvWES5qaV3W
EjuF/AmmDPQOHnvXPk+4GKzbrdEfF6zcDRczZvpgGXMPXwDfKFo7Rf/A7qts3FkJJnoDBvZ3Fmnj
RC1w3WkiUeNPnqjHhlOnat/dNi6z6FmwXinYthEYAkNMnn5jSeCu4vRCCJBvH5DDY+EGU8KtTq+t
QYnJ0fy+1llhi81wqguWBoiddFCgD45z6fiHOQq99TZ4wUrvdhBgPXc7ezicb35QA/I2kRLHBkTY
gztJNMHIe+BgYVUi+85E2+Hm8dx3U7uY/ckfjg44q+EyN4WJHTVelGDPjyMz5yubRZXcLZmrIDu3
1EEv10K1HhFeLn9rjZJumyfULFblA+Mhcuf/Sd0Now73+rNwi4dLeKqAx/0C0zLyhv0uznuztuR6
2hUOaUyysJ+VnZprGkby499+UhvCSuIL1gLKX9Nvi/AMc9+kGNL1NWReeZ9eSguPoL1/DbVi37ns
ARjHaAa8X5SbPfzwHXIrN+1uyuEYJd6zQ70KHhiydcvf8o/1M6jL9Npsl6gM5XVZYLxYaV3bIdvz
WInCtkksmqe4tZZEs2fnYj0AfLOtxfSOrEVeDCED4BgcHmggFNnna8aKD3rz7Hn6T4drAo2ZdbAY
lZuyMJZmcU+zrry4luj5VtcU/+d1BtoYz5wt+0W8hgaKyBJlAfH3MuoSYfs7/d9UAzNgr8cZoaa5
SMhUqV269kikl0rJ3MW5pogjWskY3rk8yT66nMnvj4BdZS/3hlGOkLgi1joXLuGpMHSrk236xKKI
GJjQ2yWQoRXl7uV1/AwOQPdZYi85soH3LsNJ8RFHezWfT9xc2gUn8CZ3+mhRehOA+Mw/48xr7m2d
BjoCdklCqSVT9AF7Qhopob9N4z2syKQ3VKLzrs8/uKCiSPfmBTUDx2ZJPhFrKp3TM00APZoaUF8R
f8aC12tPsvA7N+qq3ahU9C8KCOQHpahLY2kT2W/EDBk9rJS99MWKU3pOfB0Iczm8Qld/Tlup8t1c
0I7O0oLKiZlcuj3pKlm/bsLmHpKsguQBAtxkKli/6/ITGAJfBQJBskGuu1fcUFvhhEzLgbPMcNJl
WvEqsmr+RIdIVYSpqbcHote6hzKELK5gGMETTmEMaaNR1qsRrraJ03IJiblXRj1LPUTLerlyNDLU
lJzCZ1uCt/woezqVhAS93e3wYcKSDOB7mRWYq/Umxh8wgUqTFKzgQPcXsgqBzw/EudQal40Ii1ZC
ikjZQqwig3nXJnbHZZ10JNblYIw5ePCUW7O3CrywYn9M5CDUVU4oOsPJ/2EH/8IINRQc9BI5HOXx
Kfv39wifhYa6qpcxszXZucQFisE6vkPdaToDE3Hdfg8ljEkeWm42KH0ncvj4zNkWtDAKN27CaVG6
1rlfzqiHrLpT3KtAsqM9HDZ3Qga8Y7ZwJzev2vMSdkq/1qSApJiyb1I3ZNBFQ2te42QZ5q1LAnfr
OvoYCkPyuU033kX5H19FsrDsdCXrszdRQtbQMu1boPM/uctfd2DzBaWhpkqdbRwYoi5xdS0Jkdbc
GtLZIAdBe5W+IobWRf0kIQTL2yCZjHVBIvUuv38i4/kL/RJ41OPHtw8tbng1xXaoiStx3//4Ul/X
e/KJPWGeUA7Bp3/LJ2OfQugmvH4eryGMyClgCfQ+tMSIZx6JnTfvw2wHgydB0dUjbxgdcEvGCvF7
a8MDOLI8X6V4hTi+0G7uZvV+oYnzG9uZ0kjtt+qc6BLLLBzrdj5tHt6AsokBtrEvqRe2ubfDTbEQ
z+S4vBANCwk7LKNGhq9lSZEW51/BkwcXjzNlgwE/cynGXvk0E7N/z+4Qp2KjT7dERo7oCNl2tCVD
kIylTSZAaEi4BWYDqSL6ap94joDWz33XAVOq0OUHqgwgTKl+6PspifVs7PWkNeAAyYf6l9RAZe6V
tyGgfXCecU9uHs9s/8Jw1SgbHMk0cKASD5VFquOuj9UU+uSm4v6WEKns7FupfXANN2Id8mJotITc
3Sc0ua6VnqvBWayutTgiVTzvv+Brcyv0TkJT3l7egnKWDF4ISelj1lpvlSneI8pU/JL0ejgXFCnM
swWR79wAZkzsZkEz388YFW/sSGLrpS/ngbt0QdlRr+UwICH+jF+grZ1UupipBPMrQSlmMpJMu48Q
rmowm1dzZnJdi5DH5Q5SrgBEiBBX50G3wIyqTgfrqqLTaUiMTYF7ei3n2XyaYQRU3ozS9Hf+KZeg
Tjts8YIR1kXZcYA3qN+KcAZwkrDiubnoUDQVh4vqOR9JXpvedDNER5QroQPecrDnbnKUPBB7wnmf
XZZw66oct+vx0gSjiSnvge+7U4E3hDzD/fsWjCTLUdJJtuV9gGZVYjJsoQ5KcKz8+AD1ZuNoCr+6
ybB4ByBbnUwx5ACgNamIVR2zcsAMA5FwMXxxvpr21UZVyoB9WTCsBfihV1aU6NC9g7qFBRyuDkKx
LgVBif0E8Rl/SfwvTG7nhrWtgz6bHgMJrpRP782kYp0HjAnPsgbbGUvGI7nz7FMwC/JrzYs103Xb
Rfje7HWfdP+Ups4bzy4mtQs/tWepWfXYd+1qYMfn8Oc6/oi8t7pZ4Y9j0S97s1B64o45bmcjHpqN
lWRX2DxTNSQPPN5O7O3MYQQ4iZR1pnAPU440gghm+wNblb1kXQrC5xA6X/P2wsc5Hoi2AdnDe/MA
t2K3XPyoKljg3hitRCkdzp2Ivo7LwMUG8A+mJn26tgWuSk/TxL7t3QLTOLj93pVt0hmMc0igFwa1
1BeRNaW9drYqnW02jBQLU5cS0fkKpkbsbVs60r6OjUwPNEKj7S8S0H9/Zckm7ultgRyTg2rQF7ML
e0WVlSZfOp0LmZ762d2tOBW3UUZHtLnxIz6xpVBnqpkyYoHaszO9+pRUFPtZ9Z+kv2TQcOegCl1s
wtGiTSikOAABq9lmkru8jpn+MSf3l+AzzUVDcVjpmpjQbazRglVMENm4SgI5aO68KNK7zBumNDhk
OFA9CaNRSS5YNonDP18VIcFGPOACoP6cPI9rGfsdR/7FWVNtRaI6qeOUfaOMczx1i9EOK69UHEly
EKxSqqbEbJgBqGOCyHliHSMlPK+r0rNuIDCrUz+IBtrCqjzqkRpQ3czbOSrP/xHDxY2hOECSu5U+
9A7PXHW1vfJ2tOBa8BZoCmW0Y9drUW1nBPpBWX1tK2cQi+ImIt2vF/NJqhEXRYMkJU3RzJMb8tpU
4sCdscvLy/C6v1Cfdzugj8zYNFB8P3ugpYwB6rNMURtZzkFRizB+vI68ZA1xiHwHjTZ2SN20lhvE
YBmpbyvVqdJCTrWsH0Q+/JrvH4bB8hji9TFruaaZCJoFnFATr9ovNOdgicc7Vel5B8CfguUu5YLl
EvA0ASUmyEQ4mGYR7xKsgxyp2OuGtmwiRju5QouN6MVOVRNXzdoc2jtbLSizE5NfKPPOfxxvZaqs
pYodz/n7Igj4L2B3/OfaELFUcWp3hzKvm167PTrJsW2wkeV5igjLOfAQvLylI4DdptUx5XZXH35x
EtXPBquaMkdTxTmdZSNc+Ouz4+ZwfgBQnC+4MVrVaD/yEZIwISz+tQPe6SZ3z594+UxpvDjzDFZj
bE0AdvpfAcV3wQujRlLRSYTpPTNrbzMcqVFdPmrNE0PtvoGbgE0hsfybTfl0g9Tq/IBGkdcURhA4
DlFjuxs+4Mksl77UarvY2PCZZr8gXGTsKoYanBuYYvCQWmJDem+gUhfpmb5HVJwZuLeh9qqQcejO
SRhEjluKaQvZQ6FIGz044hI41Q7G75ksq6lVRUKFXCwWak4w7ipYsaVWqBMmnkk8JkEgPZbRxcXS
v1cHmqahQarGkE2KqHPI+wUmpHEfu6+ve+1Yr/71IJKvQmUbXV3OgM9Yhfcqu8tWMu4EKUzc13uf
dTlsVegL8Oqm2wvFmDtQiH91Xu/XQi3GlsnmmZuADrUKISnwG8vbk7AAnPATpJ/hy73F6NXCMu75
aYogIunqTifJFU5VtbkGuEcnJdmVwlepRolU9oF1mF1xr1IYCe3YVjr7D5Vlr+fAW6NCATr7xKR0
aqBZ7+CRaDbuMUyAmXcFL0hCm7sJOiFRCRBONRDNCDcH+fuA5tq2NKZGEm0kJhYyaczuAt+nXMVh
yKIbCd6gh4BwkOfdiaQDZl+70sxuN8xHmcdbsDuUjTX/YVAE/mcckvfhn6l6L6XMTsLDObn/u849
Dq97YFelQ/EMafMzWsA8OwqLH8w6AhqvTpPfdkDGq3TUx/xSh5bkXiSLg7gRafzkH4F89ClIjtsC
6L1A/XTXHvvVRg3j+8xYw8qHHKNuYYX0rZzlderPb+5cJHemqP7baRx7tMIZhC4pkDywZ/IAWVex
RHr4MwhGkoA01ryjU5SCLhgVwfMaVtMaEWjQYEtAh2/JkYXcuA0s9SqQlHGPBR2NLs6wq6FxCcSi
JSJa+bgIpa7GiKiTsHAEbvyxrzV6f7Ctql+0KFX+IsydjmFPt1wlpY/pVZN0rdKzkyoG6V5vokrL
aJ1DeYo2SsJL1oAk3x5gmR1wuzv+R2n5z4Z2T4L0FsAZNDhRZHeB5lcYrl3pGrbi09ufV/o401Af
8VVvT+v8lnjYqZGHXoIC5GwNtXI5T3Hp9x9eUs+Nd3n+5QQOee6iI35AtSZDryh32E9jufU4kiC9
B5Nl4E/Vm5K8394NTvjVPsbPoSbC5ixMRP+btp2ab6zFGbg8GSn/QUc89t6hI22MSWKhgthaazsE
jUn3KEmvDOKkvjpjiOU9Lu+1aflZBw5vJ0XuoonoyOIR1mGzALf+ZbYdXYDLa5IJqvrodxlcDHCr
pRQNsulF66W6K1bS9aNf1rvptiXNFJrm9MjEeXG3pAcRCmmsQCfsQhhWst91qBSJ+eHjqX/YKqZe
bUxaHkWl19Sm89YhR7Ml0GRcFVjN2ISvChLnpKMuV2H0pVBAU2gMM/0N8hIJUk/QCW3SF1X88k04
6jFaqGLn6ALZL7Xy5nsPW3BmHl08u0EBIxLkDF8QrWa9Bw2KMd+vs1ECv+OpQmLK3DnblBURCvHK
8DiUJyB85TDrME7GkZPIxQy1sSr1Ylz7NiW+8rcRsVMAiMLZ3nNvRSG2NhJXvTa2jmrLrKaWv66t
fL2rlJz+Ih1YYzM1qHURjHQpoRfss++LhY449jvPxn1dcYCyDisBTSksnEnofxCIM4lMq6hIEdtA
KYBut0FdMpmL0TytN1h2yZCz/q53PrNd8kj+EH2Elva1Q4Ii8QGN+4SAEIK1s8XPlgondVxNarYk
Uur+xmG/emQpPDHsPv8681EvCoHCFteWy6t7sABfdzuXVAA/EB3Y9TXelr+UbErH1r+vxfXUfnXn
M8IzD3pXM/mRx0qfAVW4ms9AMe+5+ThZCQk/oTU3BuTKfNSBjthuf8S8/IkBgtGOuEjS79E1BRV5
zd9AMxIFuKlaJiP+5UvHk+YJnsHr8zyCvCCBAmos12TXVjVs9H/t2RY96g/11CQh3v+CVY9WjUH1
x1RPWuXE7dhaEsSk4GlMMOA/t1PnK9wLkQcyGt875C5x+ZX1dkdwcQdBadVX2SlbH1OKp0yOwpxS
f1uktdTWdnKen3s3/GGEABAxwXu88/KwPQmgXzE06ddyZc0Z/dZTxx9IrLBsQVygsfwbvPQ1O86I
zJvj9TatyfZAZz1GNTYGgnqpN8rOb4Dw36XAiorig6183AroGgVW2kVNzQt9178bdakYYoT4A3qO
EC9rp/KxgxSIVU0agl3WnC/mO9MAZeAFqJmy1Hg4Q9nFrn1Rk9LE3nNwx3sSFGNr7y805llIPwKX
yAROrZTD4OlzPTFnfOaeXRiidvuASPH+RjRB7lC7n6RsRWDA51xJsdJzXrrRZKcwrKaD+63HfJdX
RRv04i+SYXPtJdsA4qHRO734K48q+s9y9zvU6Yv4Wb/S4BM2ag3mvY6tvyrTwm3FuoEO2gk8Smtx
NOLfk7sT9bfSSKphwVJdW/xooQlQS2Ei9pu9KaT5qfhzON8IhcqmYqN4K5E0+jb7jf84mthYZbjp
bBIWtTiRJ/nrUAMlZvBDtGxOMTomja41NekQYMPuMzyQ+d9pX1sD73XGuY/WwJQ9kEsUEf0C9+IT
NOdPor01hTqowvZeRO2ICCd+FQaF8cRbPyZFBGlZmxosv9vkaAg+s0lHZBJ6AmWLj2CKwl/46zvx
OmOPl46xs9/yaejKgy+7D2vW+NGd1M6zimDmDLMyDJopI4CS8DG2VRnyC+CANPGGHoAuWI02q5li
tSzoLHcemlbIdvX0nC4phQXouBRvOVglz8kUUiqgVJv/5N4ueGzdE8UNvZdUiK2D/RfkbvHGzJa4
AQS+HkQCA/0z1jj7fJRM5I5q3nWTHs71YLWgSHoCGxHod6EoVc2ey3r/et7G8BI5BkYnTemSrX5B
uBTONyxMZkJe8Fz3BYJ18OP3uhClpYI/20yboli0jNv5NUEcPx4kwlf82oD3AQmm07v7MUD5/+4n
Yh8FVZ+A5NLXOWj51b4icI6VRyz7D/eAQ5RAPnsUTyGGmNa00PdjiHw3KSL/5nT1OmxGw13By6I/
givQBqEDYexyoAAevtetPXHQLZeYMwzv2DMLy3EZXGv17cGDGy6aMFU+i3v0hhzIAUGwK3M9xKi8
nrPG+XqHg/83fqqdTD7/YA7g9bO0TdiuehabsQJlPFlv44o4ZIPB3IWLFDOtZJEGBKfjgs01jkD7
rcfNClDJ9wdkJ20kMfoLiOTCE75cpiQP4HDT3QrnPiM7yEZJV6SNejI7NkkdNeDGYqVpUbU2lwLn
s+JmaJUHD+7cqNXa1qnKp/gBUMjfngU9ZrzWONI/J81gFbbM1InWoQpUVjGHIDodBpJbQ71YJnHD
ZaBsBLwm/zeP/80Hkpox3u+vLBxwvRctP2WhJXaZkU6SGFbh3IPc7aIMtQHneFiRnTaBPv3pqAgd
SzcxDxSJzCWVepmG2ratdWIFhUMQHJaWz9cHiYusdRSHR0BQ4dlPLPX9huAE1rVj6OOfJD4aIkDZ
5ICvm8ahjPbLSqpDwmkjm/BDzLyQZbWO6jJyCdZcGKRK5TXk8XvEqOGA4ELV24oDkQcWZRuNAjll
b9D1dr20aWUhcGEnMVtdnUsWgeJwnoJ4NuyPEdXR/4WmMkMcLTsy3PWrhVPGbP2iL/y5iFa8g33t
3yFslb2jIa2dIE6CgIvKYOLrvG9kxZpWjLdL0DLNVV68M0WsGVBDZtmdfR2TqbuLuXyQpox0TZXe
eTfmPtPRbBpd3uqgHv9M6uz4CF2wNhtpCyJztiuUxLXBMs/UejCIarz6EadZNPOheneo2pVv/czo
XeweYXTZcY6LQK3yz+n+arZsEWL5cAklabL4NJIihk8+1A0PAIycsyRH/Y5i9lt/ceR1EFdkwGA+
PEQ14AhdR5YbUrxo/NEKtajy+bq30om8xdWaPh7Z1ATVm3ldicY0Hoval8yT24NnA9G9mQ4nNQVG
C27BcBPALoaQthOyn73BKNCOHKaywiysFScLgtjN7mwpHAgNVh5bpuz9YGVrWM9+f7tkqMy5Acac
OfiRzRlmM/CKoWxmBZmdDenFG7LX4FbWxsqqrOYaLGTNFQFxRpWGLS6W2OLLMcK4F3fuFPa5SZlN
P/WdM39AR+Z3jXSfAUp/xX0y2uC+yAUyluIVgzSWkc7PXbKuLfL4tRr/9Otg3EESGkDXmVg63fvS
5pwJQM89B6IrWiBfB+w4PJJJJ0FtmdH90oH+vVKFuP9TR4Bx3++CAST6wsS+EKpvOnWssWZF3wnO
u4XuV93ZMoYz3KLsfyx4jv2xuXGOchtpxaqOO9C52lxd6ZzO4W/HLtTODMPLlqSFjlJQdJqltlLZ
98kM75oXmaEbyJdZOZHJWzn4Fky87kmcKr91RZM4rMzgEOJhxMILKHCozyCtAuhV/aiUdXLsGPna
qqaDKs7Ul0H4R5qMqU2eytnSI5Xr79yeGMynFfbMszjvz9HQYDELZJRJtZl0m+KnSGCJOAVOmp4U
NUm52CBhoJOqDAoeJAFjbXNGYYuVtNdU26JIxlNbj6hguyfaKRnfI28NqxreEC8Aude0yuL+ioBt
akdyR/L5M2ecNdu1PUaAoPE8IUsQD9rLi/7kAu0DBeQ2BqodeLLHUt/2cUaI+9bjD+2TPv9pQLl+
dBG1ysE8/hU/rAfzzoPamQltU5Lxf05ZINHIeonNCpwosBdiNqy3RpZT/vh4oLWjkDTPlytfJQIT
X38DJyCQrui2V53wFjRiLnKHEO3HxEL2gUFA5v4XJTxHsQumeTaj1yF9hThfVK0uaa+18GQ2wmiw
UvLM8PE2VFIyWPjn5MyLV95annuX+hE+YG6alzwgb62tkSl/NOBOWKvgU5l4HKyMXYn13jGlLM3/
qo73UHmjP3Jlc6e2wGgaB+BQ/txOVhJqf4/U5xk1iwINpq4pcN5s4ziugaeClkn3cxS8mKu9BKNu
p4epSu0TrsUK+DpCMgI0h7vk8sIYyY5YzGvYoXSyyRLzW0+6c9gCAd1+9nuRfjMtfkB1LSBWGbn1
Q1KAWzqCj04zha4nw2xjAKLckmXLiOuX9sSJOndBxG4fuI9wOXLoza6O7p1RY+cAwZLnrfluge7R
r8zI+d5c7ZUZj4fMF6V+28IR4yESNdoTj9AO5qpjoGZh8V9oFIOu2luVvrlII8CaLaKiSlg0lmD/
hdByAoPZFWj+NWexbdcgbBEq/jNwrisBhoEVkkZGFCzKAT33iwkkvJzLH6naWBQf5GLD/Ib08VmK
2yMN51VPL4oZCrlpf7kpOiKi1uCbOxfeNWFggYvYVTj8T8pbgn2mkZXI2BRCKT55MLZiEuiAtyaE
ggGsC+iz+EWAt5FnAGVa8Y04wBmMgSCspKecCR3E1aqaxBKxFvZ4jTNpn/M4sjLOj7Dfe55vkVn6
tbYXLmp72ymYIjcgRGrpGQ43LCz+UAFJeWB8N0lfQRQEpR4509PsWqzLRVfJ9e6KDJoB+YAm9aOX
WpnfL+hu13KwxHuj0HnMudut4PONmRbYk5Oyd5vHAZLVvPkQRf8mxR05BaU+6ML7WkqOANAmPW5z
T9tm7h5xUMAjcgFobHBJqR07w/FxrPeqflyEqAJpQ4Bfak28zeklr99W6y4NfII67FPDdelqDGU6
Up5yr5ipQDL71FA9n50h+aSGiWO+AQ4FjVm4jypjgaF3qKYdciPl6U2Ot4FnRwhtDGTUgcxYh3v7
D5rBd/XXcx2i8L6HwtAYl3ICjUndo5JEAOKx/q2kZ88tElx5Ds9GQ1LynFaO9HPTzynqApuSjRGg
Pg5NlIJQuP7T4nANasm47SRpm3qyXZhGIsrMPMi4+cBiIvEIdafc7YZV+PBWrHWyQFDHzhDvQFye
gY4jUM/lpVI1ZlHVcptr5wLhcnrNPeUCA9l+trscWiM8qcAU4mXVrWDIs37H69O9/Pn5QI09KTiV
TLQ7J7fndWPOD2cOh0J5otbuxhl3cTmxNk9+kzWQDdfmFxoQOugDIjAnQPBEWHNdXyzcXSQSpwng
vhZO3Td41Rado70YL61mHYZyKI+7Gjo8bixfzAZc8EsQ5sRYABSCmsGDTsBkCUJQzdXaSZTPkpsz
7mFSpiB0Ols72MVRKwkLstiN259bkrt73ib31O4usbRjKgYfCKZjHSrGy9dIK2dVYeN3HGSpY1E9
l63V0M9zljB2QmkiI3H9MaRnkOeTw2ABVFmZcNlIDaKQxluEMirjVbiPnP39rEw9nBVFrxQ5gJkc
ZZ11MzZATa7uK+0vzafo4DyweT8+bM6C5P6cucNdy4Ajp+97YCw6R3VKAIS5Z3yG/heaBGx+7OII
ADNo4oguSrRr6noL7cLRKOWjIP2O94CGsylzzF16sRN98+qDDrZiffEhQrn3TXwUl4Heqs6NOczm
4Bx8gapDGZfd3Yn5akB6/nuci3FhIdwR/G4j4iKibXcT/YFFvvRvTnWt9s6Shtd/XvXZJULdjpVL
WwyvbMAe0vUrByPxLNAyIPPTT1FHMxW53Yjl3xJXNH1EcfvQOBPFx0zglYC6F+ZLK2hsec1Nisfh
vbSG8TNgdi/IS74iLj2B4OWaI/5T/OeC0jaebFddasF+nrnrjpQYTwf4jJGARSd9hcNp8b0zDh5S
O7McmfIDxuF69eezDpdMuhsej+GdJmBt0T3JYnece1qdx0QARwp03WDr5Q7CRKZkwGsfuPP4Ma9Q
hY0EoJE7iChwaQHlv+SRT3fd3GQdYKyY/uu7A4S0TR2ZIycvFlUHM3FPRoIcxwN0wMfSvcufMUZD
Yee5El6PBj0D147OJa7OOWPjdtuAfEY4uh3FKc+JtRA7D3W6auM2YNnslmQWkUllFNTJmlww/QQb
Cw3LvKud1QWsbWowgJL8Jd2ODKcKyr+OQxpFh7URmJXb9iLcJ7kU9hZlwT+nV60qwm0e9tDqTFZn
L5dd0LapdMzISniPmknxVaWU3mxqjot90y4oH+N9guufLng1pA7zJtsSSYqSgRAgJCkEUWYB2gEE
dnIgBsIXS2rIb21g/Xd8Ak1BF3eYPdowhJ7Lsw9qZrBe6uNzyBS21YTc7yz+VSADCz8ibyQcCGLx
DjaFzqcF8/G8DxqmeoW6T/5LdKY8C8P5aDUXiYpRCTpzJepSu0Sn3lKWjAsRMGk4VL7A5cg4i0gN
AEcEDhIAKk2FJ+9gjay9fDvI9JIKE2hCVyb/HYysSc72P2FxxbBX8r88ot5qFy3IjuL3+uhAB+JY
Jkv9HH9gIXUl0gY7sgHmOSZyIS5chg6lZ1ZCxtfQ/YcJZ+GI567fxmS0PrLwIzpaYjDMDdV8bjiY
JAt3sCq8mhZ3TfZDfXR6Qy9i9+ZkCwfbJAta1BR5fIL5nCBQ47/a3DPcGnK+NZlK4GBjdMx/FyW0
athBGowhSqypLjOTigIBUS7OqVAGvtgPz8bGKj9xpcsrbmubdqJ/Qal0qySHihnD21D2R60bBX8R
MwkfL7egNgFkeK05f5Ppstvmllsmr9hjI/78ClqmH+WpFZ5YY8lSQHeRMNkrnvCo0IElp1JHg+Hh
AST3IoRODX7EbGJk8PqcJp1pPWCRSJsJ0kCLwCJ2C5TqeVDYOsO2y7FI4SP/5GNoiFDnFHqXH5+y
Of+uOEJuGPa6fpRmhitMRBmySCaRmre8UksHAAVfIgpM2Zz/yJyQ27MqRjy4YGx+aNM4xhCa0Uzq
JmA6acfMn9GFwgBAWN/2YXOPx/yiJVdK+8vdjeQOicvGsS5oNJBm5Az56mAXGxk8AvDKfQZrAaIk
bTnBel4UQbrgceCEHYjOHz8nddHdNbnx0bXKQ/z6xcswZFbE4WnTpXI9Gvb+zV428C45FlfQUb3K
HUAcry5414D5v+hpEXiafosaVXllerKMURE8PVacnVZOEDzt3efRaIwnmtFv/23Rg8qrNkr6BxW8
mFsLDefxC0u0s6cCXLGvdybRRxml3Ujc2iBONiwjwK+ahRUdT2W4iNsLX/hsP3L+v3EOdkI/CX9N
N6ocEpFspHszITry7+GeLfKfSkSZ7vkO1xgTY0x5HytIB/nttg8ye8bk2JGzZPVA3BDz3HSwAmgs
gvjVwE6eKfnr7p2mxRo6L/jMTqeQ0I/3MxiJob6yijFjyETWuFM1I6Z1XmrKtTlgv4LyOwToQtVs
2iGyZPtYvqBOcJ05G6MyL3akYPMfwVLA0gQ7h5EgpIPzuT698F9ar1XMn6OKaMQOlPWi8JRUVd08
C0LpekbUZ3fCTJ6mavnFrBaqHht+iy8eEUt+i+OSgaZ9vyWoHi3bWaFspVdluE4/ofJhu7XHlfcW
FrL7XBl99yyL9QSvnn1gL29bOApLBqiWufjhMOSjIiMgyDKwgdSLTYxV4+9VfEG0xafFlcN/Aa8d
73wNnGKPCmibbFUG5cW60wPTQqUQVL1czkGsVKr0p893VyDh6aFR9k9ygNcFAuZy3gG/xRzzqykf
q5aRSia83dUF27eRQgMrSNXRfOH3O/IOmypag4v/2n9QW9/Mfcb9oAtKYdMMSyXu+EsJk6pj4C3h
yEmHWtQ/eRSqSwlk1DpGCycRr9/kqcc3FyOwUf5n8b/FVQcwIAaFe1moHhgR7EaQO7egJZc/uBFj
JIQG6L5BK/1ZPUFT5S3DX9IX7lm3aY8Rypw9K9lnUQdzu5w/a45/QbffJxWBtfIEvjf72NhHkTEL
hanvgifL/irlXNqhIj4OD4sFAuts45XmPsBV33UmOK7yx9B5TDpjwIYqCb7Nnu3S/IQdMC8VGYQ0
nKdyPCSw0h0t8XdiDgFM3vaw3+Md59doRBqRRwAKqgr/J+lzdsdCoNlBuOgpx5IROiLU+X5L0cZM
C+yVBBhAESWJBXPFCAoQsOMephwGN+rU6znzn53ghpXIzDxQ5Vk/GXqoY0SaKN5WWbznma5LaoFh
F8BL7AXR5RH31cgXxnkeBkGqQlPk60kwrjKqc7WnZfZ6qwY9qO15en3ZibfYkDlloOrFkVyj6UD4
l2089KzqDthATsF3quM3I1rOOgrXne47/l8kXg+iU4cV3JXFFha9F7bfgceJpTtJVww/WgzBT2DV
42g2iLo2lhzqkD1fct2dKXAJaoZW7lcR2JuB9m9O36u/karwbpyQkFRNrZ0Clt+XkyMAtmXxPoi6
XgugBW5eUkbDBWQH1UlDksz16sDZGVpMka41I+6MhdMEpLZakPuj/I0Jn9qdlUsitp8eN9/4IAWt
FH8iGF02IRpiKtKamulykosOtJqQPHtJCeEug6gs8wNMQV1evWd8lxf206JqDCMuPtUXU98X7Ky8
9WTJb2X4geNmtFVGQSCO0myqBXV4MF1jg+uUfkfDsLfEDsutMDQMQx6Y5oTt5Xifr/u5d95TB5ct
iEMDmUNl7H7WxuiyivvMPSlMnn+BYO0HXEXLCBN2G9MFXKeun7jX+vaElzSZ7FhS5aVhPHOHgExq
HeC8DNb+e+O9fvyQ0uMi+kh35Hf8O/lLvvWL/cS4EG+Vhr6cnbyMSTkGi8nDqsHK5Ws7cNARFMIJ
70iy9Cr8NAQxVVoJkvkm+y4Notf5kuC0a9Q2vgXS1Yyk/IIhm94NpzJhaCP4jm8Sr9pypVpGr6li
Lrq2IG5Se67Bbw1bAf6nzHGNpA1l0usfBPCSPaUbXBuxJ3DuQF8TDk/+PnXBVPo/hTxZZ/ADLj0p
0EbWu9SWK6r+VqM80suKvzgUVXC+gwyDprFwVpS+OEEEfnTv+7kSmqtRSlwm6ONpUo1foGgRdIXV
KK+3jqRb2NTDvCouoe0uHnhA27tKtqvlivL10WEvNDSY+izwhU7WtRBYwwnzLBs/Saf9tOjUoxGY
DiBmF9KLAXxJBIg1Ianv4tpy4Ag5kJTKbBaqRNmdNmY7Dhvv5zg7sinAl/ymWmzAWygGeTduKwkN
j6XKjEgAjuJRrQhdILFsHWQzzOblTOL0CCejtJ1TVY19906TjnIfh3vin16u8kFHfl6bJcj6xEbt
7LtGIbWnucPkJqem1YlyDgBqcUC/57Z3U/OHTXrsoL0SOSmBfGkJJtcyw/v5k1xjlqQQ1oCZUUNF
2HCFvKJzg6pgLGZrkLFKLswoQtPRH9OX1wsQVOEpQVPSC6lUMP93y+frztzYCkp14Rjz6KoZFzBH
XTBPXA6tKduaoNakJil0b2fKtaBRcJaD4FysHYfe+1Rezxdg/MApL+T1MqZzGhsX7pY5vcM9TJzL
ZaQYA5OoD6XughZGBxu+Z/rghBXBMqxbtVtE0G/xNVi01JgHuvo9xzTMkSbNhDdJALN81QDy5RMZ
Ip1n5/fMwPjujanstqGYkoCRCb/N+HyTpr1k3Al9FPxVdG1Ja3Nmwn2shAlEMiopo0rXoYvWutYD
abUiL82axGrrL4nnOPBSSMniQai4Gr40L8lNZAEk1ozTlHXEzcV83pm1T/Pg+CqbRqRNIj30dtQG
4qugLHkvc0IA6g+8rwUsGGYJfzDVk0nASoFZDs0ZhTmhu2lWKYSmoCsIVIn5DLS6giEGiwwlyszP
ADtYq4zZyB0gUEqA7pCgGJsvcer6//9eOF+AwFMovreaBrS6EOQMW8cXvde3BulR9Gz5cKag6jjg
11zt38ARjTl7+Apbr/R/n07YmMWKBtzEmwwSuU0lzV2UzNH5gQ5i44HrxIf8CruUeNwcUtUOU4DN
hqlKTYBdOgftFCKUMkCQpIOqnjceSCACwMZs8Yw1TtB4xiimnUn4Xcgdjxw6ZZXw1aEyF/DyckbS
Nia1O7bQoXlGPrTUZMx5Hj7zdiiuDiZ2Y0hgXzushHfhw8aAWRKA+97V6F/wO+peRqCi5Vp9Fstc
8Xhj52eKWrf6R/UmscYzZsD0NlykzATzh+10oE4KjlQkd0nIq79Uf9BNWxOyM/b4PgpcDSHkAZoa
sOBe0y00SBmIVR+o9iJZRzxNZZfrhixiUqrtdxibW4lEf3T7XOVUKKAdxbxfrNYWj/hiOStOHazU
NVKnEJYjXH5cLJpKl8biBueWSA7x8ko3rdWdtM5Ag4aBfeuOpSRGbVc2/mbTO6Gcw8CGIKhgFPM8
inn8nbOF1LcI2NMnC8irSCAcxHiFSmNaLpfc8eqVcTxB1OKZxpfmnsbJqMw32DP6+lI+8EWgwz1Y
MaddI3pBluhZmxKDBCcOT17o3iClKgpDkgMyfgfHKm3DskWc5S68gpSMPcZs8LBLulEjiVOHrRVC
e37fNZW/dp+K1L9XzPC9gI3uS72MmNVgRCoyRix63QHrVqf6/qYrB8F9CyXn8yGaxlD0mRNwrQKF
oVqZBFCo3g/R/vjSKQQzjvNRrU93FvfxKy8nAt3VV5EJ+uyULvw/0+cNWbgD25Gow9Ni5eyKb0yf
FATxAiGdhLkhLlCB1upg6bbqKjHnPH00x5V48vFi5CL5IfNzqzdvM/ZXbHP3i9xDzwC0RS2n9XBf
z2Obenrdil5Vyj5yuJvu/brhiOQgNlbnF1WPNO9UIjWz8yLcUjuRXFD32tmXcV/hqYmcmWqcmDiF
Vt/CIhHeE5uyp31hbQ8h5lhnB57dRsrMh10HfX767aGmMwAYdVLcn/LFGDdW6xtsOBNsYiI/fUTl
XqjpJ6aR7GittdVRA0W2QgkPwijrju421obkDHw/yYf4x+0ttUcVLle3CaoE7ur9WeAQGTjNOjua
PCqCttB7F35c61rDUhl9oMZRserxv+J2lQmX7gFcqorHl5fGcejEvRPX+svP/NtopN2iR9FLnstb
nP9ubqFImyfoFWBWXBRRJkiz9ufzB24/vzuDmrrji1kg8mL7B9e4eL9ySvHAYJfON1oydW/17pls
rPNfr8nAjOODLXTvBAQPUjBpRvw5EYYEHaMSmEZDN669hzuSUvQUJaGDCUFfEY1FXw4YSLLCUGgn
dSQKVPi0D/5JDQk0lCVp7SkoPiz55wCNrwt8YcSofs0o7e4WScsbSOHZIJILsEw+cDHsDLf9CoZ1
umaXMPt76cRoKPfCgPDP85mrj5mbnXcTxo9hmLm1XdEV85iojzSblC9UrDaC4wQ+T7pZzuE+i7so
mcL1K6s5G6GAQ4z1kLA0gEubWzl7uHP2dGWzPSCK6BYrtGXVLm5gBjg7Zw/0lB7QcRMTkR7fzWQF
H0YEfKxw4eWiO9p7HY//VoB+Fva03U8bYRGu1qeCsBkIYATzRDeKiBZ5Tgop3g8yDpp0O+FpyLT6
uzIcVFS4tPUhObzazGp9iKegQeGVz3ojChkWeB3OXcKOlVfscXDbAyRuUB/Wl732wJGpLMsblFJa
d3nESwSAyozl7lzdW9wpim55Lg+Qx75nD+GHrzNW3szLjg40UrT/8u4Nbm5/WQsUM28/BnjDK9Ls
Spx4/8dGJ6k7bZO79kyOQz8oqByXRhAtV9ZoAabl9wfMA0SxADvOO2FsFpJNMp3TkRy18P2m3kqb
E8DdFLNkXJ6oMuQnpUqQQL0KmzGzu/h1BbegpJrVoCMaC3yQpKguF5SqO170IiL9X5O3xCJy9ue4
rY1Mfaj/Ugx/i56NVdC7lkXARmQHj8JVUbMXusRktf307NF+y/EcXJvOEz/3iVR5cNzpIivxURnq
bzIblR9VKkWbPgbfDDgjLlK18wP/xKyWB2xPv0DfNvQ8hqgRDQP5naySSku7+11NSWnShQlJPXyZ
8WOVWtvSizwphiGYoRQbrYTFL48pA27530CZ4JSN9ad912+13xhn/vTVAA4kwjBJyYwuMfuMteAz
g6HNvCFkj+dvVB3bzknbr/Zqd4pvtQCy2cQuhvCiflFPVOrxJU1WgnZ3gIY7JIuPZoJ+d+zcBAR9
Tm7tKrBMYA3H45m46Ofaen7O4VquaquaK06T0d5JwVuBl5xGrRZjkXsp1t/JMgR/OVAihxVKnf/c
x49u8YNzH3dLgG1s5t/sV/CbNNRBAWGsNpJf8HJGZ/j2pApGduy2ZW+Ay0JXzPaXMmzPlOMOb4G1
XN2tu/cAcJ0dVt64RAmMaFyLVzlqRWMg9bTJZVb28uwk97C00fK714tS+6KMVNQ0kjiVhhSdm/wf
lnBY8d0h30JevhiGisa1yQq/8IZYkw6xfDLBySm/DQcCFS+8RY+eTTqZr0GOw/CNbD0o8m5fpLAt
Ts4PCQ8rWHSB+O/eI9JWGAfLpAWqreqG4Q4hjkddoyqGeb/Z6tqZDF58Yv7JRBWzVtxZ9T8i++RP
baoJVCvmHXRTF4XwkHNAA7YDJPvrpBAgGLquTahng4oWkIZTlJs9EtAaLk1YN02RNr4u5LmjC7xm
uL6A+eYyE5fHTGSnVlo22rq+5MmxZYqO+vo0Srvih3RU317hfhsjgiWTn0+sH0ogC9JE6ACFG9oV
rrkkyVGz/loJXy8207b3En/6u4nAcwW6RShbbSAM8M01m8yKti58Uj1aUwaIaDaq+dZHrjPONB7y
1WDEM7rjDmoyvKwvhtNwJ2gxnaVWw/QnHwIh5Lb7Tie7ncVbQAOaBZ4bgfnhfEWEgQPQING/p0uw
1fKpglJnOccD33gmLD3viRH+22bE5gU0vkz+j/NMIH/freg8XavDgSjIzhdwUgv9bF6nDI8orESc
9UAnmzz6lffUOuuuHBe08ZWbU8GG3C3oUxOdqTCvKY31y7c2xH3eUoKmmpH5KDdBFORZmUKyO0/t
B71Kp/6SMyr1p0fTJcMS27YqcA7pNKuUcgbPL7bm57M2ebuwzbhuoAdyNtyxpZIg0VZRDveKNdTu
7b0WLZmv9kWAciL9G1TZb51Sn4H9eBwrEtw/HQfWxxDRUggxD+jlnf7f60wXubzD6BdZzNAJPhE8
0TJCVfUFoPaj65BaCopksInHDf5yB660uA0TLEvkUQIX0vHDj8gQYhIbDC+2i8/A+m2WduLU9oeJ
YjnEivZgeO+B/bNUYgO5b+VT+VkwOPNuRGjCZqo+9klGHM6swGJt8ZytmR3DRShIu9e4fIalEDP8
Dpz1nerrU9kvcCpGhIl2bgjFDF5CPbRSProszNbujsbCDNk4fsCKbEqTsvnDevtgpMhWlxDF0dN4
tdDvzWcB5stcD9pB1l1kqkX4yROxpWPhICymiPhpaTfuRqKisqg3vhiI2gd8p6Zvf7i84u4FSA1k
INalUrbNpa+CR/eaXNaCtpuivxSnlqbjwDm46hl1EZA33dJtRJrKSjCMWA9oMcPSBo7CNshHFhe5
nezNgu++89MSe46EldMx44+zs10/amL5ZuxM01qdhaPu7lHz9V7z+u2dBEPyBT23fMr+8eX7pVA4
S3/tep2bYcYM/HJFmKsGj/KHJWhYfSHKMnQD3GllkeCjDbBnHGoYSLJ5NcHz5IlSEFS39X5OBsAO
tdbjWWqvzSfb7qXuxOjPYd0Qx/6ac84Neu1EPZLQEtgRD6DSzjiSn1LbxY73SWRR5v0EPDJ2R9uN
ycJU2S8xJQ/X+uVdRC2KoZ0GDLYcpclAJ8E07PSXYihUEpvfZjL5oKaSVQO+AUa9Fgfa7cYOUTZ3
Wcie87lfZYtapgS4TMZYMIh1SmJaeQSizX+UEfwnPbcMw8KOTYUEFemm6mlGp/Xrtw8taz/R7VNx
UMrHd9BoVBjG6u9Nd+Phg6wyhl8EKrVzqPBtPKDbsc6J7lufEpSjaZDsOqGGqRXWWwINpuhkF4oG
ACtxJr7xMuhndLGfVrSEvfJCGOnBWsYVYtrewVB3LvzddUlrUgVIJ3NcTNP+Sd/kRdgKcxvLDmFH
987sA+3qH4dJGKK1wvC6jOEEETOBcrHgSZjIHHH4aWgGc+xCsVlcn54VcLKTIgB1t+H23aPUc9O0
HFQa5ZGYKltrROu1N0FEtgjgQ4Uga8Z0Q6esN26aRt2yJ8nOvHnZ7IIB9AMbpwpqp/nYxG9wJnBO
IwrykDWntN2ybSJ7aooQnWDwnUnYs2BkORlgIuP7D60WHrAZeUanZVyg2oFjGKOORfyZqXT22W/k
V9byjEk+a+z+/wUG1K597pOlLS5qhuDB9p4fUG/+8ypcWr/Uc/qXbJXxS3yhCMtWa6URbRWIq6tf
oykg+7UQo4jS9zkIuTqW3QFJoErOysr/cAaUbMSAiwRnMNqcEzvEn3BPl+IkAw+v0ekdaRvQDvmh
kx7TkMb+S+ZNNmBIZQ6hfKDHi56blkBiq6d4dBYB8cdHKa/HbuPTFRdVIL3mnTpRfpe4HSYB4LEl
uj5WRwQ0EBvSfyECc/yCa3GajT7h+/aShBF5mrjU7E2ggPcNokaKHgbu3tJbfMLHvpVnapT5w0QP
rs7CuxLGmEGlJ1x9Hqs1+ZV6um6zuHETqK/2LvqhvsnBhKGusEqJBGZSTf6HgvCDZJ5+sLnOH/q3
n3Cs910xjQQoWaU6UC3p5LWw6t5CGarjSONHHACSLeRzZHpXw078iB1AWpI7qfCcA7+o8kZVCung
zLY7LK63A3xxqZ2eQlBAX68gwbOY/Gu/Ue+n9T01vJE76KlUBksha+jNKj+simE3hVcao/wzjEMi
plzdRVP1s7LisDUBX6y/JFJ5JMSlwSV7XVDOglNCtkWENc31SLJxRwTvzp2LLfZQ6OzzExS0K6Q5
fvQsLU+GuutyoQaZPXlbjP/hiFjDvnx+hAgwdPVpt+qsIWPSAnJQRjHfpE0l7KyciKgenYLFX/iM
lTa7iZxy5fguMd8vJrxzxmQX6UCyPQML3mShpaemNpOgySPKF1CtOq5quRmj3oI7kzz3va3cCJS0
4or/UQBfkNFROZ+Him8xImSYDsXe40IIoiNClEDdoDPewHZjPsdrRGRfVQvBfVcd8ERanq/wfTcE
z7r2Wqm2lneb4CO8HhOcKBkCAxErVURsTghqF/HVBNfile49m8Fav+BVPdTfp/Xv7/K4s6C4jon5
+jQG0bn7d+zTr7g5EOSDLD93so1gy+PeDPJgv5fPdGuct7gGk49KY75rH8zK1SJ5qvxBEWeFLAcd
NMmnvqO0ouEwvuHt8HeF0j94mlbyKGfZ/ktDssTfXwHGwbveNQAvKA/EmoqUZAFrlFPuUr3F0A/C
DRUIH3Kf0LX4XbZXDUCePLgGqlofuqutjKJK9yman/T1CV5u33KBM6JnJpKhmsIwqauY4uKMoPfI
bEIy/zM7QVJgVClpz42WcrMX3dm5ertzKhBiCtmHG14WrAsoWXnhU4YbJ13nbOLX+u+Rm20vI3zz
vqfrVribT4l5kHkNe7h2PR3V+0Oqf6c2rCkFfNgwhOHC7Ftha6y7vMYr28rktOZg3ZjGHH9UbXMe
HHNOG+ipUPNFtlegVW/sWmACbcFSeJLBCKTdBO2UCcVnkgHBWEcUtgaTbAwhVBS5BnY/GruhpInk
Ns1MKg0mOXwsuYeKI7tdisq9WfPa5KedtXAlJLTIbjWR+lE0jZi9aBDR/0aevAgyE/LPGi5ssgOi
IOLEPzAxR0frCB7pS+tapthLEI1kPcdheW6CBRbO/dMSrxPB2xDrqU1B/I+c9E4t/sdLdhEXCY8S
kU124397khUDecWz1JBn6d1kpKZWJ7v4rKaPp2C/9Mo2avVNZbcfzM7bPv5gPRxwaVUPJB7GDGfM
MqEtbNMHZIETgOPS9H7zLSnDTeRU6UWa2bn3QPRvgqt1pOAiyd1+S5iY4D8gUhnZwirMFcWHA0B2
6MbHfgz6VH0ticOfTRAltrZ6DXB8KNXQJmI5vnKyGC1eAzPWYuZ36FE+wCSev6JN7JKrHrFDShss
5OZkMbQNdA4ZWBhVgAvkQMfshlSih9MazS4bZSK44oxa10fshqOTknaGzu8nGJTdlMv8BFz7dGCN
/Jv36NPhCxlDowGNQh5Wb3O3JCUDUZMwosp9HsrCNQ05ALe3YHKGl1hTiJUDDgwQm/uZrv4IQh9g
SffHfbJoaIprPKQzbb2ygZw6MMnpayk+/7up5vJxArURNVjxAHVTZZQkgNZhasK7llOI3UdyM8u8
GLHOsCX/uUCjeYnm8SxW1bzRDJoM++tSpSq2/O631LL+HMtRqSmkVGpFqNvxqjcg0qKRNSY7/rz8
hsjyzsYS+ruxXfsZkraAXgu8OzXcZhJnMUci5NuiQ2mF1y04PusJtb74gyrobgVGFjmiOWHo3ETp
zgSLAhDbqOw3r4tdaQv3Mz8broHVvsRpzuwaPzwx2RMwWuLLFz0r8VVUJUGKrBNF1IRN2Ygn8WSw
sO7xKb3nplJNwEH0MzBy8k+0kJs+2aoepkTR+Zs/P+f4Up1exIyf9dpaj2VEi0i/RZGj9ff9pxmX
ASZ6tGkYHJW8QykhlCtRJciYu43y3jydf16IGu+qzDaDEXdir3CZl4xD5B7mHYE+D42adwx9KCib
kONgPrjCov+nOi8CdZVcnyr/78Rl58UvZ9f1PAtObMkXOAQYZ0IQI9iPRKbxnUVuN6o14uy2QokE
mPaIo7C/25KqffcWG+ie/djlt7FWG7k+7MVQG772xz9ubD7oahHpMdZxlOiC/BRtBHl6Ng/RTsiJ
fwcH96Pz6nrCopWKM/RdSOoPahlOtcFXw4eQSGaYvkr15h/pRy4EfrxLuMmVFWsINufO4UF5sU+K
H0lftk8ZWm1kymHPOY0aeMvB+BlZaLgdDiEHExuW0Rc7S59YQ5cGJ1ykIyFad7on3ehmyLI3M3ic
zwWGLc2Sd7r3xMyRUxLw/PlLip3fCh3s09BEpc0lMCJ00JRT1OanV1ChPXNNPSjK42OnOPIagSQJ
9CsWROxPsJF2Pq12os86/T6mxw1yF3svkLZZtW0dgDRG2AtO2pjYsAZ3SKiZjpwB0R6JUT8gLn/k
PKAmtEdk2Ikd/4kC4QYvfcc8KQ4x9af5Xya806H6L5h9qnR3UuEsfMVId9CRacfmIXBtjF6UOCEa
nFX6m6pzLVTKCyFJ8ajQB6Q1HJwEM20SclNokP4acb51V86f4EIzS/GqAAfQv4ikp4EW+vwvK0+E
k2C0pFozTae9CFc4CyBK0iscnyDbFlSd225sltvsQLhP1RUke/jd+v9f/yO1vuGeNfj5F5/YKKek
dZx48k3cgehJ8vCONwu4tbxQ4ix+OFu317Bf3K3lvOGLjnTolQKi5he1Wc/U9VExPOqTOYyjaECg
g3kWYHz7w53Apowq/3FR+rFkDkdOvT8xYtS5D3S/l0pm2MVsg33kciEsGv3Wu0Aumy8Fe795jw1j
UIggTiA3qszSWqV/tibfb/YR2/1krOFO0Wt2Rs1yD8Y38F3jQL3f0+9AmLvAV26gL8Ippa2i3Bli
Xt8Kjr0WwkgtNL8sfX6H2gVB8P3tI0BJlmEMzvE/a7TEwyj1nuEedFGwRh1BQfmsrvViAW6tH9+Q
NRXetkd8S2RvMRg6W9dU+pFlqAekpHjei+KDwVvt3kLQdB4w+HtU+Q/xb3olO6duF/91/I/fKmHd
z0bSg/Ahyd6qCYTDDTozjw7WlGKcdofZN8ElpqbmM5lLjNL5HUCRaeoRk1nhAW+iDMP5YRrNxohF
MKkrLQeGTZXuWW4D5f8Vepzzgv1EdyGtJhvAwKeLOa4t7AXugfbZc9Ex0Q+9FnT0yI6DUlMJYMAC
EGvx6b9p+79IbLkR9jXrcFjAZ38+FymMoXliBY1YuarLiwfBGvDFnT/dZCe2NQNCljzQ0/4WEu3Y
sILG3CaVPWbKjc5G5SOzAm5eyzgNRy5Rj74TLsZdSQ2rnYvXS1YnPxyY+JGSBcgyEiIHNkGTURAR
JO4cHQBFFaT9WHzZNtneCDBu2jdXnG2YiiexjjXQwJV+g5bi0lz/GHN+Omg6lJt8mw5RTor8tjM1
MS99guZyhmFXO9PyaGdL5RF9LDHTsUw8UD5QZw79TRhqSDFdRLOqkNTLpsxQG4OyraQULaVbtZnC
0VmTkcxuNBBnm4ACET4IzKlXxBJWBDDekaJ4FTE512SDJFpf4O94sYacpczND1w7Gfm5/JlCU97m
2K46EfKSF/zM8Oni1pocN6oYdPVdIhEHqX+hPMCklg+vx9wHbeQZHsYv6M8avKhA+ASizlET3w4y
TRjka4VeJBvUNK10pKluTDiF3HS/22Hvki+nrj1biqH4Rr2nipJhMre1VJskhSuMIqfrgf2qrRYC
MF6D8Ftsql0oQibvooFmofyGSdxJWIr/P1Npb2M5ZMMoMvhKJJ/JB3x776rm/wVsJH5GtsRh+slc
tISnMiVOE014HGHr0BxNPa1gjoop70WIEkoUcV+dngQDv/u771p9i5i/ONSzasu/uRRIrXMQAX1F
UiUnaUeQykCbUt3X2WjP3xfKwiT3oG0DytfXsQk7prCAfldf36Fhc2YUWza40EfXaPNHTErZjoPz
GTvs9OEtGGGAg6MVF89ER3810XteJqmTI55jyD21Gu5ASlary4UH86wAfeqnHDUgcW/eWvpDuO35
qbykCGPQrlL2wiY7sJKWJJPueQASzMIHwDr5LOzGejpLfTAg6Rq7vyoxB8Shs5kEQHQOUjO0edGW
KET/hkPcsKvvi8XzcBP5PU56vgO5DO3xsz43WD+JQA4s/kvQ1T48PiHqcdqLZ/aUD88kFOW+51E1
us4j5KDKF1utY+I0iGoqmW2cAbOcepeUtsf0btOzeXBSOl/RuLSmre1BW8QObOs1wHeFK0rnXRUx
5OLrTEg+YZ2tyzPFGQzYyQmqyqZFjTRv9PSoI7EM85i3OypjMJMRbf26rkpoH7TFVjWYYdUW6kB6
vRedNudccXsvnoRajDVxkbCIQEgryua4f0dGA9/ydyVB7X1YDELHE8OSoptrOMFZkk1Hc9eFnuY7
niQM5riuud8eQIYm9SCQxQJi3SuwTKSWAljBVpKfIU0L6mUJ6EcYOuwpqQAnGI8EW780t9flc1W9
kSbpczgcfZiINvhx/K1UH/jBeJbDu7KAww0sDKTJ1qeOH+TeE6JsuWphxFa73y9TEOXSsEg4DuF1
i+CXPs3YJWWQOBa9VfkKWJ7pznPWelhsvW0Yo0YlD7ix3o8mgIgRDj+NyRiHMtQpcK3Q/IkHExl2
1AYT9mlnc7BFjqQbGutdnFN9M9X2lQU/svKBrQRKWlaFXge/z6EGOLuBaVYogOuq9++7483AQ7wL
O2kbUk5ltQLWJudPAvzaeP1KfeI+mrGPf07CNwMuTy+zVPWA6H+CwobVvFmWNkK9uZdPF0uVLs7u
RbV3iEoE7K7jQEqtqrzov0Qxlej5vZQwsTnv9T0jFjpeShfH3T6Q6mxXkw5iWK98gt4sFb47PtQy
WOCaBhuH0hvsu24ICTYqE7prnpYPn4dSiMHziX4efKieGreooXU6AcZWcnSHn81wD8yy5GhiKS1G
QiU8ZjYgZSkwonb2/nyyF5ljn80RxGvglqtVLh9pO+REPXWDC8LSUNcpgjNBItjfF5yy9b2mbq/l
bVa8Cb2N0TbPeONoX+8sndn5Yp1YO3T07zzRYi+UWLzBV2HJfODu4ba7y8lRpwg4OzNVPpa7H7bt
5M2ywV+QA2hNGRKodlrm5FJRVSCK9YB2IrwmQ1i5NY27/qABJ7tivyU/rfend/D3ZuJAyb0WF2WE
T5RsPeq7CQT7k+hfJ5p1vk4DOwuaWKBUCVKBE9cCJ3YSjduKPfJcNtJnPTVQz739/9ezo40w9GSn
EhrlHoZS0cZw3v/LDap2U3h/j1l3cULJtwZJ5fGZWSV1N2BpdAbfdKbZPZUdQwC0lOB8AtvQVaD3
TxxEws9RuB+J0Eh57h6K+qSlLxXUiLzFoKEpll+YL7LVMm1asXCwoW2VmEOCJXkltOZ2FOSClQSU
hAkd6KzL9mqfIgVz5xDRXZnL0gS2E7/nrfvvaC6sfbaf2S0o+dj6Rw2jUA2DwGG2HaMOdf1TSFtF
d9tUlbMR6gAjzcM9Ut5u5kZKxyg1kK9o33p7ITyGEV8M6pY5fNduEPVLiajgdoccY9JHGDjvtk7Z
/xWJEhbMHXXUPAJW9NcfWrjpbN99TuI01GE+cLIYSs++yhXQiZCzwUjuEkMt7ZZa2NQSiYPuxRyV
tCvbCgs0fDuj58O9N/TdVWigPYm/F5/mPQ6qWOgF635s0QCL3CmPuBe0noCMP9b+3TbxAEhI+KEh
jriYQwmfmMjqKWEQ24wu9H+3x9FmI2dFdUM6HYh9C7+Ne8hOyxi5kmeQ4pWwsn9qvBZw9G8Ne9OL
KaZTJz8N0WRddP5rmT8AdcCbmjJUz8H4w7B3i294UKbvHyQkToo2dZ7Rjno+3VQQjubkQjNYLSOP
dVYZuL1Oql4eHiT3z4Fyv+v4hOloR5KVdGswNUcM0R9isUJ9CsWwhSQ77oLUBFUYUMhe3rE/EJ38
sxM2G/5rlMFbmia7b50ehhRb+WBDcBQn5t7uGg0EvBKuNBD4Yffpjo/duMv9c+LB59TUSFfddpXG
eaw22h3uOIJkxo3f1BdihkvLMC674z2EIhlZ1WPX7Bwn1ELLxPnFtG3sDTF5LQUzqbUXNvftrlsM
llmNHgL59HsAAwzeNma3QM7pTtV0BAIvE8sbMbU4SYGVCMcj9Id02pFcoCgweFf97E/ZyNz4fHSC
Oy0D2Cf4N8+iVXvwnddBbjAH2meMZBA7n2k3ZeaZe8EcfKBLEkPYsTW0XC9w70Q0lshVgzxZjwFg
leDdX5kmQipMredViAJAdZqmfshg9kPcbhstTFfLbDZyIgQ64KwRQAcGkw4GqAquxbgAH72HsJUG
SGo/u+lEhJjkeH5TNJ+zPax84ji8xPNZXLoPEx6QK7TvKGiZJm4+syK9+buhGXGBmJTiVFrIyS3r
OMzIWUnxZCRUOOOnHtXo/oIDqr3hhjOkReLPNsi+2qXYJG/vMgpUjdIJ8snDSi+FDlXzdGR3lHdV
rs05qxqjfkt13oAxTiyDCaXatWouuvB4zcQ+aT3w08MBmJJq6oVb4tA7InGYMCuVzwi5Ci5bczb0
0BJlKb+bxfnTBdj/Wb419uGgortwJOASxQoCENrLesyz+LqjfJJrzqekQbgFaet9DccNs1f+Mp4X
nZtSyyDSNDslRXwo009FF7P+JMusl5A8/BC/Go/Nllan7XuKW+7840plA6Ekii8biijqGKL44778
0RLr6P7+b6e1V7QH/y8fS3t/hLjtbugvvU+4KGsaUbjlUzhOq2phDN0GjV1F3G2m3Z9TKasKk4ru
PcZ93hTThpch/JD+dupWj/l4tWMnBdQNi8zbnR+JsBdqMZOmc17QYIYDdC0NDTvceJS5e6rhrP9a
eYL+f6CU9FIhOaJZy7GJlY0LQVckdxy4Ku3iHMFXRXSCk1GIxM3mp0yKL7XxPUwYkRJKskz33YtL
LHgEXm55r/UXa035lxZMDP/VInR1Df30ytrzfx9tjOAJP4toi14mHUd3K6FqJBPZdAd6meo2qeqG
lNHvTLOTl52P/iE4dHGD7d69+SP7Ck+FEK//1CmyJNVaEw1AcGMZ0q6cMxGGhIDxULrEJz/Q3ZyJ
bfSe9WPP8HoRK4+2okOgZwaGhIkUZuxdfPuUWsk+QIXRH02rfNjeqno0rVkBIeU+Y0Nh0lh0GjdF
6WO6fReFr2jbfbegvGkLFX8tDFm3XzEe6D/oPmIXPQ+9KQroAUVnApjOJJ+/dfHInByeClL4Gs7h
mu3HfA9M5GCiVzYAOkSx4vOUia5v+3TueUCukvbsnQbp2FZyjJDZ6BrZLlaLua/99S4gvnXjKDU1
zlxNpXCbx5QLtBbz8o+HwnTDM02T0bPsb1/mjnVKKj9krLW4+LtiOZzp1/4XNMJRA+Zgj5bnOxq0
/fR1UKD+iJtd3fgsFqauJvS+/71FWG1jK/g1lhWJrT7Crp9Kf0oQ12vzaSrzKkK17IYhIt86QcGv
RKQX60BndYNgFkIA3iGbqrNUCPbBP5v5G19djD8ma1HopGT5VoOaTEgG7Tfud9bu6cb81kcZl7e5
m6+JaA3X+SU/AgZ0YLFzfkahaYRCXgXkm6RGM9nWA0KWtJYDkPwlT165R1fQ+f3O4i5YTrBnagzY
FYLCoakMGZ/hrIzBf3GPstuBzddsaiOBVRmIhlo/NqJ0I5J42WOdnEAGQkprCbxc+mbs/gBnUG+F
JrqBTkFdvTdmpu1rK/pvFSSzE8WBVuisym6qPFKdrOJKpR9WO/+NCzDtaHt4nAV46QoQBea6ltKi
tyt+Arvdq2M6X5wW74oI1v/IIDrF4ksRgvNRFzIMDPdreWa4hTP9MIzXoTie+m4zeZk/yLMgb4dE
4hNtoSo8jb4u6aqq7uDa55aWjKm9dDHSn54YmkdxUD/7Ec79+0xFqujkkZH2EANT2nBJ6B8/QUsF
OAPhOuCDs2EJnt2gwKu3jQSGwsZifroGEiuAgkqhqKA5cehLHlKe7O6PcwUwqG8i33W8DmFiAr68
A6lE+8pt9lgE2LkLzj7kBpYaL5yNZCrxM72ROGSjUHFXyjwLT7JfeWZJiYa5zp/GfPJiyZ6CDmpg
AywbmHRfdhbadPutik0QBhATJqbixXcQWj+AFbOWhkFrByhhuAVSyKj+hkx3/NdsNN9hUIEKoF6g
a7U2vgpZ3psqPwewJ1fp9WceigTb21MaTbT1MFtFfxhiif8WUcubksH/HUR7tSxH+HxVmoy+pOwb
Q0kHHqM3FZ56Dqqb8u5lmZ35TjxytS4vrmGLQXKE4DdN3CY7ctWIJZczIV9E/gk39RRBXFdEw0hw
Sw4UhR0+/UHwadtfkmiFtsrVl+eH3H76wTsa6UmOl/8HJA0EVpPC4e35ZPVVgcWE5BRxHb8nYR5R
55VfeU8S8MFvFh3WqDDQJO5PVgTYNvIuei4RDgtzFOmKuvcFPW7pKUafaRd8b43pvU68cq7Jhu82
ojHUeUsrv7F8E/QU7yjCma7M0XtNWMmKSoDKPgEuEYQS4qmqq/7Yqoi4fq4GzC1YEFwlkW8nXZyY
e0tmjU93TWq+t4z3zaI9/8onHIbGoyvFgIBqObu6cBH/4aTcFbG6mjUs2ntwjOf5qGkPgVM+3X25
PoEezisKnrEq8QfVWIqJnkIOd0c8QkU5R3z1FyK1j8pD6QEJzjNkyjnEYO7/H46Zbg+WWSVq4Y6q
HsLgdxYPQ6vE4I+8upI2f54YMBQSkQwZouc3X9+8RpL9vByStMvq4IjgWaMLFwQjwY9DzUYzY9A5
OytmrsGni/PGDkv4j2g914scuGSlo0GIK/GZOeVlU3EFifSKxfN2nb3eKjuo3ApRtxBwVCzrimd7
Ig7X35f044dR+CTBtJgyDxwaSucOFc9lpfySNt5177jUTWKGEcGsCyCtahoWQwiTGMLbjXmV3B96
ddUEKwrLvgwal4IqkflOfFwFaqmAh4dqHcRWdblS64798++aP9ZjYB1LHmwP/i7zU66/UDvYUl2C
/0GxWG5fAWrfFBGqQYwayW0kZi/KnPhps1eCYwDwRLORd4/NgnH/o6QGgsJiq2f0a3JIHOf+o+vK
MUl0bh4no3ipvEvMwEgUrPQc2zdo+2pnaLyj80vqOjfr5h590pwbyMrLnb9qclNJTLA3kOCyQ3RZ
P08SU0UXHamz2YEvQsC2DrTtAbAdcVRNIbY0xnGhfxK5nkOA+hX+Bk9HUc8n3VISbhwXdSzx0Yh9
OgNllQOVGiwjQGIQuuezRM2McEcz7V2wk8nWhkkSpbtsTLqDo2rnvBQcQ9BE9M4VqewEwG1E8nYn
iqw+uvlLpBo32hEKEKpk/iGZGfXHy4+YbuooXC78KTUSIs8ivrz8/oak37UIRmtNz0m0CkJdL5YP
ypO4B0tKCsBQTaujIX1weVTTagx+moRlqjX9yi9a/6vTurmmiMPckFILaf8YICv37jSTjmnr67HP
lNBkpjrLa3IaJCPqutUUTCq+Iuaf+unY7shEkvFDeRWTjDrcdJ9MdQWJlnJI+tdmjtl2r/MS3YwF
kID5i/lcNfENlTL/rZSIArFQ2g4cHV+b37uO8lpRzdkG6cEy95ms3HhcaDLW9s/sBRTFoF0cOYiF
ddQcCJrv1ICdL1SHNdjlKqbtyQPwrxwBL66XRrMIK5uQZ5fnUQeZ9uZGENWa8dR94HMN8su+BFYR
HBBbLP9xQBdZSfKSCOmSdtfxHKb90zgII1jUEOCz1SF3ostkScruRT715uq+a2WgScpA1ojW6f22
KAKvRGV6//u5qa83gXCrPpwfeOjmTiQIkdSpF6u7ONmNZtMKaQIRFtDZm9oREXpnoMCeoCKi8vHm
Zkoy9gbx8nf+lOTUMe6kxq+2+cyTOAumbmaaooHX1WIyEO6IOlHZRMFC0+FZGomCctwg11X08egE
6ARFKK4jfErPSikyaoDmsM75QTdL+iEr+SwJ/SEN2ASLD1uY6IcQTHDcHdndwOZQk2g81evI1ccQ
otX0uKWnuFZFAAhReJlMfMeL9CjI/+iVje9PRvJtFnA0v3IlAK/EftU5KZIIdfahRhDHpkXeMh1P
3Iu7dk9f0kA9AzFE6AISr5FfB+UeaI91UdKSU6X08lpXZQlFn1iYcwhu00YJt6p0rxLG2jh/tHoR
/8zGuS/s8/rVPd8SnizZvRznRb104Mz/TFTsvDgJs6pXFsWvpd3gxe3b3l9x+tQ/iEerTWjdJATB
4/gp80GmpxvDMZx6WroMFHiJJJKQ9wkc0KeUWGt4QFvc7k5qbjyzsuuzzeHJvdOxpabn/f/Ek75z
27OKDM7Hj/3x7Hx3eweRqHeeVH0ohP4bSAPdRyC/+BgsfRZNhofk2vAqFTiZKGlhUIffXSGEDdkf
4P1Lk/+kPEDbJnBQ9Lt86A81vs0Jlq1q4lKjJhR1DeuFh4/sdU81fhT3U1R3qste9/HQANDRYz4I
JFD85II0jkTr4jt9JQYuurCUB4TTJIEkpS+Rn1wGMNdFCKVGQva9EdHzyjOXV94iGwXrOltsipXp
gNS+Yxsdcw8yY3IGfTUO9QfvSL0drS2t59zobyizbzLyHXwAgY/q5hkzu9Sx6B1NEGfzmNZmUA1V
aPTRQx4U3roZCr3JOYoe/EHSY8l5CAtQEQTVuUTpwEoLm48a1C57MBcs5ClbwFUgMOlSp0+y/RW1
pGr7RdX4u+517Z4F23SZN5Wm1i3Cp4+jd5zprIbjw8jr1t5Z/zvckNNqqiTGEB2s63xGGngzg4a0
ZP6j/uTr641xmUptVYDz3a8h+CzQw7PsQb2u5Azc2EvLDynfBEqK9X2WQtNEvBjmd4JYULbl/AE6
GqG/EutuwqSRJzNYSb+f/q9ibzxzm5T7hKA1t0/1CsBJICl2bv+20/7CAhVKIXefquz4LR8QXq2y
AxkIzn2yyEWEJxbHK1H/MigKlOMtyzHCc1uEbpRRqLGeDOzme/H81EN9X0N8j7o4C6tl7U4wvGFb
Tw3XAvMRy/n5yiMSF0V5SqCkiaJUg0R8LAgLvgrRj0SJ/Dn46ervpY+ofiOdBu8NpQU8xsKSwpvQ
3fuh6BvSHwQfyVX40wX89+waeeDYmgsVoXuOopBUN/sreFu6UFRApNDxc+Wim3BnZbmF6+VklpQe
ypNuziSKlyG41XaxAt5Lf5PXjKTuz2TnC9MZkUyah2RrgCicyopHvTGdXILdoDFmtshuBajz7HPn
BlKBk7YhLnOr9+5mTa04siqhLCxCGsq2wQezLjEKqoAaItg2hB47bLvgxgz+5ra6m9OiJxk2S4Tj
bQ+86R3FbtCkYasTwjSFwy9FuTYC05DwQdUmyps4UkK9//bQVDJrHRC7ZI6Ue0KgA8z8Mmz1jd19
2cRNa3MACs7V43KpZT2EN+K2jEWij9Adwq5bZM9XvR367AwXTznHY0Ji/0Qa3Jz1OJiqk18ef1wq
fRPZTsH2SB4Ft8tN6I4ye4j/Ts0qhYkKdDh1dFSW9x+5XvnaOK4/y9+tp2cMev/pkJlmQZEHpVuy
4L2JxRPtjJyiyzvQb650XxgafkD8sme1Vy0pEAChQ4Zkzt1v1M5eZMq47Qr0fbH/4NWYQngE8mEs
y31sFLsqlGZsri/iRxzxtXRpI2criGqMFECbAAv3LgYIi8Izsz1pOvjqIgqbH+YIb7aPAp4ufqTf
IC9ne9T3q+dgd0vX9Dtiu7ZkNPPD1cdE+IYZjMyS6MhC9Eih/7xvtOKb2+5BBtudihygoAgCuePS
v3fkk6x35ml2DHfZFRTu7fNmMYJi00QrZm6BUJRwhR6noDNE2aeDh1XHp3ixidSIxwtTu1Av92d9
e7j3WXEN7mun6jRUn3vIiTQ5bzk2gH7AMLDl5k2xFqK6Jf6vrk7MpLL+/RW3pQ6luWVYgGo6uyJv
AIONhx1dDtsaTq6cuv+PurCYb4716JLCxD4Rqfscf1Ux9xZ50o1oGmmpRgz8buMgI9eO0RXfDgUd
aJDECPdbl4hNMXsOgSyRYlpqtL/qnrg20sY2EGFe66p6u8qv2Uz1eBvdibnnV+ymvsb0ToCiwqBE
hjEwTyiXZ8vHdxqLcD9sQEGll3bt2ZNQDDLKw0yKbkOMHgOpuA0bgWj1rQH4AbfF3Vbb+eqFwXQ9
74Yr2CEW/Fvs1oJsLvmymCOL0hexnYorpjCW/NCOiCRd8edrHXtCNSJnXQpTGnyEtHUgPvzB9c82
JioSDNfdeteD7tjMfaE8SNOBl0KsvXte1mN41t6vrsMzo2dsaUptKY9bAELo2IhnkUhCVAkKMro8
pCEGpzp0BD9o1ZRANLbEQSkMZJP3if0+XfSE8CMjLuFUjrhMlZcxjR/llfMKflw6ALhm+PiwAtSM
ktQrqq/Vx15rOuswfbpt++fYx1SCsObHvm7H86707bHZETpJNNXcghcI0fynQ/ja4ZcJb5HR6/l9
FjqUR1BHEeXqK4RCq/lZK3jVvCwtP+h+VQNdfB3DVU91ocB8HsxqHBp/Eln7/J8mjo/3buG3Uray
aQ+GMAaK3gsk1YT9AgvCnBTt/5Zip6IT6R0wfd/rSGb6XPvjQt1saFxa0xoB4xF9++eLyItxXAON
LnIJ5SZIw6DgsUWsfSRAfiWCJy03+qHr09Axh1Y+EUHvdIXDR5RvVmR8sc6jO1gaq05nCRzg7Zpe
byP4k2ayO9diGBhsnzOZYxNhkaKehUgSIokbCPdfNBQMM4Ug18ZYr9iTP9fAI5dAfyIMwKlX0rHU
7fmfk1MKxVpt9eSSkmW7BDGqejLu6GZkRrLrp99ZXRnNQpkZtWH0JW+cv2xcpYC0BbYw8LTQctpJ
T+XZLwqQt+elTkl878F5UtIcJLexFC3IudOAQcC1IxCNhXphrSRwRQYzGb9Cx/tjGNaS8xsGj1QJ
WBzWNnOvm6QfKhEvkMFQtPvVzkMzkgVoKx/7OjvTQEfCg/0gdABlwev+G5YFnOOtFYoWNWUEKnTQ
yy1N4AfjoDFso+WXzc6ampJj1H/S1JFpsMfBREFJQHbAf95+Ji65GEff4apamkJ5b57PRkbvHYKU
SRPCJ7IpnxzKLb4z6+TTOvn4bpu4Mn82/xk+AFtLlWa7IYNXs9kBowKt72A5JpsV24Lm8lht/EnL
CjiyqOp/ukdnSoihAdYJkc/uG1PP43IG5QmAgPjkLVsq2EOIOr4eAbCDMcqymunCFKwDEvQrQYIa
+8dWcMRr4guIxyeAI/lvbrZiKkipFYq34Qk2HlkW6fsOIcCSv/7+46e9QfSNCEY+wnGvk6Fehcjh
Rp2pl/SVKrX5P2OnBh8TRGf3TBhWjm1u6HvSJTnhcKxr/s8y3RhlHEK10AUG+mLUexPyxN/g6V1K
xMPhRi21ydAnyEyvuD6GYMqk6Au1BE25X9k2T9X1lw9c8qIXr9pBjDFEq4yQTW7kkOXHtypwBAOl
tldZD0sjFhJQ4y+qWMNZEfYa554hjQtV3hmLG2c5zubXAdG0rgVa8VvO+pGGhCd7rGmk4PctPDjm
JnSN55b4MYNN1QYSl4LgRXSkYqNN5Lp7yDKJXOSTCspP5wIcf3sKNHoFvOBcnc5DdfbSshSJrLm8
yMHoZEpIGYH5PVHuzVhrJhwqn1TrShzbzj4kXhpO3CN7udmJB6apWK/RX0bR2TDRFQNBI+cEV8Jd
f+znrN30+tHWnM0VJNm1/vXeBva/KalzYotiN4ixq4O7vbtUGq4J4vLGI8ua6gf9vojEmhWlXU6f
oCpjWv58yAkb+HzGx9KS+qg+mdrgenqMipIw5pe4R5wcIkETVvDjr8/P/uGfIfhj1/YctlR6FVGR
hsh5S0p9FP+OOLPA5s5nT7MqGYxrv8u8xuUVgIkecms7aCH5ah5n3hVtSvNNMjxjaBa7YMNON+Hx
XEvF6yCJIwNkclxmlLboRY9eTzKiOWmH9ZAxJpm47Lm9H8exw21BQn++SRQRBhw9SdCDr9TvgRWn
ujMjd6Hnzz7wEUyEEgtgcqHDrFObcVD1bPrwxeHOe2tdAcN7awImqT2V0g+ynW24IundO6embEuB
2rVbfxqoK5t6gq8IRMrZBerz/l2iNw3/8OPM4QQ1408Z65fwf5nbipyMmIBaAMiXikjXSPOOQ6yo
tH1doOCnesEVfUEBBk4KZW5ZRJgV+FsOzbJdjiq980GenqMXweRt7zjtSZJAv6NVyvKN3ng/C5hP
/8vI3HX5Y91MniA/foSEkMg8GkGWH4OixswbSl7+6f9A0EeCXY3/zK4mwue/PJenqBQZT2oPBapo
ZzloZOAu4q4xVGPR9SW3r+C6CtvNp7q9O2JzKADR3AQhXhJDX7j9Jg1ylud5GGnaa7+IkSe8IMMM
nGaOdD1oKCzJym4RPl4nGFDvi/WKaXfYjHRqpH8+BKXp6vXpfD3nSgfAMMJ0enD/CQ4xXzxdMuLk
oLUzmzBjOvfNVPTY9kB+/iFo+Zs4KOOFPV1S/w7SBsa9iS0neFzMTb7Eg1DudIXzF8lIoEoy/z5r
A07Ot8gXYMawmJK/ACbvT/tHrQNtjZb6U3AdsC7JWsQWRfAUKwEyrJh+ytjwQ6D+/lpYJBxmmS7w
OsF5+U+CIfedm+h718eyM7bQGTl2fl67cPKewDo4w3hd4ZLObIrTWjvoCbCAQnUNRRs2VRHM6zz8
bvmnC4Q01adaPqouRxqtr1C2hQBiUg3h4W2bSND9NSlDaIzV2inMlQ+ypk+Wh+uCor6XXs7Ry0cw
B97TwEsMrBjl7XgRn8dyVO/gJBcC1MHhROimBuCfa52sq7hNs3webIr58OBqcf98PNsUxdgnFcLM
DtSvqzHV+1HWCrvt2nL/Qb7l8f7CPAOR+0s1Y/tr+tt8CD1joLpe+cGb5rsK/aKOGDFji2XRsnnu
JDMPf5bCNJAvQB7AhYMRba5ehbbB5LzquLBo7Xxc1AHzYwZbE6Sf4AxvYLJb2uXYmkBPidOQBXq5
GDZm3yrvvtncAUQhYVG29kUCelH0ZAbvGXj6crgaswmqAxvJhFxQhVmNQl0LJGdDCqyhrIISzgxE
9UJ1LHEJeoBQ3icgUqF4Oen/ztx9ThNio/3AywaKVuJPUqXI/L/2bou4if9TOaqSS/pYRvvQ6BgQ
Ck4GlDUeuaHbWk2OsbwSWq5ght/+F5kn04pF/IQkgClk7OzxWUJgv/eXh7cF1yz8EJzDrcDwLGe6
jabGgcncqTGOrbwaZsUW2E1Q3DjHTtU4kw7xVuDBof0nqU0JX14dTQMWR7fV/BGCTJP8tLjytBkE
1L9NuYA7j1DZWGaEeB7DxjANcef3sgDPrN3WMlOylTA8Tph1e+SDcC5EiC0gKGEIuDUir3OQSnAD
4kXpGZXcYaOP5Br0IZRWv5p2XUqNGYoeDq8mc5vSACM089Da4XNqfDtSQGy4nTAXqxg4SObBHv/m
bBMGQgjvyLftPvbMC+LSWxrIf7uLlCLXiCetvf7tS5Ny/zxZyUkZe1mNgEdIYbfgzogpc8q8xlQf
TK7UIU8/LGq9VXb4UgDzqb8Lc9v0ttC/mi7Wy59IiEmRblJ7yR/MxnKm0iSge6CNbogChpFVI8fa
LLnOghReJsbIGLhMEnKWC9ByfK3PEQbPhDTyO4wfSDN7InticmLX45KyimaRQjbY8TK/3M63fU6F
oOYuAODP+iMspOYDOuBNUbuyRLn3+D+4Obgu00pTEyZz0lnWVQ8NChfiVZWy9NjerLpLcCkqQGBI
mNhI00SzDwjdGZJybemTSv8jCSjthyTT2so4ohEaWAAPzDSTxpCMhMpYG1TK60RsaK0krjYBmCNI
nqRsKxvkG6nk0IJob52DT79K6KKg4x/oyae6DC8Ei9EypxEi23GhYOO8D/dhuR4It+cj2F7xPo3V
IWsYGewHQd2XWukQsvCYmUltrvsgzQ/MzLXvLk8+ot71tmsnLfajaiN/V/lI7l8eyDyTVU80UlDW
caWU+cckxV5ghc1fk8UBPPss0DSyN+WPWxfuiZXdcRAsumXaL20QyFfFlWrwFG5BQVGcYdtTmRNT
/ivuUfjOL0ut0HbVdu+6As3XNjnupIdqKfuq6Sa2384Kg7ntFpi7gTFCLxQyBbhPOS3b5FI4wxJw
NgL9XkYqTyOZdklXaq1eMHzqT0oB6/2UeAq+UqOZJ9jfDlgb3s5P3KEL863vJZe/6Zebmy1Q3NMH
rEwKiX7PYCCGRMChs3MKg3oY9pkYnXtGgrYLNOeEJR8Xp3za7/yrp+jM98qVw7OKumoFWD3oIwNi
+pFR3i+APocHzwV+cFW6IoUEnhkobi15uypYaQ3fq8/NFxxdYXygqkyGJpgfcYNZpV0bELk/mGHl
iTuywMlLsGf32eUBwOc3sWLLE93/wb7tR/QlMEVq1RnRfOXtptWx9wvOov51Ffu6hCuz9YItq6ob
R/8o/2VMDBIz/U1aRUoFLL9vMfUOZ7h+bvPt41LBDpRyvWJYfzPfFwhD5O9JxiLkVpmhKhjJ6lL7
oju924Y45MlEJmQNYHqb0hGIwvect/6hAZFDp64JYy+aVwO6r9XJCYyf2H5NF9R5iHf+cKA9N17m
QotDdhPBGWzuXsMUjkrleUrlZFg6EYcj5Ze4Tnl9/YAYs/5C87/Sr0PBRQk+jXQBKEV11P1WGd8m
XP2pys2FDOoRJLvsggzyR9qI190DHVgehonS+Y0aO/RtjG44Yzcf001D+3bBPwsS3WRhPXZWPRM0
7/dR+V9jyMU1m7cStuap+xgbmvrns3pjtC4xaoUwld/lTMFV7E3d1Ur3CJBcwj3CdH95acF3ZsYc
dbN05ymnGYPRRWXk0OpnI5aexgHTAGTH68389XYWBiHDuSKlqbYtyKFJyF7y6DoPWSulhsFh75Ur
JY1HYDoQqUloh5RfuJn3+lH3OArGx0gfYkOK8K9v5BvxBmiD+TewB/7HTU3KuUtM7KW1Swr/Bmxu
yz0YWHmFXnfelImMfqzBVvqkOJ8RVzZ0dnwVXxCdKYva6sY+HAE2oogzuSZc1l2eFVc3GRVLMm8M
UtPizII2JAryEKLY374asOvTY7mMxEoYwtIG4BrkaLIhqR66qi6yKJixRebnFGhQZwqbNWSN3xk7
f5Ddze8Zuw5P/AAbBsfzKsB7zAgcnDmlruqp2eSOjv/TZXhcMO2AAMIJonofX5Xwj2c1z8ps9b8y
DIcjLagX+o9xHqUgYN1ST9puU4nLJ8zwhZXq2qKGx3uAntyKT8uTJynj1js37C3CeshVVLojdr1S
JdT0RgDxW7uOaxwqzx91jJrxZTMdMOwDqI1R4Xsujt/JWuzfulFPSZEXDMFukKg7rVmTgvLKKDja
8nDmuef2gReSTZvU1MycTIgCjv9Z9S8Jm45UqK5JNr0wOWM+Caz3LfSJG6iGEgkIkMIL72na6rBN
CEBTAaYTXiR6KGsSVMMO+J75MRREQ/jctzVffFQ0GZMNM72kg+/jHtRs0ud5AMJU6nuwaMTo/LTG
oNg7Tj+EiTJq3+GIbuVFHHpKaxd7cvDhpe25h8jr2uUhdXDqrHIGZ6ouf1psHNMaACFf7lNnPLYP
x0Elx34h7eVMvclp/h2+CZAAATN04KD/LOSDIMHNja8N46Ou/c1gu/UrkVOCAF5s781GGXLpb8Pv
R7EbptRVjrQjk0OkxxcGKsdRE0KltQsoKPXdPe3eUp1HVDv/EjHRWqiXmiAgbJ6+dEWnoUi8CcTV
eIC6mDqKbb+VvFcwVoJ3Rh28S68BqhpqbZe9P5TcSzyZlUUo4bljNBHwytGBwsCSs6Zm/syAwV/Z
jdUReLwGPco32GaaZqWGiLfAyC7dA7jE6G0vc/2QGp8zkK38Kdo8aQAFArW08zok5g5lZqCKFQqC
SFQ8WDqx+0KnRpZXN1biYgGkn0VhiS5Ca4n/7Ey3IcnHk5Q+wN79KiFf3TrvoqVXTV96m8MlnJSW
46NFd/PikNO//yn8T2jkytft+VPB6NSDMoQkaJApS2G+2UuSqJpQV/qqjbSpOkL2uPKGA0a4tGBX
8AGJj4cYx4qnhHSkHwL7o9DArT3Qlq8s2TBbOsrmmFu0DXBznmjqR6KYV03KKD2nnNjGHxZzz9d0
G9/8/ZuwceKuVGRosDDzCNZrY4IKUe464o6X0N9990KTRL0Ea9LImChSYWkZpFigiOJkfyK77b1N
/sYXddhBETDLm77HvevE0sY4mNC1974X4Nt7Iv1/AzFbFhd4F4L3EN9J8bvqgHSOyTSn+TiTm6Ti
3VTPtG42d2NnKvDjN73rPrNXmBYky7g5Vuulrdk87uNBFT7W753UsQ3OUM3IyQyaX1T8ztVrWf2m
G8VtNmx84Ry0x1dbBell2X2WjGTMhku740sK6HsMx8a/8dsga9qAkujHkjhuoq4vgoLvSZ2/3Iuz
AfQBcdUQ3XTLkyFDbX/so/gBHQcQVKgDDXO8kLens8UrSvcfGzgLOI5T/UtOykbsmIJVTxHpn0xI
wqScvD6gVjrIYBznk6noHqurdCqTH89Fyz66cqTXdTLAgyyGyAEp5C8b2bWMXCH4IcRb8KqHR7U/
InsZDBFA83UkCiFP3Qpwh3tMMA9CMqK2ItNyQnnfrJXCwPD2/tEbCn/DoCaGiUEfw/IfUZ69lEsc
Pd2HIw5x/X/KXpOzx8Sc5XDr2z5SAG7i6BxuXJUUkDHovkEyq6UYlckCVvi9f2Yh7O6Uc2VUMVKN
rJkmO0kAJhR+6xVNFVY1sKwEeD0hTGtc3b11cveDWT/KimxWmBy+3kuwytUJd/5GuQQCPcOMrBNu
dIGF9UpTAR+ECtWXJl2JbQYR+4dDpWrbcy8LRwb+d3fbCLNSlRa73RzS0DHUDOJkshdtfNrZSw1I
NJ4MXESVmTElVcDMasG00Qv8WNVR11hlJ/mpycRvgFgJvIm9ko0Yk56Iud6/C036RtCry/ymVJnq
8pWbWZB9mwFnyqW0ComM+tUcKvp00F2g9caNQbpYNfSJ8GmZG1g+hoJ+Lk60Td7usd6PNyftTAQJ
mXWGv8x5vJw/VVBn5T2rodNdPRhJgy4EdKH0cFPHoApOo8sM9IBmPaOrBdEYkoDDcJtb0RJ9vvRN
Y1GbeujtrW+TDDmT77tJ2sOfAbklTqf/zvcXjDeC0GIXEAfbGIkXRZZPR38a7xSnE1GO5HWofr4Z
+biOFEE+ycRaxgrNCA/gx+WPLKMrOtDUeH18tpSfLucb6xQMS/qGLxAZnyOqrXnf1dbiBf1WLAEw
qiMJqNXsdUlDqabppMaoP5IU2G0JTeqRqcskwehCpqT5cvwFnlDuYiLbRzYwBybD4Q8WJzo/WzJl
AAIhY19aBH3X5XIY9Tfm3Ox/NNagSSAUd/q6nH73/zE9WIEiHkDzoXW7kAX52KrRfZAqU/YOx8wQ
xa6+PBpIKPGYg1lQopIxWMvwULCwfiubFX6shBgYEfnQrHecezEYG+b5ruulaTeqQtk3hf9b/1kk
i38BHi2hu28xhs5qi50d7UjtkM1hVGbO9SVM4mcCYi3ntoUu9jRkHA991LNPYhfL0JJk1o2UCXkJ
7cSAmxOkVUw+zy7WdDg7KAzWK5u/OKk+/8/MOtofbHJFetTRp6navauwyxDRTsBnTpjN8DHZDGje
6bek7MoJJnDESjMcbuQI/vqAJ8srLqN8aiaylrZc8+SyFf1Y+3XU6vV4WB5eHDHEXDodBFOG32h0
OfEIF9jXtvhZCd7YB+0T6IKJgWrKuft4RDKnk2PKTQoRIpWbFTyJGkHDugs/e/ANt8xZN8fg8ssT
Yubmk/WQDSENAwMOaddGyphodpFKDnK9aFgfCkwlO3QLV7BWVLwnScfKc1TGgKkVtpmebqC/etBs
vDwDeN1Nt7wwFpkzs1QPZAubEz/PFzzu+HTXDvlCRFbTZhT+QQg+gpU4rY4VfgOR7Z2NLlX8p8oE
rUTVqftMdUajx0bvxq9ybYIzBj0M7e2NDMZwmU8H4HbzFdiNf2wT5gWH6wioqJCAl7B64qy4C2Qd
sSQVWut7gLBTZ3jY3ySr6rmOY+qbUf5omc82g0zUbCMamWfxTq/klFXFF0ZDm4ESMHd9wMOmNKvR
y51HtgumsxaRa+AR+btKgPSsepTheOTr6Rf/d+ztNLta5Za++1fJapRvTgL6lm71WQWuRGqeFQ5x
NvmKdyJ5LuvTrGdAE7jq701yGifEQbw+13j6ikHrv6xjvzJ8DvybMqpTsk2GoHS5Ju1aNcM46afl
z+drhJ1t6Z67iFTHmaiDb1cSwFsXSuV3eJg+Tdm+FxOlD9zv2mpTObmskuQtrN4FtW6FAyMOhqhf
mRBqLP+OrCn9fwtosB//ZO5SGUjbRDsE6hveFtiTAVAM/yTYxbwsA22bZql/Z01/CLgymGyn4xeD
zqQWoqX8HK8EBaz3/5A0sK9qJ/qz1837JEuQwhmvzxltUTKP4lN/Vy9xbuXQFQ62W37PQdLbgHlq
Hh49Qff4uKnkRara6TgB7vJOAMnLv1fyywfIKVARFKcQ6k49nCsMWeCMANtMLzDdpvZagS9EYuc5
UKi+h1LfowWiZkQUG83/q+Tqq89L50gEUS7fRlHcI7nc8/7Uzu2gB320Ov05GF1FIDzQKTWkEZ2y
yJGR6Bn+6C3FvxGtSDSfTWgmumbXffM8l6Lf5nILmExFpi3wnOd7c9A/RiQHcKAAMP42/x9h5Mtd
hYZOMJq2RcPEX7rCidgZon5k9IB2uAOEdMGJElNGd+sxgiEDnfI86SXQoB5ueWZht9Cn2rABLS3L
b/gorkZHDT1OkI5Fkm3hMiWTnrA1L6He0YxLhlUHaSeMi1E6e10oYu/M5MLdJCx7BNN6B/Dw8zSV
8pwSlIyW1Eks3Hy1NjFK0WarrH3/TxiJI6rJq6QoaNKJPRUmoiDex46N1IYuMmjuF35w3j97gwoF
kaEJUqPoIB3prjZ5dthwpoAj2HVJGB70B0YF8zFLXUq+SwM/K01aJGHBOzo0VWGqG2EnpY1Kxo02
Y/rdHpbte5aKiHyxMzTzV9Wp6FTf6qqmMrIEEf0plV1ypsWbivQ1pJUZFJMDUIMWjB0wd0sTPJ9r
bMx/ArTlthuxaKe1IuOEH0M2Zjs8aVkuhnd0taMlZSB+xGBV222eMNEXS1LmqqgMcZpodyHMNhxj
S3pVjaBuhFJmO4zDwopNt7MvT/6AjPVaqURE0A7oVfaZKfnF3xOu2UrLdkChEYahCOFE4z3QUwsl
zG8eToNALL3+GU4UgEw1y65Ar7KOBHPjGg6kkUh6La5ZhtbVebECCqDZJBNuchhNhl4+Yg578TU5
++LZhCC3J9rDihamP/t5PfNfUikxoOB4T+5Oaflow1ZtjsPAlM1Y3YKyrQxNEj0XD3jiVHHJtjaj
NGePVQ8Hn/ve7QRRH4/v22LSAISQPYbljk+XZxXLMbycfjXUUnaZvHmFVXyHFDh3FOxS0Pe3rl0i
Gb8qYPBh2OZRRKgwcDURK5/QpVf99QPbT55gq9WEUM+6uvJ1EUp7vMawttFR2Io8Oq3rgsfs+vn4
eUm19Vilk5773fjbbuWFyUH4uiMeEVcUBv7vvWJ1k1IvXLHo91VVk7hfByOch7vvmPY/UW2bwVos
0rM9wf7wa9jB9RT5+7CYjwNT39uuj/DKNaUAN1xKgsMQL0RJZh/XWMZe1WWVDI9U47tqHj6EIAda
ud6eb2+mK3WvYRoh/Y1kHOtuwzpei+s9OP3DDWB5PVSyqQJFlk1qitzMJXI4LZZph/c3Qb6DdPHs
E7ko623IEi981VfaPb7ynrdlj+mjuetL/jusKQDMuVTOI04EkToGVSK9N0ngi1sT3ym3TgeymIRv
Kc0V5UGGCdqYpcSALS6aP81AKT+1q5JUSjV0Dk+8hQ6c/SvwTc4Ce4bPrsswbwg4vodrglExu2ag
x7cjPCFAkeam+YPcs6fuJk4HODUGgefyUBDxwJiMApdUufZebnYWK7MXCAg2wRF9thOdvbHPnbr5
scbSuz2l6+bSVyVnQxMv9zgF0XmD5VDepmpbBZdnsMwSUcd2sN9b1Bp6f/rouH0rK163B5gPg551
4MiQVpwHitvMWZqz11Ln7ydh55dsjEBY0s4+xDZQJ3UueuCfWbjcR4RilJZaCMq/M2/GX89/buMT
sLXY1fKFCZI5Pek+QZEua9YOHhiOdtBjThtRHYPb+IML/458rOH5t7VzXOxMJTabjWydrDdF4WI2
4W4CfoMHl6vCRjPic0QD1THNE/TvAtUCwMjCG2G+qkzBFb/SuGAFiQBFiDX/MU/Ok+DSLq3SLRbC
tU7LGP1YWjqnbdl5OX8kzmh1ek4iQnazuWnDmLVn4FNlOlUs4yQteb3QZS7h6W+y8S3pGZe0SYx9
ao3uckPd+OAabZtYoPbs+x96J5JwMMAu/u6SEDCNDZvN0gOmEaQl5yrDwFp9e+cCR5bIVpACXo8a
L96zZgu6FY82ioU59DFHlp87nVAwgeMjfjfW+v/tCKyjAM+y2tiBagD3g7mPIZYG106I33y4axqW
xvP/z4Fh3GKXKe6KhLTKt+Ts9zLojQRtLQJJr9mSn6fR7ULFlhLMxgIOY2Dga1H4FhMl/wMDS5+8
EkI7YoConyxXpoEGtNYcWe2NfwyWoDCCNnZLBeE70MCK7t1ef1c1eyqiPy7adsrMYnKGUAbTMxjd
2oXCCs4FS2R7C3i0r/Fzzclz1VQbPmGr6QE9XkLZxIcamgN5qdBNfxxz6PD/UpHRrTR1r/RXumAk
EZdPkfaM0tj3URcPsgw96IvDjGhL5YpwzMb5CyZgGWjcVFD1pVEQBmDic59pemgV8+lMLG+2Hdcl
jDmNPlfT1trjKbayiKpsIh70oat83EmMaTTADdJEFmgXd6NkEQOv8nwMIwUZbWO2BoWkEI9YJTuX
oami7AtX33TE7+19v4wI9AKg7Zpu49UCXr8S+d2xiT9nzvO3aLIgFGq5WiSRx9ISh6tNQQGZirq/
W6BuTLSpu8gxuGLJWWbqSHjJQCUhQLqjy32+ckOsvTAgNI7BiMAKKpZ7UzDyNqScP9ZrdlTIWEho
ro+sk2SgFIog5qBpakJ1faLJOLK8u7EjjfgccZpzYjOhU8dpHiZLQ4UbIbCVw17e6xvYu92/fZSx
QhO8L0ytB8oNkC+CfWPDysrS3fvoS3jTQow5td1mmCtotU1pbIkpKHDGuipTKspbjF3YMtaeE76c
Nm9jmaJGo7WwTwWQv5waV0m0vBaL+ZIASVI0GCWuiQOR3fmA3oU02AdKsqcyNUmvCERT91yVP/ka
DzJSWP+J062MHRcPaNoRL1eTxNsaDvlb0ePrTNL9bLacuq6ko7hoBRjnHYdqCzI4Zx5lNw1XuIRg
y0wUkeiXwt+tIToN4ur47013kwmy6ajGLzZl/i+OJOMOZawbU8SWdjHI5ugUkAL/0nyi4ABw48OX
42PcgTznOu962LRKfUVjQPsNs/209arG3I0P0sHAdY+3eWBJtNKwtuItmL7Iwjfw+98Gg7u5Zj1b
mLCnBE2Pcr05/3dpTamayyoHzDHuuKKSiX6cL0CFv/p2fg6LKQXr6jB3vE3YLNviQFSsBhRlVho8
6tuyOb/5QrXmmJDFO2aML/s43T1K1hQCufjaKvanfUCf9KcZkPLSYAYpI+48LG/iJG5xzpRT7+sT
WcLDHmkG3HPNkDIz/R8pAWkOt/7usvIOl3wX+JcFjH+dfii9aPj+mqWpGqaMnIkpbGKCvzpUGYZB
bGqzWCuowB7+Spz/aqcprXBFycQZ3px6ckcNg+6lBUS3BThUmCXLEaNd0xvMr8/MFksBAKfD8Htl
FWTJcut9UfKpBWZbhWfiKmVznWfKNSER8FXGsgOiBot5X8QFePwCYz37hzGZKxTZ7tQ7qa1r8b9F
Zlif4sknu+rsEfA9anIzUQidUgvjE5GnuDrznbzMBGCd6rn1DMZPimRi9uBokT9Gq85KEMbSesF+
685G3wgd9pxJap1OYXNPiDyWhg925VpY7xh/CwZCJKRjTFqRBL14uVQRPKgjmwtmTdw3bphZ9C4o
JphZCkHlKv85l3f1I99sArbHgStbziaTFNgZ37g4Zh+GOvs4Uw73c4sQuUOsE3Wt5Vch8dE8zJUY
tUSveBi7yod95YSx4pdYghtZkT7gcJ2vJqKMQZg2e6BePA7VMBhCqfmNmVRGEx/8kW4mpgLmJs2+
0EoVJeABkE934he5elCnMYW9DasJEVSagRzgUiy8HfBu0CHFeAdP6Zec+tG6h5cxNQOwg2iN6GJ1
3TQflQtaIw6/tsnuQv/sYeCLiPiQJvoP/K3aQ4FG6le1lmI7lrU8bgoL27x5OoWZA+IX1Vr3OVl+
JHXfJndRHuKAAy3vMxUSyi7Q7ZGcmzcPfuJRMUYlku1Y7iB1wbF/Rx/LuOXI8XByNuSGLL9UmwB4
PNWzeeuOT3wZbdL4LT3zeQqFnUm+0yoYWmWL6DPLy8Cnpl3tM9ZN8jE/VsR3vl53t5X6oDnKt3Ii
GLgzbRMBJocQ6nEtK/XiMAI59pPIwqDGjS+nsq3TQRIdFO8lzWVkWlS4RUl5aeZO8PpuWwnFfMoM
DQVcyfo9M7xDTrXmH5fICjqcRedzGkExaPWdKeNuu4vlyKioiM369kVUOrQALZskCbVxl8dUIhRk
nauaS/folSTXgBTevia3Yh6IH9yIstf1O8dgV5wA/PcaF47JUplE4h91Fpz9tUTDXGdxI/L2wT0N
cBbFSaVaRltC4UMu/yOWpUF+kzD3mNp+DU0Cgac92y8uC1DbF9rDjgaaKBXVrC2WuJCXUh0JjsKV
r26ifVLOxSij28OCyYOeTCm0k6pyCJS2tS24pbFrjT65dAmHAGu7B77CVaELZyLW+Jy2ajlAx1tI
jMH6w4ocA1fUBoYsxbN70UoXtF+JhORZeghHhyPkQggm6dILdDEXMVuJHJ8d43qGj2n6hMgdb8JQ
qfkg5WomO2KVuWEEVXfYeeFpr6+E/yipbyTK+Yxmu/PkEy4DM00LUrQzB1w1BYSeFIUgxIcVyuuP
SCd25JKJzosEwG39sw3KuNEV2BYOF7P2Y0OSbVXEYuAgtk8Vus3W2XYcKRy9fIS9CzEKe0hHS+PA
UKID8o5wP7gwXoBpWdlLc4bO+ssNznEfewPoEJrsKHs4ckqnqgRqcd2bGNTz8KKNExR9x99ChGsF
Z4I2WQFENPSHrxsGcz0dtQitvKkxrQyxhgGAS4+4cK2hyh/RVPyoRfqsiOVKP9NjgpWBAqiCD+1l
mGd7zFZNmdcMDrIwV/c2bOhlrwiQJREkw2bx7zpZz+LHLD8i/VBEQ5x7jteO/Wh+7PAESNv4YyjM
W3nAlm1yV1moakTzqDE6FQLrpmVBp6hDdbfz52wW6NaCrd0tDW9fkjpLTdM84bsTaWkB4qhoZE0v
nOROqWawOmkvHCmTz2SGrVBEjuYW0EDE0as30642n/mlFGy/Kx8vwJHJnWOQBd0/bLYzawpl9tRb
CyAgeQXWfo4KVYTTYcKep+bP4i5LQaTQEJ+YymYlAbNrkCMgEzalQcjWvvBKaYD3IjanXgNEFcJU
16PZA8G3F0siNQbPSyn9kfz26tw6vMSFFjEuthyb47jgZ8Vwl8x5uS2pHFTtQbZgdwAuRUMw+nNa
ciTyWvNcgMzO4DoqW2X5CFnn4dGKZtufB9y9FO2kCsMa7MCI1eFvNhxA9WQTMkhpXSE50N5JmOl/
OfAakS66+njQeHaLCBweoZY2N1XhJ4mwjmdlVb74/plF0U0eSYMcmOvJlrIqUwb1zZrK4V6hs7KA
1UmeXbh4SOL54yIHfIRjZi7cAxCV3xWpk6YECZTDatj/C+V2dvBJA8rfCZOtkPNspK5qmOcLBO0i
iurN7csrEqLQ/Cgtc4a1yy5ruwYNGJ8Ahs4IoOT+KENhwiA+aPSZmWbimFR+xcfPPW0Ql7M4x6Y4
WtXJlXe7cgOKmOz69BtSqT4Ve9pRON+8vv21kh/4F3p90JLbIcYHDRnLLl1kxy1Zp+rxuXqR0vuU
3+uTl+9gro9pM2ZWIkdWOGsDqkg+ikLrAvO6NSz2cNgHGYH6LSY1MHOR40SF/GH/k8u43i30Tc8i
vnKfYX5f4U7UbA1Jh2VD0n9nnGj3xxyrGAd+na07IExUDNnjFK0I4ltG1eOExsTK8IOLRGU+ksQ0
iTWnSLbvRFhRbjUq21POtDmnRV/a8lXd3H76lI3bYYK9EFKVjNzCxkVYjmJn3CxbZ+inJ6V4R3Nx
dkyLPFokGV2d1cM5rc8YG/IrQD5t1PL2y3kfWpzR5xwK5/deCCpXJ7gOZPXv1qYceHqNIjo7kU42
eklVvgJCotANDMrjKzPK6quYQt5uFrftAgNUYMtnEMmD8VlyW/DXFfVMSHVrmJh124Ad43IVgchI
WiMZBmlDXS03nZ6cM+nXEaXi6Jb7balKA7hscoHULAv7Q/ZyUgdVpFbXXIChV4eeQN/UzsgQUJ9T
nXJbkmreKmMWBksJqRr7oi+2GpV8dIM6aEVi471GdcpoAXqu+EAbD8cKYhR8jykvmFygeE1rkFyx
z6gx51j/VtNYN8SJ1KUOdxOWjFCFZdhAXzXB9Pgq4Pq5aMoEx1jJ/4SE76CZMRR32tiBrl5gQOD9
8QH5EwzlgCUDuY9gNrrQBNYhzonmLwkKbCgUHSyW7/YZOaZypqg243Uqxuh05/40o3l6TvGBcHR/
gL4I+Ig4JZeiot1p4B/ZLuWW1VNKt2mZLu6KN2VaJmXJBr0kmD5z1QUrqs6VvdsLPheKekIQuLpG
kjCtdLIf0F4YVU+L2GF26vIa4mczxXpMthSiaJob2y1T1PKX5O0gffvaGTXCYddQGD2PrfKYMLd3
loTYYtdY+3EXksyYw9ne2IBmjKeN+QoF2uFQcfkB15HiAvZ45HR5qm+X1TqGQuoV3QZ8/rurpGyo
Sxbel0AtOUWMizHmRP5uJ23+qpK1FoJCi3OU7DOcVKuTDKmdbkXEHlCfAeyD/Po8fQYI9OlwgVOv
tyyEjbUT/52lSooKGk6WZTGGcLPoFTlulFjYRPkoovWsfn2PyS7ZheFjOMqT/MjcYnMa+zEoXc+f
Y31uLV4CvsOpUNzOnWRW8NlBM1KGxbRH7iNoG1gxUytIfZjimVmmlaGFHOHqlyQQ054FsvUk3mku
S01HLJX6nREuC1Kx+lLgZ9yQGOCrf9omLjJGLhPB3yv8zfs6fU9y4YZUUfHQqCLAkOninijDb4UB
q9KDXovlYaZ4dEDfTbNEaS81dnaGNQWaZsjNkGmVAchd1ner8QXwIUwtv99nvLXQjGqH3lhaW4PL
7Txp9VuA02A/E+ILwN53FXPIHfSLHbeAk7QWgSimurP2oZ2DgK+RdD/QkX7Oaq/MBlERkR+S+ueS
M1Yx8xCSKzPdwqFov7IBNpwJ4jBaFXmdfA2FcmATalV/n6oX2YEFxlR8XztXtwhOP6WZx/1uNUBY
fgrPgfacMxKFU6uT9ePc+H2CDmVRhDWJskvaI6gx8SmWoz8IjHDls7egc0glp5nVbkq9krVEgRTH
N/8q8psY1rajT7EQIT2GKydDUFCjYxbR4xj5Y8RMCtq6sjK+gCos7/skgnu6cLgj0UrJQUGaEz2p
EGgAoMVQP3V+/fic916GvvjvEsshBAtm25xVDm9PxFJ3yrlbwGH3SmqS0AV5HKqr4l+IuqzTrRbM
rLoBKRPhtK5fcvCnNFefOTfl41RXZkpVkqy3rNil8TcJecH4GGwcLeB9cf6P5g25PcX9Nel330Ke
uikUfWM9/F8m5zfqVmGAOzZz/baOVqjM/Ec47T7IuhM3QIxpagSE/65q1Zw4AXM0bg6SoYJhvzs0
JkpHJmhxG7BTxWep0SPKW7PzU2h9A3ExXZNP78ZQFptg1t1I0xl1f0K/ZZsW8rL12rOSCo9mQxYr
zKCZXyKsGblnXE8iI9VHtbwlQriavnSksEGrxSSUI06gfqLEGDFXl3IFes6HkpFuLroxUzf3v33M
cbe+90zc5SExbsZJulu6QHbUlNRuOAzkvM/HJr/nE1BdfVzZzWzb3wjJPqWDcEvOoRAnbAayZhco
JufcAjwuxJRwidYOd01GhnOFFJH+UKyjJq5HLxrv8cyu7xdabiPWzdKUJTtY2zCN0o2/qgMWPFu8
wbxqeVWcSjDnKzJcME5dKqZxfsIjq6VR0FEtN3IRUkdFqpyGTI/IYNAi9XTFDb1yf6cQX0oEwuzS
kAe7c4Sdp/jvizmcio1N7H6f6DmVoEIzUwWAsVMkjXbPPo1AItQLF1yu7ZgVpk88a4EsTCOVamfw
YLkAsaJAVoQgokFk0RRA6gYu8xOHkNmdW5BMPALR4jP0FLZpiVDeFYwW9JRfe4MeGOTtlki87+iP
tK5xTBmNfakObTgW7ZETXNsp51EonOQOtkkGBpl9adZ3AevkUlUMVy6Zoh9cnonEPkF8ktDl1vVN
oZO3URLDW0eIweULg7avqeFUtCYIsX6iNOsb42KZbf+oldSAIwu9a+neYGPeiJZR6a6KjyVcTh2X
j14niHfF9C8crndDWe2CErL3evDe8qG/FXx/LpQI0rVtSA+/xiom44NNheul1Lqkj0jNHmQTE195
NRwy5xtha+JqPQ7uZl53X14yOQhwyQGcvfHi5et34DmW4pevq3i7VTMTD7nr0tM6WUxIYq0OYD43
z8+oSIeU+04uqHAdcP3euo1m0zvKbyPh5xuBnBYMTmr9VeHC8ZjICibyluHn7AUP4l4mlLZGHb7v
bEW5VxjSAMbYvjlcPIqIePo6XjzvM8Dr9HPQ8eviNcZ8oKGfeoDlr/MTNigYii1yI3Z/wgaEZiEu
o/TgeMz3RFZX4wDY/ZYh/fYiZRcs2rrt2e7lVFEkiq1OX3NyElAbXBBsNKIXROvWTOWmvjYTqg4W
yPXFrtFz8D1gXLnAandDlObVzeD+fShWLwc3yFYEeAFypDgTir4aC5jWj+rlaWVjPGUEkN325uZj
LvobHEVIg8nwNF3Maf78CMGq800X9w3Y920Eui/doZSdM5NgPd6hRWZ8k23xFLd5Y8s3hRHE5Ml1
eZY2hmUUs36cvpp2YxA8bwvB7C1CLLq7CA4W9maARBBdisICfRVI/5fI/FCL5Q56U4EoJvaeH3Ps
avtLyIdR3d9PdEZD/IzJNkQVD41XdBqGvBhgfpYJM100KjShcL1Il2HztHodeUYrH05rTmNMfH8Q
YE94Fjkin+Z/msrUP+LzrluXBlEum6Vqc3nOYRfyskJlrnpuh72xt+UtY9pM8IGdTLA8ETWi7hzl
wRugmJ41IL7RIePbZjs3vc7kloC/LiOwmooHmAnrdwGctSDanM4yGZgmbeAS7Tdeq9tnAa2nuvci
hBEZiucOX4FrRLu7u1lj99zJm7rLI/YsGIEx4tslUGqxm32IOgeTfQuIkuBtPU6QhJjxRwjS5LEy
efLkxenGJdfLzg2SpuEbn4rNwHY5ls5lx3I8MMT+6AewNvZxX1H4/swM9CwdsKcIt7oGw3Mc66gJ
LmVanb0qx86GDe40uArxwr15NoDvPdS+n5K0cVvL8DD95EKqxH/HMyI6Zm0XVJYHmlscHB5LxRm/
1RA4gVxuC9/TyMavk3Cdh05xvvlhuMFFOGaNlslJkX3X8SHPCtbaby1N8q95LDJI0Q7JHdH7Hccz
6ClWHo07xLXY8/8rGwGFHN4WcJy7hmi5lj/qRQ9Ri6Xo+rzNhZohKdfxn76nI4SS82KHlayTCya3
bZS9l3w7YP/Rc6E4ni6cYXOUvg+yZYuLQIuLtvYl5nOeFFBX6AEeF4MIuaxoEcdnx4xYN22nyt+V
UptBc3KzmFhjP4rVzPC2shIdrY0XXLiZtVRTvJZli7xXgKEawZA13dhM+rm4mZETTW4WnJdMyBne
jBJrHKm1Sdq8YvS7IkBYxRyGRTFFPqGbHfZYqO+oxnCXn11rIU7qChjuUvZYKRsebnySbUJaf4xE
vsv7vhEjnX78srXnsbEfq2IeSH5RuAmKuszm9gNt/YBXF1Q9/dJby2Pl69P58PmKN4e8wrkd7jNy
/oVmncHe7pkaEmNPcisFo6LFuFWEfoTjmzdEV6sh+9kliFl2DE/Hn9j+XDUTCQ2bZBpP83Xk/B6o
ypdh1rKuD7ugdvSFQOUQt93xkoulrFmFCvzqFl8+NeAsKNXH9DLE2EbmRWlk2jk8a89jt6AQ1NH8
bxAate0q6I+GmjAXhckVCs6WYaaMPI9eNHoorsPpLu45Tz4B8icJIhhdwJ44rtlyuT6L2e5m8tUR
HoSkG95KhZ6cD6zd2EBh+R1PF6KREf/s1aby69DixUe8EefJR1jRVxZoYxTcQwP9JzSDwlkUNJ08
KCJf7tmVEFM56Hrnoci2g15ru8Zi96o7/5z6I5VHB8aM7Yhvmm9c+rQ1lzFB+Bj5lPsGjydjVHa1
xOJ9ExYcdZgE76r13DNshn0p8XsGTno+qFnEz5Cdbg+fSRS6p+WbuhrvAjbGncUMmeHiNpBJYBsk
eMLa/GGj7KFgU6AtsY88N92OaTbK8WaRRaDJKH2Fh1RDKRXt6unz4yiYPaAURqEEXFmrIm78rlYH
oH/H90zq1oEnLye2pXMkyC63sMgxcq3XUZVFtmMDIyqsq1CVRa1h1knM9jaWyJFoqWK9puhDbTmo
/YyHUoyBR2hBtnIXYcVfwxTELCBtO8bpZUKi6kpzd3HDwGOHnsne0zmbZ9RNY5y6WKyJCwEv9asH
bZXLLN1GofV0bRuMZeQg3TGrBF9zEyzHRiA1gQSOJXkVOn/x/Z3girt98WF6YWM47exCpJovOZje
FEXBDFsGKGMPTtgw7HIogbhPmNqDwzgLJ/ymB6KWOzbNUc1yWMnbt1WOzhNAY65UF+5g5d2z5Kuk
VMo0LtoKygT3uAlv1R2C/GAqzTwfbfTG62ubn1bhY8QN5TVn0OZdFcNUsdn2iqn5GK9UvGV6/DgK
2c5cIMmtKwqHeMBZOK2bSGZN0uDtvy1RRt8aPnFEYfAfu23GuJjWyvKImzivs1V/96IdMU1NJOTH
Nnp0yo4P/qjMmEwWwvgtf5qaxUUEdE7hkrsjNj1q+3yYiyEVqD35e8NOGc4zkewYeI217NgtHfHt
wbCcbbMvsFLDpWdgeFrIBpqyvH/ZCFEqoAudjVFGPS4Ez+0zHuAfVrtMjEqi1Sq6hTOGnFqHK6He
KYDDoBwl1iQYXPZPz99SJaSgz/Jy14J3eTa2ZGUwXHqhKa7QUZTHgBl1ONHWGHbr+iLbdQycHb+1
TbsHg0S25loSltVUkqlfLrh3pU4h5tNAdxARqUBxpzgp7oLpAzIQ9Tzl39dP8SwGzoPlByeexsg0
saCW/GttnnrprwvCAEd4U+pQwZcoY0qlgg9m/OdJqGpleYArNsRMn/1oNF9rZDfN6I+nOSfr6gsQ
Y70Pjfqo8iLLPc8ymIeHhGkY1UCsUJoBVrvMvJ2NPI/8uxxMLTGJbYcBU36eA27kbbjD7QeJ+9Y7
F5QkBJjrUs85bRgHKX7gk6Xj1lfTaHsMAMq+58KlsmfniPX/0+5oezCx0hnyE1BeM9DZWVdS4+z3
9EI1CedRJJlvjwHSKMy5aLyZHoLEP1cwYnNARZXPZklQhJ0HgP1DjoEskMFdk/BdkyASnke0CvvA
Ek3WuW/QFDkD2zN45qbJ+ppgbwTZAWAZ9aXKbcFRzmdhhnz4Ofcl5pR1prVMnj5WxYxTrK9Wucl2
2Xu69vsXxRHDqNbt5X3kBOByUfWESOb852MMMzTKk0mYBfQTVnmIQGqIwIDCNaK6v/Cku0FJWoyP
Czc78NG4s1ktzzPN8cM4HTdcZxEfEGd6508TN6P1iCR3k5oGYHsN4IX4iNC85rWbMc3Ws/yOhTP3
qdcek6JG5RDJk39PKYDPwyEf7HCbfDobP84c24BbxA+jyZ6ANcVen9+HTpqXNAqOZjLsIlNcsvEq
OgAJXCK6WXZtYLafG8cFaoaRypwcVUn11L1UmKRlkU4yEd3ylXziVW7sjfV1ENHAqFtNxQgcNLUE
QfI3F/olf5wgSLWzkZS6dDzN2CEuNzwEmUQ92KsOQglQpxLn1rsiXUl67+kcxQ0a9QU2SRcj1Ok/
T876lRZ+bpXOo/IGRns6vd+7149blHe+Pu+tLm7Ab+2iBh/UDhz2x/yGZjnPo+/y1mMvUHka18rj
Nk8Rh8uwre4SxmDsc0m8VEUshJ/f+q0OZsM8laq/dKJNxAeT0YkgMADMIXe3bOxBA38nzEKIZDfT
CTJHz78f0V6HjXJm4VQ123qyNTR2EndOnqHXItE7VUmuifAVvrWbKtz14zAmPhHy0D8sPphaMByU
mCnLAslYpjvxPmKiBPiJUUPqScpQkO1tooCxAgXuBXpS6ipVufUN1pEE7gOjbgZXGrzFwHITCLll
7E8/8nqj7qKeH5SQr4RdVl2XXboVIh0s+CV9d/i5FlZEFmX5xQHjtPD3ZvWzvapVSHgss7FrFuUb
QdePAFGePBfliUi4mSegYJMcIgL0Bs/q2i9pYCsUglezbn2jzsuY7GtGA58FZ93jO19Yj6uVBTiI
Aw4XTimfh2mD5L0c2mlcoGZvJeNdBI6e1bX78kE6bnb7NBlWGz8wAy8XtJiqdHx3et34nZAaDLvM
zzQy9bi0JqaBa4IHBiDBJz6x/aUwTkSgR7Ak/UmoMDD1LR1IEL04L7cZ72rCvfbfuJdhY0N2rmLI
QApWzGzLAu857eEzuLgUgi/Mbj7+zlod/uf/ZZO/CbQ0nyUoXVW6f8nNovUb/m5PyP6FYb8RZsEh
8s19H6jUoOfphyv7iTti3YDdlbnp0jKZEVnuGLeoq2TC/H+yEtwD76wTGB9GEW45xSobeVX8BVqN
0GX0qpQKseNvPokrs2Gifw+5LwXC56RxBV6tVvc90sFJ2VCW1srY+fVhOdKpiUYqA3QfNnn5YESA
v1XJMwrlTvOr54fdWR9Vm5sodwpUbNTafqLfgyNobI8GErZiXtHF5uwj7WSVR++ZmxT+3BexkKHe
V3A0jUC/5ZEfXfzBjeYiHqHSNmJKA8UuisVDQYvwM0rPvyTH+TMBQqccQ12rRv/LRjXS0svle5QK
hxgTAxMlopMDRnA7/ns8uuAzyGiRmQm6spoqjTt/V55idSkS0/Yb47N7Lxyt4C/6WehD6hRVCIW2
rup1S1LxJV2Rc5tex4dT+75ImBYp1xGMEy8R7s3i5tyFx3y3TESiVE3cnUhTT9/z7gP9NRc0HnQy
/9T3RYyekWO+JbPwQPLXU3xRiBlcMsUIZWb9FV+QmMED+Xk6wHrGiMlsjg4eIqNj1Eol/aLmRy3K
/OHyn3zcImip/Oj8uT1qDb1BnzPFRUgFfDIA0c4aBapOo4Lu4DLXii1EY7KrBQIqdkYaXoiRpSVY
rX0dcGu00fuKgpzDSBibevYe4bBlWte8f2Vt/xsswSLlAXcruzFGTKx/hc3tI8E9jTVZ/dSuTIKa
TimKiHUvh8lbzrBDuDqIdbp6bFrx0WB+cSyX9GJyT8B1Tdr7I1zmrAE8GmVRD6p2vtYt/M6FM9qf
gTA5Bi5saH1jvlMVtWR2DlpY0UApZRHMSDoxEdNYopEJ8p/1t1dFv/B5PnWkFRHRRuOGQlwMPj74
QgjoTQn1yxcLLRkbI1QE7Q1p5G3xBRQQFseI9jDglCS2RqG3/p6GSFaWp/3tjTTOk3qENGDOoT3/
6USGUNDMc1mRLkvfdKHyzKpaqG4T8zz8pkRD04tS5mBJUFMwGDHVW5OoleYbQSy5hC3KSfq6+XCA
Cf+RB4OlruTtzrX098gD5Epc1VSl8lAHA03GzZmEmCflb9T/x07f1gxhv3Ttgy2q5D6Td/fsnlZu
s8+baNr+pOxw9Qn9z6DVBOmiGx0J6BzV7UfTqV5dwWWIxViXiPy3sIn3vEJNJRC7kiOwzDrDmw/8
453YZytpFZnLKNhsQiSJ/1gEp/R5js/i7UtfHxxDgeQaX5v3AIBIsrhEZt7ws4CR/klcTex1NJko
nWr0zDCcDR5hecPNYaysKlJa6XtJ1DagokhUP9e8+t2ndNCmgidgEgZBACENw5aJ1XAf8nOliPN3
rpjf33m54rnxIoW1k/1RJu3xlkYs0w/XfjWkUkkZdP1vNPKzbpOquf27Am7vF4XB9BwjLXskJIrq
OTxm42cITXJgjicjjc28/3UGKNAZj5/akqES9Y0Vk+DFELkUl9hqj8D4zhng6FQCYIELMSdHFvpf
gupA/uTNXNBwFr8Gs2HfJkgEw7lXJVLwfmQN8Agc/J1dJK3/XtCdQZ9xnIiLL09Jm/lde+AL32Jb
bOkBjjRaSUenEszgus8O1qYAzvb4ghC5V3CVLqilkzg+Ps1R3acPWB3ser7+uH7i+Vt+vxKpub1f
CaNU7bKHqxeOxxyPkoouxK/31T0vCvpJnk6idQr1yu7l8t+DgiFDV+gqaaNyI0Hm4mAItOcZlKn9
/OdtgAfgubprPryokfBfuHe6EG7xku56qbxp0cXau8LljwJNiNzea0/irqNwNe3G5hskSgNfOkus
iy9rpWCISYN+hLIqg6+UcHiWiL3I9nECQh7xQtV0RmWSqlT9PPDaDoAjwycnBX2dpmijI3byW7IK
9RoznlmO4NebQX+G54dFevNuOt1aMLydZhdW97YY/G+zH8y3IoawwYNsUb4W1g05TEx779Mz3E0H
0/L8dI+Hk01zIYQQhwp7WveYr11B8wfezjVnaQFE08DTgXihEetaxG2imdj85K/q8JBLMHOBc8pO
ilGWOKD6JfLRaifvCLy+kngbLzK2kbSHwbNLxkhU5ui48Gc7gBudJRohmWqma5Pb0Cf10rjFGQn2
v+zU0n5Kl83IR3yJeoNyN7r5rWQmlHCHB2Ebc0G2aAyPVaMnmcdtm1Z0FOJoSw6qGJ9D4jLx1TLo
PuDLvFI9MVCEBUUawXa2hzY9NHsJClqoc3fM0PhuZMRnDqnMrqx6ZXr3pI4TNJPPq42GTWzRdZPR
NvBYlrf7q6PF/haAjTC8Kyz8Kuoaq7Xfqny5hjGhPMs7vkPAlW0ueW5O1gfm2epx+OShK3OLsVLg
iYyitkCZMTwVxj652X5hM2q53aZg/Auk4wyv0pLm64QAr9rgFn1Ur5MQfeqKFAyLLDIak2AwUnrC
Gw5NjJiLJKG3wJnSEjxjIpB9rFFzxn+6O+hs8IE1WbQA486iRhEDbs9w8zJgthrWUIxuG58vlCSm
uOvfa1siXYy6e/YAtnHeyG08DSOueqdGCUxRxozmwqJ04roNAJKFBBPek1abLXRKeW7JS3W4TY98
8xLZykC/OY56vEuFzH0/1NDZcmnwb+nopOLEWKfX56PmgzHFvWyI371cT3f8Th8a4FztbziyKyxh
4HPskfu72+FV4onmjb+YD79jPUvWwwJ18/NCEzbG4h5sM/R1MVFRIVmLj4lVlSGtbUWWC6xjV/na
aBH8SLFWinWOJh8yAXfX+sfUHYwZpHxMQkkWnnlQR9xZWg+LvZ5cGvQ+Uf5FI1ZRfAJWJ8QV6YnY
DSOljoJLRhTKyG2NeaAP+5Z9YSuoAOv0e2iKXQShxgKKzymVYTg53D1Zpgrv5yr/FDzejIRcjlO5
LWNsMHhDuie02mLk7/c2pFdqAxBHSl8hnWUTox6xdlhB27VwJkILYKZBGFB/IADdC3jO6vO94j/x
RlxU9UAuz+4TVieZkMUjgx0HLowuVp5EO83tF8oWIFZZ0o1Uys1ypzdsQRJ1GYI1FYVpB9ac0spW
eCupsS3dDUawpy6UeFGFs1FFuG50H/2PstTh+UnqpXaNxV+ba/2ltO7dC2iebw9H0LoEv6Quq5SV
ldeGVjzDrIc0jq7YUqhSybQiB3wpmdmPuEYRPNpYy4D11MXSnlDVPan7Y+SAGL0hbaydJizKcWuN
2PVrN8bKzCzV6QVw3tOnvoV9GXE9t9IP/kX5QIPR78xzHn23rzR9KHg7wqAt+PTn3nYZ16WOaMEK
o8ECtYag+D1pNT2XmF0OkCsmFWRZvPQzLUsL/k4qrsTTV+s+3jCOu1CLn4yhvlopVFsffVQKIa3p
1NDjcRC2kTrk9iuh03o/JZ1eI+wUmcw540C7clH7biLKXyl4DJqoyfjkh9gpwC9sz+ixE9BMxQUB
7e1rzrOkZ548MswndFAcRbKO9rPne1c+kHjObI02IJJ6xvZaaU2hK9miMrSpZz060PlqHnobMQpb
/AAFpMqkdidM5HC1LpXk5dvCR9048POz739umbd7SXiZoTxhyVH2G7slOcqMMgNgdQXsakq+xfEP
6gFjWLBP7GurHSoE1C0U1xCehHILGkuIt4oi1aJ2QN5aTS1CZDt46SxMbbpl2KEwuCyr6yXLK1sj
eXvMBxm8VHVrj4pdQV3zwzudfmIVIisXjXCF2BMlPNTFCBtZyivC1NQGI+Vhkx9AtSljMromAKgU
NCpTOGw+TPXsSggO//FbTHAQbskYS4zaMY7ueNHHDGMeOkG5EbO7o4hW8HCbi24sqagMSIZUB6tS
QpapmP2hsXXVmymRzW5njDBx5DCuNMwksuBGptwliRQhNDptVqUO0HYPOufQ6BvueDNU3qoaedON
1XOXz4F4BBIGpsP6TvfEXbtYC+FmMn6GJq/J6+cte6Yw4iBWpvdwBfGAIHYcXbuMBm87aBLRY4Y0
SSEVHI6Pi/ygS+GwhilFtOc5WIGelpxDWzZrfHEd5LV/pmCdZ+rhq0tB4q6YH7iAmEIOb7MARRVZ
Zq3rtQzkrvjE49TIKTZG9PMngqUIIKkIuvGKP3GbWxRBaH4rPbxKg1Pqa8kjRVW/YGz2AkJcghCv
xz2K/qEsCB9AjpiK21JzC/4v+C3JlBNsABL/3PgYbXbkhhd+UGM78qLCvcvvhluryC8uPqbaY5DC
p97pbVmccgkY80IPfLTGfMrC+EHPzekvI47J/82e9lMV5C+9YgqwAY6KP2aNZa8XIiiEc6zMfJ64
JW4RMOHU0vwp9Utigt9fNV5oYqpAG/c/d4xEJHAa1xcv6Ze8ePJGrAMYOEl1WgfMnNm5D+aPHdZT
vlmawtfqeynwQcT2enYizxYD8QwkfRTkUGP97hdf/Myy67ZS76q24Gl9tYdfK4057nRjjJ2BgXrn
H6dITfu7NRiCjBYPlSutVmacSYVbkrK2OzUGSKLptIjHQC1bKYeHy53ViO2RLJgXWsm3hXnOBy+M
gTiDWgVhB+3Fo7f+ReTBALlL8CktBuPRVd76jm4cfzMscyWLnOR6yNLvqg+A5SRYYeKoQXMbojIJ
E2z3h8Ksl9GpzIVEIyitLAjzLFNt5Gtf0WprgWrtjcXlcG+Wgreu0HoRJ3DubGg2HT2ZHGTbMf0h
/8zjYv/zSqTm1rySklpdKJP1ksYMQ3YXax5pQ635meqlZ5PJmPXANfWTRtGjad5Oy4bxgGwEd6vT
t7ztHUDHaSoul8ZdJPt3oJ52moerXUPW+DBr6jaVt2CoL4FVyx6goe0e2LEtni0LD7svtFNY8Ins
uRQvWlYav8Jmu4oDofnHi05f31Q11l6x9LojrS9Q67Ly4hjKsmZlj3r+P3iUJGflkAUJoCQZGpJK
0RmzEOpcYggx6HpLn696rQdNIin2jsam0yLzM9VE7RQ24PooWYZXKnSHQYsGn36LjMo+wUUhlWx7
PIDUAb7z+JA3solhXsLda3Z4k9/EVGotYLlXGaCILRhxcSB/S8Wy579d26D3RYVdWL9dn6O0gEtu
DekbPwdHarjnDiY84Jn9I2WAvoHInkiXaWnTptBnq3Mu9IViunVAaRRd2QRdYE5CqqvpO/S4ih8V
dNhhKQBUAYIr62U9A93COI0bkMkwhZYZ0EqwfqzvEZLo0/IxMo2VN/WYs8WIprqhixJN1i2guIzG
/2GQqd3aJRZ1HHhdPdzOEnqTUz5u72Irwq4T5/sLfPyHv17MaK8nnTI3o4rAzwWhtPVcLIEXZFd3
8SdgGyetsGNt8Y/WeSKdOU0cWbVf1NMhaECSPQqvMsa8MQkMYZoJ/gMLGtWB4jc53SLsXhEqiKZq
MbOunGuJsZh7cHd6adT2Vt5lP3ZMrhhFC2NBkdZe7xZ6Jy6eq41OUIA3olCn+Uy8c/HrhAbiLRfQ
Nk2MaSAGrPgFqw6mAFG9lxxJQM+Ia3s/3R4peOw+/pYTTDoNfyqjHkqup08RgaBM4yvLsQGJLrkr
3gXD4o0MO7q9scZHa9p8CAEJQoXOJd3/3daTi+31m5UOmq2d9wppFsUcB3XCtnpwSqnIWivq9/oy
cMgtzHXDng/gCQ3dfyr9vFFHnc1gi0MCxljwN/f2Dp6cSaag8c8wIEp98/eP7N1vGB1Lc5N2hJWB
qIujxhty3zc/ReVr1hpO9MvdSKUbrwpvNw9bRoeGxHxHCm7q8zmB3b2q/UX+DaJsoN0bY0/lHqsy
EwEOtCJltY85J9BCi3dZ5w8Yy/Se1HY+SUuCrTmVtaN8rmSJtjW1dyXpYTsb9wOr4fGNbUScA6+8
7I2dLcmQ0/5UZ3c5VLS+2ORJ5G+6flAz9D+E4KLEDhCaqWQyjMlHRg3urM/wFYeKPnluEO3K1clp
KoNvTK9fQUV2xzu6MYzG6IDA9PfB9A3C/BfUlbemsGAPP8JCCg5loQyBN1EsCpJDTP3P3dssmqIQ
zXk1i9gCCiWnPzU2MLTpreHnuxhpMky8zY4dRDoW7CSf9Fi1PBM8vLyu3zAZsIlKkqRlra0GOFW3
rWYWTi3wOmRjKtcvoGR9SLfYLDWqE6mnk+nKLpNMPvyO5nV8iItUh09PW2qvIbRBq8xuu+styEpR
21p30EKi/8ij7P8dF5F2aO7iEk8JaJVoMFViyuRPNfztuuQya7j5RSZvyXXvr8mE5pvKpr0/8eOW
nLzv7kkthXMwruw+edPamCuH0uqh0NpleKj43hRXe6UM019yxe2XkVM061/jEdijFS3H6rmfRFSE
OOiy+IysIBDH9dSKIYMNysRIu4vtl6fASlzM4pKjJM8NsxMjVaHylXC0FbZ4YkQZR26Vi2zZ/bP8
bhlsCU48dKB3epiWzARw3O+5j+3UsX5fA/6A+7bZiDJG6ukyzA2cW/FCaW++qhyVmFdIQuobPR1q
A+AkOn3a0Lm1+IloJx1SDjshbqoPltGEX9wMy7suGWExXCI05bMCeFZXk45SWsOsExJ6tOR7yfm6
TNydzvzLDBnSrtApoqdUM3z5ljiJSU/SaCGDaYsJL5OU43HrAbnbb5mpSuVAYc+yz5YiG4yJ+ixL
dfpmFcKajHSdkSN0qkyKItLTXg8SKpTyc3sAeQKzgmG3IaWQhWhLAXcLf38lS7tl9iGOLQ2xhXT7
8Z2jMWnlxEQlqv7ipAJOvabQ/xowpqPr4JEKIzDl2AIoUH6fv2EHk467YkkXvn65Wr4XDa9hZZ5x
76iVQlYoQsJf1iJz5BTzXwFV2l5NH63SHLtjOcwLUViYRGkhFysPZLP1lQOw8e6qwx37KyszkUOP
K+7r7I3aQmYuzFYtPTm4cjH/lguI/KmWnGftgTwS26JsKd/Q6A13x7gfvJSiuXplbWBXSQ804a4I
QHG2YyH//ZAUwrAaGcgAIh9ZdcmL62RnFOGnUO+2boGfJifFhpvTQRO403muQXrgrzsx3ZRFLTDN
6SL99ekVp8dEBXINabC6VmwUNIsoyeQu/hY8XFUAIqTgIjwNSqv+FXjzGao/LoVfgGWxq9vlMKRg
+I/Yuh1IxDQpDVcV0ITFj6hpFdEp4CWJkOtOjC9e8hA3AW6ayDTkCM2QxdO4NQXCjk/JITzPC2aG
EPY1wMIheu/6OPfW5eiJFXqSeBpdxtbJ8cxMNqBlPxvKxipMdAkI8wtS4n1EYWLLfjomFD2E0H9g
ycCvmt7dvawRTXW/3H3HbYt/oIiRGHMapWmapu/7fmcGNHL7KAjv78B/IsmIznlQDq9fAU/iX/rb
89+Xrf192KDeLYusV4jgl0kpmEARZlMec06aAxwSOskVVxcsFD2Z3U0Hf83rOIcpIt4T0AcDdL3P
kAYDGSVut+3W5IYppM/aFUKO65mAYfRAkK7zZzbaUiltOVKhwfS70TgUB9sxb+ZqlaN4gaCbekMM
ycEpdGrFgu+v5UMMfc7nxZcGxSZNAve2maqdGxzynviCEfLDThKuKwrVJUfctlA2B4bMbgvi7K0q
XRUApDOCQ5DCrjuibaLut7zEysj0UsrQ+7GDlEbpg/RxoQu//fJhIiTNMm7t99lBCMRxp6dq9p/Y
UE7n9Vsg9FVGYHmqongwyM7Ly7EJLbivz64nlw1WP6Vz6OlLVzKuHeS8lZqr3gya9Oj0/keCWv1y
o0umZs76rgo26RsnnDgvuxLl+B9L6yg5crvzD8y7OmuP56gWeUIsrXzfpvLud6RPyRNLXEv+QYsf
fKOHg0OvbPL0htIZ9lLy7PfusCZcOOsuHC65IfHr0kwAiRPqQYWqN9z7/EJGVzhkoLo6ftuqPVxA
A+F4GJF4tir4Usd9zI5JGOpf8wCrl7fUDr9mKeA6/KxCGf0oPOUQ+uhCFmVoTAjt12cAGYN4bQ3H
MUkgyJ3qLOKhWzNnpLwW75M7TKrW7JkwsC9t5Z0xAcLiJ16/6nvGcS7oavJzZoAmRPzfGoPUiqXO
Jgb0l0Wvhsj8nWp7Wy0BxiL/IJp3hG/7PepYWKA9MpwRW+j1IxCvthdrsdwt14N7y4KGR3x/jXjx
q5R/Gd4mDgQUFt/nNhfpEYt2/uVCxDPvcvyhUVEVehoQcoYgYHL49EXPkYKi/aBKeqsRcrW+OQcR
EEfsc1ss13h4vhKAl3jcw75aaUZSf0a8riaB54QeSKuRYQ4BZqejlbZQqAoMqyFuoJGhQEvlcMSt
pIScr86xwah2Pjy2K5dSAgsh84ohVXwGYqw9XjEhES5EIdeNSeR+PG2KKQ63545Jwyl8LHHeqEGN
hyCw5zHIKty22cdsfPgUhIZhTKjdpzVKSXpWVOcnCKsRMW9/aulFv7x+0TVHFTuo2pldOjySJEFG
v3N+ZKQXTpYoAgewrhllP8y6Ze4LxrRp6DoiYXEif/6ulKdm634fFhgOpwHbOvRRzyU7Y8MDyoxe
7LBTghupzjDByWks6v06FXyZ9obLNvxSkZKgWCbNm51NQJAXSdWEd0sDbVZ3okheFDui3Kn9YGPH
+RIoaq28+QHGtuldGfbRMfxXNHvqZx+0L+QzqX3ujWunVfnIqCINXwH5erO2H6+FcqS1J9n7P1gM
AGJ2TJIx2LqiZIP/OKHu15izx93aVOC0vA5mw3SVIZ8ZMbWqAVp6wt9aAtJKnFnkRmk2OWN7sSi0
fpFVHLX7FixZ7ApLH6f18d2JA5es5NP+Q4J5MU7yXahrgcd6KKTNQx/n3TK+vQ0RneHLpMUdFSYT
gIoTCSxMrEOEuQay1A42WQeoX7rw1eoNqBWXaSqZmzSzagryG0NWLWEb9e65CEE0H9j8IfBho6rj
0q6fSDtREVhlk5dBUqBf65A/kGjVd/aRVV6MVrV+VbV3SAyUt4ulkQyJVw+U295ZIVHkCY57DMmb
zu6VWNhEBBrSKtfaEwvzoHGojFwVC9TXtlxVF8rrOTGGY+aKtr/kFO2Luj8aE/MYALCE7SAj2D5w
RmJVQkPhQfbolJCVXGHYEeeT3kkASm8hJy9eZ+z16FMatqlcKXwXXJ6PNC/5xBUUFqmrHD22uCIs
+6JUwRJrTiH431zb0ThJX9ywbXv3DdprabIpTDGZqqQdgvNwpyGUF59vc4346CPr6pXSKjIOTRKJ
FpMqee35u2rJbzTyDCcKEPduN5PZiyUkLQ6N2A5TrnXIea7Bcsnsm42LamsdlsZWItqwJZ76Qy/k
QILDsq+oHJ/HENXVQioNAybPs3JaCRmFgHj45S71+ovyW0RuKUoxbi8t8KZM6MLacgtLH9J4ozek
XpMwocthW57QV7ze/cNuMDG6lj6eGMM+IdjzCFwHRzx/ug+xDto2fiPD0I+OrxGaDiWA8b65FI4m
oni6Iz2C2SD3mGHkBRyT9tjf6pBcx0vDGxjbO68HmTzktzbepljb+XvopTxJcL5rvJOQ6pZ8L7ik
NuIbaLv76orQJs9trlbwxXrtMP1cCjmZV7FMXCJVFkvyzasY20kJXtENHE3eY1yilzHcycJeWBmk
SHEEnogVssGin1RykQoeHjlk0iSfZiUoFTd7k6ZrG8p6whc+w/Vnd4yilxSjR1nRISuBy90ev6qx
SPihps/72STDPHHh9JHLb7g9i0h2wINQDCDwVXu8j6ArWUq8GfAUcrUBEkgGxQYounV/BEZpxjns
KGrmLSc9pPWkP7YjhqH0rMZcWYmxzDqFBN3HX+9oNzEtGUDLhrfjexeRWrfIr9Zb7b+eZVh4Mzo3
oA24gimJqoqCrluzgcFaAWZLTIJoZ8MZf8AJupEu00HJUXo+hAbZEYvnC1R9Az5dxl0V7PLQsufd
PvEdPOtfrC5yYojESIPkCdH2hBWAxRroU2Vrat6Y+L4Wy+fzSGvA5DNmdg9YRKfwoxY7jGQYXGwp
AohdW0N8hfMYKkRF5EPy7auiGVPKcv+h0zo3MoC2vfmx58f4je81czj4K31nK4nz2aorR1khKSUL
SuRvrHj4YIn8vlCWhHea4pLuqoi/sQDS9U/3qS0eRq2XxTmCcT9uPgajXP+pLS34Hnk9fqk8it5L
Wa/au+zPGjql/pEtldukzeHua6RoJNuaiWyS/L8qGG5SWfUd+gwvAt/II2erLvRWt5p7g76isbSY
72QcpeiEYm5N50VoJCNvb+Ay93O1TYf8FG8PgsVLqs2nuSGy89OM4DQu2iwKhZjIquaRvhRRUqBb
MbshCfs1uA/JL0zUKqNcFRah8sYkCwrFR4F1gKqiDdmh8xVsgrmLC6aliVsb4f5uLKeE3tH2jNY0
7arA0mGoOb3CrLVr2ymjXDwrQoFR3CxjiSQjQIf798ntbCOLjLDv9e34hCfKwUWjkUwe9X6heDmo
W2EIp2oVdLeSIGzdRHAYGbNAvXyP894XMNiy77UEDSx03D+9/h8uqK1Ii5iorm5OvuL0pPLzXsJV
5GNtG15IXktB+fnVXlLcQRU8nUX9WdnVccK9gD4RciYIf5WtzgRcvEy4WxjTH8AJG5WcdJRdjlhd
ggfQpi3KO5WlKmkWfhe59C17BoI16fpyxkmoMofXVAZHr4RhqGFm1WIH+XhuTNfXj1ZpMC2DPJLO
8xHyjUyY9gqd8by3tGE69WZj/AcTVkL8ctVFrMNbo0U8fAp6RbkmwYdjbb1cTxZyk1PKmZXnlSSk
VkOgbx2O1pNVUje/bUitPwjTjXpOD7Uk7eHt+8HGKV7spcCTzG4nkeNeOgAGCnFrqxzsIrvN/sTp
mur1x9C0B9/c/iQhmGqbCtWJh5DtmO8uzYv1g0ilXmvB4YQtFmb83BuYttlWTTpa2AJC/YqASKcJ
70ILTOhzK+m4jZck7VwhLxHKUCy5rvxcB/qJeJChA0HyhX3Hu/mxTwcvYiycpXRRP3imB3/WvQMI
KOvh0uDRj2qdWVtT5THUWYsU/JNv9zJcQ3GJvts0Ie/sIyUgcjXNUAda+q2OBGURLr334Klp/LDe
orfgPW206BAD4wFsFBdpvfoxhWJDNIlUqTv+8geNWqzFAIkQ+wrcQzWgcvbFXYxeuw47QmBKqiYJ
J5Vns+0F537Y2hVW3DnveUYDLR0uLNCaOEtKr2I7+zKHyyEvnKz5Lb5GwE/cutPmoBD4tLWPIodl
dTmU67h1lGSy0ZFB4v6v0AVJmoIDyRyxK3vF3XfFbcgspOl37eUyCcjaKf1J5+MH1BMJX9sj7/r8
lbiiQM1TKehZtgMlw6vb9/28+DIqyuMt2glrgcgVSZ+9g9Ke7S3dZEt9g+M+Nz51uIY9ScyE3k8G
FcXuEsaUT5UOl9qPG4spQRf09DLxBikcd/b2aeOHJ2E/7DQZJO3t3g+iNoRwnFc/gMj4VFEzEZqV
PWU0MWh1+sU61fuKCSF9UjjPfVgLQR7SEg1IC37z2WRAmzmrmE5sdFi/vKs7iapNCtQ8nGu2iFx6
I9IJfCSreKJoThPnDHtDxz6eEbqKjG/N/U/KB3ucTapZCj47fwamDj1b+G7O73iW8YvSSIOoQu1L
9YB9KbkQla+1FqVkXwZxP9GABvJ4oEgbUlrS/h8vFLUVSY/L3Fkl7zbI6/Qn1WlXIOoOPziwuoR0
MGX0JLJcqlxYXIzZBSunNWyGfY8/3ah01PkIu5xpch5/ZKJVWTFhmPNCJuFYZznovDgpU7tKbFqL
KfD7D1ifiPmq3ABPV3waHrGT0/IRWhizdZbCQ0dhf9zOS8y86Psl8pW5kteXPmQ27z6loAc/cpbK
ONMjmfz2tNue+DNfhGWDxj/mA7lsDrt37vFT9zwz1aU0VEC2OFcbkJRZOrSBCZGYpTJSV3kXOw0X
kZmQGmEYGqSSoDFbEA6XS42lPv7H6CUFMuK4ZQ3j5QDKHJ+voom0OAdTKFumNYagFwYylfHzeHFu
9QptCQbzweWnv9yFwjAktb729/1MbG683KgSeYdkclATPUehGioE4fCFCunjVx/LxkWLAu3saHor
1OylUERec2wSH09PRgdc0nC8ZnPQtM1h/XTdqUM/mbc7rznorsdmNmyVNjRQ5LyRZiFZ3i/dojm0
uKEJ2n1AFji5TOER89c4gehIrkHgjyVUHmIBo6p8PPR6S+xywZiA8o329pHpeSsBckJ53ck8Wyvq
VjzWARykMtmmrk50y+CGrDepwufCOfLLg/qo4REqEV1R9HiTM2Tgpj4HUvGEs0K/VSxCIP+JmiIz
XpYlXFNSIJbhX3hmnEhRDNpNEMIOdoNLyTGjGzs9Fan3fc0flaggBwVwceoVPDNb14WqIol+o3IK
YeCxqxg2EYMXi20IpZEjxRV9ABPDRhsGd1kedDglpT+xNI537BHafg0v3+k2lbTPps4UjM4ojjFo
BcK5mwkUzvlxdJnbzRPXrwJRNqNe5NQVkvhpVHv8QkaBApjxwfb4ZUwnyeq5OZpEAYOPeRravNA1
qwuAQ4t6MhGWvi/mP82OMF/UDEdFq9Gr6oy7tqS1KctvvFibyKBV6JGJuIG9onV+zm56fua9jhfB
54D+V2RH6gCtkcg9uMS3xgYIxv8H9osr7sCdtLFsSz6ln3x40eamzx1H91FJfD5O9AgJdkCMTB4l
VFHtCYCok0SlEvYOru0k4Ts6D21iUamIx0KJcFKayCRrM4YWJDlN8TGVOsgzGVWnpy8J/VZ7OPPb
ZM6BJmnvoJGL3Cl0LC/7fyYCLy5ospr3IjZJwEz2JVOcuQMG+UxqVoy6d5PFGhMztXhVFrdTVPps
sZC6P1g9fnqB+tidLrGomrZcv5dVDaG3v6Ds+jMRTGgGQ6YZRcdKhDz5mPWwgbV0D5xQnk1JtrGs
08KlZwPP4xGWMcvMBV8xnh1kDOLEc9nmsLhZPCgUa2uHD+ODbd2rHId9fkKaa8u7IOkSM5YC685N
0VM/s2CumInxW4vOWUyGjz8eTEzGU4cDA3Q+VkNlLvMzNTcnoFdOTHIoNIqZJj2TCsw81/8nLLRo
9GQtNNJenBNxymXzU1dRWWg4e159MvMcKTC4d0ll34J1+XtGcT24qY7d5/pDLTxwlpcLl5yInBkn
5klY8DbXzLmgcL/NooL36jZ9hvMwu3Zv0tYLm0VAiuvR5zBXZAzupiVbQTmzhhky2Hh1bJuL/5a/
TxfYbceOBCCPSRJfSenemsIUmn2o2sIrUf54cVSbvPQrhbXeI7WVUVb1DnUkC2cqRcbP7N2grpLZ
uxfpFJrx28SVc7X7x9kgmcvJE7WFZhZa9IBQwnci2HVMVfIEb7klkhg6D3jYeOVvgMqqAXUdpF39
jAZDx0WEYympVoQyjlA0gfF3L6GiXqk+e+UJ9KsB9a+pUnOm/a4l190R/v34wyKfGnq7KytUwQwL
tWzY/+uYRBRuKOmj94LXPepRlw37UyMy5zgb0Ik1KN4TdphNj7Ohd6ulpvc3oesPRyJZl5IZeYtR
pePtcd9VlXzLzR7NeMQVAB4f80iFYOopWuzgkxALngRnD7A+U7j0j4PWefwqAfpd+KburDl/Zevw
kJxrkUu/lhUcP60lUJK8rLVn2YQxmJ2q2MbecSv/Ho+vJs0mViwq7nUcpn3YPJ0HIv0V5hnWq1wW
7dox06dKr21Kj5rUrwbUSoPjrll7IM6iDE55vT8JqTEOs6O4xDswWc3ZOXmHXfzx97CUMw6uWi8B
S1LvzIw5EbYfeHl3QkhMNjDwewJvfen4xm5h6DvITV8JI9zL30ep9kjB2jCui3cjuF4gaFr/GJux
MU5V4ukwfEvyLpVaoALMVyOKLwdgmo1qB03bi5ExOMos50h+OwbJ/qySGtMe2LC6S10tgzMQ7RY2
Q5q85cxkk977mEe9OdgVLFRq2U6D6lwLmmcQ2YfpUcermGifx2W0Z/N0m0Q6slz3VB08/6lp8vTr
Ew1BJyzVoCwHs6uQ7qUkoKEZWVrsD3cfKH3LWoFen4B4extgXXlljNFY7nZOLTspNcA+87ZtSDkM
tA3i94BLvaf7ge4sJiO25IGlyzP5+AoVUrqtvO+T3jlCGvTwP/XAmCL8VLMj/wXmsIfAdOXOTCYf
EhHP5EFephHeTgg7UYCybJyzI5Ggx7ZmnCE6bLi5g1abM0O2+9d5865K8lipA0nzsie2GOEsPnnY
R9SIEy36j6ILBamkgwi+qYJ13npSL2EP+ihSWCwjjq0ydZEZqtTbEUhzskM3yb+FfnPPIGEtd47y
Ya7uSg2TmNjp8hEZhBOAuSzP+LtnO0NcAEW4Ca4rMUzF6Y2QKFDrljr1KOeBxpvso0eZcn2rplhb
Ypz4Pee9p1lthN1cO8MF1c9Zt5SonwTP1Zy8Zp1xgnnjckZSIcoqDB1nTRmmW+f02L+SCqkigA0h
qWdrJxa1DjmnXbJ17fOzuqUNSknFb8KXzHU2Q0oeWH+eev9NxCjY2ZAH4++U5uWf7Rw+LgROzOg4
4VWnIc9jCoNj0YOOpY55/qmM7hCoFujgbXk3YW8hVmF5v/bIZXxjgOl3o9hqbnF8s6lGfshulj1p
xCzZ10rLa5vN+k1Gz9FySq0L/vftrdjPYzwHADyi9G87A0hbvIluW2MyMO2Ld1dGj95CmkcTORlS
VJXLcR7KFFMCbj8uWOBW9npnzZ5KNdp/IeJeZEvB5pG6flIv5ijc+OCodVjPwGwHi+QFQp3ahRVT
Mt+jyNDeAW9qhFM9sHHT3UiVoe6KiOIPC1zRx2PK0WwT2DvG1K0O10p0qpURErDSJabGMvrTuNhD
be8ca2dCcFOofDGqLABXKRpDHYneu5QW2JuxrOHTJqA5iwdMFauorN9BEksnCcqNYc2CQWagAAiX
kViXMeMqV5bzYmA+kZ4uu3SmneKUbZ4OdKL2BZyeOtQK07/gGQq33txnANO/SgnVEm3bgdAWqLlK
pr+vhL4aIZhgiNoUHoJ5stCCDV8feOr7OKjaa3OtBhJovoA5XD6E9lCCFXmWmLVtP2gN4Ri0bVSL
idq0jPFxTU0AqzD71JE2fHzwPd5e5GRrY2d3E/bIbVH7JcuYG9et3iCCi5v5NSskTSF+wOb7OnxR
u7vU9ty7oERue+Da6iBY+T9BMVoA19+XZtj1ZD29H03QMbIMJEJEon9VoBOR4NkRgOg9N9vogwfN
DldZRwoNjkb3SlhdxZJWKYFj1XvJ0FYZRIzX2cJNfUmwURJWPjwe3AgYEnhkFwA49AO/m9ZkZuRW
W0Ar+RDP/MaBkiV9GIqXHjUHInqo8DLncTwsAy9kJNWSDtw7zSLCSPIr1cKD/xnTxjOihXf+xiPd
l4UZ0muo+8o06KqFQkI+G30dqjJyaX9srdNiv4qI4feKIP7oFgnWeep3QmtclR9KUAzyXRlPVpyp
xR7J1byMgOFikIGlPpsx+29KC/mKrTRbvUfExYA+vPURO1xQKTx31D2S2NKFZsFA9/TUvJcqr+rW
pBde9psC6HurRhs57kDQa+yL1YD8mXmUmS5quNyE6YquNWs8QezXCCoiE408igcKC12YLDxnUddN
qMjmuX7rHIup3pMpD0Fyr5AntLjzMtmlr4nXwHH6zOlC38p/3xW8kktwCN0tIKjm5dQK/rveBupI
/HFB1ce1aL5SrIcaD5v/OWymkC66VVCiCB7yiuAw9VecZf5R9tftBVCBgd6Ub3eGhmT6n1RWzYGL
vQVnyDcaaCyU4uJERIsIsz7Y5p4XK/SGQ8pDnXEsRL9Fdp0cmwgX8U+aeFVwRytrE2sGbKnUDeRS
Zo1aWL9OggJtKexNvh9Dz96xDIW3ihEbn+KNTRcPLEJaBQ9K+XFczSirtJsHVRI73WrKXSDJ9JwO
6hmfUKfhzRtkRDLKj3WrEnPU8PWWHBhHvd7XC1n7rbEAB50hlzmNmZ5aDskA6EXf1KjASBYxREAx
M3U9897SkA7Q8KFL0VKqrveNSZ80eFg40S7KMPsMjSkfNyAih4GIcCCm4MVB0/Sid4ZSgnbQuA/V
rk8PxgRbAb7ClSlLFsd8k3uC792ttoR/PhVAncNbVJGLCr09A9v9QSYlACf0nspmyzIy5OUYoQsK
phk5ffswN0ucOGElvqEx4Eq8RjgwePgs/+NtdGTAPVx0kvPr1YrZ9R/NgrQpkBohLrpz68l/NfED
kos60qAbY8iofhFpL98mlLDlkl4ETbLRAwXKqZg37LzflN9bVuBIv1C00BXdv2uZoXdxcDkYW8TX
TfrOA2bBV1wFnQaRnGsfjWqyLoqZdd70qOGGT9ijJ2Q2wySu+nRx3RrQSHAHlQW5fqUNCAIBQkvu
Lw2BGYA/k2Mo6kVR1QXxqHPvcWAWEkr+TxkJrkTRwAvqdLNXGPXOUucdsg0k1EXMFgFUJcCd57MV
VpGY/M35VsfV0e9IuuVolkQ5YZjh6+c0F3O7EPhHm72NH08hBV/aAyaSTtSvwX7q4kRtmw4+6NWB
9ZaTSTwcwCSGW6rTTBE/0PW5Vf3WkKexqJkkNq+aEZnHnYV5zhZHjLt0+QEbcmzxEwX3oG5qJzwv
b+a52s/9lZNgJ52Bi1bEP4F21DqRgSI0/t2mAXEFxkJlJt5a8R1qVsLiFutW+sbRWXZP0EyRXYvn
gJdpyYK9IBuaPz/leM/L/9Uu1pbgZQaT0LQkTolvkrhGmVM6x9wUnSTt31d+bkN5SLJf+u3GUjry
ZcxDoWTiFY3ZzNW2lkXgTUuO4qIn1ev7EW6GFO8Cz/nm4JDYxnFTKyhXSc2quhnywdukPXXI53pB
FgLzKM/ejJOOR/dPY7EKjn1Bb79VCjHvS2NwYLVGySb7D/WGwk+loHpGpbrf2PY3TxslZvgsJZHZ
dzRmoeLXBLmS+tmLg1igw7nT9J1AuOYa7dhOOaizJLRMPT3HMKlZJQgTty39c9ueDTU6c9/mgCwN
+JpfTNrMhonp0AgtNmzw5h4BrnTmSAI12zJB9eHg/Oa7j4lnIeyXgT05Bqxm0HNrmvp9lOQYNzI5
SDS2dJjgxO1/mN8KreKzPK/mij7NsflWR9Wjf2MQg6arohn78ZwzUdSzRouSY6+fpQTqiJdEajct
ZXkJAkhvSKWAhV8x2Nb7WAgtuKOjGqOCA33q3CN4tsbc7j2mUhWsafHiHetJnYctBzenvYI7j/Rp
so9amG93YCtqt3Ea7ZOc5D6F1TZ36cbItVM6S2awcXuGUByHbKXtbrraLDBMLQxgjrQUgd9oeYj9
3HNuTJQtj8kAWw//zo/e+Ukyq7AnqU2Y/VcdhMqvtuMa1m3qpLnxUtortWZtn7zsmN4/KrcA+49K
zLwkdI8TByHi5xpGx2Fx0ONXBUg1JvQjGpLnzjml8zDuzF/u1COYdEIYwwX6WGl21IMLXHFjW4pJ
O8PeKEmmL05v3JUeFpMrFMSfYPEVe5Ahex4EbCXdiqsTgLCVchSswbbYsytOG7G7bu/IL5GZAqf/
HcdJPO/KQ/k/Ck6BGiuav0q61sOIHcBstpnJLpSe+yFttRckyuWfLBV6o6q15cGJW4WJfRbRsCOA
KQbDDqhKQihvAVsC3B/+6FBXq5dnxDLWAdjmptOPPVKSswPH5Jx1ZRpTX4A2gp1BgllRQkzVfr2c
rxbPdj31WoaHli2H1eUU9GOjioff2QeaU1ELZZRDPCKnbNbxMvRJ2o4jwrONtZnhO6UFpaVwKqFm
c577zI5gqy5rPzi4Q+V/c7WPocQr6BF+RtG4Ky9wYiJeVQKSm+FSO59nSlKj1hvvNBRAzCX7zdkQ
d1fRKsWSAmDeGOGtXz28muHpSyw8gKEWbHvO8Su+UYNFRzcJuR7/M0HNZYJjxbAbXBBVqsiCIMdA
AneSKQwFEpUy6r5dFstW1Qc7qQIIX9XpPA0CYapJqhjCzEFxLuv0clN8Z5uPRCzwukUJrC9r16m/
oCpViEYP+xlCEynIuYwUVRf+4NNW5b2lzES/zrL63Uq/TjjgOzUCjrajULwW/64CdQWcGB1a39Oc
NgXPdKDiBHaAadd/6r1d5/74A4m3hs+Xvh0v1FuGErD26Ue7AzQ2cRNys2SOgHtBi5KNsBMF7S4G
0HXqhLqx1Y1kFMGfTTVwRoP9T+fhkyrNEcCDv6IEx+9Ln7AH0RrDIauotHSj/dQ2EEwVreNXgrBY
76+LM4sgb/6r+qAWl3RcUHGVdf+KothVpRSVm7yeeLM8s1LBC5M3BjilA6DZ20U45S8N8gPNm71C
KpteDAwL2v9K4naktt+glN9SEKMzVwG3jzjNTbrcpEXtCzst0ytFEAMmYqJtIhMfG6tXSK41YvIi
Hdn1Y0GE+qn+I1tOrwnGPTOhFQyVY0WDUg19SnJ0eRCFFmzPQWBNb9WJmu+7Ta0JoALOP3KZbt+y
d4s2g9LYmoBblU9ZcIArycubGj9apwHnSY0HVJ+d0ZzDc/cG7EaKI1OCVIbsvTmhSNDzoKP+uJDL
vewmvfoIx2Ez63xPl+nCNQY2p9Qj977GvlVSr4EM0al0rozuyTnqyvV9IEE9ah8N641JDJpu1UmU
zMPzEXAx5v/jJQZgH0Kx2QhHV5acAYu/zrrmzWeBXWaktxW+X6RH7jssFt4NJW13QhJr7QXaRmx8
2Y9aSvtAKrEMZYqyfXL40hlt4jfwn343YdGS/fmg6tcdoy/Bq04vpKZSef7Zek/BTHv4ArDj9U3s
1/2qR8ePv4G1vRrZjipcXSkhZy0t9HRpFuOUHvgEODWqrVhcHTIZMnm/ECAhgbNQvWq/goFgI/uD
XgQzKL/9o/vi1Te7n8p1xXBGnx6SG1e+tMhXXsUlJrkK1M7OjVGGZqazHmIkAGvmA1lxg2eyBG8H
pP0Zgp+uwuf2JZC7qolvH8qDsXezfyvbasGshU9WKTgV+LY7AAGrrq9fVCSBVJdDWZ42ougALIl6
sYpjFKgwOUWaREvmiY1cfECFNYaHrGcXqGkmIjqb5RDYHEo6+mRDVtEiXIOHMfeQ7JEA8FlMMOkK
5J+jsNirm9ld9YyBqA97XVMAobvGTCHOnBGLMFFPAPp69bqZoRPGYccR5gLRNXWE75u5Q6BADqYO
U0IKN0mIyRUC62CiS9bC15idT0RuutMASihQ9wJmM8r6jqP96vpD7o4lNNjwVIzRuebpAJGAW4x+
AwyEWwfLONicomb+A7fPepCqQXuxD+jun3y7Fkg1UqBjQPrL7BW5SjmTd1SVbSJbVskHo43I6aHv
/A+6t3x6dWUDwXyDSnwDUW50X/vmsKgpjynnECteQkKNDPBZqIsgN456SvjG+PA+arjj0ST18jde
Yw//nwVwyy4sfwxffadiYRUgfx3lsv7KW7I631eTFYcqY9PtZCFVaAfuCMeZRg3quGcxrOo5a4Gb
gPfLwFlaUWfH1PF5X3rhXbDSbsUgoNSMjxGUouk3aTcdSHEn6paf5W1sRCZCFOVZPV+37jFzwAV2
e58NoyilTlKqE7iabdTMPDfCguJV3KXXike7iSJmo1JOBeuHIV8Rbj637P5h1xD93WP+68coFo0U
owFl9CIHKZ8/qrQ+J33NCpfljAs50Q/D4UbA3KJZ5e7OFvr5Oy+gM+TNfpUH3LDOT81MvDvqX8j1
eT0WpdYoNxda+CBd+SKPbJMQ2PxMzyUzG1+15nFwJG0DusO/hoA5tW1sTQ/86u+fCrUBgTljuUH4
Uu90cJaScGtDS7LznAKZ43GxL0hZlvQeNRbm163/in5ZC2z8YXl0/lSn6zdGLTndq5abrq4zG8CP
4Ysy1X3MXuA4G9uz0uoE63iaaj1zQlGs7WGXRc6Lw9GtNi2myxLS/ayXbzXx8Q5to30BxU72ycxZ
/ZksUsLYMc5WwOuZucRS0dCpxGTgeF+Eu2VWLaDJOl3J33npdcmkkiQRdPEL8R2Y5iv33uYz1xvl
F+C7fR1EzjB65vtypC2RKwAyg4ICjBOUdSjxi/OF0VQbJJajgXlrnacG6dO6xhkrdnvvnVUQGmZe
7nZidJNYIhJiyBTx4B0EkDyN98f4nTxEu564qsRjTBid4wR+ZvOK8mhJzD0a0VhbZv/zF1gpFQDA
kbnB5aAw9sxM/EOhdUvdQSdnBiufw2dHS/+qkrL9yrpGE+2x3RJtDZLsKL5uMeJ1oBiFp7vOT8Ug
XOyihft/f7vrl31kySx0La6vzWK5lUzzyCEY5O0V1vfyw5cnoVgYJrJoMQs9pKyCOCeV95zI+eSe
qeAIWm9LEsw4HCPEb4TJzgoJrCaw78bAtEcsAl46y9pMLm518IL/EDQ7kByMptkJ0WUDxQg8jlWV
Z5bZFF/1vVROBbibNAkh1CpWDXouNBJFg+U34rVSiFYLBk3yVKZ+ETFpnMY4TzmcGqgg/DiMXZ+A
w1vKinR9IR0GlIEdBKvX4EGeqYT7/zbNgL7Us4IRuhUqT4OeUiktssSEPNybcYywt69svsvVwUx9
yo5HoVYE7tG4bsuIS0z0Q4t6LvGxBsECcrxougHfi87XjGsdrZP/l2T+e0yHJ3LoMtoMqJG/xMcw
TyqC5/8qwviX/c97W7F1m/DWMiWESo5yMDTsOfvPIWDY9yy3iQ7HQKwH/dGtAKt5PU+jpak0fKNC
vj6pNMpBDvPVcSpItRDK1FHe6Tmsf+jAvldvjDTF2tPauMJ5PVGebGIwAVJJRKSlxZkybA/2VqGW
rY2aZldlvOJ4+pDd23DVxcPJM36dYmwAUZg+k3ttXLaMNfOZNLZbRUFMmMem/Ew6oIWSaSwY27f/
h8Xb2AWGeOKlBaYBOsggMa+cMxC5Hl9kZrRPW2tRrwnsQxSeRTxLfaLGzMONLrUk7rJ2HkYfss3X
saJgLXBt1vo65J13lWtgofphcnI61OsRIgZ8C2PJku+lmvJob1E0steY/Qcz+uVTlCfNeCRjyC1e
uuj+ownfXKA1CepgZHCDfeUuicU+rfjJDI9AOvQgvMMnFoOJ66lGNswSuqlvdUEts1aCIk3Rp8kG
VRMTiYtqesI2VArL0CjUpFhowrQNR9Jl62pF1InnzsfNZTM7UkQpjQDd95T7BFvgurENEqs8v5lF
jm+uPZ9u/uAh0g/4qUlNdAGqHdI53uwrlaS6lDGV4SrgNzNZNYN5zrzAkpsrb+xvqnsTZg77UobA
k4rk5DX4q690M8Lr/FrM8vxyNqDdSwu7Cynv9Xv+hQSbYn9/C0b7WBdWiKnrjXQVIqRmD2IW1dYN
3dkFd6+50x05ZDbjTRYdaSi5fo0X80QsEG0oRvxwI77ZnJJ+3cmrTAGaNnake2QnSlIY8xoBAC8p
lKA/k2k1ToX6qEutvjHWca00AGl1nJW8rkRyZHMB8G1ZfjDYdqY4cGobO1pzxSUJtGnBBFXtG+31
gPMv0rvIss2Dgu5R0X5WF3l8xvOWim5LnRxA6oMQT84NqFytDVSxj6/YJrdpmD6+/rwkjhKrUvY6
4bFpau3XOvSTNm3dPE0xqhhsl3n9zuiP/y/1ntLvrUEPiPV62XS3I+PUrRk3g1pLodcvK7CPMeBA
CK1KS0EDOtHcApB2j0Q0Kc0oH7868o5pDO7//xQnuEHmlHcNje/Ea1jtCLGTyLC6Fek7ovRW7G1P
WZ6h6itJ+0XIwLNqMN41nspNgupi+s/d1fYEQrTDzKwvF53l9tZa7OVsFZDsOwHg5sWOmZmxzefm
iWDi5zNFp7yO59vSdMH+C1kXE/zWftADU79l+vGB2sVcbswzYmoTPW/wbCBAMBEMNyLCHmA54ihq
lBtf8EBUmtb5lJ1RvpfazVwULz35TVioXwT6ovb9vSTgv5I9FETiIRJevHn1m1IMNrrJj2R1z2tF
uA9lWaRsLQUOykxBnPAWounK4qA1+lESbHm2tr5C755PqX2NAhMCfA+/GqG0W/gbckn0pwg31hAt
FMuKSr8MmlkTt6bXz94EI3q+Ot+qR1ORxRfhaL0RHfOEQldhwYAYIJ5mMNMWzy9NFrmJUd5jkrAC
D70UQ9Ur0eEf4XLXoubA7Be0VQnuauYGuMXlgnCFLdVc6DPsX7Lr4udc1wtysTtJ7249+5r2lqZu
zQKZybRfhMQtd/CUppDbTh18n0UY8xVG8bNO69NjMrA1QId5l6vlJJtY2zNYeK/BwJeopkA9V5eM
7tbsY6jKncWsxKYZ3V1JC15NjEAOQkA35OG84kCe6T4PZLlGvwMqy+yEw8welscjrTM9Wq4jzReR
Yp7SFp+KTrh3f91RZY4qXCgeEgROhsiCV2RP2m+5ZzYHrTnP+SPdWEKn3xQVME1wpSU4+HFS0khb
iN/4VSQcX257di0Sa7oI4ZbSc5kzgna4kN1mlCnbjKP5SCBVXZilNzbK+ZvPgaaMCAutqg94IzqX
pWU6DsDnjvz77LSNVR0xl/oHwXUqgEz/ClGlcQIeIWdYOyqAhIkR81jR+mQcCnKG0LBM7QO7ucj/
E+y+t4h4yodF2iWED3klrTTOlIxE2sVrMctakBdPsHXZPB88DdfUBPE+ohOtd6HyUxwhBsizU+MA
ngrfZb3AqzMLO8h8zlAr4AZysIeoIuMtN6ojMD8oiLDj+xKjm7pBlVaoZZ8vITnpoU4qkCxnQYGm
Xo04t9MFuj6MYsHAitjKs28n4rakeEEVIteJP1gk3WLaLNjNRnRK0YhEWowVpiUHDyDL1kYAMB5H
qOubUwc6XBUGqRzu4b8VNI4JyL+BVDkFdHfiTIKg/ElIGfXnPOp2XK9k66QCLOru15O3qW6Ys+85
EEZVe9C4aDZNxPz8nb5nEwAB990qSawbvsMTGFZMHqo83RUJMeByOPUJRdPHy2qEkCy0207y1z8c
EQb/Ihm5KU1rBAIU1qJaOaJHYW9/V2/2yYqwm9vkVPtSl1GhwesAPwE2qaNeEC5yGM0dqQQI5HMA
i8jcmf4bkGapjhdTtDFVzggdv70vBcuStoKSWmV5h2bQ5iMgVKKu14tlaGCvsvmiu+ryPWZYIf7P
KF6ybYOH5S0ZJdl8X00KJvMlUuFk4i/BWKhC2SE1mx8Mk4dI5gcQds1XCw/Eh9v6Pj6U0MghfqAk
IXbaLlKmILyvcadCfXmU7PwnO6CEQMaFt1d7bZSXYd/8URP57pl4RZunMAU5uUcVoXta1jvM7RWO
Up4N8HKN8nSM8IC1S2i2oPiFcMRlOkabM24Or5v/EzU9cfUWvYbGM/RWcaXP2y56op9KZY3IFrxw
ZnEBEBp57ASoIlBKMUuQQFCNb+o0cmsudAPOY657D0HOxsp1pzgM9SxOhts26OWQN+yWRrtZuZhR
nu0HKz9qDhOeL3Rme6BlPqQYSPiNu6lnh0M5hKBj4zT5RcK7EgJR6Dd+jO3W2rkD0nBpuD4AFOKb
XAw7uK07u5eVoJl/lUGRRj64lqnbad1bWUMosZG4ihsrp0U63hi+8mhJKTl4zpFM5+oJ1kQTG2pj
x3elCTnOqPMXsCucSbg0q4ezucMIh6GAtLH8HuJPCOnCdg42gh6Hk6oQ74+SwPd0roiHfu4ZqENT
c8wMTf/d4ewxYwue2uxUbhYRhOetbE32Vh/zjJ5KSFSDP1J0UAi9g8nmpZwIlIs68mzm6PDP2cyD
dUKzTeW5hnNRnVnNP6UViJERju4Rvqq3Ndsu1lhbsgHC2d0pQb04Ma5heIJ+dxvW7hkJJD1bIHzO
dMKK8DUj/qacOv+Drwjy5PKZ/tcFon4D0glKuaRnCAat6PXrUqy1teCD0PRPFXHIUa94k7vRZKBn
TxYPD3FWGTQOPAzqnQpIaPXDlnJqRQNHYCqPuJsEVuky9ZzW2Tu0ICiawNTb4J4R6SiHf8A1vvf3
6WEcxgTyg5qEJAGPjtlPxOFobSItl5HbfluDERn//q6OBMzSMjWeSCQmxvynvEaHcAKbvszOMEQu
2FY/H8xJ8UAZFMQwMSRYw58hliWnmzddGNhaA3nqYhureuxQt8L38KK+A8gbMQ86L48sTXdlpYad
UXMr9tsScwmdmTpOD9Mo6Tqe/oQ/exAt8F30FvhemQIX5Y5q3LIg6VKVd/xJgMZhL8Q/xat40WbH
TZUmY2UlCuz85fI94aa96uL47XeIS6L6iL1MfilcfJVZiPKAfkpGcTM+JdR+R1lYvjmbULo6NPcL
Q46nAU0crK5sLAThvgF2rlRlXQNV8FIzGx5gyUFFz833o6qieQlAhQtOQNI3p0pxhrL+AnNTa8h/
jYJIa0EA726rMLTR8UH0L+5OKC/QvUBl4G7qDvhEY5AX0HyH0JRnTJecydD4pjRsEamnleneN6Kj
0ONnZ0B67eL0f56Z5iqVk/5iLo4abbbxB+IE0jXGBwgOD2/qktlnxomh4A9ObC/HXQSfl9OasYZm
HPWmyoMf7rZevedIS26oxSE44IAUGn5wibeSFoRxaYg5E5PZCak1IiAJhB+eQFBCg/sizpRI3nyw
brwJWOB7kP6NtOObH7/DmenlzGQiBdx2jpuxU/r8RWVKbia37DVSL5tk+tg4zG5A9BpIFXOLnGdh
DMQxQkUD/OTEjqnJlaxrIUbjHjoQoGnUXS6bolqIlHNq4LjA3IQWnt3ajiKT3Y5wSkRANUa/zj79
GgyJBxrpp8gladI9C8MxU30DjLLOpV2UYAerllp8t36wcasxYT0Dh904ScrbyKHzQRGCWkLaR1dZ
MRCSRNy4xcYW6oqe8feQrbWhx9aJvCmffutum2GLvklUwWwfNZzYvBF2RjQF4qZAsRw/nkBkrS8/
o2Nl4077gFy6ZDdXkc/oNuXojwXdTRPwgPv2TUfbzk6IdQOS6Vg5Tl0XirrnC8H7WlGekM2WZ2gR
/d89Iez9UTV4PYiK+I1Cqb6gG9oGhXzq79BBv1HXPtqPgx86+WfduZRtscu0vcgcj5Ar4pwOPeHS
3ZRhVyFd2FsZtwzENK6xJxfgp5HbBLZXdo1k5vwNxmU8yafP5bXWD73o5TnDr838L1rD8RjY5E9R
covJw3bXONIaYEH9XUEBI5AXjAGAGrTeSiHDjIhvEy17bDsXDN316IlWZ6j1XYVX6DSt8oxM5jdk
JtC7IzesVrRlGwb5JIVR6AgaEqakylOe/lUMB1JBJElh6J3E7xO9xnPAAC4+a8LJ0aFZbHd/cluG
sUnLAssjajk8911oVMbwGVmPgLGi05rmIY0XCqrdZhRpFUL9YBZocsOxcquMu6K0C8jYN0i40VPU
GXi9wh+IxgFuEBujPSblzisYDDixzf0wbValcp9lnsjC4O94F+3OhtinvdLFAiAlBMVx2SaWmjO+
1EEc990LFqnsg/U1OfeWvkYg5vCpNJ7lCRmzltVGItwVlONOP1xn2CRah4HTZ0hv8/K+PID8DbLu
h/FzBLxxEv0tkdSJQU4LTMzkZvBWuL/mO/13Ou4HD8aQLg+TcanPWNfGH/XJc8+/Jtf+0nTEZaXN
4Z4367driGNjRqPmBLeGauS4CC/yienwIRdS/MZbI8b5ZHAySVa5Z38XRu1i+aeiocVZG5uLn5di
t19QLcuiW0imW6eWA/eZCe0sBcglugpKNCy8aVCLPg8B1ucA+WByOii9ILt/0wPRN7DR0rLNuuHn
z6BsXtTrYJDCxQIBKo6RJPVjqa1CGYUnHBmmW7uTMVJK7f1x00Pk7m86SssXyk4LO/z4ZaBj6lWc
kneiFSeIR7F0q7o5WFdRtcUEbxjxFnFQH9fYaQ1bs6hwsh0q9kTZqhDmxGR3yBXxfgbMKUMTTrhc
E+qbH/JiAXeG8167OHOGQepY9p2sFmpifpw366XAuOnG4iD1PaLoTsywMDvOBShoo8qUWiWJxw0b
mG8tduJw91PUHFaqnQ+tN9ovoeaT3q9PzzMTv7I6xuAelwTCcqyeEgDFSOQVANz6GVp/fMcAzb6d
zdNzZOoNATZ8FXAjJPKdd96Lz70vvNdX2OLRDNgwO14STd2a/BLbz6LnozfF8zV93NzmVgWVivpP
uuhvxYYLSy0o5fJpSbPeJZlbWtR5yh7Z8Yz1AcNqqVvYAHrR98XO/bZIMDVRTJfDL6pwU00V9vTx
Yc7v5gwWPnvecTlkSBn1s2Cnzee9tLAzMgArVH+xfxuuEelvRlvXQu0EsCDGi1IrmP1zq18Mp4tE
170TcBIgMnsstEAl5a6u0LvFtZn85lgQ3zVmlXSEln+jFhZxyGa+0K/qZpbGDfzA5k50NilXjipq
LJFI907UaFsXoNXmAHAa6vkXwwq9idFRcvA4b6cwmejWgbAXSzAql5Kg0+BJpZv79shIuggPhdwk
/1EODmA98WWkgYBP176NZoutex/4ZSRH/zUsVn1t1onIK8heAh04P2z0Es02wpqgZRXtJ9cEMlZn
4JKBKj5xapCScm+YvqQnBi4FPxZBnkK90A6PGKYihJqJGpdiXRZ5kiCnc4Sz22VLiPVFvTlb/P0g
K3PVs4Mzb2k3p4MS2glXAM4F145hRFwBGFtDLvOoaNqXGkgTxeTjnIyhGnYaTz3gfQ+mZlaR26/O
Br2RYk/wT4FNvO/NX/J522zBRpuP3HZmPuUN6rOt/93FIyhQZ1QSmBadx9QhJ6yBgWcqXsrIPUQR
8DhBRl/YeMfgwYpPtJdre7xPgDnfeJLeEjoR3sfhdECSL/ZNSMgCcsH4I3WvNGAIO1qY4gOr0KrI
Pzhc8lmwU6dqVWtybJijHydvzvDUkEQ9knmZYfeRyrBuA1oAb9iUpkAc1wXElHmb/w65FI+soGVo
bjYmmJMbZ7khcNOPuKhO23C2WeoscGjZqNy8g4pmMkgdBayhP5oBjVz2ATryGXPLnTXgFdNlbtGk
Q+rl21NCqypK9js4LlIU3FGrQH/Rt0vo9uxQ488AUaK296pluZwdTHmSe04puYMnkZ+ZmFn/laLS
KNQxs7JPdfK96vUtQ3XQmHiFg5BK5MrcPPT9swXt7oX63c9/hm1oj2ISAFqJLfvpWOyzHPt2MPAM
57N8gRg3sgeNfiJrP8rheMnSHzvOPezAkOFgszTCaps0gd8MCK6BZVSYSrfpFtT5OUFl/4/WZxZh
8yvdR+c2I+PuRV1cZWEPhxenRyNYSg9BXEHTDmO+ZV3dEv6vwI0YXj05/n1CNGYKBczYkfaX4X6V
kT2RPxl6AJz5S124E3UKiPHR9vbOPW1TmwdLSYpdQWf4v/y8zgpx9jQcHm1lCjZzo2B8cDbb5m0z
tSeq6QCTYPUbjY90OaGy8AnpLBtTTDs9tqouE9/v69Mdnt1oQ9ypZ4Q2QljQnBhKzQ588lm0DNy3
8W2TOFaLJS9L8Be4BnkG7CjgZIxGpFhxpigeRq7Gb6jzd7/uC1Vc3qcw3VIfS/03IVrJ8gY7M8T5
ZSEzIGMXWv7DbqtmVEQ+a4MXosygQlYd81c3nMG/pLF6yavbq0hZ27HNMxnTRbRHD0tKdSsSE5pG
4J5H1wAabualPd/w/UlqBPUO8hXYTPuNfoGRvicioSUiqT/ca6AmQmz/99ETQpoeYW+4QxLJ20Pt
cWlESuaS6dmXkdQ556TaTym7AtHFqVcneYkOA4ja70m27t5AAZdLt0GzGzw7qHZEQ4B8nxPNgD37
jmR/vt6wENc+841ShrmPbaj9k72DIx6IdDaEWF+1Wc1ryo8JcE18XwPnSfnrG347Wy2ccqfGyIKy
4ONL0+cPNUpZcYT+y1bAakYtJ/aITWysTGsrWZCUdCIbPGVZND9A8l3/MW2u313PWxC2IyrB/ePT
gnNIVJDbuzWrk7GNvkwM4pCJZXbVBRv853xzQKpkL7IW8hUZPZO8AxYVGS5P6teblExMfKZzx126
4im8uRj7AT6lC5E81w69r99E8O2KZ3/+8c84l/ZNBfNJlMqS/D/e0AJ7VRmJX7b91Hb9bajN+iVl
znlaM7OsvTxWTciWZ52WpmJK2ifPkNIzN2nlNJIt0ztplG+slDurm3ztQ04CKugxWh8Wixkh3QjJ
1lutcOCB0Ga8GT2FQxQUlY3KbHTKsSN/hSI4aZ/kO8kzch5wEpYdKWdegiaQu6Pmw+HyO35ZvU0z
ZihEc2F60w+Xbve3FdCa91iGn7UvIGlYkxQAfyKMi3e9W9l6bc0L9skhv70TR625GdN8Yys1UkGF
ZWGXGQZCNVOYw2TVYbF87m8P/QJ8kMhSZ8qkghreujKdGfFyQ+W/unDZOBxQ9GektKDq9ri8so++
+NetXhrASO0/BGMTbqX7qGsOvqdIIutWXSYOuF9X4YXmPtBX4FbAYnbZAEaJeF0rgd4E93pobWPB
C8XYXNdWmQKeoIHWQYt7sezy1xlP8ImGgOr7gtU1NR5JaYMKNaWBOMWT5yiE3yRf5/Hqr5kgm1XW
JhoU1V3zzwCRXDTWgc+yvhQW0QRrUTj9dxErSwqr7eoW6r7yJwHZLRRXqipWwVKuKJI5OjU+Y7N9
ab/4zSNOkSltw68L127S8VNiQGXhV67fvnx0krW1iQAei5RaJEMblsusUlTCqJ4ZHlfkG3UboU9Q
7y6MjpmxwmNxpA6q3q6nsrPehdveXGD3GzqZ/Zfx8+vAYMoGzpkZvfzM8wgfmeHUvawI8caJC5rr
j14vo5iEeB2LairOYSd/qFJQ0J/l3wCmESoAc3vrKBnRVCxJGiZEGnpnkSrFASQcMh2a7cfpK8gC
giL5T9CdK+UO0e9m7CAfHC7hO+79e5TohcDvqYSi2eJ4grvdJtTEE7173LwAgb+Ci/wIE09FbC7G
p/OS9bmdnQYmJGVtn576EOTpxDrtBON9c6s3FkTSrkxi3/4bc4KDufhxrxXG0Q0qQfFlex/5XYQl
jNyQDnaGc8KOV27MOX9iCaUJIytgg7SvSsoZpWH8InrI6Rghn7Az89tnzAk6GvIqWW4TBBPigpod
97JgAkJUQgxkRPXrRIu8kOYTsw1JN0rRegdqJ5DZ3tctvfg+OA2KA/rtw1ps/XVgQviGjcH9bmy8
U1Jq1frOQ8rkkB7rMAr7uObXYDqpCND5uGE11xSXsD2NvJ0JKA87csIJaUtXAYYed/Ln0HBoalkE
7pVw7qnuEKiax/fBbatkAkAhX89x2Zd4VSF/lbFktapY+jb/hoAcMhc9A2uukikhjMyPvOAIEBnU
rhENp4Lgb2kDMGJAxDLju5ojsJXXfpNX11hDwjgA7SiPeoVASg06AX3SOuEbDZ9IsDMcDWy/43bj
MNcAt8h2CZCoMlIuUHEC7kK+8a0hOREUlCp1Pk7PQaWY4cKtBCh9livJL8YOHFY3H8snNt5CMUts
V84hCT9mB9KM8/es5nrJpum6MLWgaRWDeBeUI8YF906JgLY+es3YIJ1m7L+Nk+mQUjN3xxlTr5iD
hm4dIwoKH0h0CADJIxBGS20PX2jo2gqRBNbEcqG5CDCS6QKtkT1wFn0QC8mue6ORljNQU3FJCjih
OEu0hEW6/f36AqmjmBEjnU1EuKQc4ifwU2kJaYYMGGtXOuLEPqsJ2ajjtbRB9OnI5xs51qt/VbOq
FiAd5modBrWXRbmICP3qGf4L6ZEZbynOz437e0TufSN4o04dK4KbhOmWRnvl4p7pfKrWjqKtA4Bd
P3pLsAns4FDfS3ZuOrOo74pHxn9olpJbt0RwJ9jbW/gqQvDwk3lKo6VhqrP42tOnA7Smu0qiPeTq
kITrdi/t/rtZVcpWdRaOqalsL9b0Yy+p/jXDEzS7Bvci+BW3X3EW9Bv/08Y7qUTrubX5lOUygeh/
hZoDyVDCiXiUC78+w+eWM12+yp5WRYien2X7i98v8duRuVee9XGwzbIyUaLzgO92/8nhIVAzAwjF
dngx4jL6pJxO5iPCBB+rArwBNIij+kBY/JBGVd6g00m4+6L8wAbYiZ2Kja/l1Xggh2zTAGdwmmXi
Fyotms0Ypx8btVcHRxD6EsjhySB9F5afVYcH1vPPEanO1kjSnpbzuSqMQ5MUKW2YbwzB5s+nF8+Q
dbfeuvnjYDwVL6UiTlo+As91TBCVcQH3y+jra+O1lI6dSJzU+VbJmUXNGvcVcZoUNA36Tt0Td7rV
PryXdueoKDuWcoUorNiAGojINbOqPVFPsi7t56RCkp+kPp7JVtG7tquGpsGReNcHY7W43/v+l7Cf
0TYR92oWScz250i25mlMZ1GOrH2W5jGNkC9+ZrhS5LZDNr1sNCzPSVzgQh6eDLWq86A1J1GA5skB
k7KUz9ZR+ShZDmoKr+KOG8WReayxdSd8yxlMEBZ3EKCT/oLAXg4qgIpI66G0xc5YHcH7HH6jKXmc
ToBbC64IkwO/OtiHDyjeRvV9Vxpr04hNgTooB6WfiHrDTr00YHSMwx2ww2H7Xq/X0gYy0oP+XLJJ
zcUu4I5PE61y5Yb3bZqQNIEE5pL0k1xg3QyoFw8fnxFd1OYUsAOftxSRpINViBPZn6qhwBwBc2lc
gpFuH3ByacKMIdqDGe5iOEjJf6ufM73SfjFn7yI2/oTz+uXoBhM4ripVYrMAqeUYwPHMRLKuQe6o
98S7Y1xJN4XTmPtWsFOGNLVBbdh7UYN26m+qdUX++hAxjL6p6mYhrcO0uHz7VEKTdN4lAGC7fSA9
qPNhBupGW2uOYFGXDGS9RxW8BlaneK6pFTXAIllnhbY6VUYjDa1hvugVuo1xuUlXq6cf0SeX1Qgl
DM6dXQwokoZbm9d3toQD2jcKF6tH6ElQiKRZ41eW0RAAeoxit+14gPryIYhGFfuP9l8B1rEPYtx2
PsxbPi1r0B2P8RbK3Hg43xsGax3yoXouYhkvlkZBbb7elajSGgb5BrWQgYUY/Xmmkz8EJMoyGCTR
ZfDAbc3rnA/+1h1fnwd0OYfiTt3M7+hgNXrGeRe4ezD/lXexONNgl3SiNp3ktTYLfLUZECfizLRd
KwAR6r/tybYDR9cQ8gQnxZfXf8MyCff1/8sxjmc4QBpAbkLGj0eKg/jr8ttOItbYSjQj1+pJwAbf
PHroiZprRxV83qclihXhvLI1V+/mRhmkmkzPhZmA3MZinDEHmkgn5OD7tIidDatgmWldxoruuiOr
0GMoY2w6B8FIsmdutYmlSN6z63zGcuN8db/ir6CTpmAbs1qYJ4/N/e0sDl96s0B3/EQD4peFQrw1
9nlqRDmlNOUpXqqpyDXLFjKmH7GkjYqDVLfWO9BME4yhSqiTUCZcfmz/+Gae2iiQu1jwD6uXKZZs
kkXRyITuy59SsWnRe4cg6qY3zLzDqhgPcY65UbLmLr1rEKHgqRrDP0f4+C++heftc5uI9JoZ2pCf
TE8Rk12R9SZcqc6DZj7meqD+n3L6Qsg/E8nRVC2NdQd5h8K8DfPo0x0n8t/NtNyvZlOkiw9zxJ+t
s8KtA+pUwuzKS9z+DsuLmulVp+hbvD7EDtHq00CP+ajVWuxXTVkL69yLW2NVoh6psidcVkJwFiAn
YxAPiqRp6SvG38EydQgW0AlYJj6ULuoBjOARKwHJMUMwU6V2654OuM378F6ywKcszzIh4Yv3mipo
A5I1Vk8Rjnd+xYfhWtqVJnJLPGYdvvvPbpm6u1/DiReIOp2ZoPGIFlhEsmwhDMBgaNzy7DSuj5gP
CztjxrWKhZf0vFWfeo+wNbQBdSZiqt4ovseUmGbN3JxcsoKmMgHebjvjlSoSFnJIOck703m9EpiN
it8OXQoDywfBEKJ7gsqbEuCKMHLY/rtlG4qQfNPZ9ANEfqEVLy9ubxuqWrCteJypd00CgM8SXMqd
xmSS1PMo4MUwquPr/RN55uC7yr/IV68oXLCXkqm0iQDwcotuhHHBLw1xMfzRgrMFzopzXQasYvzj
cKZxjYaE3dBEyBdVJsuMvimNqXH8y2PSsF31guE3Ly+lx+wtUXL8O/Jvk5dChIF2jbtWTlBGCOyD
eYVm6T78QuNltVSt1Gfvz4RKiq1cKS0WKJT18W5ZIhAeGlbSETzGtiDypB+pjRVTE5V2p2bD9uy8
bUxYzM5F9LcOFlqE+gcTUJXJLo2i4l0Cpa1jWwtgg1LA3S4ev5ucteLl6IvgM5p3jgby9Kx9pfs6
a/L135bi6obCzHPzXTFerdctT3eTIo7XMzrvuR9tnfPpGMVfAIPoiTaVTLDtsiUlrhlgdE37urEO
9++NUdiMLVXKrjX5cMubs6Kc0hm9rcI2aNMOZukB8HGFhuH+8QoItLc8u5zWpbkDgY8yFUMoUSNN
Ny0ASxh7JQytPpAxofEHaBtp0MUzARvRn16liCOtW3OzWwxTWiBK3L4tTVLZX5F1tdsVfyMYPDZi
W590nh3OdFBBSFGPdoV49WFavlHhA7j7p8D6Qry1B3+1tiQtn/Whxy5XYiiwK6kRhlg7Qxdq0kxh
+b4h3weXtyhRltTuqwgCm3QJq8cJ+HYf4of0QySxYj+jEgKN9Q+f620xTTYBdB0elkANxaMykDwk
vJNkogsRMghIxskldkSWO6c9cMlvSTJngHZxzivYZVDd262gyFofdv6srLuw16gR897Z+7Q7LR4o
GxTIdj+aO7P6qxo83OfBlEhf5cPhbMsSh435VdgV0+9gwEjnoJsxL6xIHSv1dI1PexqPptpEe+Yy
lSWL6KxMxHx6MPggWVLA0ESgdU/+wrM3++ipyFEuxHJ6GbIXmodoMppmUMBH06x2K3LXkLdNJDqd
RHnXGLceJnhjw6LqjXxA3jlrZuChSrpXVVm56sqDHmJPKq3JNz6Hwb51fa3o3dv2ENHDbnrmgXna
p9I82a3g9COdiyUF3DqnSmZ1wMYmvybrGMywRkKzHKre6PSkmkSip8ju7j8D6zP3/zptlqjAJ81i
y1wBljT3HQLrZum8bRqpcvySB1jhtT3+VOpge3X+BZM5uqsbil64PMAQQxr/xHdK/ZZvOjC1ros0
AXXtjKppiXRPv1UHPJDQHlMaMQn6nRhVLN2pnXv596nB+G3/O2JMcHwfPMX3q3hXtWdeS6p2DLyY
NVPWP8w5Aqjem13a3+UAnd6ixPOEWMm7JMzWP1VgX3DYMghwhzfdmmRtSPfkC6BiU3IlOuO5jH6M
akHdJKHeMNwiPRW10oP187YBZcBelMrhBvisbQDYEgkeqotnH/yQooABlnKqkoqOcJ3Qssx7ROZA
41lCPyFVPt5TLDgY0UctPHR6vnQYVnxqccwzI3s/iGWS3R+01m58kCnZjShurfnTjLSdLpkp/o1I
2p+sdeDSilS65/shTnU7Nkrv5YKDOcDy6wS/pdZRqOFQKN9ZeaACbPmHf20z8TKK9xKeQtTPsVQE
DU86lAPlwDcfov8pkeShTIlKcJgtvaHIuN7aqAGxwRcfPub+rDK3zePuZ0eJmkOB3bmUCTcdYjsu
uW52UKBcUFVpFtTsoVgigU0T1KP5LIMkYTMy0DmcIepq6xxdCjjMgN+c6iFtQQKbUGvWXGDs/vM3
GN5ATBClzed0QjlZCZTnwl9Q2ArKQ1st1Y5xYZK2jMn2I5aON2b7JvCDQcngcsbupkMHq+Jq5Ft7
IgsteYq1xQHJ5SqgfqwqVyFmVJ5EXh2nKY9mvLgmwkNYwJajH+QVBmmyWtAHV9UZ+qQHZ54gEJnh
Ph6IQC479NgOBx0ra9TvKUs8Uh1vPC3/K/zoNxkoqssoLV/8CoGl9OcL3f0ZOo9mN412hv2qo8qB
71dBm2rKoQ24IWNfn8W9Emvk/vwUVA8850f5l/bwNF/SFrrfTlCyJQbb55TrDMXbqy7pk74R0qqM
3/RklQRl5Ps7nLBSUT1bDMTZNe24hKnbIUCwQHC/W/z55nbVe8TxW+2NfyH3zcYM0VGET8ppJqIM
yJCwAoTKtHeJztBnEyaEuYZ9kOBAgEg2sNjF2zDPZWxt/HgjILLxcywol+7RlDbA8EvgKpugTAQd
0Hulwfphqj5+d6AGRUzHQx0SKyRPSxBJL9t5ra7n9ptS6bM34wFV1lmcF/WMPKOr1y0EcOSk+zw8
Ujqvg2yZWyi3+fcXI0YM0DmQC4igsT/KtngjA7xtP/x61laSAMsAjoP3oe51M6Gl8sWy86MF3s+V
1u/l6PC99GV5ZTMP7O1wJAmhHtIyoAlhD+MdYLOoyXob2pAkLxjFdwqRSTuErCm9MjMEIs00db56
jDmKyOwxubxplYAfiKmAWzqZpmNTkJHR1F1YuuvbESM7I3XACi5aunT1sUI9BXEff3a3KFEaXsoy
Px33VB2AYMNIk3gqBwMFt/cok84L/wzyG/QodDCJ9ZQUPQwJmg3RjJAGt5ny/6UVvNjcb6yoR3KQ
vd1jAomt6g6OG9UI52ZX9u6pRfAqAyfc0SL1Zjf02MaJg3Ozj1TdyWoAjniCVrfyZs6FKF06S8yr
Ae1fUovXDFigxYEQkFe0jI9PlxxITpJZJHERQrkiwdofbs2Mn2UBmARW3yQ+P+HScK56cxhChAnA
JB1H3C/2r6azAguh0VOFQuegJDw3ook4/5IG07Mg9V+JQvRPTKeCH/H3mCHETfsH+NViitxo0cc4
QgGwN/f/e4qrrtplga0p32227lFXpcWjME/kq81W1BwwcP4NEAm7hS9ltA0FRReZNRkRTaArj3EO
/WS9dG7T6uVe1QF/siPb2VPeQKSm8O/xlvlAvFWDk4QndPwFWyxBm1pEPop/CzsjWzt1RvvtBKVG
U/0OQVeyn2S0WSHAexgEToJ72CgRaEhTMgSK0OUPvve9T6qufgmIR7PmqU4+6aolT78EOd9zyMKO
cKfNtEtTQ3y5VO6EJiB3eXLpBIq1ggNCFh2k4uP5q4Et6IclSmLOypW4j1F3yg7jRKqTGbVvJrQc
WbEWm1CxEhrSzGuhmjQe6LmUH0BD2JsNCikofCJN/srXNll4ehg48AD+DTcHtS/FEtfS1TEhUOPC
o4x/qgjV0NY3yj3rdmBKSjh0B17NzBk6L98Fyxda33o9F3v767LBZZGu8q1pqSzKiSlLbz/JtQpY
Zy6KJ1c/50J5p6Uyr0G+byjFSYakxkTcXoLrrIa5Medn/o4QKrsUxvVNtYOMTFNycc5DaNIwWppa
Rds8iJhuVeJMwIdqGAFxUwqJWa+mIp+6SoFl6SHuiszq9JB1QP9xrnZqLko54yCLZ/HXVkI7YO5y
lMKtlSYFYnrJ/kNgfvPyDlW1j+wMr6j/uB80hZhEtQUR5jYuAogwBrrJbLSQwZ3S8dFE15f7KOR6
sZ/Xq+asK9bPMHEEPVZUXLyUdftz1ML3+0doVgrH0XeRb4aLKcZ/BW+z8DbFdrAXGQBksO4/+7Mw
liT4TuAoPkqkPEMhOSxqz2S/9QsrH7W5KFU5qN6437+2AXkiAd173m7G30HV2FnKhIF6YXFEpvxt
P9x+A6L4LbWjUkaD+411e14AqVvO5Zwsj0G/hBtbQWw49EjQp4mPybuofGKaU4fm+msysVVmwrPW
6cK+AJiSGLMIeBc+O2fKlX9vmlGvgABV3dYy2Yts1eLsbQrkXosLxy2Ua6uMFXe3SXeTNleqGqbd
kW48Fuc7ojhbCe5KQnfW9dXN2jFNdEiYTwOXdjgEjg21DShy+Htq1CN8YD9TB0STRGBUrAHNbDxN
A1nkkQJo2LzjNwgCz9XeSFY4BEr9l/5+YYic/eXZA9+hDdzuIfDCjxsbLBpK35XSLjlBwe1AQwps
mULrsS9QrtvEl7usXTb+pCWxyMl3c+qjd+5IkHsXuaY9NelWSIYb3sJy/1OfUgZVrZhGt0QMZPgD
Qfn7Ck8q+hBe/RVA9azHHbLWombj3yBPcyIFUjoFu+s0WRB14R0H/LQ96UEhF9M2UJ+Ie2YmhmC2
usNvY+1sD34x+2tp/7y4Ou0RkneDXPdYOFSPz5is5b33BBGsGKngdH23wbBP5VPHYMm/H+iTPhb0
wQKu3Ti3LqipRX8nrPRnCTIT2aQzFD1NNx5M7HsrHVcWi+oYNWg8BqJ3ruLKA3A+7nlXMybcUSYo
ab/nhFqsKFcLqNJN4yA3rljw4D+7mHtUZYPI4xwiO9Q7ylvo0wQwqFb0+3fQCCxyvkwX6il7BwT1
9aScJilOl1Gr7AIQtxzihwN4vjlSQm+rChrHzI+KYPt+EEoubZN/U2aPzImUfe8qggBfqK0SNUKD
XNTKeKw/x5xVEqsLBlCQw2Qmygo6wR3u/VJ90RRaWwntqWJ9JdEY8Yqc8bGMOur4K1oRhXVdTtS4
OF7cWq1BL8Kx4URFBYb2woXyC94Mdec6UpG38Io1MobRXB1tp5EMSKVIcm938NQVjxSJPCLvwhVG
ECWW8tq25FcvJoFRL4jgE2I/ODYJBr9X0Yt9I1gYHKlkvi4owcaoNcvSFMFIqOg5Vw17XveDdCji
kerLpt+E1ZVpTLXyd/kWqKfcAI8dTXMIIuaFcn6OHIShuyUpro3vVJA6r2EohO/VKcmWEWfdMcAR
9PjJw/8JjLDyLYH3AND4ysMpXSoi9VULpb9EFkwK+qFmiBg2A73iiOdMIm5McrGC1UgCjgo6k7G/
feiTgMciesI+aGbXFtToey+8JhdYD0OuoQtjYVPpOiGeXOZdCkbufBDoeHTFVtiAMtY52vb2awhw
rdjo4MIM5GTh2yn1kYYWzSMX9BHNhIipkiKdoAw1xbzLFB+Z8TlXghOWU45+WiSI7j8Z+f0ozGs2
SqgoD29q9iZdUUZjPXiV/viWCTFZZNoMec8HWy6JY6t/WivYNxIi6Co7edFHx2jNrzXe7RXolnoE
BzhNiWQPm2E6nvYykDjqfAbTztCJl4pSfYHyGHZj35gsNcxETQQvWD/77jhhS+oqiyy42j+IL4gR
Qaw4e5FRUri6NHch44GB5gzfu5/pu7So43r3yqZvdgQwbU3h6LxENl2GHQNk0kCLl/89jl+eekiT
X6wGaacbuEcs8QpaGQYabCvAeQOL5QQ3xQKLUKn+Sdcor0g9IAKPYNtgM+r86Ccgi6BGXeiqBW74
D+qjeIX04puEezDHjxyKfRhfABuANLW/PiqLdxsQio8x0+iYX7jVP5rcAW7SO/znpaY2kV9aZnrn
m2LWQxCDrfb/oErGdU4+rpT1tPZtpCvrgakvK/1/pSXYS3vah7HBorHjFvvK43hwwXPkINWNDsAT
x8Yw9Q3tJ3OzvEdzZ0n/yeFhsK6qdSWnwnL0qnMw4cb1qq8gWvwzPjaCgaHXHj6CLnhDPENu4zZa
3U2EpuMXyWggnmXuA4ufBnCqPPTsHi66Jjc8oaOGl1j1DjhekeTw0BbS+1B28oS7lp+lpWApwmFm
PAYUt+CqHyIKAqpMdRs86BIPaH5C1Jw5JSp9ia/84p+Jga06+0ZNHKZ6PYvpFYzyKSBdYIBx1rNt
B9N3J/3kcfZe9acRskh1/9cwRSv0is/LndP2fS870TnTT1M+vGf7M77IR3RJYy1mTK3eWkKjn3f/
qRzAjH41eLWG4oH2y4TEffjAJQbeXebGwDgYJsjjQCL3xuzuycrw1S0FJNQbaljhd+bIY1enA2nX
xNo0YZPKQ7lkHkdD0YY1Xzvrk3rlFfQP+19K+wElyy7367e0UPYsWLlTUWiHEHM5Dg6NL4nqrevq
k9TjJwzT0nnhVhSHVg4lHSb82ivBJFSH6HlcgceEiJfYaLJNAtua4kLO4vjWWPV2xM5kxBifi7Sn
5tjoGBZ95a6HHeJ3ihyc34YOzEcGxT/eVfieyxTQhlgeFevkg7GFSMLDS7Eb9t9cXHWRkcyJgxfq
sYWJ+43VsSRwZAJ+d3DYu+udnv8BOMFw6COZIlvrd7WmcsKTySpnWfPsbbBGx+3vddnJdj/M41Hb
eSAzkELfpAIfoTCaMIgVT3PmOcGO4jjR4SpYjcAAr4e90AVXdAINfQdzgi4CHb8/N5qnov8pcjeJ
uJoLIvTn4NdFG5orZKNeKxhqadsDT7Z37YiJ4RQUnLT4ooThHtG29HIqHrezhQ0qdq+f2oZVH64S
RgOylYJWFACxg8xZGP9iVyTAhK3pN5iPf151wgmobwtVQXnvPgrFZck61gxGkEcUiBK23SdSCAvZ
xLOpzbrQhW+QhdsKsEiPZZ2IFP6XQQeRQQX+s9Bx/4n2ddL/7dsnFJVAjMMK6OveImWNBRyRTP0J
s3M2VBHH8jpm7029i0Jzx8xwaqmMBcfDo4y/dkNvDgieWaMCRbzvgxlL6EmchNOkxcF9vjNHdFln
gKDyBUlzJiVsb1w1ZhmKlcZ0Y1A1kN7YosQXPGVWUEg8JXili2CNYfK4ifzzG6WOwP/WwkFveln5
Eu7QaKSROBSvZ8fu3ea+lu5HPFt/2D0ksznkOwUYIPvsx+Ad8W9puC39Oe2qRHIPVFzHIYD6prot
PEHursoHZaXkmb3J1kiZEt7ikXhhHv3qaXLXaZJA9boz/FyS8zpo5ht7eDf87IjOvInGkkMQ0wKr
LZEfqTMN4g39YWYECC++DPWpLK+wwtyMgHMvhN9hsukcbjw9ZYuiB5JeNMsPLTjrFQgpbpnwy03R
Ahx84WS4KYN0bqp81w+1bYU7XS/89tjDDy6hgW8L0IHMbYd7CNWiemqOCHGR/HE6FulQHmvazVg1
wj2UDqfJZMD4/FpVD0G+VV2FE2AYmE8hdk8TMfiD4ukU2H1L46tyzPHDOCf5eK7/XoZwVzITCpYP
znTa/5EPsSdo59IuWmKJrj6v4M+vbvRQ6g1wYNKYRKxxKUy/YHsOlO/iU4DziEUonGHvICqjv/8K
vQJ3JIUqFzCUl8YIqBVjn9G5jAq+dn0OsPejvhm+HnrodfAn8LP+TXT6RIq3JSMCRsTZ8fSG8tdP
GsTyckyk/ce4JXJs9TTBvaVhAtV5alx3JI+PNeUuMCgQhO2YPly3n9aWh9MegpWDyLQva6CqoF0g
LENWJMD7pEvuBtO8A+czw6Ru/LxRkiR8mosorckhQ2csVD9x2fKjdWS/iX/z5DakixrbTtq9VEXa
T1dA7XIRyzti15fnBeyayxIP2zzQbzeI18RhSF1oCMR4NvrzXB9py5jTQR1ocA/x3+SbngG11MZh
RULo4VMxlu1L4F2vSyqcJvpwJgslGdhDeT88rIewY6Ku2caOLhhvLQuvAazzGbHc7YuGOoMjj9YK
zvN/zBhqM3QvUAGxUK9rZuk9Q3IjTIEJSNaUCihJ5yPZv432gLM0x7ABWvdbhPZsd83LZTVYCXjc
MTH3mvKB+oosJgbY7W0gv1vSMiqJQrxoS4lzaTWXGrM+2vg/2uBN2hA8U0t/TqhK4Vc2aRjBo3Wi
1QdVTIJgKy2BnEEfNtePZapUiNnVl7QaOKHBw6H9IKUzZBvzDjIykjY14eL2PTvu72w9nNJlcGIU
/bGt1L3Mwp53voDTCFp31f/YbNQdfcrTsDPDF829ogK0yV8eB41MyvIg5j0Oy7Z1HPCiwhMTYH7v
tAsiRB253x56JtIyY2IIJPGuq6CLm//F3gz1SKRSBDvQD6wZlBQvXBSb+D63evrV5LtLusgXy+OQ
DZtN5NVhxC3zDm9QoR58JYVvuKKxoYTIXKCXJSep4hwoXpXLEG8rnfdkWhblTpEAOzFRGwFljEoN
Yho4b+V5+/szgixZ3j9A697aBtn5ZcCBsZ7oW6cQfAzCa/l6fY80CS08F9PpYLeed8hwyrvcOOjr
rMn+YUthf8BdffKNlTNpBFab/piTOjkJKS5DAzVOhkzlDrP2ct4cXZmF1Z+tOLq6MqlmA8QRJgTo
sJJoV1YGs5LrZBRGwBAT3V32D9JnRuosg02M8DTmwOKpt7nv/vraX+krLTudsw6edqjw1elyb8aF
xthl2wJPWMAT7yqW335V+J0OXACfZp6YGniQ+6Nho+SuZxvt6WYqgIYT+nMPRCVYCTqWo17D4bqc
AOdZdkyhpLU3xqj3tNrBuNZfV7yzSGWR7yaIiyYyeji6CrJSMz36jr5pdhqNQOoPptcEVXVeMOZk
hUZw0byzOwcVTEkoq7+gS7ykYU6lmR76bAaWB4Oh9x6wINiC6EyNxTDWY4rOa/c4ZPO6Amersoce
eTjHvlwi3WR66i5jGc0mDm50Xox5UZeS3Z2njFvFAYjLze5DC+AzxtdwT03DnPmia3CBajiDIeek
r8LEvfmZVLEgGqdVt/wLsXQBryaWZwuG5OBhD3Mlh1TpJTr8a59k4x9A+tv0yg3yY7NPxMEG7Y+P
baFAYDs83AbUiVUaimoEy+ERjMXJ7PWCNMJoX25CqHUGHALQ+l44waEwN5HJYWHeWdM5CtZaJLAv
ZUPks/g2AIPraYtNw2riwYrexIMV1zjf6T/BxHrJmvb1kf8AaUR1++0QYV3ZUdP5S9pcDYL7WyRX
+uOhofzYnKKHkUiFnApGcXYoZGp9ALXS9V6sMt4413Ry16MboOsRTeKg33fVMTiCdra36yQ6uZ1b
kHcs71C86u1ZAwyqKIBu8s1SiWecX4xSlaapf+9IqzgtVIY1xOz2/esp73fpgPZlgiTD8d3g5Bjn
AvsIvNqPTSUZ2qJs4iJccWGsqljL51miKyscLpjUwJ+HeCrhCXACvRr22gtLLnM/QcUP6wyR5Xqt
rJydtIKH4sVWnyoxgCtJxAAjdvvJrD33qp7ruKa/AzFnFdc4WhbXhlfxa0jj/I9hx3j3ZNnanzcV
k2c3noisUMv+lvLTxD3YkQGR2LY63gqOAaY8viwnrNkg9QSJb4ZdHrkXVSRyRt08xedWL29ALifN
/Z+9XzGQHk0CB6+S9Nqfs4XGfYpV+6BFRC0uJ7PId34SqQmu/bHZEZKy01hIF9OAXUQCFYyZumsp
XMAA2eSc8gltsTe3uW8GhtPx0rw0QWKOi3x0No34Bst/Js99s4udZB+V1AbLTzBb/zPH1ZyHL+nU
clgyE2Cx8+GZkfkbaGpoJzZlF17CdemSriqluJZ0pVELjXBiGwlahI7ITmVVctOuvmFFqKIWuTUz
arF3reSU0hH9F9TuqUc+t7JFQL8C+YvcVQjr6LrxrQjH+/NDL69ofRioWU7PHvxPnpbZDZiBdzem
r0hK7JKstutSFs2rlbLulGtbatvLh0RqqbPdfWFbajN+rE4254/7jjMT5woo4TNjhSIXcTdeW5hG
QSz76P6ab8pr+5F1Fr51sAnRa+S07OOq1YCMuC7YDp8k3HjefrfeIfNBx0WCZDgPj0wuKnY/d+TK
QMfL0VIjLbq3IKieVi91C2kpHGMSqnztpV7nYGM36OP4EW4TA7OMmI3H4B42/NTSdM0nG1stcNcH
Rg1/Uw9lB2sKgG6orhdKq1MT7otsfgCh6WZcW3UkTxzgbAy7apDe1Uw3IWcX7rg36wBVrIDoSxUk
+pICTcpwyKfm9+9uE6aGSPscBFHlIT4JXhm97Yuuf2t5mQba4SNoGjO8BGZ/jcnSSjdiV11kmIZo
nTNIpJwDw2NkG0W7XndQx5r7i1LjFKVnRD9efXDye6lO1lwJjVhQj/G2Q6Cc9/lO5wEtE6XJVVrK
lJyPtRlkdMD8Yu9/PNeHdRIybxkU8E/GJMSMEA34VbebKs/xz+iJz3OfGLtIw2EurTSXMOd3tyy+
B/tNsSxr4pVoiE4a0QkKAzhgkU9yi60zPATaSnIbB1ndb93iBou63Au7ZbcWU9YRLY+BvrXwNvRY
yAr7Gt79nIeWXlfsq1ti47FwCSAUKsqeCRFTtCzM5RVBz/Fkx42Bes5tdkgDnObtYsgHwe3N5KN1
HEEL4VkYESuZhkvWML7uPuSIYspmx/nrmsvJ2DzaPLqHPX1CoQ2dOnFMhfRtuHmIAxtGtFUmbsqY
/GW+BarPNcmfZCrhK2NWAWjLEscPlqryEH5EWgQsa0XGEAA2cBHmbY77IjK8ItEkzZWbCvI7SOmk
2uQOtUFGs2a8fRG+7/+F987E7kd5sS248WIi7HwUj7sGnhcC87GitT2bWVC7pbSo851SHlSCN6Pk
LxHUXUkLtvQAtXukcdRTvZiSlxxvz3hw6ZtoKhY6ksB220w7ApvntI/XzheTPc7BUmlGmyA2yxhs
wOlprqgD6HfURntXo4HA6ya/TEOJaNqYPdm3/8V15S34SKWjRLLRLkMVwC0Dxahxstc2EN6oePzX
j/4cgzT5RlLpQsdBIgG2jfzPV2AjLcdHw5ffeIA3fYzbyT2jJiugT6hdDp5W7N19/lR6xCRUVXBc
q61UD3lCYN+YF+EKqywHeWM4X8sxXOwiGVfWQuB9ksUSucQvTUnvnjw+BQiGJNLkKMaCUSwtNunW
/+V+rN1mfB6OsKmzJhn5LUy5nXjOtMbfEqzIVS60lY0y/xKNciyAMQN0cot6VwTq1TsDTZNLNkn8
h7H+OykkaB9hR1MTo/pm4T5u9a9HlTyIUfHEBsGNyecUGBGhygzcAJLrDpL7djubPAr/eb/U9pBB
4k3EWOTGJ+QofWN97Dq5/Su9dmN48Mvc8vIU314AvUKNAGd1zUy8roRDFssZK6rnt9A24PcWdXqq
nRxswCPlZjbk0qRaoZ8SZAQApCsQnxJsZv3zAJvJSvsa2eQR5vvzPTS5lYVHl31i5Lz1RhZcZkYi
pjYT0i9QPK1XiOgBhLZ7L90FRDRblg2xCc+L9eHJeWAB3AkfqckGDf7hZ515lsrv3b6j0Qks/8u+
mPNZgiBgoNv+5a1lOhCTbB8kb2A6J5KaQHqtqISxG6k52RZJ2Qw3tLPBWV2JU23bnfCRJBAJKSO0
W838TZ9ak+qmLScPATLsDqkzGj8nNwpGNITpm1yZC/FwXcn2OTPTcC+hvswJYno+Sr1Po3LUHjJG
cm0kO1PCzk500MyKL/pJH0/MPnGqLSg/obagQ4hl8FEQKWzwE2lFSFaHNzGYZdZnEeq5LQ0Ew0lE
ksJurfE+FZvTPYqcUF+ZrNT6D5rVMB1+PDqzie6b1oyTbrzuXwvxRk3qpyqOUInE9/fbQs6+KrSm
s3wC5BjCsdGkKWgUiA/ciTqyxUOq/mjFgm9S3cXV+YTahtexLyho1c2Y1Uob826Yv2Vxm9Vtm/6V
DIC7jVUDaomk8e4+AtyHHl6GjKJj+JpFwrgyB996+/epkR3aqNJl5mSHtoU4tv4o/tF6ynGS0rYj
AsLTDqHL5SytXGC9tN0WiQ307Sa6hIGuHLpGujZdS4SjIHZrDWWm9YyUridGs3VyHqdSIt4/hN4N
b6mu1AtbA2/lN4lSiJH1ArxPu30ZHcJm+OqEBtqutn/8A3VhZhCFj9Wey/hn82Pt1Pn5FDLqwDV8
k9R/LzD48WsVNkwswDv4gaYvAkZoseKFvz1UYnIQoHA3YHot56Ol/H33mKSA2ArADYsYfpSqTXSw
6QiRg8SDf6qOXvK3wqUcs/BkE2J2FIcvFjo+4SUuXT5TAc3kC2+Y2CleoHxuAdX4xBxARNSeWIaC
5ezCR0hapQHb4YCK7WnJhjkcIuwpn4fFZjr3u8nTLQcU8bAFx8dyWe0JKyrnYugOrb2Y1VVwsKIe
mNr5gwgMETdv1wXrfjtrAqBeCAzvDazVQVJ1TANW69jvZwRPLDI6WGspWgTNDvHK3+iGLuoxSJMS
fDN6Kn0CMTRZY+y/zuTzjddwNcklvd7gMEu/06fFq0NjICSQVjGhTf+Szz4eClEoTlIsDP9SVPXH
zctahe/gWkteFZWFnrQp/fgHeFyk2A8KKK502jtg6wdsTzUntNqgBfOhC7bBJNpvPvXGA6xUc2AH
pKIWKfb9/yqFvcoMnVUsa5wtIEIvxWBkI2QTTEI5ozqn7yhpuvkbb+IqmQj7El/fCXEQZISCN6KQ
VCC4wISU/nlzAiJ8OaXzNehODSUJ8Lansb1HUAnWnZlbyk2Zw+oy5GCF0n84SolE8Kb9XmPiYj6F
k96+v4uDrcbeX157YKLeXWF8jRm8H1ce+BhKnU5NMpkzYxHyGDXPNKZxPswMdLXX7nJTXB8d8enb
G4L/Y36mtN/xtwIT8L4CBoqAh5TN9kFJgdAwDkSGO5smJdSPgmHnwJ5FKpNErM8WGneon8/+NaSY
CUqT9czAem098OsYfEsAW4oQ0vfjAaQN8lW6PPgzDdkWh6wgQaNz2RYM5bnkIUt4JRMxh4ipKYFH
QC8s8R84yLhyudjDkTtmwFgzuVdtEVZbRPzetNxZEVxnihqIeoTHgpSOX5X4dRHdPKs3C/SD21qx
tkn242bEXqBCfx+KSC/l36qwAvH6oc8WC85O0pRaak4lTb7yVAP25xM7S1lXGnr8WaU4McgT+CF5
Rj5MA46M7FQy/fbp1aI8+VcGuQxlv/RLOSOvUATqWfmw4sp9NpttobFhAIQRKCjq1GikW1BrZ8GO
luhpjqMGLRcgmc2qvcWq1AMAS35WkkSEj8M/sVZoKfTALzsVht64D2tW6rF32X6LdE6LqitIti5k
yZtGUpdNyZ27Bz7xNioWjoTNVlFDFmorPz1EQ1tla4VgcTLNnTOq6VDCKLkmj3CGOEATih+o8uei
EH3TxbVrbG+bFXR7SiI6bfRr3LV4aUKwT8kVYy+N9VjGnzsadEPh7tAXNRQjtB9Wo17gGlPp2uv5
TxyaaOhlr34Pl6X/lAqXL6iqVGGVL7wHgZ7UgpwbXn+FBO5eD+iLwGkhFC11ZHhWNfS2uk/NzK5e
3GAZZV7fn6Bcimja8VV1cXG11gvBDy0pgT6n/ewN4kvUN0hjHWhQEHuapTnty0kRWJtzqPpHJb2c
6q+sH4uuu+xwQnwyYP4z3gGjedgykLFXtQ5QjV/HNOIlbQ8YNJHFmusScadV7aoLE4Y/Z33349OX
AMh7PkqANoV5ToAuxWe5FmklyyW7riL0KZACuidL+XDRNp7GM0WbQFFoaNGFKGfCfSXZNQV46MAE
i2R9oPO7giDT1actfvAzbf98o20lRZRmtCrFaLfLQo7o4AzpqSJlABxvidRLv1Iy4p5E8pwSV3J3
TJJh6w27gMc1KxhW336KRu486tFEmzIfdM20EleLJL4KW4B9GHByM8Ob1soeH1uQl91mEQevU3Dk
GC9JNv6YKpsm1uv2BC9FOiLfkEglXW2gb5/iBpjr8mwF9on7DngtZ/wafGXdVKb+8psryecv2YNt
a+HIvMBZPWtEqT3EzG80+FAQtl2wX60hLFjberbJmJKp6pwTJMz0u/zJYOS3cgSpBESZLxhoBEMn
xS+xKGgeLfGa1GHXhaakVLLCDSELpI/97ayr7xw51MwdCLsskg3b4RASIZIz/SuijwCzcMVYIkbl
kUtiRPa8kOO+Kzn5ZuGfrTx9+rGv/EKHy4f5943QEH0O4qcq3LzHxdjl2kZq1I7oZZxCCANyy0v7
Ako+ZsH+9mJnDehBvVOYMod/VmdwrcyZHUstlhxgIzgoq0zldkMBt3Qc5zJXFN6ifAmLEEnxhQsQ
wtuOklOZJwdZ8BAEfwo6+MxXHBmtdxO+iGtvwHckaKUK7gPq4kTnIVTHLoTEOK/0dG4szLi/9+MF
ozBEoi15RtbceuqzWq1uOLSyJjYtRIHUz2HerM9PtD0iuHHqWEtsAksDDxnIHBgMoNZufSRWtbnr
Op10oc1z/XleMNfz1d8mWRevpFVrKSY116wpKTJK7HMiZwOl7+Uje/bZrkmN0vThGHPBoxHz/3Sx
3peDvPHAZI5qxUqO2uBGjzMW02FTWKutTppUyvqQjHJ1Ne3weIB0x5UF1zoA23R1QgYSocHewWJ7
tzfFhcq+imQ0mqX7pV6UZrNbUzUcqevFtXB31pWrZIZ3EnsMBTFGglt/Uuh+jM5stfGvIYrskp89
3+TmiUbfSToVIHhFDFIA/P53LjV/Zi6szwOCwpi73rEpW6BAqmroBWC51LtH1nOdblcj7ySKT1BC
X+p4/sRO+GxWQT/iXhQ9//mr0Ej2vkyvzKsJYhM3mO2D/THV6TK6O7kUdR3HvWxph31ot2UkFlUk
zi6W0zwKfP8PJ7jPPctK/GD7P0+VuQPSpE/UlI3TGwY4rG9TuvU+Uw6VTiVG1fywJAhaRTbcxdaA
Oc/AZtd0Cng8GN/uIuOBRXcJDOORVbXQoEHRfoTYbX3ktvamsFvQCTX8bKow0t6Nwok/KAVq7VB+
eq0EIjD7F2ahqOP4vn9/3KNKSvUA9uBuya4+8z+LzimYJDNSFXVoKyZei9Dnha83yr2GaMcX36ri
FSJTk2lzDcv/bpRUVQ3Jc+xSK9uMNK0HBD+cl8tnN6NlKoLqQ7wz5I3yPtOznTEQUfFVmEQnZ7LO
VQ/WMgDRWrz/DExTGXP267cVOkbUos6aOOzLDYLJXiVvCPC/T9VU42pTQjeM3wUw11drw0l1NUV3
6HhvLa2njJ15T0xgv4i+D9D6TA5yprMsjuVOFNFNgUASrNu5u7CQByccco2oIjPgbAIjIK53N9C1
dWIG9Usn2Pan/SZQml/2oUW+CIgCE45IEk8G7lWq1DRPuXhcb5ZtGuyH/uYxs0UgG3zAR9nUKgtp
mhnwLqjN4iNeAKlKd89dnescFtsWLUtoiX4zT8dr+i3CV+JE/TTwvG0q++qCfMvQA9HZxhGw8Vj3
wpuHAV0mikgA3gTnHKTMBhFhjTXgtDXb41vVVIYDnJrgJtnlnZgkLl7plfHhAuW4BIhHETUYgAQq
sW4T9gX8v0Jxthhthdva0qJK4gvDVHtgdKB/Uu9u9j6PnPusLNIhiI9ce9BfMUMLdV9qPBThTDou
9HyL5akrXfzaHQ15aYBhp3sYC8DHIHwmWeHnPSl+EA9qGkgA+epcVmS/GlgJpBjyTtuVp+FRfKfh
TpIGPsFMNC6U7jc1KXLCB6WgfZA0nhESZ166r2vA6Ker6nZ0wewfMHqX/VjjJwHcDDj1//kZX4lX
fqyzUsbmgvkOVENAvX1gnfKgQEa5URxXa3kffDfAEYkkHE+juVEndkW6pGKUrujjtQ5zEIWmPflP
53xtDk7guBfyAV2tL/KGoiMZ4+5xNJrQDR+rdygMxFe5pMexKn2VL7z/h3A5z66LVwn2WFeLHfP4
P6QCs2hFENgS3tfh2qyl5xEMs7WWQlkLsXmKN+cJA0YQTfJFqCMw1DUaIHwTI4Q6gndGl4yCgw0U
p+OcfPF5wM5noRFL1IVHLXo03UBfMkC8ByJQP8t2/fuDMFMvDzUTKFIJIH3TNdOM29Jt6ADavqim
jtxOf3G4OkgqUJaL6tS+Kn6usRwSz+YsZPizXc7Us7ajokY1GGnFYwmijt8jK2XXczgajtvqgibX
bY+bQbkRshp/Yb5lRMOrOgMBp3MoX4eaokfUdgbWqr2YYuWfmW9mGcBCwelKB5kstu2+AR1Het+L
8MGePW+lxK5w7KzyyHHiE4EuKOsgj77d0PEwucAGV+NSvS7osx1IuP6Ddwfz/5mT3HtAvVqedHgq
w9A8kYR/T4iMbdhIY5doinh7dC6H+Xnejc09VEO7JnuhwcnLUMDiHRpeM1AJDNtZCBHBsKyMzpDF
RAZ+jFh78CtlWy87nCesiKzFXF9ViRPqMOjWmYcYJdCcOAGCF3YkZTVdMR50604iIaEeMOnLEa6q
b0PAT5xOlmLiRho9EGMluE5BpmAnh4y1mOWi/uZjmP4LrUaExXaME9i9+kMM78iGGAXZA45lDYqw
txmEXNiKAv+9tZ9lp7AoPNHTdGCsdxvuP8c8Blw6AZ+Z/Sa86bZj4kb/CcdhQ9FIHDk7Q51dmWor
uvTipZYfqRyo5hkR6yDsDg/+quy11sYm0AObqbdmkU7c38j3hXriDl8YH96cVvhxsr+MSteSfk6i
uUuReeU8zxGee0qvtG3W5KJ3/NTE5uvcgxCqqYDHNWt/u8v3oRXb+fxuvF1QNPcZeEQ1eZADzruR
VMUBwvi5JzhRaOaYuqLXBZ0LeenPl2VmbZJlKfaav1at6KB4QyeqG2bTpxKlLaY9dd6lFykq1X5v
QtC+3QD0QTSNEmIm063K7vIYdvtc7AE1SGODW3VDdCWCrR9C5XchM/1GdKZcD2uIyldi5IYqKUGE
vi+50VGNjKXO3T2s24QHG0j/81LAtKXyLFXed22Hu+szbgM+hQomA66FLNyyvN9wOoB9H0tztFlt
PYpqZQES1OXX73C4kcGX1b1G8oeV1u8oCjAa1NoIQr9VSWRbnRHnS3nlthAuDRN8tIiEUp0eUzqY
ZbOKgAhVKlObAxU88uaJsJhpyGT08pmoTZHGMGLdv9Lk8jojR+DhqmbfRwjPwnQTkPMoRsKdPyFu
NrnTjpt/XWtXBHE5wLFqzml2p66wlanjNg3frr52lBppSfK4B7jW6VvhCfbLiYTkMEVToAli4OtY
0BZBdotz8KfEEFbO9loJJw5JNLmx+meBd+fIK8fUakXB7EeDj8MJJZFw0jaqQ+UrbxO80/fsZJ+k
U+WZAuJ1cKvu7bOtUIoxe9syRo9FoQNPzl+0m1RHZKFyBIsu5EHhXnGRhN6BRHom+xV21UucpyIP
3RgIND6kKzrKl7TXoKozLA2icDuMLWtIY8AXhgPMt7qtq9BWoIvoWGEKCwUfCL7BnS4x4+2674p+
hC7tSYnsBWCYIXno4X0E+2cpXeFtFHMP9OY/JqDWBIwpiiJ0Q1Y0/scdGakRuo3gnmIYQGhdruMZ
JLWM4caHX6VcQaCG9mhlFkwbGFNYcxBbqKDQzCqz7wHtmCu1sQS7rmmYln+zYpM0wB88zsjqrmMy
DnlxAIkkyhxkUlf6VJdxjt4lKuLP8eyKyyaNCWuTrdZK69RzvsfN8dirZXTENhTDnXKgC5P8AoSM
KNsHFDUa9/+v6McMLNd2oS8WhZrjwabGpk8BeTYDRqk4QbqadpJHmbe5wVpgkSUAgT1fng6NCTDY
wFedLqXThL6s4xniWwGcaY/k+M9ARhvdAASlm3dv+AkuSbiC/P/X66sOZYx8NQBNEDumXGqZWV5y
uIbw1w17LTZz74SDRlLq+YM73YxUNdCrrfYeG2LczWlYhlE3sCjMpx3syURNuLjfH/Wmz1lb8JnD
hPZgL+L62i7SS35MwkSAoj83/yKDPHvaB4Kw6krD/zjljp07CWwWljAbbS/M4nvpI+nbEShURrNJ
kGn62SfllsRimdhZXuuwTLGSEeo6mfpQMWEe9D2DdU/EpDsTa+jPWbS7KNU1DrJCStVzKY1UggUC
2a0hv6apiu2K7E4sk2I9aVEHm2/mcOAo1alS2upXhn8DDxmdABFOH4g8nxCNeuhejbqMM1cVYAO4
7hryhQYIOsvbdeol1uOaubF1uBFKGb+nFScTbemabJ1hUgT6qH48Fa6a0engPz3e9WoCUakfTmt9
V80KNLCgT9aoBzS/SCWujXjThHHpc6EpQRt7E9BgNOyKboPgtgy//4D7VhbriXZH91RIqF1FCSiQ
1qQvOxOmypS5chbIy6GaEmSdvDNgQGSydBBKoaxou2CfcV1zWJzt7f6HdQEhyUUeziTJKKByInmA
ZKGqXoqeW9gva7nGa9iQzzUXxHX+PuFhNTEyWc3JDAwPoKl+o4PxzRlgxaWMxQ7CfVQJCZiuMgxd
RGVk3LYykpIGLjR6rT8pUFZED+KfjEAsi854jJs4V3fit7+fME11nUdHx9UmJygUxZbcOL8yHywd
pUIJqsYULYBlWp3PcOQdLmRmnniS1jW4cyPtf8HT9j7cIhSZUitaVjzRs3mUOPhOK9+qfGCri0z1
3jPcfldkRBzLrQS5fatsROuP5appLGl27/yxeGoStsMvi6FB7g0Iqfdgv6f4J4uQ2zORDdIYSKSu
kUzDSDR+NV4S3NokNfPf7siwkaoSdileub5qj1hMVIXlb+lmlzlHkpRrkyZMLcYf+nhdTRliCdsv
uplb7c2tNcRymfh8arnW0AXrptyQAYs/xEXaAzosUNSQec36kd6m++KBs3CK0j9N0NZEH+Gh0pVw
/EQQawHx49q1r+djUTmjXhlnne40+4UrrN54oRBDnuMQ3nq2X1LlIETjzGjy8DKc8bk4AXHzr5i9
gROMCYMfvI7rybuxb4yB6hSnZJb72xDODXFyFtwmMuwFq7DRBbbkg9WZs1P1sUc7JvU+pIMoOlRj
7uhBuWX7bAqbAAl0ClOinrrCWisfFF80T5gWnuaCkl/bSC+wwpcqepFYZxJdm3a599eT1BDpGXwE
LQ/iJYg6X792GUmI8kiEdyDhfQa+PaGC98i8HZXaz7Phpt7BqmU9GK3KfIjPfb2Cx8yuY2Nslh78
DHSHAYYNswObl/mfPYkpXclXHu9Y2f9AmDtMUhNREW3QQ9nx+LkGtngBUPxpC1Nay3ZSA+r16HK2
aUtvNjzgQ0xUv8uaCut2k2lxfLdymyOnSTf6PCIcK8icjY+ag9pZvyxUcMdX6hPuBqqljXNXSQKp
ZakgCIcMZAeIbODg9EZDZPsoMV0wQNS9c/MDYO88KcpNrEyohOCNMlEmtOO0WScDGER+9XEKYkPW
n71qrqeWt8PX4pe5EnzXcgZ1Gj/3MurmCfpzlw6BO3taE3vX8DleIBll+J1jSUX9FXT+nZ6eqGZ3
tjVcqCY5MLEjgvHIt3ZoN2kTeq82Ib2+Pp2M8+8Jgo5nPOgasqQIgzZ3m0qMNy36fseETmM5rxaM
gA3fq5Ri8d1rKIfisO16N+GODEDHzar4KhwDjmn71iQQ1tm5D8AmOzXo3mDRFyDUxcOHAjLydce7
Wz60VL6uLEDQ/+KyMccUrHAJHG3rRNDGcnCVMeijM/rrMlESgwWSf9UJe5dkhxOqYAwIax51cl8f
jTgaAtbAJ+1LZQ0P2Naqc5YnucZQNEAi6RU1Ol4P8G8trdWdHJfxhJ6pHcCZzClID0dSU4B2+P1K
Xo3ByMfnj6EqH70wHS6Z+CdHaOgM8InY0O0V1v9giMs3IBWivrDC7A9HMXIBVBWg7riYLIt9YGa0
p5vFyLdUXLsCYuRzpfg0ULCzyW8XuOq/woTiVhdKthMjQy8MsuVLVH5W4/XIwGaK1OO80kgiPeD0
6SHfxq8wtnsS1G/+4m21Q4b0HG9BOky2wDWczbJk2vxghXj+ucbkC54cCTyxl/2tsYPEVzSzicYP
t8g8fhZLV3zKJjDNgyLwbyzDioOszHewb03Yug2F2+SDNc9GCEW4OILxpGI7APhkkNfKuQ3JCrqG
0YMJQs3kxosu58m7kxBEpxDLaAHIghBamKHoq22YFtCvgRyDdD+tCV7CJ8TGZYNhzwayuzF+I/LW
49jN/ICz5XAzKD3DS/rk84bLlyhaq+jOOBovMBTNSOwCH5kD66jH2TnxRzDxj49/+VrNcU3iNtA6
VcW+6xScVjiiUyVet1O7RF7rTASgahjAc7k9sOvRkrJFnIJD4871oEPMjouktKYpNjKRCaTDJl1o
/T877tZs67mSr/Y2zCGL1ALDi8YERcwufSNIiJLpoU2L5zsf6+niNSkr4SSby528ZXxPuhM00Pau
G96Ryl9/q9TeIeHpwo+F6Mc+d/qdb8k2AoJvt7bYLTRlPQ4tzoulxkh7ORmE/4xCrXtg//Ln/gEI
Bc7t+GqgGZrj1FGOnEvxY2ZH50/w/MMoDiz1C2mK/Pujf/yJvFMATbCtNl7BjufbYWXicQ7h3mcc
OZT59VeinE6z3rYLANhd8p4bUoQx1/Pt4hY05WcoQW2o+5EgrsEst5z6Ycl6iXGlvXr9Zgrp7k7Z
51Ou9XixWHUgxLxo+KDm0PCfMKEVVM72MhztH/2ELui7H7LeDBD5IZZL1BObFXzPBYn+AvYvGacW
njKa3zPESLoqEQJ9e4DREcATNrashqxNUfynEqT0/o24qQfA1TBYFd096++oPQNCh6xLeIsbSAYk
ZcpDC5RqHi9L3B0h60PtbeDjeOJptQiG7xCFHkCxJW+CLgPkE8JWFBqFKGrZvUfwwAizKBqLInsy
X5jcmxRJM5gH6GTVnYhjHmDuwuWNz1nRFVG7sSo1HQaEp7ex3ya311etf4lQnas93+2yi8p7pCPe
IijbaMmBzIMNtbe4AwHdw38gKcBxj3YF9NtdouMiKaT5Vy9JKWXN4kM582kQVwhwtMCcZOMlC6Lf
tnWP8/SZMoM3j/2Hj37Q44BoawgnQ42asmlH6+jBFeDxZeYfkLZ9IYZFjNzs91lLxANMihcjcz8A
pq6cjKiSg+86y1CzdlOTZoV2RVw+KBvZgIUtqJdBtsBXADnk+pGb/6dGRobA5xuunsCVBIBI6Yde
Ltf2ebVkS5zzR/MKe3xpMsCxr4An0t6uJy60tGFUk536ffWhgD5xI85+kJwng/W/AIrR27poxmby
je2H+nbq8AdlGYK6ib6LXIEuv0uj8uCcWU+0WPAKcnEebaH7cUNQmbbT2muWq2Rk4TliwxVn6AjX
b4gFH9nP+O8FbVngHNudpfvyHWEzKgBuwf5So++H7mI5I7aH0oz9larOGqZRB/I4U1WWdHKVDj1Y
2m31CDhfQI6YCaqi7DVfnb0JF/j3u/9KpgYBit3+spBV3sVRTmg5xN8GNGK3hIYJcrY/9WtqWlvW
dCfggVyWz8zU/F+4ozqTYh2mBOeIJwAzTmS6xM5ph/RuRa2V2KNycsJNLevdcutmtvYy5ADCx6ax
CZ1nkr/1+Le+mQZb1VNWn2J6VSVkTK+tTlYeju+KP+5GlE3sw65kinhDn2zVcSjMLxnI1mgbHXvf
jgODyX5Vn4BrYTnuYtbUd6LOI9KXAFeGQBK7p+/zJQf8UuuNAhObOht3yVS1MlwfHP/f1zwEsBqj
pZ5nUSjG5ElNl1OWrISZPqUR3GJiBC0GelmtYHlAd3agdCfRi8V4SeKYz224Vcjwsu5MFVV5k+OV
Zzp3RMpQm55+ogZ9Hs+ZRD1P0Bm+JZYsToThI2+6ZYpdhJXJus05MwM4JP4/4nEsGGDPBaZT0Gmi
La4oJKyt6a9SOu8DEjEadl4Y/wvE3R/IcUpShcxFGWT3PCJVCspUlwRpry+5m5SFUm/1yn8WKneJ
6cHUQM2axoO8X/kGELA5LtNwzkbN5oV3UIajJ1Qbg818PuK0gE4bWU4gzbCutx4IZDUeWlO8z0Wm
XCk5RP26YwRGQuX4uqhf6prePcsuJEkq6gd4JtwDZPqSwvQrxh/sjl1uyoKpe5YT+2z2fvPcYVd4
hDmbhG9aLK2EKcftuwidolknE3rXIHycgDIY2xZSI7onQ3ScO7HU+wKbkrg4zc1CPZWTbEvplD1h
4kPIYEN5gnOS0jMrYYEK3sVfJm7+CF/UVjWSEwLc6NGJEe0xoFRtfqQYd9VbglZublvDhnXmpG0P
kwltpDJPXNLiMWpE8rqXe2dhWPbKrCk47yhB2dRiEHd+2No8Mg5WwZLTFh+hwidPUIzC36D4fPBr
ZZkK5xCKcilQOi4i5KMS/sItVPFTN/wqEoE4P/CQwCrUOuOt8NdlIVpMVtPWnbHGu223jZ3sFBIf
OJWWysR9Yfqe/Yfs5rIaFk0LHXQbTcb3TDS8QHXVW2BNxsYDU46Wpo9o5xVkoHwRQVfAHzBe7Yne
C4Bgm/6jjqCiSFD5WbBt0WjzhWu8+FvNdNDP6r6QfCtczMuUGSLiLYAnE3w5O4tlW7UN+p7HWoEX
rbjmsmwjf45gBKN1d3O1pML5CZjwFLdUexRci772nGGYtVXlvf9S4AvGlWsaT5WnlIL8eD+1Vmgl
DQHJ2074jyEJg51BRzNXV2hcUq9xyuykRAogORXhrXP1KaVNZsBZxcp/H/Qoz2Vstt1Rp3KAAMNu
zeQqSW7SCHjTBuFjxJKWJhFNcaocDXoKGwqZuV4HKpNRIdcpsWB2poRtpJiLjr6WRvstJVDCPcva
C1O5/P5aroJHfYL6YYyVSR278151Z/GcZx6M4ZgZSV367b4LNXWaSVQ2Ht/V5u3bMyDaVJagrGJt
DvkoEiNUyDag/xIhceeSOZmyT/prpFG9hJfNP7hn9XSrCEa9rgSFV/QSWUilwkY3Ey5LXJkHyanX
0wj/KOpoCEwKnP1Ny5K8ve3N3EXuCoQg4i56z0sRa1pmhRmTJTmaubqNcw4OlTR32dTWPpyff34s
eKAavN82etXqE4zGw9keZtdmpuagrNfWUPnWradStpcIWHikOsJ1dRze0IVD5g3ACAh+DaHYa3bg
hACc3t+0vZjgtg/w3oWmQQ1TRunO8KJbKFVHEInfgU4u9k3N4of/3f4ED3AW5TN+W22UJHg9GlJz
wNH/XBaG0FQHCnX5s2TezgNpQ0h+5Hhl+HLH5RBqck/FgqySUwwp0JrEmpvePuSFxbimZ2sIUT3j
oWIVcml7asCznRuozVmALz0zhFAX397mCe4gCFGkhVOM7XlXMUA8R2sRdyxKIasoqs5/ZLmdWO/B
RK3s7EmQdm5r+8kHKHS9qVw8ZMuyUhoDPjhCpbf9qusVfD18l4Krl7IITUHF/lNkx5DHt6nsQHjv
tOGykd2vvzmiVdcoELs8KEmVwtYJoVxil0hRd0imP5IwaDQi/UwsBol46ZsYilhbaq/8YKxwvhq/
q0VobU2Cnqy0dYUh19KDkbxsyxIIeS6Uo0XFMcwdYUTEDYGObIQIL/cmS6O128C9InBjAV+o3JVB
WgTj4vEkvUalhov0e4/wQW70JS22nw8c9YJkrYMGeJk8V80UWeiAMed0j8QrQJ22a1sKfVYicObJ
tJHlnMe5T7YYzvuFuJ20yDp8lytpwzbFdbeFScmIAlCNasjrWKsTpGjbtzu4k6k8KAfQNBpEfh3+
DEU/R7zQdFvG11qn774oySN+oXA21QLDzUzufyIGVv7sfK2p4orZp4VxNdYEujlAgndS51V6BxHN
clZR1SXbkNAR1guybT0YFg1C5Si1m87i5Yylrahgydw9WUYkDBgAk0h1hJ3pOY2aHtr4uyBGw1Nc
pnW6+W0QvhUrHa+6BfpOL/VcTnuNqH7+31QlNRURrW9vDp9mrA0eZSvao0feHeFaB8oO0x8K/q5y
v+S8bAxLku/2e8ml7x/jBzK/kGdrcpuTLj++jF/RvtNdZwGxgezYkni523BvVnHJ4vsMCh4d/nLF
2byYlK6cU4PYebImG/Oe9XTJ09Z9qDvP/u66pGxs5q6xIKWF6WIQFq+Y253ItZso6VAnlpmRy1N6
/1upGnxRz/Nfft1U+NJnB+JXXe1t6GEhGoLdcG+ZGBdDWKVgCr9oT9UfO57sk1Ep7fSBnYVcMA/j
IVlIWhfTRmFgKI5LXO9xSRNfRPtKyiKZRmuN3hQi9HgyV8iXRdu1knu/uR15NcPmzTYiiAJw72EN
I5OwBvbOpxb5bV3wuovMbQT7C7wVtSiZNMs46YJ+ZCTre7VVCIDK00fuegQpZPtaaJxtRKMpYwyz
wTWIaElCHowxnAFU7as2nzpNmto+hK1YoDRCrh7x2WS85nYVJE4EzxTqCPKeTxB/UNvrf24w0BkS
/GsKHM/U29aGeFAiCzyZ/htCRtxgvPRxoeYDdbbbJkygMYfkHztXQBhhWJqpXvuGIfBZxs7D7gc3
ylP56Z2+2RP0J2llG84xzWUpfmHVAbqRB6bMAhZ3asd9TZFrHz9lZ3lbpXL1B2wke/glsb4wzj+Y
7jEFbeXJd/opfp7RUZS8VS20393qFoAvr2tfQ4fRKT7+XVVpj5om4XBm8RhHUvMCAFvBp+9CjG7/
ObYwzq/MrMCgnRH4DVluDZw+yK0EUH4AagwHjNdllKtF5iKvHkTW4w/oD4NAOCAcdlakoClk91IL
rd1YBN6yhLJh9EpIuU4tKk9wIKbdwY4aBw6vh7/nOtwKQU6C3/EA5aQBYVl2HmPdzgh1FDrvSf1S
tMxw7QU59SjU887cjw9qRbqbqMQuwLs6n0y40/U7tZ76GQx62ZE66Jslk4ldmUqh0HIfXPTLkDBT
YNSXxonr/zZl+TNk6fF2cAFa4hHnn6oIIr3D/6ZhHSjiRQQgMI04s9rwYk9VKV28ZKVbmVoI2AsD
Jf/qkvlyxaspbvr/JEW/+QQh+aW/KLNWdOEBucv8xNw1g5u7JENjFNCGLtir0IKN3g7UXh6CIMqS
94jmUQ8aeSqYX6rcz8miLVC1CDbRzczCur571zsAtIEpHHO+faGkDp7rwth3IXjgrNBd6dLzzCHx
510LQbBygv8AVG4sWiq8o0Jzei4UnWRTK1zRmQaOUvpKF7DWRSLC8rZVPG0Mt4/2KTDEOQXDF3FE
b6+70cn7pkeW5vaTONbetvQF8hf80BLrHzPAm/rYOWfQus9bvONSnveaEJ/uXvQt0K369bpq6GCB
3pvLe+dqZtSJ4Kyskk7lUqQYIkMMXoFRO6nfNbTvXqLz7EtdlaGvQJ/v4oARaZHYPRQXUwEQGJw+
Nw++Hy2expEqkitMKzfHSaYMwteU+TfxeWnXo2A53tsTmD7SGZQZ/gTuNPVfOf5p1is7Guh0H4AW
bWGEWvRhApeOMSaLn4KmQ8Aapjq2Z1hPIucTgTAyJWxVsZKGgGTH40w+/OebJ7L4OtXJ/RGNdGvh
E+ErTiyhGAthRaWPHPart2hrcrDT28RcRIqyQj/tD1jKMVcg0c3mukO1oX5MxQCAqy7KnTUJdygs
Zfn39UIkC4+8P6eQE8ytu4ziGU60buk5WBgBnTrXS3yVuYuMbGJRzZPVu2h4YBcqSssRGkF+qzKf
8ojBsWvNMTzFxoT4S9AurVmIIXCqMyaLbXgJHMaerUm73/X3a1CxYedFEKTdQBfwjloyHLKXiUWT
UP2+Ei7esREikllAg+wei0bzwqeCG7GQu0jYLSx1jZsAsDt7bvLiCXotyzKmGoQwy2fysKSgs/r0
X8V9mWi01jFSWI2hbi+u2VGC3ZCEq2uGuIC/j/+2ossOL589yh8YO06ySPWWxdObbUrT6HcTEMM7
a5QH3bkczr+pYOY8+4cAWOQZFey8eoDSndu9AnnBlW0Es/RRVo7GmsLs0f3P5bPtyKYI7DvJtl3f
dRzq9T31FkphIzTItZM6w9zv3ZYn6nWJNnkE2ea4SpTBs0X5kCiT/o0zwxGgovQN8WdgFNdEOnLu
j5rfH+lP2LOPH7a+v4j8pw5nqtx4MxncgwCH+GfJnZrwqscDyIn7kQMhhEqn1yXI93Uipe120eOY
OBcnCIMS37vv4VaZkvMV5382MGxRwQCdQw8C2j0f86xjHmaE3aJW9rZBsJSDTlpQ1hyGck7/8lYa
2oQ/1Z2vSyOrdr8Y6LKer/paFsn61BuuGTYBkgdaQiqAZ7sYEMgqn8nlfkkW3seT9NNZ0/P3OpK6
ggga8VIDO6HFrxbdnTB/8AZvr5CqTIAs5ONrxccnJqbgenaOmAxg84b554qcca4q5mLXjZeS2xpP
fti9gDfvy18RNjkMlDzBmOl4whB0axLU/HvKTKY1GCSWtv9qptuFwKjS6N8/mZf7eIA0/VjiB/iF
iOhjRnEX1Py/OH2PMCDIILrkPMS95asFA/+UEXZgtqunc5BYeRoG+1xW+XL9vx4Ynhtxj9xa0mDk
zc8PACOu1eXD614SmVkN89Vr9NUAXM15Pt7ns8fR6nm9Rk4emI76t3LIrP9AjTjEXTazE5il/G5/
6jBa1M8w041bsGYaN3LbOQUrjL6iM4DQRkk+0RgZ8nXmzl3nxfPmR7irWTLTYlYEucdCaZsxHkeG
w4Npry4su9f3G0Scfsj7KwbxFo7tc8+ALopnKN+ZdI7nWXIM1QhNS0o9Gu5RS6Jj4sszS/v/38vi
eBKO0z+Ba7JHQL6ExNZtPKLX2uu+A7bhTwV8HC85xo+6pZHE2OCC1P7zEoOlL/xqfCmbhnOs3w0G
pijn+McSQ8q62zG9pwhDNgtqhMo3gjy3iMzkgxq9iJP9w5+HkbmVsetSa2rViMGz3UNPrdyboitE
/wDoNxy4N+PeDuJgxq7F3Asr5TGM4i4vJ9fMkeTLZKwu9dUlSPvE0+R3U+Dih6ou22tlwJduc9Xz
zfILQhsilafvUJHQQ1t/Oy9V37heZoi0CVUfYEGSA+iyGXmoUMUflCs9EFUHl6RZzgzDO5bRObQD
cjVipqDjwt23uhCgIaHPhjvcMjG/f9AzKr58SY2H7dl86AO7kw1l/cSuJrqBXivt4vMb9c5GmcgD
JkGtqRQBmeina7jWMaYVSAFWhcYUKjmiWvOtJRDjdEkeiKhbDUiJThj3xoOlaX5fzPWZ4/AU6RaX
j8BSfvXJDjidGbXUswCKH8iXERWFZ/ZG6Q3XQesG4cW3jCqVtLcZd8IpLDNJ04T3OBBbxFOWFhI3
tI4Tx+oi/kinKLrkVr0juVVRWpE07FKgb996ap4rGMjj4f8Sf/oABsEGA19ryxy1jxjDq+EcBZro
z9GcJTs7T5nGR7gL0dcD6kuruxS00YdnsL19YfpAVnya8l3/6vxc8SBHnBEy0qwXm7u6xPl8fU4m
ZYVLLhC04aB9J94knPjWdXFDdrvnO1G1xu6aVGKgQUU0dIi+ifQ69PwQGEhU9CdzJgBmgfJahWrj
0V9w+rpYdzyj3sUi1hPnLftg9JdU28oZ5zcpWkKDzE22vkFuDoF0wAV38a93Sp7tR+8GWz49/JPB
e+lVl4e1uE2xj08aQ51afDH+DkmPPVZY8PRY/1GOyBIFS0l5h3VezyIpoSffxpfPiEB5Y5XmEqQS
R0OHCehWWYP6NVxNd0oaYjDyoG/YnN8foQuvl5VHWbrHE2OtrxJ4/XeytMqNaoHMDtxiiYBxv0T5
QroCVunSTCYVrWNTSiTY20LMTzmXNGu5x9XniC+xqxU3CJDYmGwnymky/A/czAZqAJux3HrRIpTV
tVsgZA4vywuaK6MdnWmsntDyq9RA7T1gBnBbELeejII9KLqGU4FlYsnp2JP7ihlcddGT/GXkgHcO
DrElXaleHjQPogEourgsmwFvEscNHMj+pFDi7atVMpm+PMv3iUD3wohI00K5YB878GcfRcdHnx7T
mi1Nh7Of+j26ghuAfu7+NItOpgOZnjPRannHvE1LG7rCUbLiD67Ruqj1TgPeaFAsJC2plPFWhphf
SAfO5w013BpKb3wc6E4KeDTQ9DyVOBpUxkbc5viAAIMfStF6VaYLKJgOE1v/oX76DwYFN7biJszt
5xUFtUoPTXaB65S4NQDDmop30o02UnoENMYpfPilZf0lDFrwAtMf0/pB4qVEGdACQWNCUbF4EOU6
exQze1qWmmZlGkJ5r9MrcpG/01vZ/CkPW1KUpIaj5dK6d03x9dGrZz8oxYfawTt0nXziMx/PC7vH
SDoRCVbIaATIaowz92IAWoZK2kmQ+QJqbvblzdJa4VCIKKNovey0msSKCtaQWQM1xwqtYv8un3sU
iJGa1jJwD5bvUoAAA7YFfraIB4c9YNAZjZ3qobA4lqNVAd4jBQxNogMIsCbF4gsfIB2DCAoDnBP3
SCQZzTCCgJQ7vf6r+XizP/NGaHfi/Iy63p55vNeNBUGNqEwtu8gUsq1+X0Kn74xgBEtObXG/rsuI
o6GnS5GzwijXFWrUxHHkb/BhVET6vR1o/K2staKRsdH+EsNCUiKbtMyeugXbubIL5DWcctmhxFy8
TLlBUyB8Zg2lq0fPz1tnT3HKKSR/+auyO7wfexmGeJa42klr8mwxRiHMt9wvC6PUu5f3SDgYAyh2
StCbz/VtCqgzaXrFcr4YUdcRyrIdiek96fdS085w35Rti3bbQJ+STgB2T9ub9nLcVNNFmw0bWck8
cdmKxj95GNwr9aE7sOBYY9ZO48WOUh1M/GCPTnlEMWgfgKG+3+tfMcGIpRUXayQlHVGThAvsPTH5
qtAVF3yjqqk3plWZ5pebIwH1C2dywksLDQC73ijCVRenBYZi4lrBtxeP+q2Kom7JJJvMMoBlq0fA
eccRESyCFO7gda6ggBfpJ52oyrt/sSCz3mySfVWAuCPmNmQYDhODAZBmrKs+ZBP1GypS6spP7jtQ
lz79RqPElfvyl9lqSf99FFNkx33TYQhnW0NwmgQu2tBw+6U+MxxoPVVVdIQCt5r6ILreYVNlYECv
WC4/bNnjUnvrGX110RY8mHaS3BM4/QTHpdDazF8P/ZB3zhnVXtEQQgqA/ETk9xrzMDtgrYZTqy4x
LRxmKebrO/aRjhikzhJp29Y1Q3532XLTzfKjxhdOXWseiaW30vMr6U3q4I8R6p2okKyLFi9ch6xX
iLczGil8DFawJaaX7nBUEpsi1K8tlmNE0IKgS5ifPHTSvn2vyrJKG866JBDPzZNzAP8qIGAQXfSf
FucD0Y8T2SkpXKEZYRhPWj9qWtVGp2/zJFJZCbtYKD5O4OF3VLjKgmAhSBuOxSQ+xebpcK55ku2y
+oOX3R40iUHmXfeJNk/R5McTw0t7oI4v3pTEaW/BxfPe/G2AqCvLXaa6oMadGFX+fhQGlN2I9wrh
FbbtxuUL5RCr1EEYTflW4090VkeXFIDrZeK+SuLXZElUuOx8xIf6w/FRib2wQ2oP1O/ki+P8xICl
f4G7iTpvPbUAHysxheubYWMzx2j4+2sMEu0Ob+oskwz3gvXYvtO9uiaNaerXVg7fUYPe1hGneFd9
UoHNfJsBbyCrO6xjhaAZQw8k04ituzoNoTyKmSCbdR5H659BLxPnkDuStwvd6IQJfvxMPcW21K3u
WMdikm6Wa0fZsSVSmb7rFgdqufkCh2RBvtQHwRy708DLq3ju/aYTfkXWoQu/v1KOK17rfctf2qM2
qJgjw2ObkkK5wtbARxLZAN6vkHmvHDdn8owhmTB5+PGnLS20liYfiZ9wTep/wq7kAP/mohkVEGuC
0skRg+xS1maxmTgYTMeZLmKl3Q/otpz15KjhS9xJBOIE9gauPV9FdDXeqrV4O1xQUk1smpiKlxqX
8ZdZ+DcJs3KkPJokmExxCoYrWxvVx63c1B6mEmt1Q5pvKIoFltc3ZTZhs7RGL6NQ+r+2mK+7fISD
78zBPqaJqGH0zKGOrfqve7/JmIZY0KkVHPQGohBHaYYLujxFg7R5lLQDoO73GLkOEPEAH5LhROo4
pWIW80ZdPiGpe/BWCgfPXz+QGqabJbWwLCMpj/2Dg/X83z7TJ+AqUsj+HmVqHq2u8fuK2DbudwyI
dMJCDRGpw6qqayEEbH3zE231sHOagtVygmAFoV8ywnTDbgHkn23FYe1Degh48zdbTmV8e3s1CFeC
EwEKQRVAxRwm4khUMppNdK89Tr9o65Ct4FxlHHEQgo8S44f0vtuu+ALCjj4ayAdFsJBMMKjN4974
RiDpZjPNVHNT6Zi5xUdQyvhwQE0YTRCcDSU6lV7UhZrjRSMK8UZJY/jY8/oDEKdhMPN9lyfOgyXs
zLbo/1ruADMkmqmAV3hbF8MHYze6B/Z8+s49WM94StDPQFvbxrrc/JFA3yjXZ3eNpRwtzO1TLCd3
MIVIkQbtUkDgBajpu3z9ypDRvQD1QLw2Euvoj7aCKcvx97gd34SmI/b7siXs5lwC9Z4/ZALsAlYP
SkoRKs+9cJ+aDzW7rhLEMchLppb1Cco88GJb86V/8bcf/mO+URv6QeLBwZG+VKhA0PztEdUbBhmk
13s3sKXWfcG6ucCjr6mRSuJ3LCizV3m1nS+g+ytsSsTesufrgOf9a7KDirGGDr107xZ2D1J1bPTS
9RifjU2guRmBwUXHpAN0l3Fvy74WUtAbcKXbDUxXKvumTXfnrVFrwXau4tMvaAaUjLppn2u7If7k
mSdF6CEz3rZ23RBE5bLCiI7Lq+NOLERvTHrU4I8tZy8hioXA5rYOyr7/xgsPel5RjHPXMbeJ+Wjt
dtQ03wB2gaewYg5sDEc0mwJA9xsq1MwawTG1/zUkJtsO1fuOg69VUh7iScCoEkAgjM9GUBHA3y0p
V5Wp38gXrdv33pk/m0c3OYV5d73UGkQxBDWfMOTRH9+PLdZA9vDF/d5y+Yr0AibZI2x/dRK3VsAX
TPS/p49/JIWWzdgcSRyJ/G/IKNrnkK8Ea+PYxDjtTIqYx3JntlpN9DPArJkA+eoTLSjr2XmvUgOc
F0WTUuE824IZJbK8n8iL/JYV287XD8zyCiyPreFKrp9RRfJ2espROO5tew3VRSu2zbO5cWoaEQar
8wCWePr7MqJtjQP7ty4Y33lrJE28pSsjmPclLWmEtor+9irXGHilyz3TbS2Jc9/M+wfgf0JYaUtO
GzrIcYlTZmAns5zpMoE8qdtEzpuhKC6FzdMLaWm0yZ8knT1nvqZ6YiW6eN+mdzGFRdriIzLEcDXS
8XQViOfuAryyYGu+BVE69ZF7wzkCwZzCVpcnrrDr41T6+MH2h54niR/FtCFp9OYRIlHiuI8sf7vS
2vfQysOtzb21k+qznJLFesVa/dLoSAjoEQ6rbVqdzHHecBVtsqXsYaVB6t8DR0OR9MUCPueYOiBW
sAE0dCvtb0mCnvMC5eN2sFmEKxvQ4XSP9YVwaMEhhww9oMfb8phjY1zjAvy3/RPVpEhiaK5JFcmr
WwmLZvSatHeJn4vx6ldyU+Ddlf7ICLUHAbJ8Vvr5zPkCKfBtRfVUbXDbxoaIY54r8n0SzLKuSjDm
0y8frVMi2GCBe5HoUFl+QTawbwWP3C6jQwJ4lmvlfrijc6JaVoXrMkpn4csZRbsIQGtnWk/FkrA9
/J8VxFatgLWS/l/4RqKuSpIc3A1fbnKUYe0BvnPlOYVAMQBoHO0p0e3pcUXUbrl5YNdyueOx0y/h
s0+YtdjePndHf/FpRJibzLL/iRvjxojnE5/VORf0fzJ6sBxwL/3IURxfH1YEyRreoHilXTBI6+cK
rDQVOZgEBoWTmU/L6ZCzEYYws4J6c5aSirMIL8+q4Q6ZI9EhlqPStgqbxsL1UxPtpNQBqGyVoX++
FljSWtWkM3Hs5vO57loKI4GQtPuZztaBZ+QV9Mecoh88LmDoVofWzfg/rIJ+yyZjFXnuoiv8Uz07
450/jx0qNLNoFVgt1j3bFMZSPZ1rUMPrcOHWpIlZhpU+yXyMEpgN1t4D7cDNBuvjGLOOzbQgc2ch
NvaFNGRUooqc3vtHR6WGUQHcTK2hSaqrAe8CDFjWvyKE7QnxNKtcjBzFtXeSWmiVh3aVnO0XSpjf
jsS3kzXLy0c1mtt9WAwBxv7ir7+BxrjwVfMKFOgZuqWlc76+5MJA3Ps3o7YQJrjsMnq5byLKN3C9
u+ElAh2KQyGLBH7fbGdPpiAttjn5vq3tLvxw1eR9JY4OB4ABApB4ausrqLj+D1wmfq86WVckr9UP
2jp+uc0ywRzsVkoMmzTMiStH3UzHsHPJPQUzRPSf3mXUinnW0cEGm0wYLbKVxA6qrTEJvxPhJuqS
R55dVmKliobsfJrO6njtMPyTWxjZFptGTbuT0A4ygRRlg40Zhcm9H4z+pXk/Tnet97TIqXbeXdqK
fvxoYqCAc1u3hmnWShw2zj1uwkhxavpKnSxDXw+/Yeyp6h/myD92aKLj3hJn8DVimh+n7jaiMSRO
RXzZvyrpEJHTyxFVvkcHf+Ns8Hj3HSKgTQuluzoNop8XJePuBCeQlnO0x1qnk0at8ry/5VCmQSp7
pPcu76/K0ejYLSHHKBBLtr77jlOB0O68GEjGjEmSXhz+J4VEbo/xWR2wLBsN3T3+OFLa53mgwmWl
iuYHW3/SBixG5zoEo89xxYaRN+znHm4yyUh6xM2EWrbHRCYanHgz0tgRh0MUpvnfPJlhnODJ/NU2
y0v17mnJalZIEq93iNdr1RmsWIE2JRhYu/AV5D+DJLgU2rQUocBGMS2tG1tDc4Qibq9HuqJBzCWu
wKmNI5RWddIS9ZPqLwpQu0NQuN3BPyldMcE36+y4D4WS+HAxo9oKcO4C0A1glnTp8vuWDGxNyKSI
87NcXQU4dAHs09wDsVtNAgUXwpfqnebBAysPDyEx039goju5eCpKFdUG4n5t7JSm3TtuyF99ID9Z
eGvr92mUssakv0VwnhOFNJ65lRcLilymEMfWZQoEIkcMgGXLBovuNy7VykpHT7c44Jsl1Dqmm11S
tMFnLxM0VrUypAEjVpmSNqRcvnm/8bDYs7Mgd1Aivsl+iLnk1EV46BV38OXY0fKHo49/a45S/J0A
ZGUsPdsm6OilhacWECcfflR5/dAHWLEOjH8IPI5TJ0EFjxO+0rzrHRPtKyhZGWMKtIFPODqDMc3/
ORCWDPIl0Q/CgiQci8OrJU38IzjckshumkJy1/pvLqYOj1k8nujizKYqnhqdfg6MW900ykIFi9YR
5Cne3B7m9ZIr+7M/dXEQ/x6ClzOyA9jQ7GBIrrAiXMqKs0sy2tBHhpmBjIfqLX8nMYGzSczMvjFp
E7TQ4f5wTHORp82i0wxUkmvfr5rZ2VDRVysgAtPZTIaYCdqy5K8gnu88RxgNwXDxy7FNYyxTtGrK
UCpn2CvoFqARoO9GD2qQGD/lueSYeDAg0HZIk5qdMsRnbCFW+9TLiqlj+ah6a5nxxVMdZHncWBpO
kiK5EO90F1iKWomYTRPyz/pe+gnFMAJ0/IjJ2mWTXXd90FzxPkWdaH5AasTIbMWISHZxX3U8oWxQ
hYZG7C32gJrfBZALIiBLB6G1781mwKwkY9hO9igbssvYwr2NcIBifNHaYc84tqcaPOWXWwwe0Ow+
93p6T7nHmnaQEbHAHVEjvnKrmb3vSxIkWyypjOASILQ37ui/claI/nG4iAnyduexvOz5bZzg1kLU
kG3qNTff7ulmLc/NJZ8mo4RZBD9VMpuJXTHZvX6OYsyeRZcSPHB462kGsH9gLA5UjPgotfl86o8n
UczwRYM8NRmU6QO+EX+M7iQMBM4AIfSLf0fkVsM+NGOBWTJUtZwvwazI30yBoDinmKi9hSnNNEma
/CrD+RQYKKspMCOvuDiGLwtPg/g38u3jfqTGq/IAvCyL4+Gr8OfCczFX1zmIdCkmxLnwtEkS/Q0M
rDKeNhgQzMP34HMb/t7XEKLWG+pdVaS98wkVjemgC4kqqnp1pKLQIjxORL5ADuWiOm/H1oVBrqtQ
2SKuEFwUj8XAbXtDnEcowz4sHPIotmy4+grKPclf8LirdX2V6I86u5qofRA8TEHHvD6xVrJPflRG
AZw6rp8Mx49NQI0Zv7vErfKYQXMOAFHxdAWiybNQi8CAEkaCKtmT5F5F3R2kBTnR2BhqEaAeimc8
2/1grjB1RXqylyOInvsIRgHBkegyb8zO2JKKiS3giu2CQ1VD8Q48ETCyzJQBG8efJkdIf/9bgKJQ
S1SeUEOgzVmbzZvG2U6NoZ+lOwpax784xP0i92BE0GLNGOSUm50XakJQUIv0uFCHfFY3OijZwRvu
KeQlrHo7amRm0mdbUTT+S1kv8LQJeyF4qbTHTCvxHezbNFBw0YMNRmV5WxzOyztpBD9vmo5CjDzi
MKuQGU/47a+02VRerBDanVEwa7sfAHuI8tv6qvieeVO2BqoWQ/3MA2SrzevQFAVT95GBR/jd4ZWQ
8enygTpbo3ujBaMHujHJWc6PhHu05xnWtcIvOA00wJafLep7TdUbeuLeucymBdWVDAzILtG5EmZW
4fnI+tOhCgY5Rq+nfxb8AKCzJyTsLgNo2wDC6KRjPaV3G3vKinakTWl7947omh02o5xIm2Gab7z/
UOV0CLh+c+Z8FTDC44Yy9ZkDq2ZITKlhgzf7NkE3W4iFdxwDoVeus1mxreDnfBQAA/Znij6jvdM5
iKH+pr/DEBEizH489ZtmHmN/6EqvKiFPW+VN4VgVqPuxdk9wm3tDJstlSmIKHdpZKlCPNQ0UhWwc
RZgqsoKjYlXr9fCb5BA0FmWNXh0cWd909wWmWJI5ee1i9rUbtvRmHCREYpzANuJ6VQyPvn3uCGyI
y1h2HtCt89FpZjYJG1SaEjYsZ5iV9AP1GpzAXcFEdCu/Tds8zAc3JeU80pbDHgoUmq/bSfs56Bzz
TsUnkGzJlcBx0UWsfSfr11DpfSQaGiIDWXiQY7TEeU8pCAoIyxhAAc/ZDaShzUdNjzsZ+Pqt6rw3
ctgkkENhQkuOaOayIsNIDHerMGkmKw68uORKwICarc8nPWsXWZqocHuvX2XssFGvDfA9m81kugn+
N/31LQyhosTqtlve022oORWIIlBM14S2BmnNnL3+9uXp2wRA5dOCWZYWj6XNF337D+hUkO+L9OPp
8Wc02xiO0q1PdNu9S0VrjoSSp64oeNTHBqXAy3X4CBcaVxCB+oaVArSD0IaV6fBJ1z4Z5pkQZyAq
zzDvQXPEwk2Y3/7ObP7iqbki0odRrwN1HOhHw12pVYOZftMVAYkvxP0l5PDtakMNohOkll85Cb/X
wgr8k8kNl55rcy1JoCkA8RhegyVz1TULWHpJe3QUR8jbR9muyv/rMOJlvLA398CukMKbtpxymut1
dI5KnXGHkqT1B55Ufq/C14QEr8akfQmzzNVQzL6C7bfYfTIw8BFT1h3+PjqJzbdUbVlsq2fSQG76
s+uLWF+bYkMoBxu1vxqZmriIy+EFwm6Qc6FvzAO9mNa1KiHjHwwNOcpZl5eSRyL1EZR0KU5fJclk
aIQ1m+V22HTTo+azz3vgBIUHUX+zuIt1CHFPTICt78e2sKhSvK2DXQq/bV1dn3HHtvn1koLKSQFz
mVMFpkBsidtJ4VABrQvRmYwzjtwEiJNMezeoeXwffdmhx9B7LE9Vzp3ghL4JHeh/t2/FvgJE+Qck
rcZiaL/8K8URJmV0XPeGjumTn7ZR2Sna3qlqMck7ArupnaGELgHEd1t7XLXuF3nKSird7cantqiI
t6rYS+OFmtKufOWluLBuUfPJmJ7xFkRbKp3wCEj/pvNb3bcuqmSxKdDg2uIahM2zggmrmvMudy/J
V3bGL0bmn0BBX1Tuy/lGY/QipIc+c6a24nJVOgqdArS4AIQMRD23rDuS2t+6EiivaF57IH1skkyV
8YXvIrJixLVqchCXDYd6YFC1tH7VATNL6PHRqigHoRpm1m1ReG+JWZW92kDWQKkMHGO9l9kw9vlL
s7C7nK4V2xDlhBJuVQ2EWLMCpfxoojMBS0PvLY0N3a8hx2UIiX5PUxPwEXro/6jrIbJlB/z7GWFX
WGIvncHkCd0JqDjS85/1H/dyNoN3n2VNxIe35YvXgja5atLrRmu/zizYivpl4VWGyNuVbZrDpIZh
AbzarET/98IVA4smhK+Lt0lhTdzsWEyGbkG2V6xjnfrXwKVtWj2xspPMCQ7pUaUHDCho1m/3WqJC
iySgoLLQiQLM3LkoP4LgmXbev0IIiILyu0NKQ9BQmvGm9DdE6JbAu6cq5z+bYin5UdKcLJ02Rvzp
DmoUkN8xDoXgx1v0Ijrjj6hW4rfaQ+u0eZF1Sb4ppyl5Cmnmqf2sjTxDsZAiLQ+JDZqHPe4ZDkHv
0Z5Sf8tS75eBqEoMvY2a0GuHsueqiYbj7ZP8TqD/NKnwDQAuxepGpV1gPNB4/sX7tWqR5arO7loo
ph5KkBEfFES11XbSHTL+WFTe/TdU2knXxCfTEF/btrcXVucajF83VPNEs3h6q1MxwEJjDpeFdqze
WkprK83RDmsqoYDl5mjk5scaONUHvp/qPaWy4xUT3UJgIwlpYITmL3QlfQ5tEqe+fRTgHCsCnA8H
ctunuu97G8ArudpQDPD/abPXfo/cvnPXacSZ9WXyZCw8fB/vq/Q/i1cbDWntZNqnMdb46SaIIVy1
Tw0ZrlLqartiQ07w77fW63mr7J8rJU5d98XN/Bl3qdLd7yuIxYKVpH1+xapSP9/8ZsTtzSVarU7N
za8EvJkTnyc5bsBbuiTYww1Wx2FH4JN8zbzzB7632pWoPr6zxxoGW63GpZ/sq+E6q9UplqU6uHLJ
v31SM5rGG0+3owsLTC85yGugC+45kf+RtnD4FB+CHmYpImjy93rttTvK6GqymZSkVRCxI99FKU1J
GvpDvL7k+no8MRCCnQeUb7w36RbSKc4CXVivLGSmIBwZ7+3q8JuhZo/6YQzCMXERaIiMBh26W9y4
oPTqUueACX+aGobToD3ZbuoCgiPaE+L1cDcfwodISl69DCH6XPNnm/lES2cFWsctBJZ0wjEnfFs1
CyTz6KyHD0LZGCpA7XkeY12c2yw1LKDZF5jlIkZioajb765RGZGW58orS0Fu4g/YXnU7b5RkXiiz
v/5EeJ3XLt6RZqNQx6NI6Om7jjXv+LJ1Fkiw/Ttxpyo+xw6AYPv1JhpLN5MhPnWBvgDQ7o+iiLBZ
MezMqpVyyvxV/uj6vyyNVrZSt7phCTbZhxmPtedvVYWqGfuolOasH2B7muayyLvuFa73wXoQ9/w1
6c58bm9aDzCKvPHKgpv1uW70LCwNTbzQ5gz8u3Kdi59BxDguvPlvbI0mnyiGbITSAgk+p1Wy9bLq
xn4m/8eoFVVShg1l+JTELX/xBknGNCJ+11WPmSZFgW36wqZKbOLtQwva8Z8E0iDX345Z28/pVAoX
JFKKpvFOpFZW+zTRzWW8B58c+PyUeUkPNOszY5oT6ylkN2KJzSuVmCd+3R0H2KhjsJ5SAheJqy4h
8cSq1zAisaQrIExHXHOpJrY7QVbfVP2Z/e89rRSi0GzVdJ6wceGp/E7GOpEQOCKvCTGQRTzQhnt7
2zxWxAkQbUE/fwgJ/+Nc2PQAPmi6sKBJtAPr54+w8wtjn8RPpKgI9pd1qjvym5g6t/+6O6bNdshp
HR4l33shWI5FmsQf4fJggOr8QfjJDgH349rGb2vyoqZrw+/9aufDzASlfaGZuVhiKjPTjFUGd6Um
LiRsVsGLLjycNW5va+2Zp26twUtebYTNh5mw4C6GlO1ws5+j2bNStrnfUQ7F1gAXod4U+Fz6b/V+
l2pXR+Gqf7/wh9IPpXOhvaRFTDdSXxWXBLOMFp6N76lqMk/1bSwMHv6YtoDig5tOj4ct3xg0nbvg
u5wvQYs8tFY2I9a7jnRAuM0narBGW5an7uUN3eK698fdazhFOGNx0r9q1n0TzEwa5Ki41gdVMAo6
exAwusfXIKIgEK3PwYo169v4A9dMNn6HbfDGqj+qdyMS1EKs7oChxd6EQl/cZjOQoHa4jsgQUS9X
0WPo/FoKoIE5aapmpUD8KKUqQMYzn6ajqGZhxI3xv1fHUDGKGR2aaSDxS1V0xlB9x04f/z9cmxH0
LKDZLrvs3mOrQYCa1gag3n3G+73IInetx+7xTlcpmospz/2RKzonjkZILhHvZorR0WBSn/11J48e
tSzQdGwVCs03TmQDyVvi0jjfRbUNkBhZqGaNFwqp28LdwVdaxkbowsJlEG119U1ePU0dSMkGNxgX
QalTL1pk74gCAHkNN79sWENqN0nySO2EQ2uWcAYes6sTUxCSogNsx0Rc6K7UH95W3XvM2xVjMgnO
Gf/q27UXwVg/IhlcvWDwVW2ihiAOm3G8mjqWy+wC3vjPcx49nK16I0N/R3sFyQYHdOiOVYaRpY/M
aImoixyLitKU0dEOs8DTfvAIEdv5/mkWxOba+7aHd0bvU+9gWsASCxxrP+PWiF4X21jvfJcQ9xlW
Pw10bOSZf4Dn8QHD69etNBqzUnB3lLlas5x25OF/F2GSUn3Oc4H03eZ6d6Vr8gjXTLMar4zPf80G
kRRya3CG5Yx+mz0ft9xN7ywvBUuVdiiHPhvbG9arJHR8dT9CXO9jP4UXbGyQWk0lkeAlmjtSwiYq
DJfXGJrTFt0NsAXnny5iFkZlTfHOUHxECUe1WNtoNr5YuRWIkjYYKYamTYhzi8rSLQMqU2cGswM9
g42r4dm60xR4W0lGchlEDOVEXVYVvrzijmE/TeL+FWBk6VP9xzJaMyjsZcEPtthMf8PptmFu63mo
BUf9yzo2UGtuUP1/tfGVgHCsXG7ez2bbaqQtcYyg+qRxPFz/IDA99MHs7qciJuISD3VZtrg9BeHj
65Q4IU7oImA1uoYBL8VIpG3Qa25cGIEqxnIZOm0h+ZOWxbWabzGZWsLWJRcdLQ8mu1Nq0ewEIoRN
dj46U7J1ddCteXLZpXjYzol2zrK7tdCLKcktQyiL18vP0SBHLkN+yE7kCUMtt9hxJ3elObASswpo
YgUEKZ35vsCBQjQ8e7Gi9wiK+rX0r43hURJlT6FIKnl2Qofyd8Oo+lgIpMSTUkGTg7olJ4DHwVci
pOH7ivv0R2BhpB821wnWGUd2NtcpYQn72u9vd9ZHkdgSZsc+x2vZJY7blRkIPzE/278J4xPEqDim
f3n7nT78/9cib1RL+uTUzMZX4/Fm+FhlWsUP+OABlbA0dGSl6xTPvMznqaZlnaAUwvZENGgFEgdc
ap8l7FMLX0DO71+SK8itySuRzc08TVlQPvUytDg3EJ+mtM5sH1RwuWX5KoqIA9n9vdsy841by8bP
ld9lb/8pEK/HsOJOu/jqkl0AXzfMOEGtqIAEYmDVW2GrobViS4JwodTorTUmU/PMR7/qbX082uVP
yXkPHLapsINbTDlHOONgN3GCFlZL5RZPsCzausV/ojqbE+hDUClheceBdnEr+J/gQCHzhKU9/kUT
B/tVD7aTANHIYr4yah8ij6t3gOaZAHxsoYP8ElKWrRqVXNb4YNN6hd1oq9T3oXW8PLAmbZKlVcX7
GYQobBhJZyM2glJikXDSU2Z+YM4Su46nDFrZZplxpX/u2bWZkVm9BYvclbZdR2/1sQqM4VEzJSWW
meTqtpaOmxvw3phxo4nfPVLg092yJ5WKcUqvC+7LiCFxhUWvaI0MnpJebNnlhs98cd5a96olRUhv
GPFUXcs4CzN/Et8Mi6E8sLJOyXbrQ+/RAuaWh5T300z0dyemKu2vDOqk/usfgKoFJq9af1fIHlnn
JSFpyDJNQ3iyOtfHlLbIjneUCqKFLcwL1AME+/QGXk4CSPEXwZNp2g4hfuroUK6gNBXKFBzhmZMH
r+EzxXAacmWKjMofCybvyC/H2di28yn67oELUJV9h159sxdTm4lvVkTauTjFcVXrw11qL85TxrrP
UALfoGAa/Z8G31bnioPkupzhp+LAse6MBmB2WnU5ETO6tnGFxT5KC/bwDKQqU/kbUjj0w/KP8rj8
YQux2Ll7MOOrzI5BZxJkGMpfP9akvCjpox6drSZw5v9lVSNn3Sk7i+mHABgTB0SaTUUqzd7ANrKm
14+FqJxWNP46krRDNxbKGwn3YQFO2CYc9UhdckYOHr8mzIN5mkdwHXF0cu++hnBINDTLQZtKrb4+
zZBzQgfqmUZ4/Jvn+lr1VkuqIAUdsFzJ9vzqgZyWxx0hdq/jfridBgew6+n8i8chizodEhPn6vGj
g9+k6IED1W1SFADGYLkvXH8V8nFbWQFE29r7cQKkx5c97IdGWrVCjJ4pwKY6AAo1vrOc7hosqnzs
a4h//XaXP+1Oo+tLwAq3tHsPEoZIxnLEhFdDVQ+aGZDyMny0gG/sBsh181CEC0LlfTkE710J8kwj
ZQvtDdtscFWM93scItjl9qpmxMbQIi833iEO29lnCO+K4MhG0qTRJu4Kjso8HTKN7Sx+cEBO0DM9
ul3lzsWOv40JCCrcbwOTCtCPk5GtPT+Wq9R5mS2fsLbRtu5Yphx4r9jVsePMaWv4CrGD4jp/KBWq
mEECm4PWcw1xbz/BuTujqbf43thrGmnq+ogEelC4aINxVDGBkpFtNwm68E0z5BJ5FUEO9vzbxpLd
/L0bNot8T79X1XE6N2QxY5amQT+jRSUpnFsF1JmuAphMtF6zSCNW6e2axAJiNoElggMuRIp7p679
xDqn9ztrgRGCUWQrake2lLBwsBExlZMQosO7l+I9vx5/Elj/4pZBEdQhMWLkWGpymwyn0Mvsl5uM
RTY22SztthF8xEZhwhIzZeWmdMhC3bhdJ9IZDGv0HyjVDNnVMD8Mqe9tU6Krp88LsAMU50ruPnGV
GWXNzMFEHgzEWTPiF79TjQosp/mKsp2zQPti1IePaVCO1yUuZ8FPXXR0MsJne1BuF0BuYV5aPuEm
JQsqVUkX5CFhRXmgdBHnSqWc0LTfVdP3Ag7IW/EHgpEDltSwHNIt3oJupHOL+o1WPzvhLKdhODZz
H7bVhdWM7saf/2r1PEcqMOivFsMYB0EPRvLsAV8jUAzNUgNZA2CKwGsWLFHCWtYOO495nN8r72Zy
CwP141V1PHnFnLIYKSf+10tvpwhMocUZ1FKYhp1X4odHIEm7OXGgl7D/nIMXduNmNJJFS84czlxn
XnfLOdVcVKZcSTzyPn38pVdg2EFqkRLakjozIcHWGSWZo8xYSzuvAZWDC9ta6s1sqqGs84lK+UpH
E262N+dc9TMjB1Lk+N9e1iYMIxXjeHcEzydXMUWFh2u8NjYGSErzL8Kuag028GFDX6v6rlvZ2bhF
1emKOQXBArzqiI+X6N1HXAmu4H0CCB8xP+e0hh2Ai8TqWde9OwxWEYWhowOFLMegf7rllyoZZ30A
QBr0/1vOaWkujUr8i7lpucInUS1IgRbra/ePS0QpgvnjZPg+SzIAfBLxMJrubE5q3C4FIqWp68vB
rEV6X+i+/Ipw0Jk7OmeF5/AeLsIr8rrvfVox3ycJh0esOiG5gX/1TFwI19uvGypXBPVHg+wB6UbM
8o7fC5UODxoKjcp51aQDlP5eiSLPyA1aRglDJwH3iddOOWzXZnePwtbhxrdKPgX9ntaLMlNCGwqy
joTZZX6pnSDIcTldEeweRw21i9KKs4L9Yxq68B1KdC/oCS64dTlbhrE6C29vXW+CW9k+4cQ0+f1n
LNiPprQTeZ/NaWgKN1iftW0r6RBbHgKf1Shl/3kkuERRfed8p5XoSQhtDK6ch4OITnrTZVY+gg9J
yrJqYNmo5sw2HdEuic48V0+KnDSOeyBem/2Hr8xbT6rWzpH4RmoGsq0Zy1KstGRISkBLu9U1VW3I
VjbQ6+LYTEBO2AAyUPzoqrxOt8xlP6of9okxtZqa1OMHrHaNualA9eAqjNRALMdL+YowppM0lKnx
rxeNhmdx3xlK41c5+IA/km0R0D16hMjmbiRYi8fWL4dRgWrFQZEO2r8+VUoIyob+I9wY6epWcbxn
Z2eez3xW9lvQGBywDQBLU8I33oXNMdvvU3vfEpccyIVpZMEVZY2NjAgcw62VilydNbgEMNquZz1c
ennTq7dNf+W99yTQLnQmCkvy8WJewq3hmZLzsyPJK31HiZSs8bIA6OMSJ5WC01TgPl8htIrSB2s+
faKdvYndVQ19GxwnoVp9gcaBl7MSK/Fm0F7PEO3TcknGBJUsbReoSzSMrch9q9G3Y1oFpLhtfb/a
uRo8qdXZcXjbOE4Ggzsz+x8wAKiJlNe1W0G78O1xM2rse/gPsbPPwcL1IlAQ7L3V6KY849DppEO+
PY7A8bDz+j0Cac69KXz4kL5GwYpn3WTDe4CzqfrYuMWAF8qaok2L0jN3YO3yChoNI+qJL3lOj78O
tFU2AUL+a0RAQQssfmnLl8iAd8ilqrroV1/Zmrjrkkq3sMQs53TdpW2epmTpgiJJ3F4zbvX5kNrf
sPNrTvF6X1djI+faNsIfFtrKlXOC7yFpGpDIkIY6tm6qRYL+a7wcWThTBBbKeR0ExkEgW/8ONZUX
/amyuEG2t9Qqz/BhlGOnatZalq7N6QFxC9CRf3VyBolLzDET6VstvMlJxNBWuJN7uh5gyMd+ju/O
vFIR5PwzuW/EZSkLP+KK4OtEMhvDpo+xYACCMtzjXEofCbFvmxATnDiJ+FBzeVG0m7sMYLyMtSNK
0s63IOK56qV1hea3KhdDlwatGzY43SECLUbdktx1ktWTU8saMTiLGNhNo/hmnNVs29mqSKO6zC39
9fBKPvkAE1WSq6PtZp3nEKjRKheAtjXz6a6en5jSuAIME6Z7yBcxW785jFuactY4zDm5AVXe06L9
UXwpDorLAeu4ACM+whtVra0oGBf64pj4pXg2ckuVhAAX2/SCvvx8vDt6kjetoRrK8SsONl+zsgZZ
WXiE3NgIZCJqzzgBHD09W/V8RAHit5zLaLyyjk94eXUS25jxJUDv03qJ2sKJpRqUQbn+uQAkmizl
AO5EIPEIHF10ZoaayAAfNi9xwn5Ad2Hrq8cgbA8tCsaeu6omwP8MwwtWta9N2pvFptiYfVN9H6N2
XN7S6+6D2hbnkCy6kqtypXgK2MWe7r8u4smRjMUWpdkLxeVOIrP/LYos67VkFRjPYwVrp6IRpRhI
GKzBK60GnGWgsU0p2LU1i4Jg+b/nEbN+NS+nyceYmvTNhXhCTdMHxlwXFHSdc8sExhOpR3/sRffi
IrqaFcR+yu/Bi86si7O292FZUnPpH+TAN1Su5TIIz87RzFTd1NWAOF20njRQEvFeYgIrX14KqUSP
Zivaxqjg8kpZs/CCT6pug8+vanE1nr6OsXaaOFzbPt5UkFeAzbnYvHK/os1CChlGEGlV9ec5ssEV
x30HoFTrY21ZwA6dfozU9hfZT+tqrWsM1n2a+5ds64zfJIYeKB5uc+x2XygD5FjUs92a0fR5EImh
pWV6Sv5+x0sxjpprJqcH17qiNNZBJCcawfWg5f4GQ/FQwAe4SOvJSG33D/IhX2Mex+ljOC/MMeuv
dBqYFRgI5cZNxQPnBl1jxen8CA1F6PHuZcKDyxIAC/yZQovo2LTYMUQZuw9TdCjLdvbovIUUnrMz
ForaLBTmN5gp9IL1znQBImvr3IAJTKJKMAfEH+qxaUl1ngAPJYjYfOi0sNcwLCKs2OtX+OEXcpGo
H2g4cWg0H8h4L+b4lltBZYkBGWe3+4/W6zXpkU1e+1sBio8sHaa+nlVfhZKTqSXvq8UraHPnpkGA
Xl3hsILomXEXJCnfUlIcQBbT6qvVuaFw1HxZzeeR3/1iwsO8BseTKynIeok3s4yLb1fAVuMQqnte
VoYE0ZniQFYHtr/jP+rCAl4rGFMYDo87WgUYAZBSSEsUf/tYHlsssojcbNBUPEMgQ9rVkJBK6DgI
L8w/zZWLh1CyWRYGhXwjVwHbchSrdmP8eJF+NJNlBUIYwZbt0POSDxcPJ8uKN+GjWAVGwIrsiZbR
lJwPX81sVwbh5mBRvQFk5l6nN7xi3aZy30VFf36iVUuR6dp5P8OCUKcYQmlpZe33GlN/tk4Kp5Vr
c1I0cpZEH8kZM/kl8sksO/aGbeYpYFiGowcY0g4W0M3KwSC0ySiUpSkyoZA7HArtqu32gbh51Fi6
Vxl36LtLgd0YobNSL+/t/CNinsd5SLfPGIhTNiQmKPmWl1ZhqOjJ/J5C+H+JRb++eP/jOyXdgH4z
pTp1TJLxdRfZxhDTQW1PqrQ3FNTbk2eMFZojNhs35Yq7i/0KDnB0zI07hq68qh+yjm+U047hr1vx
wkj3BgIX8BuX+/mZQcG7B3ZOxpQVfhNBvLBdgtaykkrbS+ehc95z9CPqZSylt9A44Cn8edTvdXQC
1mr7OLUTeb9YKsCWm9fH+gZ12JKqydlmQrgj5wOcsUyuqlH/Ue/7f/UFsg5HKOniIxC4qXsEmsLh
R9xcnCIvPxR2VWBAr8iRp1tv4fsrYJO+o/zuUw7FItJcYthFsTCPLCCmJhpxjrWqqDFHihV9/8+x
ghkrxBX7vH1sIqM0HuFJUzTe0eAlFg5y72lF+KwDeVS6mcATf/YjpnoCRE/Kc2IOK9jd+fXceb9m
Cuz22IBsif0SHjXHciZwZ1b7cLqetOi37+V0jJqA0rfeSvfBxWNYCyyvU6agOsDdESHLERULwFDd
+CatuG821lDKZzTi3FfQDY2+uAUP4+sb4uxqpIpSqElOIw2SBt35HRwHnVJTNSpuV0Rvb9KTk8Go
akbyUSweAuKMCS5EsquCUA6iY/AvY68EjJGUXq2i4iD9KO+EUwy5MFUFtQyom7y81/0Pjny3dPI5
S/g8+lZewjeqtoFuAlpMn3lPUhGzdLLJqehpFnZ/jU81De2yDOuaMo4F5LgJKRVVrh/9HRYE0X1n
JI/L8N4iFsboIS+riCeDSr7QFaAFn5fm194YGixhLWT5e0Sf3k/WI0htE239Ritz/Eu9AqWss4y2
ATiBbXBWQ6m+4iDKAtc5kiGmmPPjML9tJ0G4tA3efQjasaFAGlkTcQ/hk6CjQKGAkikcyvBmNksL
yxobZOYRGtC0kud0/2ztdGUUy8IInFrRv4cLWMLmlIXjtHUUNkovwzzwYdtBRVqJuLcmD/hmzB+B
jqVamt4EkQFD0Ay4jDTKuuAnTmIqtoigQXrXJG/kqXtPtyblv4yNQ/xKm6aCmYmrmqZ7hOJ7bEdb
JFZA1fKX2tXMXLuq6tDXYFPlNVrp8mwej6vdj7pkQwDLQSI092FbBJlrja055JGhNlcDOU5JA8zL
i5CuVJhOydigaKFMePk7zw/+xGhmMAcK1px7/j0dcybP6w062xhA1TsvqvSn8Z005EUMLAWr/2LG
mCi/g8W1jRXh9S0gUxjnG7HP7d+jRrCI71E+VDbVRKPYKJWK2+5WQ42LehbGuvJ8vQ7pIA64u0p+
cjXY6g8iZ+Y/4WCT2m3s4VMb2de0/jnlvCOvw3lH9hJ2jigSINadpW3+Q7nY5p/uVe0vxlGc7juK
S6elYlx/tu5O+zZSx0Z9pw/qdivyEwHyaPxo5w5mtbUvH+PzBQAWRKk4VE3Ko3wYJ4fGFTNp3hhW
cFWsJsKm0UW8xUxW8v/O41jky4VXqXibpC621Wtg1QXpEk+hDXRe1nhOjYme++Tz6nOwjfzqANND
ISVdaXg7VsVcvOZ3LlVyNxsADAomYBudfpwmtjiAQzDBYsq4eW3eWcwlEJzXUewXwQxxgnZHLfE8
Orhj1SjHXdKQ1kXBlXiYmA7DXN29xQ+NTmXeJOrVCX+5jUcJr6g2PmTypc+2beXw0cjihnhY2dDX
IpxFRllx6qOmPl68c/n8K24HxSPofVfbGAvFACwUbBgHJ0i+TmD+fGAMzXkZYTySABg8J3OoCur1
Z4GxNnbiFVOmJhOtq5qc7joojwqR2J3ASmnhgmfqYTSA+MT47nwcEHMVSigOL2aQoOkzKyTRpY48
v9qNnwB6SYqTKahj0QMkKRBWHtvgaPLwGsrV5cLYfPYPC3/QWeY1OP6tNGe0RQefSTc+9zQd3tPI
Aq1pHUTWnpNSqmsrKqbHtIHhZYO4L5yT6y1pQ+YHTB1DIzddS2+iApFVHrmgMgz+AqoynYv083HB
km7x/magVgxbG9NDW2Gqd8RbdSKS4FP0vq7pn8ikm3CiiRCYyX9qokB+gMffkmh+CpeRyhZMbh8r
kLFiNxyftiUXtUym6gFfhkHF7MJ7kWBMkrNOp2hMropfmsY6ILfO8nthbNH7j52IfvbeWWLeEJmy
7rkANBteL1V8oOOfZ0O++3xpUuIFwnFyRkdpPsbypYsF2iJeOBUrT6NsbTbWJmY78ig0ODhq/K8P
Zvr3+xrYABQiTz6WqXX/j4wq65kQnRvAKb2P/spxIfNQWuvbTd3sMsM6/NwCftcfTTVNAviP03vG
g+ZAToG5b6BWyYR80IYqwW9t/Ec4bPgG9jS2wxDHMQ3DDcN0k1agLUjBgDdqhIqDLdc+ovqRb+6u
nwnB8JgGo9axoziMNwcyf8PCQ4wY8kDlPWmRHEjDXOfV+bfziKh6NgpoQqD5TRvHkpwqs5A3pRRl
RawdZEO0PMN4lCFZBMdcT7ZX3tcW5jPT6aE+MLH6T/KuZcltL3U9ha6mPdKka/4uoETc6OSx7LtM
E+z9Ayk1q1qZeJY4K1x5QiSbByK1d+8dZLJ35vQJJ5lFDELRri56IyeZlpmu2FXVvIMD+NdERJ0P
S6E7ZusetTcL2E00xEGvIlfwz6yT8WasFIekkEv2kZTYq1+1tQHjvJztpwgyVuOdUU3mht3MgNDs
+YRKWHJ8uwtQeHevhFMz0pmCmwOUGcXYZFTngxP/VncArBAn3iW+vENL9cS3Yfj7hNAZDRfDL8Km
h++bar2fcgRcx8D4WPgVYybIT71L4oZXBJVYopvRL0ShTviBbLm9yqQdo799U/wDNf7O5uDYFqke
Era+mR5gnk9WObKqQndz9Lum4xDe6uASePMXuMpBcBZwMf17RXlNEdY7WyM6nPQ9dt7+/shNdrbP
9/+Z3XmMWXnshMB9RRnOlA0etD3ui5jzcOspLsod3UJUkfknGDtvxTUg/61vgQcHhRPK4VlBGoi2
rf9CXsCVwlXuqPJcA+e3xZNvvpBKnGyBZTqJGWG7teSIdGFLTrg+PhmmRokbVyqdLpLxMqhmoda9
mRMPn7CBh0CnrRCrChh2fUpNsVDhyQ+esix662WwrBrTrIAb4RpcWJj/jtmR2J+EytMam4nBkKgY
4q5IqoSf0+SiNoYGcpzP0LFwi/QsXhP9GbnoW1vcuaq3vvJWFtAJeifwsu7eiY1At4UN3imNj1Vh
hqXhbu+eV91fuMTB+Ci9XScbseLIdxlcTNyYL3AQtaxKaKZjvHUgELNxUo922WXa3IzmDRJUNE1Z
Tmhc0gVvxVy4XbqOd88hBevE73eBBDsGYbby/0y4YoOPu7ee8Z6yBCXPT1q4Zx24p+gDfzPF6uI0
94KQCU+Oh6WA9cHEcs/v4siYCNIqriuD7G2xWZ78DDnMr/LYmgvBuSM92Ez615wUHZIF8DUCBlmU
N4dTh8nEe0L9mFqtql+U3TAzDL81Fxwa/vER4XGxA2n0h3HojvoaVmjYVm24LhxGfipO6ZZyDIjw
CbVovVxNVd9rS+/GpwlMr6jnAnYpJE/TmJ8r6423VrRy+s1yXZQ4cKGceKZ2Zh/rUAGAN/IeOgTs
6v3IIIsk+3ddgtk3lRpVyBw0PUKxRCZIKFJWH7gEJUF10m6ujFCnnpEgMQ62RWRBC5ggqvSD9g55
IeRlMLSKz/jcDwc7ExDSxl7eMlOXoj6kJrAcMGyjit9j4tsBRUmGXhckDwdxtPaj3rvTYmFHArFK
26+s0PQkxGpkSji7TWjRgcEW2gumAKuRblGDjMol6EpRtQRDNvfs+Qqwic2APWiFx2K3IbuAKSA4
m8tA+f2NBg+1gawKCRDXwzaYX4J0YnftOCIidmXe4D0a5WkoVCBN/EWD4qutjrO8SgRONAUbboQF
vLfluUM4RCwZUSjj0JDdABg1PzbcTRhQ/ceaTAweGAoYLMKsv239lsDeBHGiscll+A6yVkbZ842g
o6iSqWJncSic5E4ZPmBDXK5+zsXIyBnDzmnegrL9gDSaT2KJlEtHdRZ0fwnCLWLxv2TJDjrxKVtp
w5lSnXDhsH1Bh5oXxrPsCWcJRJ3/efrcvX4l/8hJBuO4IQarSGDINQet+11R/xisNjN6ziWYZjDg
d7gfAWdpmydLaQGE11qWMj+i5bFN6O98q67z6UJUqRh66/tsIrrNAqCns6EnJr7+5c9PhsgSp91P
JzSOnkBvHiY0+ihPoh/tY3elws8Sv0oi0TztS2tSiSICAqJyzPlMH3grUQnnmH4mxO2ejCsamVow
5DyiGrxsEL6Z0UgoQsB+cpi00ECC4irqecbxOWkrAJW+Kgw8BmkvEH8oQq4v0fdJ2BeAuUpF3VoF
JSr/teGIRP/55oT/q6rZt+b4h5X459CRSsfa+nM0Zs5iONnlSXWIL8eozViMzLmeXT5XctTwziqx
gbKGtoB8aBNu3B9B91SrU8wokqZ0Pohytklpm7iDnBzfIgUpBifUTA/xE+kQlZNh4Hzye48OG8nW
HhesPd5BgmreZtIbt4R6kKjW8yhv5DV83VuK5GPd9A1YJYslF+yivkV3UUJGw3xcjMHaZwqn0R41
VBV0Pgf0OomZYwl+Lb4a08XK4p5u/JpLZ4PE3LS4IfB8zNONkzFBsZpc//Nyy2TBnZfH8cYQcOMz
jexcGKNFhgwRkEliEdOI/Zdv1HmvlMKqP4Ldj+r+ZKEQKSEbOaT+sStQkagKOA1OewV3DkxCNSdD
60zqEl6EozTWsMS7JF1Lmcbs8SmLPFxdGjhb2WVfO5u6S7lzsZRzqAfeCxgsA4hDYmc07hxRYvoU
E0jhXmWmqwRJenHh8t9N3Iw2XjDif01zHN6fOdUGpnCyYoCVYGGJZAVcAly72R6d6BkUbJkA0jmo
sVKioFs9ca52318IQJhV3Ey4OvY3VU1saUItR3qp8wfMBFADS8Lek5LQ1Gm1yNcE4YoMQ07+x2M0
z0kTVRK/xBP2xlU7N9JczCFxOxVeqiLV1jzCx2cgy8xwsUGqZi7rroxy1QFlImbiDWwGDeEXopbE
XXXuQoIptnyXJWr6LhyIZNjDj8x+ACUCZxWNfLnP3w3m1Cyy+BPRweSFxsinn8Febx2R7TAWDKTW
GhrGKWbb1LyO1TVdmmYQ1UFrGhacRn4ZVYOiVwlxEypFEXw4RrLAEAoOLzQYRs37jHmZJkMY9stt
2rroRp1Pa/4qJsuBFift/seilP12711Ulfbyyd894BxNvm8uSFtYK1d5ta+fdMsWQ060IkTijvl1
wt9jlw6TaKM2cPbWPm4qSshT4O3A7ZZI0RbQyofjvucIt/1XgPO6dBxmxkcWi6/GZQxq3QSSxBPW
CTZgjREAvJCGJ7dZnOVrv0Z1OLeU2y8BB5MmGhhyBeIafVvc6CJf4apM5bmst3RAvKUcKg/7jhsv
9XCBVnktj0bsJ40AlWx98VvBI19XiJn6fap+gwo6IeHqOv0zvwhDJK4viJuY5dxY8xUx3yoaukIt
hSBtY/M0B/gz79qIYUArl9A7TFxbIyPuxGWHKyhbLPpbY3dp5ZUteQClKg+jpZi93YiE/OscrLVD
DasEJxkKBZgZqRPgxA3jNpWWZlXBbKa8usequJ6tHrJHpvewTMYVUYELuyDOFIYPclKs8hyFHqdZ
Rec7lh4NxfGnjtyBczzeONIhtx1AA70wJ8dfhNV4o3X9yo5p4Zqvi1iTUKKSAC1hZWTwOyqYkHOl
/yEkCYwwjefb+O0OnZKGZnT/ut5V5mQETYPZMrDZpiQKCUZtgsgYfr4E7vWH2nd7o/rHXUu1dhB9
MP7lGYx1n5ufkrDJGptLBNt9sRsDCvwWXPWJI/dUzsTI/vPjWgTSz7YDrOZeEIVqsjthE6VFf2He
4kDv9qPT3QTenBnEicJW+lk2L3kRVmDt8zucbDIyim8JgMTfr3q2ikr0amhsh2qhE4RkcsmuDG9p
QcT97a7NH7/f4Osnz9LRS+PVVXpWbqxGHRS/fXsVuftR/aT+GKtI7UJPpWzOIzgpWnx3EH2dtoqY
tqAsDmJNnro8MJQMwdpz+P/PZCNJ62yr/KxI9AkPnngczoVR9OfNMEwodNwbPFlavCHHBm9RA+Ce
I44qzZLLGKePvd7o5BObfCDsgsBCAHYa+NFLV16LKSsAHLjl3TLvRU4hGEFUAKNRzm575HRuGQUn
+kj8M3+Q7dp7Ie6j/+GRiqxrlHo/Yr6c3+PGYbQcBPGT5/jqIrjuJ2RJIzQG8FsERUxlYztCgaWF
M6OJpmuaCo7aT3TZ/BsVwvREzdo+JisNYOaVPzoVPLW+gELnuqM/rTB7NwRh7XX/2bEfNzSE8Syb
wTWX26Bicr/3GYknQeUnsJdNPAyjjb5CzCGgygzgamS757sdO/7zGBX0ubp0zHCMKVMc/vfP7h1z
xRqyfqjAP067JNexR396p6DOXCWBYvBhGoE6yBfR4laqWi4TBZzyKJCwoJNTgETwFF/9LiGNmtzR
qkOZP18dH/d+1JSrBe0ogUVoLo1xmzSDQaGoRgfTtQ3x/XRX/WPDRWyn5Hh+iHiFi+dXVBL9WaIv
kl06lOMkf4m46pJqXq1qUYBB2UvBdygy1LQjJDbk1my/ZBrqDj+Grsi3dRjCb8+8L5spy+ytWYta
H/Eoek7A6C37rJ9SR9g2d9Lrf2QZ7eGRKF2YuaQnLaf5ilfwnIq3igmsx1OZZWjHnqU5RZC9D/Nd
EcpxyTYaVoc7XTHcVWM6+J0Ek7aUpnjmnakU2Gdd0r4zDwicfk6lR524/dNKJrPFnEekKf3UlCxj
4S9E6RIcYRIYXWqDRsfujuJ6H26h3vq8yrbnlc0BhHu0u77h/rJ/U6/xkLoUhRKHOVtHAdGTeLTZ
tSdY+pI0LFy+PKkP0b93y++qYiXNxg+J/UdId4PL1d2AIVXliwA3Be2VJ2zLzTbSusO09wL7Tmgl
S0PjbYVp74+JIBBFhxLsQv+XTrePaG/+vkcNEM/+w5SU2qrwc1XmwLDWT3ywkvo/1BpnqgGHRI3s
KZn4O02RKYyUZCWmo6fBqMCsFunEAXsi0r6ZwUp+sTrqQdg7V9UNyItwuv1YR6VVJpTsy3iXynNH
oB1p0/D12HhXXQ78YI9G1k2zOD1dKA/Yi2sC7YZ7TFQEWrnFyqbfSnRGW4i/MP+jzdwg2SUUhoFI
etET1epguY7p3+MCSQ5+G8owFOY2zObWjFqV88e7LuGONBiTYzwOtN60qdVDNCzETJg8TwQKabEd
hqGKTpNKmyJ2QgVyOdPmfR17kYk8yKouMO/ityHP9P3d8F4Wy8+QmF7PAi5N8N87nQefKV0CEYC9
zxP9A9okQHkHrZG85EW8ocIi0cSYDoyYGZwuUP5gPdZThEPow07ExmzgFYntJLDkGIQArNou+naK
ijtKLhbQVydk927pcDprp5CYTej/QR+PZT4aYAbycDHrm95XnoV2b4QifMcLvkDh3J/SEU9AE7nG
v6kcpxmqnZySKvtGnuTkba2bN++VRt9uivTR8jHaHwo1xwZCWzA8Rzcj/Cwv4SnK3nr/2xX7XbC/
iCphXNBCF7wZjvB8Z2r0ngSaVHpjMJhWkIxD+dhGe+JGA58XeEAN3wciMieU8zzMSsitTPPEe57K
OKeI8teCsbvg/k5KVamhEzcicyT0npXTmqo/GG7Hdcx9SWN7r58aqko3/wVdrStEKlIXwVDgiPYq
0x1295xwf9uRuUJqA0B7U/eAIkdLf0B792wteHErNxWKpqFteQPquRZSi2tEBlBKlJlm3T/uU+hO
kKoukHGW1UC3BZ561VYXXwFE1Q/HugPOuEDEB0KOgNISxuTCSydp+8PdmvCgRfSAQWycawKPCrsq
AXBp9RIm/CkVLL+I1wg8435Q8/CLQp8Oioxs0ZIi5QQkYzWAPAMsNuVioFXjqcJaJDQQrnle0fdQ
915Cw271mfa6uuPl0h/chyl5/LPqxXDMMxUYHiXQwQssN6Xs0SmEgtXvJQ1tIrIcyOXNkHhS7cql
SHZwO0n/rOURfVMTL3cfVv+7uwXyifKLEycx2mCtHbuW/O5ZqLNWiodhkSrJTzUW8pDkww4rwjHb
pL61gp+93iTGbu+6CYgpDoYuIoUI2gZDx2A501u0GFIAhs2u06526SeDN6rZbBBArXOeUcTPr/rL
wLy56xMlwnCz8ZJ6h50H1Qsvd7ESsdWLVj35FYgb8S4O9RX7P+bhckZ3jE8MgP+Sw9OJ5/IEmJWx
1HODAOQcDtB3nKHMvDSquT5KXxI+ZdSTEMp3YdsmDTy5OY2sypwkRj7P0ubB6D+2YjM/RQCSVKd7
kchROTRru7hz9NUL/9X5c9N4B6tyghOjE3HxlDTek7MrolGXoPwtXydfZtYYP3W2PW7BrGhKZxq1
BR65IVxTW5nG+SdTS8dY/cbcLgbl8XBpsisHdaHLrA4gPVYxIFO/2j7OyxhMVapkFsGCxqpNJhJN
cH9glzlta4za3crV02y8XLXteZ7ftw6pbWZBH1ix8ZNgrjvHoVy/D6X08C/mR3VxfltIQ/aBvfSp
7ZTIWYNKHPNXHEJonC0ExfzRo4h1fXvqkqj9IOtaVikz6MyoDJHgff69WO7ZQo1yXaYek/lbq8ss
kv3RFW4y89Inqhi0qjBJ+xH/Kzyu+JuFFcusgisc7Je92nkTaZKdgoCGU3hYul6QsNuMMeHV1qRK
UddlGqzkQSpDj07QoxnFVzi81k7Wrj6qWuqE1at/RgfBpcsj4PxTmZpaFbq37YyCZFinCsP6/rEu
O+yfBB+GcGpFiw0kuOMN50f2G1ibh1FDNf1HOUGx+dwREEeHWZKRQ5EqOjtVQH+2wl/TgNP6yP7Z
zXQWBturLs52LwBvM/QyFpcu4pswzyja8b5+ZVow24DNebKH48ueXgq7TuCyCyNJVMq/bU6bbFEF
nBO4cMS39DE8Yj5YMsHtMEoK4VWZF4rGpSy8STLOJeu8rVyGXdt8xuKAZVubKclbvwDlhQX1JWU5
ljvfZnjJFbRiEanHBOpzsCuq2Z0GqnhgXN4oEsuRpyASg7fboeJn0KXeTSz0aEwGNO8lhAHflAff
pb1b1u/lKACsUxJEtOgBNHoRLrA5ndcoWUj4w2LepfpnPeQ8Hl05rnik4GBdg81yDE1o6bbG6GYO
Td6aS7qIEV5qJR0o2r2mGDYnrwCQDG8zbx94TjZYeKGGKa4pEx4fcFpezt7o9GUedRiRdVLVUjE5
jOB85f2o4WiRl5l58wxJO5bi+YgXdGYIGVV0Goa2RF1ScABBxdpbcYPRZE1EA718MJQN5/b9xQlz
jnHQQx41VcgsPUXhIKXc561hZlUwWa7ZVzC7941DcTYzz4QZF6+BhZSHf8YnR4bD8e2UHbR/FLnb
yWLvjSpb7PaxfBCpG+6ZpxyDX3+eVg0U3p7LvcdmxGJQ4kLlr9OxBy7nLa+4ZhPWrPy65s7W0qda
3KVmzgwulqB1ICPep/C1zsCpBUMNuPh+bFjyz882ObEEBiBYHtE48uK/Z+u8kYLKg0acFfX0DOcn
xfo5qSekJc6pEpmD3lBOaibHWaqHfhLWthrilhZ0bGaTBeMB1OdMx2Jv2MEJlaZ4iLM+0MuAY4A+
SwfbfyYqca3JNwWy8ObXlUVfwUkQwyfY0p8fc6Qe5Fey6bR3rA6BhdCjPRseRHmqGh+nQrSH2d9V
9nJZvOXykBDtJnIAIPmON1eOL/r9TMelbEO/kZpXV14kVhmKsHFjzaS5Sar8V7lODUGPrtn7OLGZ
laRQUepVP1Np9i9GlcR1+mxtkjXvQDpcvPT48f21i0sTt/AfEc4nz8l8NMwkgforxDohAG9moD28
gpSchRZkhEkXDa48cvJQLS7KdgXOM64DKe7XCxGs2xJ7PSjUlF4YKVIJP5zdOLcKystZ8/LFOaSs
Z59dGcS8FnLb8CZhP4pF431GRgG/aB5SDlvQHj9wkp9VqLU7OBTmrUeQ60RKpTmqteVOSIJlsntr
ihtCIjY8xD76CktJAy7xfArCq+w5Hq5MiWXg//HLT3BFTRWeM+rHmPQzNeAeAn6ji/FMpPIwaBek
aSuMIVm+pkpI6g+Oz16YxQmiPjOTrXJgM3PYKkXI4NKWD7CtrfhCfTH9NDNbntdGXc3B+P7PTn/Z
krGVv8qMH0Hfg9Xm+nHH1DJ5/ACAyaCsA+PMjFmcDIOmLH6l0KKaMvXPEbX3BhojKKHITfkyLSUN
/tfsV7cCu4Dk13Wg8StYVkFGn7IwaxbBjeVgXCpTofW/Snjq4pdysUzVld7fIe7XN8yO78xBHnI0
+ICpeDvyNUmqb0mAqO9ats+yqEwbEHq0HJBHaPyp7L5gB9s00sf7DkTPsOlmt8Vhpih3n47tNnDI
0Yl2nv59TG7H09cNv07iQCTjK6xVlltfNoeE6w1lQsdLd9feIWwbxwEqHB1/r/B5Ill1McHpJm6l
DXBYJLV4pqR46r7y2EdpeJtQdlrejJ2qaznx1N1Spj5JUcx5Zv7aSuKWGZCprcjATlnmxjS5bv1U
VdazFOsx+y79XJ5A6qle+8KfDzuTSTfuvwMiD8hobXsW7+EtLoq7ttVHHOeAsxamjFSOL7UDweQ9
EKKJdUgdNsq/Z894U+W6Rn/46rv2bssj0OC0hyhcQlXT7e4wWkoYI3c/QJRZN10NHArf0c/6BxL1
G57hyV9/hYznlbAIsYz6pFWDWJ0tRqoTmB5vctmoxW4DbLljEm0QUb7VBaT41AHOe9sW7fw7z4OH
0W4fwDvxwS3t4jr7IPf7fb+4HMdC6k9o6C51Tf0f5o39Bq8p0EeFNuztkxhaDcNi7CkksJTdUvdJ
lQt+XKf8L9ECxBHS7Enr9X45Ita3f4Bb+gScxtEcTwHzzpeiBfsCDLI+/5b2hSSmhLnRmvsFzXOo
G4QDb9BM5StEKRexUEnrQctUMsG2rEJCFTJwj2X7ximqq4CLDiKa9+/aweB5XpqS44Jhe1oZKfHO
v5GwdbTwYATFLV6KBwg2eKZs9+m30JFBJkx1LbzjLL2W4p41Kf9UM+KQEIjEs1E5JxBIoD6+xtBu
A83KG6HxpG01zYvxrnsenrMbNly3A64P1+h/dVXVlq24JtSTEcmrvW5wmyrS+vkgzFODXrv90MZI
ltfQBEwheAc68CQl1xyzDtE27E++2T1H5y62puKUBeiLrLkC3x7bRibVaKVWu91iDncJb7DkJDn+
8Iw/o5qe6dvZT9ZlOWosVJfarhjaT2rG6ciDkTw52xTaJXavtYGI5KgAq5hZKGKZvrG2m+qefjo6
prWhcLqIvHndh8l7OkG0SvhR63tOiSfFd9+V6FMGpgjy5hd0EVVOL2/knVweHE8kxvazxsb0XgYg
S1SVRZ8TFs6z+G/uj+dn8Lu611e42IEYomafR/d/82wORr1ZL03JefcugXdOIFaMRzBsJO4fjT0X
IMqXCW03mcSdR5tKpoJihhDNSq0bnTACTA1v/vMPd+2r+oyFoQjUszxg0CeHmpt+uTlZDxm8Euma
O9MYiTXZwD+xHuD0YPK6MCqvFXEy9IgiYnjrflFiWbDfPFDHFvtlLJtvusLmDJdijdejWN1UutPI
+TzUG08T85zFGvLfv0RvLTqgmrS/gxfkd8+pI7EplJ2QXU6wNDUcNt+pGSqduZlvS/nmQov1DyvZ
62jHE1TvS4dwqHm4PM39XhJssct6tST8wRN2oWKym0eZ0/Zk7HjBOjrp0SyA78VXQlsfdktwTeB3
IfQlKQSzxLtBlXxZapIOqokMP8ppz981mhnii51JxKgkuSBIJccq4Nj2u6PH9KMi2ssM8Xlv0Exf
mqTyfqgOEdhuA653dvsKDtb2pdTo6cE5B0fLEGAAvbxRWzj2pBkXqlI4T1Fc+bJmPE6TQMxtgQOt
Az9R/NPeJzYJ74esFsFtjXT4UsUD53azJyud3XHCFw/5X1v5I/39tFOgUXl0dHk4a/uDHjfL+X/7
yFygrznmrDR/yfT5Ti748jdTp2/qPknkjLK6EM6vjbXR97SC2Es1odg1hiS3hC7VdrAbmzgIQF3w
1a7ZkF6ykilt+hRUjLIRv7UVSjYYj/YQztSTO1GDkJ7flOmwBLgcT3HCQ2dL4oyiseZk+yyn4HqD
x3Hgc+OaXrd7c2kybwrqLMyTZYgy2Yt7uP3d8mNsZoYrjlzlXBVLrKib6PCtHga2hxpEdJ/s8zZe
e4pX3PVEz+c/Hn/QgY9lap9tEXWJZXvXuMmynEqmvQJy7h2RwaNwOcnkMv4Vl18jS2paPjVI1xPb
vdUWV7EXYc0ji+RU71zixbCIQzMGZAPE3uEjigd/HBTegjdhhAjADoTnKHUYhJSVVmn1it0HYuYy
VcHVw7tC0queZqy0kXVwtnMymckiM3n+UrBQF9PLfnhSh+ReC2HCE35/BABHrpOzPWT1N2Ir/jky
raMzpgWAdKkj1kbx3+YElT00Qx7hBE21JA4JHlVetbguVq1m8MVDp+YRH8WehD98Shx/ehGj3s4T
/asbyUGlyS55oIlyakIIVFNzwPBIZ/s/oNfND0i6WIAaXlbSFMRP4FgdxyZ68qkl45tXo719n0Tj
wEKmpsfKsTQPNaCda2mJmikLbPRzCShwb0OVeViZwCPM5IccOK2PX/jyMCMz3UgaSzMqxInj7g12
N16Pt+/0SUPnCgmzRRc+5yDWf+k03/pYNkEEyA1RUdLzwDxpZiF4tWfylF/7b8I8Ngv939zCD1OE
uDvqkvXCwG/8aRKARLfexgWo5rLP21bRIYgw8vm9la6auroqIeWfwvmfaRwKtl2DIJ6KLhPLbwL+
ti+khdrLpsRxTqYsbYKSA5ji3S+ggKBiPj71fPVoDFG2EecsBNRfyQn8bo9qzWpiqjA5VHlkxFnU
xptH4JhuFBHkIOP4i7NpThHHTE7OL8biCr/SDKE89OA0Xh09tYYthCkgRbeZJ6dmjNOHgJRY8Qt3
Vc6wWze+d0U8AO1Q8W/k5F+QlA4DmpktEL2WJLzJyn7TXl4Ct6vCzJqyPXIZG42wvoiCvo8ruEmR
IOPaunsG3yp0ZgDCnvphN2o/vGWRUGi2hNV7XDogd9jjzyfZb1lPjWbSUam8eKIIp9G4V3IQyP91
9bAeoMK/k6jWctD3apvAXH14C00L0A6lUiOvYCmSrkucULM7jDzUAYjZsV4/2unmozYqg0AXGJfL
LmZfFqm6h7a7uGjVtjW4Z+YwkrMLjhC442SW0X3bnQmoCTy8RJ3z+hcCvVOMWpShM97l/9fXsYx/
awJ5Ucc+dP5J0c3C9SZKJC5WYW83mjlWysqg2sMEzwqAOwW7zFx06E/39Tyyz682fokBd8pDOhMf
K/FFJj7xafW+UQS5+vIcXwaSBi4vrChHPItX2LuRNUEYDoG88yr52P+vI2waOwwqLpkBlWjuAFj2
vqnuWf/O9Rlx2Tv47YnYPVpccSJH6ImU0Vwo7tDyYcCL6Iy+kdqzclGdyWJ4HPT/CSy4gAdSq+UP
AeyYef+h7LU+Cu4cljrVCJ3AySi5KJJTOdS2SeZi1er/thBNuI9o6o3+FU0VVcf5jmgUfqTd+qsw
iFcTPU7ne3nL3/ohrCNIvcNeJY3dk9aTCAQ14xLTOCUF5k7B219BfW/U8LDZsZH0EqLX/foIxDmR
1/Q1wI1a7r5k5s3wXBexCgwSZclZD+IDbF7MYNyvTGm6EY3KdNFp/aoWcFuSGa7wo3rnvZQFad/X
Rs5fW3E87Ny9/TBvn6dsad03QLxb22VuGzUIKLbu8l0xlgr6NSsiqpHQZuFeIV9sqAGmVoDDD/YL
zQORofmIC8c6JNvVVB99avBr0VQU5lzJgrn6PkRATMHw9Wrm3/mIa2m/hVoaUJIFxIhFcTQ6wF6v
dQd/wlt0GaPSUYmKvBykKpbOVf/q/dJLWG5RhIlcRm/UxBO8rIdgDKe2q/KTe8HBZtbgt9IXh71+
L/leUxlg2MzwhDQhtKIDds6QI7Aj1aR+VhYr+PftasTgQZqn5+DIlTqch8KY9uYf0gjrwC9oXpAQ
y8bruDHOS2e/coV2kL2RADZ9BGoYzxiPTg1Uu7+2uU+hUFad8oQGRknS1e4YIJdKehKCWZYQq9tK
EL/0DfUCyVjaJx56e4aCr7XaVBsaRm3WjOIWzhZB5XmMHhkHiqkb2YPyIJxcJdYP5jtYsL6TfwRP
928hTNSybV/TAmjxD9fQs82N8XQDBdV6sz9hR2p5B5vPw0KohUSpDkYBXyMpoj1VhRUpJWeUMNDm
dR6dYrgKLBCem1n2vF8r5lrjQGmtq8g9t4o6jrR7nJ3+VnFw4YsbPDQYekv8jfWZl6V6czBR89Qi
ee9eQw7SZ5nu32rIVcRFVMsnUge3SwRDyojI6o/AO27MYc/O5PlaxhInHiogZVqiiVrTpCFIKckI
OxkDedPF9KXZRqPqFJP6kqv9WOOMfhtXmgjwfo7mFHOeXmuZusm+7s/MZWLxTqHJsleQoyMlovye
sXmd0XxeRUNb+fieOcjmD8JowoPuS7028QHd5ci72uqRarV3SZCRJtGp4c9tLCJeVl8/QRNxUlRy
84VWeatxf3Fi3+iRwfvPV57iQW1Td4OyFKeVyNEwPkd+r7ulqlBX/nc8SDNjFwuvU0CRRfsA6pTc
sI7vv7Ch1lFz5GtSwlpmVT634nhp8iiOWWDG7M3GAENkoOcqS7iX6a7VK+NTX/xqIZKlajjgl/7C
8uCzZdJ41Usy+pGE82R7gaUxKfCRQuOfr2ITcEue7uwTQtEQlQWjiowNLiBZsJKCAf38RwAZQ+Cs
7c5hSV2Lu7eevw0LnMc0DxgKjVXa7wzs8YpdiMRaPfnHW9hRvs2EJkE31EjUOqwm3Ams2y4Z6TS9
CTZLE49a09LfWLIFqv/l6cCuBX+KXAAgU6zQhZHD8Hq96sob899bftoHIG6kWnt6WxU5wabyH616
FEydvzR+EHwVyrK1c2lUuWp7nkEQ9TiCA8oOjssOiztpN323NQGGZ7oCcas2U2n7LtTWiod1ZvW0
EaYLZk0KGSzUUOGecGWYvqV7oEWk8PF2ySofC5gLgGqQFmHYkZsc7m/FkyouzNLc18aEkTCndg2O
QHJcadCd0eT4erA18PFkhHnoGbkvSuOkaFBkXmzn6Yv97kEqe4kwxR3aEFDBElNxfHuSv1D7c3iV
XfGEPNP86AgCvaYq638xGV5nuYoM/zT7EMKaCPOAMZPRUpmsybXkRZ7dQPSMWkplCmQKpZNG3vD+
r/kiZHDyuAcAClvwn1j0e49ubxAjk46F9zRm6tvho8P6bP6xbw4SqKRtrnArBPIg2WTvQoV1W043
tluTKZNCCMFMPm8oaa8NyACrw+PAozkasFHgs/4rMR07x6gFk9N9Rn7tpZhR8cPvM2k3aW73L5SQ
XxlhluSm2clfrLU21Y4uQ0FrJexv44TBXQ7A12rfghLxj3z1qxBqy8jpzodbTTRs/YIoYoIJLTl0
6uFnrlxD20ivFDar/Nh+//5L3QHr3u+5SsAUO16Tou29VCWrrWR3sBR8w2BDvth5p7aFwnxfmTLR
Q9UCsBk927VI9xDkDzZuFZHUvL7LtaFlofyrTqYOaCRXdukv7kU9f8rxeUKv5oE1wlR1kZx8W1d9
ZA5x+JBwigqcl6NwIl39Pf+SngMlsjzU7lWuxSfSARYrsGmo9D8Ab8KbmWcsu6axtGieo5V3JeH3
WimyF0YkwPhZZC6Q3v52kKGk2ycHY0UqIzeHuCBajZ5eCxs7Jd9YMFtxlNKrmDWeq/amJGM4z1OI
1Vs2XFIXEHGJEhq1LJijYEUTGty/X0KIJ3OlAiWyt7Jk04K9xpiY0ILnASzs+7UQLs7A43pLz4zy
xAyU5yhusv9Qz3jXOdqI7r5JVD8Ech9V9dorLUL8S9McRDG9AcUBlg0vzObaR8P40/o7xQS+BQK4
27T9fGU22sBduElnqqoRvSQ5EeRGr1y72rwxgq6HJ//O1AwHGFFFjthUVcNGxFDHPM/uhv0wvo90
+2vO0y15p6Wsho/Z2Zyr6pOCJJNZeElpD/ijOAowTlIjSvNDUtu+dcL9xqcQZqUOrYWKpYO0EsKJ
XEfYnX1iwoJEaw3WEqvqeFOeMg1nh67dbZQK8Qr/oHcXRnmg3x4ktyypX/ugO5PuqVTz6y6fSq89
vbER7DKOMKlRqCPdopmYw2AHdOPhnZ7joM5wOsyyfqzNJL2fD+QE+tN5QRJ90u7bdgwODVFAgvCd
hf+It9lr1MieXYZQ0f7GrafUeUHGKqRwIHwp1/eyIdneNFP2l53HNTPIhARPHIqyFgZZkxoqS/M8
8UXT3bUsex2sUgCGb5fPI7Pe0y452wg7+3F9jF2/oLMsgw5HKbCVNxCtGbWgeqbkYTULbni2sAcz
LIufeFYF/58iIJpnfaUcDQsjRjKAoZ5PV+qSvg9cplz/LZmXQNWNCsb3PHESPI+hrRK0jmlSrPfb
z4ZMogCaMUEieTGx98UhMDPU3/6JbfbNjFHO0QooAZ5cHXXCw6QA7RwSWoGTsXcYYpajfzwS8IQe
83RWhdE7xMc5sJPiB6mqSSOCd+udi7dr8KPGJk2PC3dAzXHfwHFZ3S+efB0fYhVFfQzFjVmVgfpj
V3LZE42JZ5YXN3K4GhypLR2q/YzQgtNHhHF8FQYC6dYMwQVX+4choGr5jwVqz7LRkmBdw3Btr4Gk
hRR+VTctqysFFsSLkMECgpACoeE8faQ31t0sD4a8MeyM5G0JiQqqaVUOpVIrlVyhQJAie5UYb6sx
afchWpyw6WGED0Vg+e+thZ88++p5dcJsZcGNF8kpuHtVY+l1nuyFX1W8WlX7v5QXKlKDFOcT34OY
Tu/gQ0q+8helDU9Ji2v7sPZgrLeU9DG6/emVvHXIyEFOaP/Nbp6Auyf7Jzgk3pUkK6GlmS51G8ut
81SlS8ItqWkNHd2J2VOYRvgo0/o4YwY1sT2JY7HH+pojaChrs81PFh4jUFIFJSPHGOotxpF2bi34
tSlo/+FCMgz2kEOisSacuMabYjAIbdlL0xH9QbwM1j9xI1VXtJdTCaEYayF1L7bjpjSLK9vylcXV
zv7lQ5+LKnk7RF1TtYyI99ZLtlUVOnN3MfcvpYbNlCgC1dyX31FEdbVXuBKwXDl0Nq/wwJ36SYBN
aQHDbEWZkLp/djys5XT3u2nP9WD4pue+pW2DF2WwoOM07iK0y92D6tvU+bA8d3AQfu/tnVXPbvyZ
4JIV9rc5KBay9pz6KtrcOV+QPPVWs2LkOiOfnxKhsKW++2Ks+mAZe5rqkHrLNwQKYXu9cOtjNMNP
ZHzjp6MTdHqJUYWp6tqaWUgiN2eYGH+xNKzcsIEV5+Zg59Id/wNQ2AlKMQKxCN+i+kQbTQR8x3wq
rG3B77hI4nzphkYOswTc06EqqjET9Wx1rpIgHNdzqUEsicHW7xP1QtzFC09MkV4moBwaosWsMfto
1t69bdzdaXOxy24t2sq+CRc3Y1C4GD1X7xuTpLXaWrXHYPtzTvIXxlSfEDKuQE5Hh/kqqPiU0MM1
2fgr4QzqJNT3RkS5PvGxrAjYwn0u1jWKfPZtQ1GFI2PsnadcS82Arg8Js9EgCCHsASg+WdrILbA+
XigMPkBkmkBFfjIDWG8qUHWGccUL1R0Ay7gqKEjC98MrioznfF/FnEVcppxaN58N+uDsCW1d14YF
RLO35I35d5e6aYU2PhcEXp6Q7uAJUJKYFcY4wQ88gsfh+dIxK9om3LBdETvSFQUqwoYQG/HUD0UY
l0pLVymuYG2DvG/IAAO/Xnp8ubr6c3IehLtzPb+CrNDQ+eXnTYYJU/gc3CGwOGfcri8IcGRaMAk/
GARAXP266m+9CdCO40r7TASVK3vOSIwU6XhRxx6Qe+jENPN0g2GX7eoxZqLcfeXsxmxk3Ws3eeYR
UE68EG+Rkd60H668fZ50yP0ZX94oz7WHfH77Myy/tSUvAEK3ARPUzRjFfCL5YzKeGZx+aFsz9mZe
tV+gVao3/4SK4hDA+Bgy6D9b3y2rDEPYaL/BYsI3zTiFuMv2tTxomP9mY7xieXZ81jyVuB2uQQXR
v3hwdSakyUwyVrhz8Ql2/MDjfsM5u8DKoF9/WaVvdIQ/RV4/n17DP294xLIFSlvS1l0+JGPogyt7
Ix8gpw4DhOCw4jQMYoufjzuLjjb/kkQ1xHC8goN/zdL7e7w3kE/Ht3fKgFn2MDyajXbn3OF+7eoY
m/+CnN3iPHKbiYdqHj9enAURAj141JfI44CYDnu3c+s1VzR2tVExefNyZkXkOebi2ZV90j/bP1g+
RCmbFbU1Gk3vMc611yg5nqiKTOkpgpLO7LhVWAG5qW8+XtDX+SySMJJwL394aSinkGCTmTYOv14x
BbqjzsuxuPAlu/EIGWGfW7ddFwCOohNWslD4lz4bPGHO1tWVtqgeSbQw4mJL9lNCJF/Ys54uLRZg
bZBKarV+FmB11c4yN7k5RFfl/90XVSFvrDMgXybx897dtt1MjeH29bQlPDJqWhcS+8AVg+LbjPkA
779QdzPQ9EJv9rqAYDqv5F2Cnl+1CJqDGNAu0JGmDKro4DLWmApa8fs1ULkTw+EUuu+hrnfmflX/
GiZ4mfEbE2ZT7p3TW93iUYPQU8t4B7VGdokuoE/6GsGxf+PpWDP/nimu/q0PS7wkm1Sdu91s7uJZ
kesCUh9Zxjm4EOzNZCcT1zTD+tGrwwVUxG8z2XmGdQOwXohM2h8YGNE2PJQnYIjB85l0Jo8mhWPg
SpQ4pRh+pKpzOZoV1d8HR6Up8toiKkpzya3zHhiuQoGTk7B8iyzagYmI+OhY5lWvmMF7cXfB8Byc
oJhDbUrkgwbUsKVw+55npbchUIfmDoPp/zleVWcEPp5RbtnZD50CZrEcJ+Aunzg2HhWiFEeSLLjC
byqBpfZazSQUKxF8OPFOouChJsFdYIHM8LUpZELVcTeczOQHD14tGRrzQd882kECO2V0+2cMvixq
I47aGA/tZYF8pOP6tCl+t+s3/XhbpyUg5ZdbFSvyPGNBHXAAdxm9vrY7mtA0jFXFxWiI0Lk6m3PL
7pZc4Hj3JJp2AWzrZsIpu3jXPG4jUhVSB2iL3arelgue86LwiiFcdaz7sSwSh4ghVnUB6x36gn0A
UrCRRN2diRKenJj7PVLhjBF3CSRl/2MD2UX1hAhMOQV03hBO5Gi9hvUqZg1sH5+fCcvOq3HvFRJb
gifQdasN7JDMxenKi2WAw+p9aK2s0sd+TB1+TLkNmtMzyXUCVhclfPmxWf6KCT6GAxw8+w6lpH4T
CeiKwHAKhdx2VFIut9Cc3jKYVQtu1V8K7wN3DQlncnDUlCF9d1AK2J6gTal1/M0V1VX0D0hiWfTS
TAPYLjRMlxBWZyZq5bYyoeewLEwxnK1v3l8X/tCc0OO+qd3ZHtLKmEP7qoiLtnH/TcyEyluW7PwA
19orvYVOBU3mNbZlS7sQOLaDXqeFb+sdrRLRz9OL0fq14dQY9wl82omBSR9Hv766nq5KaAxY+kve
ckaXKiSkaauIBHPu3Onj7d3V1a4+Nx3TljDFrBRqdo3H0prKQNGUYe9870FrxTwN70wooojplk9Z
RSdfS94fcdGldMokvxa3JS4Kh8M4U6jpMz2UpGy7zbr+8esKb2j5fkwlv3eZDKPXR0XZhz/jCQhj
WE4oqIBg4rZDK42VDTUqe17/Y7xA4hCKfKBt/i4H+iMG/eT5D+FE/Gb9fldnwrFzGXCuaOgc9Hlu
aBQYh6VW1ee+/NAj9UgpmruLkmw/0fLDHyNCLeGJZI2Gwlu1CPDIV6N+Wb7MO89FO+BMhBgnZ5hQ
MRsvk0tQdY1u6tPaBktsUFdh2DZpg3vwzKuD7QZcaRwgZBuU2CSWcVkriaKuAqu4Ek2+CsIFHrNa
6Fq7vM5ffyTN7FYZ+JAZwEc08qEimOTieCzreVJ6fSb9Em6MmT83Y+eUvQcsqdG8kMyDxwsiVl05
9aWX5jqlEkuJCp5VlaMhESgj7tJfKGXL0hmU4+X6vfmtLhRJ8YsWy0RDoSmPwhtQP9mMhrmMhM6e
JJP+icQYiQtan5VJYAEW8QDUzcIpu9wh8bC5VcbSwlczyChRhGzCeQ2/eIOjjB2APOWMhWI/7nuS
50x39GwlImpWjLpz4qUHvw1zB7lBfEpeVxIQSgBaFNDZszten0lz0GzuDhCS/4Yyhy5kdXXatw03
20J+0LEbd0OFTRHMo+Hz6Ww680004WjV/ZR5zUizyHevAhkX4jWcN6wqmOflnxcQ7A87COSkI7YV
X6TvhuK7pVoPVEwcUYtksHOhg3bPZKGeBaBCCGnIZGKsYgKOUMT8zJYSrEamed7dm7OZLSfKhNe9
3Xu3j9tvuc3qaZjC3FNkTb6JL2lFkrnjSRwIgW2iFedm4/KFUzI/AO/5JTA2FiP8lejV7cw6nIo2
5/9HmxBx6LErVpuotXIiAzQsi6eP1CkxvV5Rp/A/YVewzC2RdMx3/bfeSFbJQ6140Ied+lmhtW5J
AFrwuYubuAs9Oe7nSFTs8xOBSQllp/yhXw+Du6c8v+5VsO1e9QpPWM7PMMTKIauW22r4HRgRnH2p
Aphz7oKwYYUvgWZUf42liOromRHWOVW/JOJoG/U8uz41ewAIvzUcEJPB2eYQNojdNRgB8Wi6qoyF
beknedCVHB6fg0zQgqX/U4DDdTT1vBc70hoYRpBv4klU/FhCeXVv9sM84VkJEQhd6NyI/5uWxy+/
gTD9q6u3nW+FEgb6G3AJLkKRKfkzqRT/XT5ri2hYyhPg0nxorCBCGvZFacVu/4Sa6me2Y9/+h+Zd
fG6LVcLYP5iKGSSFNQuwSOHZk5Y3rxZ6F2hFgPLozUaXlaWQkDQJ7Ea5PrJxIkxOEiKGi3VFhGkL
j3/nSfM47/XKG/w1YBdgHhIKPtTCr1xieqNaJB7z4Jb6f7BM0dYSZNilGyUQrtf0wp4kueE1okiw
hLUATd6xFWfegRieKzuj0792WZ9yKjwXdwV201Jgq84nOCRtzkuqiHuIXT6le201EDwS5o1HaXlB
sjtZ7b5+SUVZJcu74ofI4+2D1BhtEnbAPwfoRFE12bG07AbzqUJZyIjkbx5cshFabpMq8B/e3514
GqVTR80k2xPqO77ZDTO5WxnUQKTNqI4I13hJmtykkwqwxIlizT1wFoJCa7Skra0ObUNQFRbb6rv3
7HOnYF5Ov3DCa4KJl4RMvVuOsSSTuKoQ3twW5/8G73ON3Det/7RE7Hg316QF+HF6TlSBqi0isvSz
WlNmunafp11ymbrNhkLesFb5HGv+6k/uej+q5JdJ+YALczKvqVNmQbjXscOBJ1J804sqa1jly/hf
PT09dhvrBmKVAOALYWrn7UzJd2tnZsZc0Zrk9CXwpKJFBCrVRcf9PzMEAuLpKI1PJ6ytb4LooA+K
mO/TcH7NTf6p19feLbJ7VjzB1LAzwxBXpSNK7JMEm1t6MJEZPpNqTC9AuALDOPjPBxeBPNgicBPL
szcVc6lR9yI5pLtlnCCsBizkxivFB0O/XApXltoqwKAxDJx3vQAhNz0H8QeZ30eNxM93Uao607NH
B9gJlh5i+H7jX8xBHg1dwpQ+eOBqU4gVTT0mlq7rbfKy47CRZT3Lr7Q+9kAcBXiAAgjnBpKxMZJj
ZrxvUli6ILRpLbp2EcSqtQlCbOU479HmnVxA9LPnSU33vM1YOyaLginXxWoiDQpvcuoqyISBZEPU
uNF0rfH3MmuyFgWosfhC+pkvm4MJPFF/QUkZI/Jg2DhpZElo7Y0vSnsNWqMIk7AuxOduFrRleATs
wJKiLZbt7HkI2Gj0PNRdfDwwRsghIAEjKTsBFXDQfMgtoqT/kitjx7Gz0wSz/sjG+ZM+pV8A1EJw
SBikbCSjfxJcbF4O0nxJ5jW4zCu1F+5i7laeGQkcGVNC8NqncDbn3JU9hQzccS6b1qMZdw0bZ7/Y
oUl0MheJxLKOz9gbYVab4SzJbOaA3nM70SBBPCqXIh6ER6b2jic8hHy2eeyml6y8/AaLNDI1eY43
yRhHVhVccMW5bqU+8MFM97w49sm47Vv7BlK9Jpd1ltKFzxZITuRkGyVg50IgKbMoRm2/1BQHpMb9
vDSCwCKvaTMihllH5q5aSy1R14ACcQSRC3RZFDYDew/gyFYR9AKIv7f+MIcPtckIPNn2RLlKoKBI
0+QvQpma5SRfLHuKErk3Kt9/WB6VEQ4E9bqJXLzVyLJfaIdnbwbtBC8JXxDMXAYioSN3DyncRFDo
pJFi2yu5hxjDX1OD0H/m0o2fLqWYV3VU70599EvO1BYQMD09XL0dSki62pPG2sOtPC9Zo5ehYZXs
rQrqcHtamyzOh6Foh2DV+S40eUCvycZgRRA+HaxLhBI9YZ5aeNmoTBHJtvYubDW+sbAA5sW8fyUY
X2HM6LR3dn0Xkv3jRSN6b/elryBvATvGHTEee0ZbqOqgAHHjUDPKIKLYvA3p7noytFx9zcFxKIfh
ex2Am/5o/9O6vgZtFiYUkk7UWqPeFgl95dqfkZcykAQHIgWM7KAIFFR9EWEMM3qCuk+hgzYC0TpY
Wr5N7roxfZnaeFfWpWNNsRid/fmVXGEsJ8xIdQltGdspG9JZ55xAZfTutmoJWhghnIcRhs3P1u45
EVTq8XvcQNm50PT2MGpVX1O6R6sPnM3CtCq5R5stpcHm9qAzPCl7V9542LLJig+V98nyC58tiR3x
DVxnUcVV30YL+Q3HmQxnZMHrGQylRlHBIzHzxgTp5wxlEcc0mFiJEfOdC8yOawY6gIEUVie4ExC+
+9WIPGgt7W/UhWGAYi/pzSs20FYTdEho7sbi+PNA7KcRg3L8Isd7Ig4dj/L6/MSEskhu9dcOGbye
PI85cgaBGC1RUIlFQG1FhDeTJY1oSCT2irIp6EuD6AVl3WOP6dnlp/RKznDI7ypVCR9lTJ8GIjKS
JkiEDBw76PSVeysHCZsmDU1Mp1PHrVLGV0YCdyEoKYhqBBXlwcsOLJeiwKaES8IbkZsz8c3Zq4Ug
K+6ELimB2CMXxVaP1aMtdg8oCHOyIkoXcKPBVcRNYBtgn5Z2h/MS5gS8j1t7rHxpjfHqcFc4rFZ5
AIlHps/QbitFG8MShO4BTev9MzxMlycWqbePrx+IHsKo28BzUnAgwApH6RfqNmkH9lNbUnspvsEb
Ae5pNz30sqfMV9M913itlwhQDPR2iGTAN8vMl/PxLay7ZmHOAe5xkpWX07w0LbsaFRFykO/mDVah
eQXFxUTTFXn/qe9SMs8Ol0Sh1pZU5GgpK6qAoz6um+AeCSpzv09UWJXx1rLwH+Gg8pdt7lI2TxWx
CNdQ8/PIArwSuD244M76obNtgWjJXbi+0TOf/CMyRpx81t0QMGITZ22EGGP4LLThQJnaFynyRala
CcAwcpVQoZ+Xpm8UbYMi0eIUCqoEpdCdDXSb1krlPRzKEF05c0gVwhlVCuTnxNqjE8CgpEdZft7x
adeBfBbH5PtQQ1XXGv3KOehJLxfVMv687g+KdDeJlvorzSPkXQDm4UHrDptkNzROJWAOxWD0+mi/
1DfSCbTmQPp4+TTKvVrCqbf9QNCln4M7fLhU9ehPry18IAbRCnRxJaoaIy9rqSYakdZvtQLZ6PKU
SS3Vm09glIBY/8a7yKyteA8xWCmyQGcI1eHep+ta4KCgjN6sMzuCW0RK5qWt/FIKE6gckipD7lou
eUCb5pAGnxCs4xKPLehpRCpY7PBhWDKGuTy0bU7kTO6xCzlDhup7xvCBtyNcQjrzalePtUByPxku
OCS7W66OxHf6MQHcmLXxZXWP7UafHLJVK9FTODn+92dE6N7P6o/DXgwRkofakCuvpgGJouzu5U6r
3NgyyOjlj8TLl/WgX6ZVk+XmEZPQxI/Rq//hd8EquKC5xAylLgQJUDL+I7MCxvDBjp8bIotwJbBf
02SQ/1RFYvsQOhgHwUY1JkC7upPdV7hH7sxV1waroqDuWGvz2+n7o9fN5ypx5YiuMFRqOLypgg50
AzeqrYf0Je8D1Mlk0y9MlKPb1Ukmg/nf+f46XGSa+HlU+gEQA9TFri27Zcu/+mvy11bmAHnxVErz
OazQhv3SzeVtk7kAYI2iJlgFY1BwB8NVQrc6E4wOl7DdP+AkvEIBLVfDnlVmywIEOcAcR0aEJ2Cv
YGDeHXen5+klFxKV6WPd14kMMeMSEMDQQUz7GGLqFiyTi4HD39277+1elq79XlcnIblEhan6btCt
tmkGGae019G6YmBDU5JGvWhvequKl+clDO/BICxlv2Nhu4kBx2A/HeBgH6b/rmuQFxWuqB1BSv7D
CA8JYbeni6N0QR9BhhwkibVRTjUAfSTKBzMLKzd6elkIKLPVMPp+QiGOPizBmEmHP6fwMb2Puvc0
N1Mt7x20kiIxs/KNKpZZm3Ri5ihjnEV3mbQllGaAo1zdYNVW03+XAbeBcGHEmxngyfUmNVob3YaB
rS5Pjrsx/FAqTA+8fzxKoSrrAqGxq+rFQgmYDelpIc2fn/d0hUODpbzHCUDZ9ayyKnDs5RlkSibI
7b+HWtrP1/rkQmD1l01hQme7GwcLfUa/cRPKAuvPDfY5f5oYCEV10GO7ejfEF5YVJg0hYs23RoNv
H9rRARfxL30BV50bVFZPpGILLt9+/JfcOtmUX0lTkXyneKYEliYvsbWEkk5SxT8znQGX3ni9wdpG
PKD6ZrOCVs8zHLVGdjtIrTyJwIcgd92qyloutUasxKXhkB9xFZOa3UEX3yFTBr3YXM0HKVXD2AHC
J/md/yNnhQY6dsH0OH1Ixn8CEn15elPha5kn6qHGn4RmqxlPNTAPPE661HsuDvF/nr08oaD7OwaL
zfCm7ldu5rn7vc7AD93VCNfG+teChcokj3Te2M0WLj6ZxYixqEH3buVgy0dcGvNKHGZn5J/Fnp5I
Xrl0VWDBetwAz2pjy/EunPMHjjBHW8+/3nYE6UpACqMbTOC2LhtC6GLWHx22KgdzJeEqtKxe7e13
6IXd8IHUB6CqEDdBEMZRXN6JXNoVzC0fYQrKphXYA0WSUOOolUxNRVrbmYcER5fMpalD6Y5HdnWJ
ymuJhA27+5jfLUgG6rn5uZFAQCkiT249AxEDhLgsvDrJ+NNoDcFJXQcafEKZH6xtSAzs6UVLw+1r
1qMxHzn+qx1bzbyD1azgprWPIyKh9vsrh+n+N1oCaT31Irdvd5KkHHLh5jxF6H7WIhX0kylfs7kU
mrl+jFFE2NtX9W4UR9/ulH+JyHOMHCU6y/tzTwti9v/DcjNKCdVz0Qm43Otx7FA94UDmh6mzxrHK
E6xxKuEFl8b0eIux0VEeZl4oT31DtUgphpeLBuRCeLwbLUfcP2Cl6lkivqoW94Ma+5EhG4o0wTWG
h7Fkf/S7srHCKso34iAc8Ub7+XCJk7x4MuATkwie48qkbq+D8nyjfcGISJx/BDSsI9R1KVNUqCq7
Y4FvG31/weNxrRIn/mKkzgP7pCyYSfnlPHHfPv9alMZV+kywsR11B7tMK/mDxOblCJ/gZwyrr3Xn
RysGuG/YdoLe4diISHoqxg0WgUXGyFVEt+lgoJvr5P9/a7mMIla0ZjkePd+LMo71ghW4GF76zBkt
zkEPBHRGt7KlGLbzgclPDphYkCI+NtaUdqft6zmAjqKwgcma9WmIS8b4tRXEwTvxpcEpuBjS+7IB
+6h0XX8tZYnSfmKGwedTPrqG5D3jmTyur3uolqeWew4E0d7OFXEBplsAjWf+xo6UKHbPNzyXp/cf
rVZextwbhealYKxN8vYlPCMzhFAJ49GN+8R4a/LXb28RJe16u8XC2gctG4ZlQFPlK1ZJmXsgmKaJ
4XZFGfL2Mt5W2Onzq3tF+qeq153O13oJlO2R/158VU/66++J2JFYvyrP4FMQLJCwvd59jkHcFtoV
Wdthd1a+p11iQocZHVwBsqQp3yfdTBMkHviSN7eKXJ+cGJSB6m2ux75ToJF7CSEtlah9gfgvPufV
HuwX1OZdHO+kvO89zBCbSUf7dNGcEiwS+tebRMOyGdeFECVUzMuj+B2A2MaVwz57M/FcB5jfe/O/
babmsPjMNig4fsZYzytJ/01aZSr3PX/gcuF/2pqsVad1t4yIwODqpPdn1TrRwsenMe2fLTN4Scim
5gskszPuAmrc+YtBOWBv1lAuvc8T0HVGCORFuaiD6wzPNDEXXWWaI9/I3YogjCAl40PZBnHDubGT
O1MLx3jgeBaX4iHiSenF9vYiODidn1q9qQZyJVGxcLDPcPjkdY7IIAbHqKDc66w2Ib5inm3/xB/k
hkpNDhQ1ioY3rm5nObdZ24JKi/F8PGO9ohPQONw/1eOS4DjdofrEocRjNyd7obgDuu0l4EERIPfX
3i8aOXFLV9s7arSiF0mslSssDo+wf0FlVHaMSPOahLMfcIALGBg68tAvFzLvJa+gWpDWtc6zxCow
qpQuCnBSQSzK4H6r07oXrq81ykLm7xjR/WTIMWzpMV1sszGPkWyvdNb1ovlKC+5hpyhEg0/bsLqO
PiyvtQ/Em55Ccdj0o9QBsmY4YB7AIYFUwo3TmotbhA/SgIXm7JLcvhyBq06lSI/KySIEthPN5OWm
8CBcCG3PaVbytohmX7fSlnoJSbKy/y7MfdIpoKJuh7THNEfAhoKIUfH41lQEj72UXQ/3pUIWCDIQ
I13vVvgrqCBCO4padY4bEykk+ftoN1XMGXMy9c5Z6bbpXSa5pr78BMe3Ub2a+apcrnNtG8X/e04/
tZKPrNS4Rvopq9DIbcBl7bzkt25IN1isBy5LItULjcMjNIJS5aNu5hyAcopwxntFT/FiueYT2A1m
sxX7DJHN6MzMCy6PDxhI598Zku9HBZ7gu4vYVcK2m/B+kv3ggW5TF5ShCjgRKFBF0pTkzaOEFrVL
XebgHaSo/kttO9j9R8r4NTNRpReH6jXmEckk8dgw9p1px/KvdkXcMTkCOWI1I27lNOqLCSsTJSGq
z9TB7RZL0d8thj3qsUkq3Vzi7GWUMqVhaPH3UcM+Nf9nQYpuMdzcQUhYJ179DszSlDSD7/YlJ5T2
TlSeEHyE7k8wHa6xgJrh/u6k5tkaPbim577sIhU90vlM94UrsX6Xoq3WYO0RL90LWt7ezXRPTowq
b0sXo+RAG5Z9eQaxtjHjLkPDV7udxSzmgBBPe55iru7DUK/rcZFigMcocGUGyEMGVtTMDMldPuUc
ae/RHejxdDZe2xxcdD7CaKapJrt+NcJFHxKoO0M8ZjdvqhvnRKgVTUYyVZ+ZaTevTxhmjrLUX3wz
d5IP6Dsc1mkPsrR2lIeEaQC+NA4L8T1TdKK4DfZtsYwvCy/96JBC54HuzI0jHvW+T/bCiGDm+jd2
IArSsv39fFwvzHAhGeyp/tYgNkl7AuDtUXEpKMswDD8YBhZnvZYwZ9Y1uzMHl9C4LsTL24CPIEb8
mpG/iGecR6OIX26Rb+1XfL9k7CXUjDxSkjKGJPB/8m3Vs2sAZianBnZawul/jAybDPkY+T62Rz73
Q1pFlblV3YTeUJDb5Dqq5cSgws+BLc1TA2S6Ia+X6TwpWsUKjPwlVs/37a2PPROdyjLFtomjhrAs
Bfy+oD9qW9ody8ushSddOkFRUVIlEn/Q6UlnvIoE79vY0xAJh5RWupTNLN2oyviaHG+XisrX018p
QI3jOG/LI2ZLSLdCSDcuIHSPiFkgl8DGHJfNmUVQ8rj+yZTdWQq9WZHcw7giDUNa97LlAO3Hys7x
G8A2Cf075Qt04VrXKt0Ye/P8RlnnWzDsSSmoTQG1pEj3YrnSmTaiWpr5CDzyO8S1Wq1KnJmU1M4z
AvUMK6KaJH1xuaqvCf1LhcrWz8J+9Jh3BIs8wv5HCxCb0IbizeK1hVg3ZXO3VO6DDTFaK3h8pxg+
G2+CfuOR/Sj+IYvSIDgXzKNbRxYrCZFo2RbLi4lDD++FXKwyf3vzxgJr7bBxjnzCho+HklikoRwJ
WICWEAauq9gDv9NJDLaV+yzGjgzcLFm2w4OlEbpyTWOUgIPeFlzFRLh9vHWyxt2KwaOvcHR9EXew
zzI3TYr5De8V5xRuKQGbodGrOKmngpkq5mJbL33hSNA2/+YR4ccv4aLpXxxzW1Ire0AG4nXJJbTt
45W2ooCAQ5IaKVJGKVOHqX8BM++sbzW1xrEox8SrTKmatZ7gFJ84sff490Nsx9IRN3PGNOrzjv97
EYDrzxXEXtnKwXVhivz9U4g5Om/b3X79tilRhPzn51Wp8oGqaBntzD43BBb2SYrQ9PNZkCEgTDbd
OQ+qNiOQ4nMkEsVvJAHtuvhTVyINkQo9mn48P1cgsK+82xLyUMSbAv5de/5pspwRddd/ADTFzsnM
pFr5BcZDewAiqOGTNLegcotGoi9W8CfOYKqWLkQlSFczfIW/pRKJ3kOfaQ7WP1uYNTYLE8JqbkIs
RbD+8vd+B5F9vLXqjUubQUN6mJIy48CS5uPpHIctTomdjB+5GPVnDbTxqjijygnxTUYUM4CHgZUo
qXnTSfyYrJTjh0oQ1J8d/PCRUUYQp6saH6rlCXWJwh32oZzgIVFgdcnFpc/yfIsSdtjsSOBZ1hcb
8jneTmuwzdiKnfWnOKjkt2XOcaYg4SgWy6jsz/U/8iZtIYBGnu5Su/VBmOKQXtkcFgICwjhS4OmO
S8H8tl4cpEoUr8yiBXGHaqsdcjPAdqgdV1gQDzgXYeT8wdTiyKjBCD0WckJ7mvBlHfxctHeelLgN
mPNuoxuqEGAM5lMBvS1SL1A3YTCXt22tF32oO6jDQ6MarG8aVVEYx+TH4LUqXb7tjMH7upW21nII
VqHNjAH9seAzK97fuuQQVjmx0VmwBuGd2tG00KvJnjkoQP5SAOhMp8USzZBIIWhOHBR4glTAoQF5
X/+MtROz3IJUH2k5Mmvhsj1tC7icxJR57bNYe6l8DdCUn8KTCUSNc4S4heSIf10OFtb/ZsaIwvqU
vM5RncsLYO0dcQ0Cvjz1shyratkOlmqTQobuzodCo/62z/O2N3w6HCfaiKjVhvsFnTYOE7p8kEXM
jHFWFCsxpdh6jio8/JtG9FDQ857mzNH4Fge0huhG2dyg8QAtquaBhCWEhATR+cGGHIIL5MiTM5JX
3gYEpsaxvo9Ss4p9+oJKRcoYbP32A1LIUKAWLU2olX7sYrkqmnIpD4g8OBnYCPZUBzpMz87Va6sf
tFaxz5rFlhSdsZapZv/vQzYlnmDH3lfwX48aXD/Q5KnNdZCYU0hENC16JJSR9IhS/qsZx+5Wv+cQ
PyE4zqeFA/p4iKThvM6suDkXueyQSA5r3AUckLfUwyiTn3EI18SIvH/iZDdUSf232es5SnwhdaTF
UrgdmiekZJ9fkT3BZKtFzCbRxRvRXbX7b8OEDP5tyVaVu6nYHIw3vsz1rTnlRjaFkOTX6WVNN7lZ
mCoYkOL1O9ra6cIH0dLYRls/te40dgTHfbKuMKIhKLcYMtdmeg/5iakmFoP5CadbGjtg9ems7jb8
mIqnck/zyNnF63RTffBXUy+74MOyfPwlSjhgQMGxffARQ0JxrrwDxF+PZn5K/YormJyZn6nKDII8
7y/ybeW+Kbm/MLQH+EHrkfQdG3v2mmoVAmZ/eironSonCqvtpDYqh+iMVvLEAWSCyh17IGeocW3O
9E+VCjR1/3xzpJ4ZKn7OVVXDuWHOx9S86rxxywbD+5vYvOZ3kfq8Ww1qrGy2Q3ZspwFzE09w6mdt
w90SKzNhDPMtnHbyhIYM3h0diJOW0/37eN0a0LFJt4gLGTPWgX/LVaF/RgoeOwQ8+VW1LcewQ494
nCu8VjGcza2GH47rprjkTxnKk4oRdSSEDAYgQXgRidkETF8S37c3GFSEkvcNm4SkvftEujYbB08T
soDDde31ho40+sCeocyjH6g6pJJfZwf5sG+KjjoGBRMAQhGbketK2AkRstmFJNEldmwWI6zHhuNm
RCmFLbqEVcJHPSPkemzb97uW1B6nq23YXL2Kg9MksrnvY0P91IYeCVWQcUXc74oSFM6h7XO7P1XB
PrDLZH7IVHM4P41bBlhoIg1j8bzVO60NeK1alFMHSo1BQbcJKSyjLAd6mqBqpq4JhHw9esdlUlFD
kETg/gUrhLUlFGxJNcPn6dN2aeHropPzupUftLGlg9s5CDwJOqsF+DR2RfqPxrsb1NezKCQsFmsY
1RaufuMUg8CuzNwIX5sOrs/Ys2Fd58cdeXQS99iwFZ3UuZFPbXOiViFcppYoMMWkO3GdtssGjeni
GHkDrZBymvsBlpE3aYY8sUE3nIyfxkcUIMzM1s0PavcQqegHM5QrxvBVFW5dwVIC/Rq1XMFY4LXY
eeWD4uOdp0U5hHX+XjbNhVx/L0duMGFLrsaqCMRPV01YAe5wETJIYJnwzhTlGYry0G43AkT8ksqG
7vRwG6nIxvalMKTvd2VbBM39IN7pqZSVWNVEq5lvSggEr9Qk3whoR4CaB+RI4xYrHgOSYkfSGmUo
82Yn9kV7J9ttj1uf2IJF4tJTYazMFLYB+XJMwtWTTCLKf5JxF5DBOfRvMdGgHdsdCusuOlczaNb1
RS9r25msArLk+k6CcnErwohjM/DzD5R+9XHF+uMCOJ2DoTtLBFnsIIpEyZHdLcqY8TmQgpmvGnD7
58dv8IEQOBs47OrPXL+siOhC/0RLT3QZ4YSra/cMKYS26j7exFI47hInX9D9pPydZEJjNtMmhIXP
tJPb5sIkSu41UC2veVz4ArOpQgtTLcg7tkhKKbhP+WS98R5iUBhid2J1RlCm3mAo7yF6vF588myZ
BeEkCQnJGFQp6WEzmU4bCGRgmrqVyDn2Zdmxhu7pVPOdD6f9DyQqFkZJEU9AMZAIjcJXR+FCX0yS
5UaobWDHRGacizr5lRn8JZG3Kbj8/5ZKaqB6i8FhkyBAAFGMKwZ/maeK6ys0bCVuabQrTs4ZrBta
xBHSJiTT9f3/34ltgQ8NqTptA5oZgKhDhz0u6sit7oqbwZeWLcPdW9+8zie9zQrlLMT/myNq//D8
SXfpveoafPYtayXS1dZRpgtLZ+H+2If4+QO+510HHiYPOEViCT0vloZk1lAPptCgN9dObQ3fyvLf
YAtdjHk09LnAhtVrJrXJYYiHT7I+0JKRyUxyRfdYFdLI0OaMj/3h03YU0TgE3OWC2ov7Z9C9+3cc
3nwcHU+M98zUC/HQ3kBx9fpuPR4Bo2QmfIDmeh8Flw3WMFEL+9LaMRyZ9cvxSCHh7rLdePzIUyfz
oVeI3ZzQaTcVrb0oNr55KpcpwsFaQ5+akq8irQpLv41zFW86IyDweWrFdNHmeTAdGh24guEZYHs1
Y0sDNteMpUxn5PDDik/UBIxrTf02rruMt2gXALzCbbdY54rdP5r8mn0jTwB7RJdfyDhDjgvORUke
B57SUw3g2dnNYXubJOxX45+7d/Kf/U6GWDIw/9Nizeapvxt2N7Kw6hvVjy39eiV2qLTBC0NWauCn
z43qrUWNrAwU2utEKK9wbW8hfPqNEqIcKVIjsAQ0kRM3U4Ru/lLY2DaskgGoLZjAtN4kkcRpGYd2
1oF/SRT16und6qP2cIotX4U9U5H8jrD6ihgPCGUkjUAwHTSkuHl5sWMQUK4z79tk4Ibw3fxcKYq8
Rb6Mpc0Zt73y0nN1KJyVb3mJV71vB/6VgB8mTgMCfLgcg1VZSv4v8ymW4zqqpN6SqyoswwD9JUU0
L2cdVdAZVHkK+rkvOI1DCDwbK/q1E7gjnSV4zZ1oCAuXfW80snHJjeHtRgE6pyQx66EA0yNvji3m
v33CP82JJu6vVm/Sa1REXVuNhw6GNTJevNI+HnqEt9eppgtv9Rc4YUilX+ZPpnpHvZzYdlpW27KK
iKtBN78MT16oljrXSUi7YXELEC4ZmnwzHn3i4Qvmp1If1a5kEXIKlizr1wRXBVbq1nzBp2hOy3DU
zL2wpaQshBJ/wpCUwxJV5wri9V1uKu9NRsZmTDFIE6+MZLrt8Dtn0DWyaAoIa50vFwN64asC0k+X
eH/wvyUR7nVTfkTZ0xErE68Rv4ZaNRvxjMBDSYymirFepB25ouGAku2Qkp6WA2xMXgVuJrG67X8/
Ih6wwT3M8fJz1tf1t8tphyDEjWEXSQknVo6wQomVqzPx3zD4nNIt/If2XWEnwHqiYAttWm4Ul0c4
RXHPdcq5iKoxewi30vSBemKj5WatP90kitw+O6ADO95oN9aO+YmfSINUX/Pu+hhhcN0h/m/V/fyb
pAYiNAEa1SnqTfkPhxV8Q24ZJon7eGaxbTw9UwG7dg3xMjuvgmLxTucE6TiBdB/0tCf7pc83vOfz
8MvARdM7+mzuj6ce/NCgF+dR217mU3BTv5+ED8ZBUyQ6ydx89VmvlxSxHuIK//CvZncyx3vkOzjl
VanfJQnjFCuwc/sx8lgQo/LRjpKW4emSoPsBZq7eR4dt4LEMSWSVde7Dei/DD+0a86Bn3lwD2ntf
6rGgwSsBSeEWaO22KyhNaIJGpM5g/Wfwlm0M906Yenz7n7dIsmOATyzet/wM3H3I5cujLMzWbOKL
u/L6+eAfWBLET5KGBGOWeUrUQyHpOsaIqZEG23DgeN9/XjYSKyihrA0L+LD2b9t3RSbn5zHXzh8d
pVUnSw9eJWV5IcrN+V0nw+95hMzjeJCEL+CnMqKcT79sYTVOOQBKJlDTTFAhZ866Sl/2+mGrtkzv
1kTFtXMyx7WfZkIba5tlo2yHSIMrE0g3qbTvcL3my2oHkqCQhbOf/vA/zY5EGm246Y6stb47U5Ct
2u9zYIO4zibYRX2Pf5ZW/p5laNMjuSdOTdlpNvZcxQu0Dmqq99jT1hVWBC0T4P/P3oV3gLKrAU+6
6dKMf5XfhvXm9cOivjntoxlJMAoEU1o5MV2n5o7lQ2CECL2ThhjtX+JdsN2z6WcIWAGc9vHXdi/4
w7ehb3hq75sXn4CxK8DxqdlFV0DDlZ5V4fK4AwnZ88XSSNVVslAxgHhv9lprjVoJMnNoXdTVTzwm
jtU2c6zoOaW4ZY36zje2P2NYHkrp9dEmH3i1m8RNT6w2IYHJrlrse9197MxelImS8xkNIMDfc2IL
jLzKTpHXKoQ+gwfuQa68BNNpcprndp0Yji6W+X/1IIgBSL4OkCb1R4OLGIHIUop1e22MU4PasZSp
kINOQ+vfzfLmj+y7JuRmlrmSaojAY+DOZ8UayHFzcBDn0PY722tJvIUVlqB9OYS0I4Rao8W1z+te
6W9iNtDyxajrZI+t2sL87SWNHbgYxjeraxba43D0Mr4puK5jR96wsUT7udMa42cbKG18JN0SbjMm
sqaUzL0Zin6HCyRKN/RRKxfH1zK72zaKDFzXpGNO6gvaRvrBODzcGoyMjvuYrSiVfg2AZLVbMAdv
oFbj5cJRuortwtHqqa0bksEtz+T4OCZrDICEXdQ7KQKh6szNv4LEUZYWQC41SQDVsCFykcENWUx1
2J05z8J4Hg3sJcbbXj1/oiL0MTDeZ1hNlwjW6/32kC7vN5yNqACASiyKlsS65wi7TMndCp99o/P6
z6Nx5UziuNmliMOthHcaSVgTjvjb1N5OFq1IW1Ytj7D2NNGHuu0n3LR/aEwx5/y+zxaKCarM8Re/
AdJYMXF9hLzNSsuXXAqvKbZxcOY2oxIAw7K/R7eSTkUEdujC0gw+hRMbSC5TsrAmt7ihAfS8oMuR
7U4N4EoLymIbdTe+vvHOKxW0ZaxfsSYQWmLNgAm5FrI/Ua12CmItnjf4JWt77OfTKfRLYdZlzsxA
TdifpTs4UmKD/QprWhOi2gOnq1TPMDWMYqcVlwz5HGgab1Ui/IQ/vcEU5fHaw396MvbmQVntBAWU
gLNpOGkqJa0h1CdP3yo/8hPBKv4HHKwUdN/RM4YEud5R3MURe0xV8MU5oo6GpOhCyW2Yfr38hKhm
N/WQOVVAStDBxHVF+ROgVfdyxJ+oYR7fa3bdv6AniEdQZRGbpJ63ZIqKI7BhDNCiNSe9FqdUgUBN
ZbjhdSBxnYVJ+Xef8IbIlESyOWSjFU4MSOFXlGtN1yTnFd18Ss6DX2WtXc/B3PfMehFzMCKgpFhq
UpYSq10Iqexe1yWB47zbslEJqAn8sfnVyiGKT7ErFH2pqGYJ1qKr++fAJM6Nzq6mP7hGiI6W2oI/
dxuLJBZ0dwjYTbIEewWTdj2f2LReHgZ/MsjU/iJGC1OOTkz0+m8HIkIHkvUbmvUPV7Ma1zf4VLbj
739IxM0hjDDsk6vU+0HiTzyQslsPkJB4UvLPWA3V7Ce0K3HVpRBUFL4mFtuC4r4loKJHef0J3Dl4
oAbK7K7l1Qcvlg2wVa33qB+TPKenQuDnbskfxmNPkHyZsPDaonbbItLgPq4GMEgJrSTRf2Z/L1u7
QQdIfLUI/Owa4m6G2ror3y3OWO80u/39VAmox3GYHZQY9ayZ3Zykti6jz7vV12xhU2OXh3Sc3D9M
y3OEmd9HtRh+Tji45LV9Tirclgvs3CngoQcwjzOwzOZykT60m03izvHUSvrBbw9QpLxRQW4BVjkk
BftIE2Sycjc9avMo/ai02865GvTckXzBSeahrnd9a6UVszgZEp5qzPmFke3kAC++lLtzbMfPf1IY
23NBZSjhFu7dr9GftFaYD173yeh4pY3ratlr103lJXG32qYszD6rrmpjpkFDkE2+SelHyuZQxCAo
oaHerGihtSc244mZTdXGP6Sa/fyoznpfHDQcuaic0/nLgxxNmI/aRDW03V0fXQ6lPapllK1o9coV
6ieSHCjuj9Pq6rYvh8h7u1Ktg5k7mpyE72yVnsnThVoSbyEsLkauXsdADrQV0aCHvDaHbJgL73m/
ad/2k8GRTulej8S1gBVysgZUWYhCUtOqKlzVfmQpwOGAdsUR2IKWO+s5VmPOplmsxP9njsgtuIJx
a/DMgnYyvaqPRnaFW2gCqVgadnpT24qhGqWv7w3sdm4KVuJkqvp+4XlvOK+sBWnsPGna8GiRkVEx
J54JW0pMoCOlKze18dZZWxZiVDnQdZ5TJILI2KkMDXU7NJq096cjNlCXMyHpBa8EjI5kXYMjfgqk
4kD3XfGY7l+zz0IcHlrKwKzg4NLodho/OZcsMfqqFmM+HjpSqIfOJ+jWh9uU9kF02vgu1IZ9zJwG
JWa4K79/vG5YDFMbFIeDWdz9+LyXAJvnABNTSxQhYLhthj9U0fsNPd7sBjnwaopcWd1Ocx7mAu3s
f0f7fSSMYnfvRpALEubTLfIDbM3CVcV76CesFj+TMDZFqkQuNmVZp3aWIeclw5iEvO4928rbtfD+
zvTEBUWw+gihDhuNXDtttpU9S9CsMGcdxA6QhKErI1awY8SztCVtW2qsUhOFcpedqpbc6AlwMbCT
Ok1gJ7fHZSzZpzvYLMt1rx6INkhGsqd2l+XXSFwaETGu54e/dwUXB2y9uWGifHA33yFWHZIduSQk
iumZ8bxgWK2W4Kvv71Xrvqh5RE+teLedjwb5k08aSJIrdsocVkq1qYEl6rrPqFsEmukd2ioYrBiS
M40Q2Ghnyn4pHw39cCxCyQ+NX3f1sPJNw9dzRVH4DqdmNqzmk5XH3MyRtZPoWwx1dLhiUJsepfvS
Pa5OmaBAPDbu+3JSrcIbW1bRTb3+JCGIdX5dMDZ85GxizUf79kiXgHSGyvqS7p6V9t3XP0fqdxQP
3Ct5XUX/OgPwCnS6EN3h8mZ2dBGOT4mNXAi84MCvrRCBpH8Rh2ZZ1JsJECwrMavAJJte/mVOnbxw
/cEC+od0vnQjx7sVK9BuEuUu/agGE3gQhh/MtsGGjydYjd2FVAb5TyuvASl+VjVN+93nC/uXg88g
dSsQgcjKIOoHt+IwfhwzkaZfE5pYGBIqow+t14MYwPlpfl4qJky/sVaBFeFo9osJnkKrF0qifU/o
FSObzh699iufMc/juaPMh+/ZBPLxDj+7GuMP2mGKn7mGW12GonLnXctekwoFZ+V8DTSw6bm9m553
0vApnyTIjE+kaEtyUuteKz85kqrU5HRN17RijtZAlyo0aAfnfWPW20zjyafc+eJntnPpuBFP+c6/
6/W5kXpADciSfk+qBztOte5hNVZLo2oRRaZSGWKWTdqOPjP62emvL6PlaNiN+ZuHzZfPGNEe8Px3
CuXgwGlV5xoGExDr/rRwCddzK4KI26qEgjJAWQm+0/aGgjRu4umXw8NNbW60A6cNlkQii17OFOyD
+KjbH13P5SlzYGh7XgzDMq3/ceOEIomgG8NxI2GFP/NtQ7oEaCaOKd6vCiRyg2lMePEmQwEtcQ2J
dcexNtKuU5vuGON3rfw63uwyi7+hPV1vWq0nBPyWnZyPkmbv57xy9nliBmX9O8LC7d8INfwQfwDf
jovycuZJDYwY3buBzkv2I+WHL6ax4yEe5MoAdk+s75aJH3PazksHjoPhPwhmzu3QqTHCXPWDqi6o
JhSfKNSgyn/kD2qjE/zOJNlQHDpk0IYRCn5UC10t9QNRaihYAaCB3VF8UkPXuYhmccLrnvnWfGN9
EHA76FwCt//s1CDGCPoLgWImKtiyKzXcxbf1jEL2sQ2Canrd+ig8u/hN9rCxOvsWfXX8wdMB6PcP
qXiBfCdaG9BhrL+tUlv1JFfJf5ShI9Y83QFtDAKeH3LcADekqEHWUtuAW01EPj2+7CzqM9NSgy0B
C/9u3lzCSiE0dgd3do4vett0HbR/bGPMzm+GjjTJF8+A6yoMG+Kd719iUPlY+ovYSqKwk0zwOs1s
gJL63dZz+KHdGtsiJ5bNC3y0vES9FgKHYmGQZiraHPh3EB+rd+4IP7sckzlNYVuOZJ8ShOxhT5mP
MXqu4djHkJZcAFKxkv4MH896IvYvHlcA/IKBD5WKPQaqcJTelJhdubo0H2Jon/jsRLEZk8NHNqY2
wjgUDl63GqyewZBeVqrvC9kHhCljiIN8kJxd7T3T4PVckDGh57L+/e+hKp5LDzzrkOA8s5iCjdaA
CRri9jK6GEEfuOsGEqP6Sdg8KzILpg6/GR/vYQfQNYXziPw3W+Ob+s+WPRH6NzyEZH8lNu3TcAlQ
n2V0AWOr7agEt3ovyciNjraLOPiNV/4ziXYZHL+YIrlTekrp2q6B8SW23UaOcj0g4LCb2iF94760
FdEcMprfeFaGMy4VHTD+xmRVs035Ui+zE/5rEZM11WE9RKQpRs6CA7yWOCv/xccRzccbmNJYGsa3
OkK8wCatqP+jY4v79kiYmS1mB6R6Pg0VlLHNMq2ar9fvrAV99IS7hLjGDnb0swLrPWkJErSBAfoE
zM6yB2Dm3USCYd3Auu/L9KKP/mcYDs9N4z1Hbok79ynEA4dZf7/lvYgZQhKqkmj8vpGFbKRdOtx2
Lj95IQtMc+IWrveYldIFyxx42EiNsWdpGNMdOiRjJ6YInHffhD3p2Zx6qqrrlMnon5czjx+UUtmD
7NUkUsGy6/74GNIk4ylXsjvOSsZoCe/CJFfagHc6Bg6AIrQGKbHRSAcLvY5gB1YbFTTa4HJXU9uh
oPXG9Wfq4A0hCzQGWAnI2/FoM7jBSdoecJGhvfZ14K8B7kqX9buxTRrTL9REIEn8ECR7l/jU15rw
40ORQ7LEWKLqb9u/PzUzJs7peqXZ1gMcqi0fn7Aw2a5dEQhXlKdtGclOuxqsakbYD0Oiw9XdFYwS
PuamJVi957w6+BBM8xT7V/dLbafsx/SQnNuhx1jffatU2thLc/gy+TIzzbiTxolx8JZKdpQEalh6
OUt2ZOJyMSmF15IF/DDrw2/gxZkWTS86EoauyG01BwH23puErlmyhCXd1LSqJ0pyrc/G41Hswoy5
LkP5EPlr76uZK99Yt26gbzJ6yI5BtRIThfEchMv98hXRLjxgO16vfpqCboRzD5MqJprONu/p62gY
xxxwin8juqz1BrL5zWj6NLXgaerphqjvux1+SLGE+lcj/G4WvSyXPTHc9rWFvR7PNXbuE0yqYJhs
9v7xGax4Fw9cuERoUy6RvgJeY2RDxuRixIhkm94BKeL7I2gaQ9FiZzT/Ei3Z1OnKdws5QyppV7bQ
BpjrnppaIrs+RaWMV5KepQe+dGGLbD0Uc4B42faoVsrCFzJkDxd4UvHz2k04XzumtPDOyq9ktqVv
Jd1vFjXX47gIAuaURg/D0TZdyHmD5aWUick1ZEK1cD5fTon2HWC+qtF72mFW74MJ+N1NWfpEyei7
O4RysgIkYUllIXnGtsDFm6obUnkqbROXL9ME1Q6ByG4e+VuPhTvf3oca2rlf9tHRzbokarZzHhcP
vJGjZyMP+1MZ8fLFIeBiQD29VMqMC82u7W9JizRMzo8gGktYgnnvwngR+ynWy/kXSEVHPkqPLvUF
z4EReBUkgYZDK8vLJWrhxyd7oElnlRKftZKRZwBBeeELzupFJF7xNUV4/hxDLNIkp9aTc4O93yv5
B4AxCuJqZirIJBOP/fz4jj1Wn/fssegkjDorubtTQkYFhULQATZw/n3Ap5dTfVfV+DRcpOp9Thll
RWB/94EThS30TLfVfRNQSqIQ3lABYEmcwStkmBadez0WuOzli1C4o85s+ZA39on7B+z7cMU71XTg
4jZzsoezsvhmUQ6ErFhoVasN2hg2pKM5cfW70suSNUH+LGHYyLCW74GwOFySPnP+ZQasRoNWvLqS
YcCYcSIRkuzt1hxwz9kQrAVB4w6wplwpOGwlQSkNOdZ+DjFrO+vd435RZIErQU/kDsEYmtNuv3H7
EHmMLhzUfX7UmnIpkKVFVI4Mabyfd+KbOHurGBqmVTfyeJ9c+3fYKNb/5HAiI4UON52IR5EBDs7z
r1EaDyBH/ezrHQ0mk+2kvLeizGhghiU5hqK40iRXi7yo4qzrHqNA9C24/6p3HLMe2f/jccSgWnGK
YzEV7CvG9UOZwBtiWN0nZs7Ylgm5U2jEZgCoe/yL0KceDIv7TTV8UPgDVZIBAIZHmeeuOAr3Iq4e
+SMDlm2b/C4ldiwH9IY3QlLje7uiO/hnVxM8MaC4eOmO1B5OMmq3LoCgVQx29IcRY4yoIO6u233U
2n9eucwg4rg5j4zonxbXS3dDgUfeFj97ExLMz1gqtheTSyO6cVIFjzKNain+BIqyk59Da0uomaYq
qiPMQKj1PayUZEhoYS1VRjEJTwFzXjlFe8A/64faYUgJ5WRKCij1eYh13PoV/VtIobQFpzyJ3q8f
Q+/nUqr5kBN+dcAglR1XVWCSTkubAD/mGTQXChJy8yyo+u/iNDhvFz/gJl4oHMcO24FU/ChpCQdo
nJvo5gnVgoFCQYTFCD0t65Kz2oIFXKEJe7qH/JodWClT89hjbf/dvKKtwN7+SDEI0caZUujQylTe
clytUe96uJLaIX7dCSVs/TzoN9XPYXD0UtH8RebrR8jRxxX5nOcaTUpoGIbHEHH7nPsUr+ox4h71
US7Nu1UHJM3NCOwjI0au5hbyGEXdctQPYLchSAeH6Db1V7gE88m5RNTPWOTyVJ+3kNzbG1ocM3Bh
a1gGfNn9VLQtJ83vOjGnBcx8omGqN7T1EuUosNgI2IFyqzQ74zvIrbRuWWDEUTjB3Cs6TYm6S66Q
G2IiK8HFN6ariuF6O05lEZIOiwqSvL0N1+l/vAPEhGRiPT2X+PdO6yzsgz0kQc8oCt7FHgrTiofM
JdF3lFqWCL6eqUZmPa62iOy28fW1LNivxbj4t9AoXAqthjdDfs1Ky9LJsoRvKNxjQ8Wj07XgaPNc
NjmUZKDDvMsLwE9vvTAIgZM3HyvuU/2Mk6yfMafjFSN0gfI89ZFcZ2WtslOhej7VlVMiQPoY4hEx
BPzuOMAjdY2kyRwNY8pgk5QdEd0taXMpA8qgG0mXev/5PEVVXM/CXSU65k+prVSnnWwGB8tDfPpl
2ks+ZpSdJdbXriMEHq8Al5a1FC/DLwSxLY8bbBk37yG0CYO7U0SVVuxxoUR8cUkUpOOIYvaeUymP
QhCNTP5paClHt/zHS1SKFF2X8wzL+AoLbi3TFfnAjsy7UPXiaWlEglXUREUK2WiQVC6UlppSyNwQ
tDgzsOGPXdVmsRlFKZCrCA4WLrYDvVPVYEkKdXLw7BAbMKp4IDe1LJk0vbycnCrJklpMyFvq95IR
lGDAf3CazWEKQ/sZWbvza1EOjwe2wkzodb78ifuUg4j+RW7ZioOxW1JArKFeVT0M+koJXsYYNQqt
/IcCoaDZFO+gmodggG8XOewQc9bh0jl+bYZxb3c+7u8mwc1rAJk51xHLXb89Dvcaasj9GqWhH4MN
i6gzfeSRKWSA+cxA3/wTk3FFlZtjRQfTSXBjsLX6ZH6NKahKgpfauJowXX5C9HTRGoCY8R1CGXYn
hDBhxvayqp6JmdLFC7vjIpYqcrIIyM6Dn9BBI12cXs+tD2NDQu5kt4/XbDA+y5YwH3ZZWiFSh55R
frQ/08Q6qosYz5KtF2g5PnnTvhzWXcYYwO9u99w3eI6oKXMZrA8F0GuoYdUh7kF90SdJ4XwcgEhp
MG2SMfG/GGw6uZgac9YYrszDSRRfNBvsrebMxeRm3qj+qGusk4Cs69pTyRgEyZcbGj8kqw0Wup2s
ok6AjQnRwLZg6a32qFfPiRSjjQfyH1pq/Lqpitz0xCIkEudwg9uZsqHlVzK+NpUHpDRxLj0MgkYB
1GdT7bmehcRw1iigXNi7+wIOVCQnAjtkgeBd/RYGNIHbrRpuW4lVFQpl67xA+6i5yeZs/T6huKQJ
PBMCEEnEWAYpJLawBbwkAx9UnZwkFhgemFEkEa6XlyVaawCjdU/sYOnH2QetH+x+zuR/bfrecLr1
dFOe2kMksUq803qcq4zmr0zsw4RsKgug3hd0emlVZjDPeT17Owv7Tj6z7keH7RGZcGXCySmlMp1Z
rtfZ8jBO/QfXE2/f4OpPvttJxpwH/V3kbGRTNAjtKXL7odMTs5p8qXmIjSt0X9/f8sIPTe/4a003
IWiRTB9rUZPpgKcGiMm1jFMWwUHeUBHq/Wxfx8DFWsSkOJwObYjg13oSDnOSYIq0lB/X3I9BfYrq
HQfTey8VJUMAehi727r+jEPtvu2OiP47eFZte6z8zQLz1TU5j2ZjEu4Ro+cyUBcz6b+iEe+2g86V
LLMQ+Q6YcK019DlGmUh3fCa1ox6SPijcJFcVsXnkLkiFTRUHcbY5ET6sGiYvpQOUWGlDMQigF/5n
d0Axh9c1ADjSbtfXkpynrGetM94kb81TsGTWsEHpphzUeg/cmGrxAcSGZavCWAoUFnHczmNxWg5B
UOUhnJ6HGFRdfijPWUc1EecvbMKzYRuZe+K0zDuEhHAab+RoWuDhalhWsAPS4eSBS7R913tNqcZS
Ax/goCI9fZ2eA+r6gNDycwgxLqbJfIyfb+/ftoq+MekW7D7mXDeD6S3+ykMRYc6qHd40DomoaPJ3
DIKqDxYK/4YpJTi8D2qIzinXCBntY490JMZAucYTD7TYgQLZ0ENtPprs+01Fn7Gw0VZBxf14b4Rg
eMf9MiLEo5+wRFd2TMMf5OXvT6rbks3WQYNF1XWgJI2UtU5GOmit1uwrfU1o0AFOUD0pQx2kv6Qo
GAx2f4yjgmlYBnHllptcO+L75jEKQw3M3wst+nAGrozZljjbxd11bYJE6iQ2lJhTPvi75ijrYks3
3Q3rkKrrQLEiFXDFx735BjARDXe9StnEbdGXXmvMe0zfbvZvQQ9k7bVUDGCNs8jPdvaCBWX2aHBT
iyFrDkPjImixipmzRHpWp/Z+gPKejFTdyJ+TklPxKujF4J+4Mp5aaSRqrMbfEMMnd/GSf3O1WjFQ
GkKGomo8MHYytqQ0rZnREtDco6kPjJiPIs+xsmhLqVUoCukRX+YWnMzL1rEMyfiFH53SHoI7Og8I
albpZKarnTYXm1JRJ+aYDX18KxftbEa+MLGOXvJxRpKbSO8qog10XVAiB8wDGVQzaSVoZM4mXIra
oNdLRq+DqFeJYoGQT84GR0rNdFv+L4jTm/rfgBpy+TTRNfA9bUFGgx5GxNqKF8WLltGo7hB4XYNW
5xuT+4nt3UQmRaKsHbMA8GxILtcKAIydhFVYATyN9d6dJe/Glbi/Z8nZFqLexGdB8xQJdJSiL87i
yPShZdKY3ET2yf3CzpCVchUHEHhQCKBQJHiIMIJllwKphoIjDngxrYdkFryyCA24RiDJAi7J2kgn
xzvdSNZmXJLwiPrt+ST25aeZC0lzEdye2NpzxjTdDGgF/LVKh05rqNQ4wKOsTHwnvxCCe40+IRp2
a6Yq4mdJTWQFLoIgHNbfYikQw8Sy+FWspePzSjNsRTttUksX2ys6T1T1JjtuAoAm/s0S5xdGt9TZ
usgl81wq/tjJpOnKV7CGz3g+EFFjs1ev8hIB2Q1MueHbSQKCybuZMcKf7akSh04YIUEi6YeKWK18
yZm3Jja/oxEjmmFzs+qCRSCTil6BaFDGTDsfuXINw65vreqGpBl2ShlF8NPYvoC92VH2gv6ByvbX
gftGWnweCrqy5BaOO6wpIMzP5IN47Ieu3s8RlvUI0ctOJhaZBxdO7DZqqn967/98EOxNyAiRYcks
C0YsUAvD2Aj1Mwjpk4gaFhhsYOBpqCiE1ZhEzE7pPM6x80aEvaktcHlZ7cxbJjG8qIakHafkQ9rS
VbyPwEs7U04IdRH3h/0vKLpcKBEthNn9Pdua1p5CBCcc/EPCBx8cKOxJxI93QYYDQ0Lu3PCHMr98
/nxRTuC0QOycjBEoGhJGRhl1dun1bSTRpLLXjIUAdvAK9zzFNlIlVXgwfSCHJK3Ewp8rCtXYiRFz
cWoDzb9AYMw/MQWVX5N9m0EAaQuLdGdmjzS+WbKbh1Uy4AfQzrjESYISzutC9XNy1RurIYe7YRzs
V/FB6mfW6K8m80ilLoPXdtU/L+dXLZo5UawSHaC4uSyFxeQQNLsAnahtqyJVEs79u3OBKgE6ZF+v
TgMDSPckbY/OR/3vrd0INAkzCjTFCUNDbDowCzd7ZEdVe9220AFjfKxhE+O05EtaFeZ6qIacDH4d
kRlCtt+yWGvNa3fT+QiQew3oYyOMHWIq0EDVx/SIpULOrjfXFg0HMiaXfNWbEWGvsOy2CbUNn9Yz
Vs+TXvk2brdIy04YvsEF9UipmNvFZC4ozgUYceat9k7qvdCdYaBK9pHhfLvrVV90Ff83WuqAAfNb
reofnl8a7RkKrHteb25sAqTp5vsyJ2zlbF8LznxT2GXBGtXcwe+lYV66TzmIn/kpAJWSM7GGxT7Q
17govOPDDtFq0qge8FqcruLXEsO5QG0qiqUh9ScTsOjBCV2B35vqUfc3ezzPoYPtxOxQWY1/ePKS
6dAvnqOYI7pqTNiZozi4KBz073+UYinfu7dj+2HFPhJHhhIIB7M0mWygraA1wCAqBsLfWFcgU0/P
e2NMPHx+SM3eOkfE0aRpda6/Z681r7sNZK4Y7UjS0aAPCOgNleMor2PZh54HSppHVcgZhAoqLoj4
NI/WK15dDrkIuOmLo8kmM/fR1omHFKkq5RIC3MVw79YJuRFTKqdF+d5pU+mkqbAOfJ5jDMvnDAs8
+jyeq0s6NI5+sBacdHeCXl5AcW0JjmaPxS5In4tuPFL963zMUWx6I2AuCwnENcSiJa6IuUwMCOY9
B4BNPN0pbx/oE3GGhtXMz7+R3t0CGyf/nBt708xOOq9oLLi85J4YxUwKKJmRN1bmWfif6krmFnf8
R4c6mTuVsSv2BmUScNOYAbmeCJ4kNni3HidpoKGvkv4AvWHfiMmDUmSdQPDf9/uPn6t1dUuA841+
HzTLzSQRm0dc2EnhYdprkeFpTOnz8/3f1+wXamelhSzhOEjtPja5qOy9GKSOoUZWfJglQmam+tq9
wTHS1gKZ720OS5bRLGSnDfUqYf7NfqVDkG3+35EX/FutB6avlcjDkVQw0W+tQoE8PsLiu8ypoSv1
4I9ApYOOuA9sjAKhlCyLMyvJEkG9E8J7AJv2sq6njqVJMLt6Ns3ypvCW9M7//VYfyt9fV9dKA54v
3r+jwdbh5Sczz7OwCXOSoianiIaMZFgO5Pz8IPxfcDY0ZLt8mchmjzdujNunLOD6rZv/UwgnmkW0
F7AriAE8vG/1HjL1jbsEQBKCxCCAsIgap0vLJn3fefDiBcVY1fWvJXca5YmFHLsTT+F5zAJzStPc
mwPOsEK1CEkTSU8ftISruXtQouGTvuY+Td4KXSiDXQPkdBk+QeILYGPdIRZ8PT0ELLrWdbWbYIFy
zZteqBZ+mz+IEOjyYKepDoXD8ssCXPGDYJIQLK2hgiRoFjGR8fZg9jRACkEKiYoUc+CendQo0nT1
jR4MCDTQY2E37bTHaSHaa+G5pt8I9TD/rQBf+6P+p06CObOIaJA5EvGbrmIbXAKsuaIp1qPtvkEq
zEnYlEdow3nBr8KNVWSEHXJZxexMfLV2+zpL1R2POJz7O2a7CPliNwVUpuJQn97qLujBfI2TRuyN
jk5D10nlMhI9OGyoRF/r83vrYOc0vkGSENKR1669q9Jt379ShX3HqivSVwwiX435qkwUegdb3LGJ
+Ji54c+br3XQpTE0qfgzUhv37pKR63TmSMfEiHhHVeHXmdMh7/Xr2vdL187r7wfvRL4aZgshWSMs
82r6zpyrhbSULxojblOfYSEAYtktSXIrierpW7WAyZqzzNmcEA5uLQrjOfVnzJktraWOb64aNyi4
bhQIMXIPT7XcJeS2GJoFdxC9w58BkFKIMdv+IKfxU2HWPwLvQOz57e0xpvjO37DaahvCWcG89reZ
aaQ8FkSa3EWO60arZKw1jeCXP/iYmQGrOvH0jTzAylw2wnMc212mqnp6a+tZJ/7H8qtTzn/JIYWc
HFkwCEYnsEk1BwG8Zd95xqC/HqOui+e/8KEvNI1EIpatf7+6vXM0O4m9++X3BMxBXrsrTk1Xg+Rk
wPW1bTRiG+AbxpeiZJMXl3dyQNt4/Rm+HawquudQcxS43/V7jJIBtCujbos9rjMw/N/tGIf3CUXn
vegBGrwf1fFdKBllI8fJRLdJU+4qtjdIUNIo5UdZcL0h2mecoj6DiADCBHB5/w+BtCc9Ogn9o6qg
X0zRDzqAIDBwhaMLy4T+46KfdtB5+tI0fWLnkTQtBPxGF0tISV66tQylWPeVX3jyzoLwHUNvFN6l
VfiSc+1LNCSIWUaXDM9tOmM1iesLCP6jT+5PXcddMMTAjbOt7PGxJsz+mi9UsLMwNF70npe9BMTX
+uHXihuroZEABCmkw8MGmoM9cL5B22VmmwF0q3Fb5xCTVcasxE94gCg3OUh++XzsSSUNVQnB0aIn
ixjR1D6/8RaRRgIzt5w2GFFCtadZs+RofpPDH9+HG9haG4SseLAdS+Q3gYd7EI1UV7WRdcyyCBkI
UZQt8TjqhfJU7MqXkWhSOKcfmT8SgK2iM5jokoq6OlGYFycRTk5MXZztmd4AHB7/7pIGS1BNi47k
dJt2iT4jaMviCj66nrKU6lXNdtZqLdKZD9S2oVjhSIECheEGvAVCDgQpH5JTKJ0fYFVAIrmxcSZW
Yf2vZuvJeLzRMT1d4dZBj1/SARzH8NRO7bCB9qeG1JIapqTmVVR1sShWCM69x+JN3Xoq6lB4lfHE
YGnK70gKUAs/6JTb79Nq4zdreMWOw3SSDF28R8GIj78zdXgz65zsF9cZzV3hiKIoT1eHqa5fljOz
CdUpWhEIVwETiOnIDiiy79U3KLFHJ8pv/SWNmYj0f71WVo9QFtiaVRqPkmjAIY14+HI1UllbWwK3
qvQIaGF+waqrP3PqjnlZSDTRVSxynRTk+IXneQ98PHT9IgQP26L4oneXmUbvM7W75L7CrEc2yevh
9JJrWJkYfgUvvC8gYTzCwvGfQ6Z0vu5UQQax3FQURF+SzRSD9LYgSwEIYyPIcOOxBnuMyO5Lx4Fe
L+VGAfnOuffsNxkfvgyTOA88ZDjpfbnW6O2UaCG33CLx+WWiI2OndLvF7fdbpSeTlJoBmw/6DTPD
Flb3CvnvZXYlSMH21hvzofkGsjsxAbVyEQOUGYuC6P5bcGbgVV8pzIvZqwNXI3eh+2H0rqg0s26/
SQD7qeUyX/OiFl3/fKrOI7uEzCl9zWUfjZsOmXGjtEqKN05CW3ybpG+Gdm3yyDi6T7TlHicfNR2r
2TmyCeVGKfzoQJwYJIiG/qY24CZg6k7aK5/PpFceNAneC6tjPKv9Hg1e+S4mGcMK2mOKZwtGoqWS
BuYWRbzEunGee+YxormPgRJK6po+Q8oN8IS5vCsouzUBYdwqPTs/WZLWJWPXnmKTBpHepsSXQsXT
M4J0jB4vCpeDiVnPcam8aGAegE2iSVNxQ/betMQwmvTkVoDUHO7LT/RXmZvqAUi2ziyFLEK4A8sA
TDp4AHtKvffsNe9sdYSJ6ejMjeou4mvWonWD8v/hCitx6pRjjNd62PUFlTR0E7hRrnLoEipgS7CR
MFOpMTc+M8MT2oYO1+jK97OmBqLwpCCPSGYKPDa6jYMZ9MZCgbUXQD8mtOwtcu0aLRjwas8N3FWq
xQciN1lUqEL1s9WmsroC2sp90NeMWzkFsvCVzSDPQptr/N7Y2oirL6XqQgPxRX0E6/mx/W28NsAs
ZlFsx9NB/lccmaatYnD1apU6g/KklirFzaLLLvj+ejl12AR3nu10g/Wb19gQ6M9yrJVH/X5OMtp7
48/pfrMVqakjVR2CRor1/s3gL6p0qyUMJO81tEMQsUABS3JDV0WLevmsCyE0GVmMOtBXzHzo9Bjn
WGAuzw1NwGaiRlE/iLPf9vejKf9TVf8dDec7mn3ipYCugsDO59RUqqVOCuXEYFDRbT9d/88RQpyP
b+UaDM96qaIGbT1wgWYv0/TT9w3xiy8wIOQJKPbjZawwRct5361oXX8rNIvJCI2uhVcf5IpQvpcG
DHRDRL5IFpT5cfa/7ocjwKM11lxWnlMK1f3fhLUeVAOu+cYvHVENQTFWLWOIo/dTEQ6YqFeqczSd
WTsaHIBEad144biIFp0ES/156x0Cec51VSMZ0s17n/urBxsES5ZmVwhLTmNwysY/NE3AWGvXZF6O
KIJe7A09gKNyNFdvtKg247qhfNEM+v+UiDX0RKne79+st6RHV2OXxkl6nVY46yOv9zeDUEvWeaG8
6zH43rYvn3Owy/I8toLOgWEKKpkjkqlyi2esejSYVcARfjQVJzLf8Qj0FCbW8BOxZt6yK8TQfNED
MnSrszxUSmGcKJ5iGC4+8Ov/UADywPmimPseMF/JU53YeB53Enyo/D+ZWBUr8o7ohYUuhDB0YpNz
igahph3EcwoZtEBsI3KCBJZMVvnbmNGr0u4yj5vsTuYKZM2ePNAFXslqYa/VB0KN/1qMjHT6VFDG
3qwITi5KqKP7ww5Xex0+ZI2VpkuSpXIDDDrPA8HY8fJFWNgcOfEmJz0SFhIRDpwMqAS/LVajbvBg
fXKlo2Kc0GbnvgITU0TzOABFa61TOtREAT7AAxv30wOrLf86GFNJ8FrDozFJhLJsY479oOV+QgtR
JRFrLPAYNKKgkxAiqKR6qVGM3K3d4bdIvHHs/1OQWp7oAvniYVTlL50y14QSY4oM/Hp82EoKjSS4
PVhJ98PL6qJIZy4+UUrAQzzuU5ZpKLB1hU6KoBiD/QXKInp2FkTqTyKu9x8nxPp1pQPy7QM5nfsw
EB02PcqwDhbpBe0IsEXlZn8KS6RPK1f+jur+3zQLQxH51Ey1AhXKfMMJEEf7hWsfiuJ/tGA4Fn3F
pB4pZfdK83RW78Q3fLf5Je+C6aGZj14ZMRHLT02CvgalqdD4xW3P0SX+O71N3PecuSRCwWmEJdrP
A88P75mq3IChtX1+TFfqgspeM1tMSHev4y1PGLHqhTRok6RbE9D8xlasgoGui3TSKkgDKExmZMjq
xfpgm5Z2xbuWooplBtX/zUflmQjudbb+M3c94Sq8pWWPdolwh3xt9lz3skfzAJSaNapRQZhS7K2H
GfNjz+wFgc4FcqJYsCzdBexkk7j2pFnQCwWkOu9uDf9BP2yD83fNreR3a3OUe1ic/sb9GZoB/zDM
BcXRXYVSzDRkBDI/BL93sGOwutIPX9mHAsbSYUnxaumf7UEENDh0Og3F4NbPgjvHPlpetCjsk+Oo
gvqcbl/H5ydDqQ+fF6MVB0gdKA3KWmqX/5sJGX7hEi6RYj/f8lcVoNxFpE2QL857/Rl9gPcCK4Sw
n1MQZPIGfxjXn8wb4lHNgjQdD3unsiYW6FaAn6eqKw+UG+Dm+ccLrQZskkHZ+PK7ALJt++GIyaLP
9/n8Wv9Kc2NDhBqgDSq1w5bJgu0u+mQJDWJck9MpMoV65UaksL8TajLjCBqpIZ8F+OWGTiG1zGdU
R/+77rJyS2vawlmo+AWuRegp8j7CT5x6dGjzExVe4wxPLm38MU8ajUWxljXqNZLbOg6iu2oVbi/w
L/iPBoMarxs31Rq6CvW0v/1pijTExrmeFklpgbcRoj3WAM1HlugLkY1YXYHJ03jj0592R2HHomg3
r2N4PmFzNAfeQ0ZFAMWyM7q5Yje0Ld8JXNl51qci7Z2MMjciwq+j/Zh2igAt1cnvzIPvHU1MpdAg
vJPtZh6+OVtoktP0P/nA71hyFUuNS6q5M5FOJvcroRQvcHloPcYOSuLwdDPyh1uIYR3h7vrazSMw
YFIEIqpDOeYDWkLA88tqb/wkgD5+SHHUKUhjdpiE//27zi5IGTvQpF71/FT74zx4OkJm4dde59IG
cfxGAfg4nhzIWyg5kqOiC1Tgmykp4m2GbjZqkzUeIm6q42mKjemymC28a7iSea+XHfte2TRP/oaK
u+4RwPBaSvwM3VOoDm6t6ZyQa50jgLfiu+6qaweIJOM4Bh31jRgtkboxmb71NRLiYBGBJN8ny5eB
yYaTWuGRSYXDTAHh6Czg5k9ldGEpHQHgdJb4UZmARglh5DP6n8Ww4weM6AoGG/917ngq8OuMUIBC
67TMN/gxdMc0pyXHe5sHxweEa1Uzp5uDhc7Jn8SCsU1Bq17jTtxeJc5eL40mp4ssuXzMlOjQr+B9
O+dp4J0EOCJx1+Ib+IrkOpcXSGkvXq/0HGqDEYUHEPPgddY3sxH5bhsV1t6pDb5MvDCV4Pw7NGzq
iC+W7ewnbrFogOZUaQGJu0la/j5IhvgL+sa9Fwt2MIu8RS2Ubw1o5MdjyvStgnibDQjngzlDutct
GXiLQFvaYyP+Fp54YjNMTtI290DQIxVkqT1sCT6JfaxWckZ/rWTEMkWkjyX/9sy+JUrk9ekZ5Ety
XAdixkFYiie+4d/pKK3z+GQLUabkz25PHPYW7HMxdAdSkE70wjBxq4KwUfPDaRyye+zG9jfyc21V
5L4SRr2tZAultuJk9Dbn6gllQrPdycmfLDPBah/4k6bjmLjYfjcPQ2z0GI9QsauAPd1XpMK2c8c3
nBT1vytnSueM0kVz1eVLSqkys5D9sO3H5Uc4zSh99JsOxh0O8lEjb07NwY5gqOtcOEgPy1CtUwZe
9KFI+sAj983zLobbH9QrREnUwuWBMfb7YGraBqXc5/JQbQsqbcW2kUIMaIvbo6yjzfeYNOE5Q21S
p3k1Y845P9bFSFQLnE44EhWKGOirZ9Kjgvs4dhIbYECvUnnqtBkA/l/RexY452meJkLNzRiEAwyi
3VwfBwVnrpo05aXaJm91dAI2A9B/KV5POEQStdWZOcMhpjLusXH1NcC7QcPI7Pv+dVwy2xzrhTEH
DDGAFSIv2tYrbollRFpP6q6AWpB0VDBPY8lCUZPeiwQ/AClJThdCgLIZyBQ3GQaSSTDXb9OT0dEb
LEMPmobESR3dHp2T6l2XEUcGmh3WjNrw3qbroVKP+RHabg8pe0nAZJD7Cj86pSHdiG6dSFRu6HeK
ry99HPAgcrwEnuRkfRY65jeSJVeNoiIwgwZOwccvrs7n/twgI1t83PDSRnntV0X3KQc8RnLAWVgE
d0hU8+8gb9KzYXGlMHG9OO598SUh2Ysis8WBUq1pNPGBEHxFN1XumqNmPPzUw0xN62gVsjcWAzPU
NuV00N9j0dgR81UhqWqntLZUWt0sq7BBlZj+GdBSLaoYqDKT7AoLXPzedMwgkBcpFzZSfpAtWD7n
sOgInHtzZudQBYAlLZTdCsb4gZ4SuSenH8HBcBfYvDlhDoj+NmpMVJYfGueVpBB79WpYRbPo/9ay
+FPVMnoaqm7M+en+Iv4WB4B49XgV65FTmCw1a0jR+eVEEv56D5Xv5Gs/LthmzCGWsCJhZZ/VKUtp
E0O4T0XFbst2AyGB/xFhPW5GO9XUqtT6T0cHVGZI8dp4KFFNskET2jZ3aa96KLSE7yCTfuaE8kdr
04fu7P26lrXoAZXNOHMs2niMUUIGl/OeoIgzroeC30fvvG8cQXwjTubO8uMCSfKm9HEeDaemTYLV
69yqsLxBHpMno3k5iV99jk0rCg9sqzyd31y/Otoyn86LEGoL15wIHt3xBj5XEaS1626+TA3zwsRy
d0KJJThWz6RtQWx2uZjQDoZn0AGRwEax/9BTf8X8eQwgd7NUynx2PzfqjAlPPLcWc9iEfvMs9AhA
z8MNLwFWTYad6P1PtXsvpjtoSdhKxItb17vpk97ZlqUPxL2TkiEKx1WBMa8d6+7e1ZLFDqkeuEw5
De7GcFrE6dUknnxo7iw9ApQDwawD5yTeMi+znj1R3np+ihwXUq7HEayBwCMAGJPZTXHPbGVCMB8T
AN5XoyuSlkSYkbLSHtrQfsgQ6CH4tnQF//ePqXSOJYheUwEpc2HfADCswJBd4xl9Cx/dpz//bzBY
A/9J+bwhxpaFXGxTJobA62jAI0sCcpa4aNR7izzYQ7eU2ITTcrDjtIXYQkWNkuaznm2tLbGaoMSt
D/gzzsCkv8VlhNH8HHsQhTjHh8m7goQD8FdGRUDLrb7HyyaRkgi+rTcdig3V8nqyWwIfUWZQxMYx
5I974Woj/H70OKjsq8kFMdxefJvTqawm8gFEo452+yejSPCbXxoknpNAb9L9Ikj38+/BDstjui/v
Me1S8kr/r7KfiIOsYI3ueORmhOBafdZSUqjSfY/vs2ytT+70+rQtS2WB6/r/kQejsAIsps3Q3grq
aSd64elega83n6UippnU2QCP2ikfKOlBhsAAjTPI0zT2V5RNhBQyX+YTM8c7WUOncM4MWFRUgTI3
EFv7KQQmZCnZNyj3+1mmRHpeEf6rV5YmImQoh4dnJT9ImgAcx/OCxEjZkP7PZh7u9j1jYNxQ8RmU
nZTtrgGQ4pCxwh3/d17cCGom1FWZ9gKc8G07XIHmwHJomKxHLeZ++dUfj7hk32m3aL3QTRqO4LO0
cDlTHC+SxSJza9EjXNppAhjgWPa9ala0K3UQJrIoT8QQOShDc08m2S0x95fy2PMPI/YUAWm0SmNw
P5f6kvm6cq7L4Bh4b3tqZMafa11MWyqhztZ9UybF2iUaevKpSCRvy1+dQWAsLZMa3ysFfqHc2dVF
A4SuCFmZau62hPpc6RTTAJn2XzyI0RnT+VKZrswqKCQW7jZcP/bte2zLnm0sKli80JY/hKL2+de+
2YENBaSJq0i57Aiu//0hy4NgT2JspBiag1FknMcvZfLN3CmA5jKuB82HFYeOYbWWjtDuYOwaMB0E
1Xur362vaVSZFHOKxB/IMgTHrRsmmUPsvDGxwgfjyJzHTKY6zI4KKUuBWJPL0j/suLCYIb+cX/dn
XaCPKK2286pnPehaH9Xn/7jEyZ9se0gdAGEI8qWerTI3lJJnTpnrAV5hTFbMZNXVtBpHiCPVXLmf
mbpIeqlpStRXhKEuBsEV8QeQerEcCj2f3iHCLA9XhEI+vSPAJfu/pLGK43X1dlitrXq7FxqNwxV9
5WpitBtR8PLiprbW5/U9+FK6vmaK56eJmFCs3xXFZyFildjPvzjhN5XDXRNkP3g0mNYLx29vDF3e
TV7oCd90UsCWRh43Gl+q5uIKlwMT7yj4jMcI3BW1DiQnf6hukZal15ji7KNVqE4sQ7RyjKoAdsro
nU2PgiuTidddWTBpW5hC3mQ49Uk/KA+o0uNNgQ1ridkQVmQPFhmcSlbchBPf5o+nYv+ku4YrQLIz
EoeqDJnCmgEkW89p2WifXsi0zkxQ3OfyAhovZs087WlesUTHfEWGVqKA4Y4bsPPY/U2yB0P6OVoQ
D3Em7Pa/SAl3CKiLv/79yj9iZWV4lTVra1dRWahcbl5GlmqCfCc+/NFjgUgp6m8JmhYIY0ayV3tu
Q7O6WN/nlOKSNMJZQl8kvAa+hON2Gsykg833CFaqQl17hBiHBheNWQ8sxlxTGAD8ybut0lV1MAEN
pri0IlVTxozhDxtSx5y3iW+pFGof0+9RziKBEF16hxZ+/vgZAdUsriBSR8khm+Tgv7Q/F9UFd1h2
eqT29jbFZa5zdgyYZU+U7z4st1hQFMc+Ntcpc0fArM7GvHXUzY8jfMLIZUViHfH4j8YL/nOyFdKl
4KHasRTgzSh9rCLZstiZign3MdqjqR9ivdAY/Wp5JgYNSfuEcSQ3iKR9IvRGhd+gwTFNrgLAUFEa
O/ZnTrXseO64e5EaGjOK3xq0Jpcqm481w0fmlW2U/OHOOVDO5D+uvvv5/zWX15pTMs2Vi/WqEqMW
zYdEFvkf3MH1XB++/9HtZxttLDT40BUWkrvNDDYE83cu8qcAfxTtLmD9UAKEl9OteBoEIjgQUDmZ
E4wDa+1HG2TEODeAGMCn4ZrJRXapUhqrZhsSAi3snVDSMQxSn1pai2C2C1/ctKiE/bFeuDdqUS0b
KQ7TcMO4s3C3tuOd7KFaeNjJ55aM+ciQUrxBw2RrO9i1I4of+RqThG98rt+u/V7oGp6FB5TnoavJ
oxWYYxW5i4amQAUfJyL6PTBqDwToxP5stcc3xlDfijpPGUUVzS5v/2Lw/FmpMDakJdheViL/VWQv
f9HtKUyrgFGzEr+LFsN4huca5OZjwfYy40RSQ/VxjzClQ4yjnGCTproc77tPBpjDXqs8laFtRAkh
Yv4l7ResrYXlGQ+j5bTe6F45lwLVkt9BdGvhGhEAxeOmAtlMHyFPLYzt6v5nMJ3gdlYkkWMdM4Eh
6rrFh+WFqv7hxaNESYWW9AUH6bIK1s4Z7NdEf8LcW9w/dTqtbiNtxu+O2EQIlgPl0Htj64kBBNX+
S71QF5A2gQsgE1j8LxBTIzaypxCLO+RKXMCM7+Lpeh6wPGaG9/lILxwCOLRNvgWWZRZV3it2Kl7l
SP/asC1Oig1VF38QPVHANYJDk2EhrYZXUDtxSpC6F0IA1mvKKtoPjMVrm8DXVPNrSXg6ljifYWho
tu9lGyOzKYWBTYbigoirNo7bZeOtw17tQoeKCDH7HSRWdd6uTpAOIPsu8l+5ewdKJwcObM8y5xk/
DThLFREKDz2E1jAwcI4o9DULEQW44QPx9tqNv1APDyIjpSHFHyy+IFTeXZkwKCaZHiTixhhL/0rH
rKlq4L80jJWalHzs+QOrUTBA1SzkRzT4YclQrUGkoqLrWxUTNG8x9DEiS7gOO3ub2ho0plbqVwRi
41br2qzNiOagC2+vhP7+a5OZ+Cojrb5LwRtvFfxMI14dau42b2dKXfP/QyQQkb+ZyBrZ1JMZDhrE
E8vmJzRKMDHPrzA5H4fgEzAgEFU96HMhE85sTh8eAoQQs+vcNjUgalKKl8i+DU43EbTdzWiNCIH+
0Mg3JUBQO98c7ZfGW9gp01wVF3IpCnaUAZZDiGookbZfbJrwX60OY/4KutvXzXGj5SP4OTfHyFjg
YgsDCTGOEGw587McUELQPasfHU0YrM171IuAWhKOzX+MZFJD/qqvh/9HAypaD9ZLQJPgHpQTEGG+
gZtSjtY+fzGwYP5AW88CuDlUoMt0DQSuFxA4fzZVAde2ifm8Rn9ni794lHbOQrvuVdmK9ShGAs+Y
VdgyJTyXsSFgZ6vddiPOpm0nkkXnGEaKCiB755K4zsDKfoGbqgeBjaTzgo3MhN5ZsxqELyfCe/z+
BG7KVNYltQboqZaksaNyQewmrYbB6HiEiMPKcR7oX7ZprFTWEqFU2CqwWL5ysM4/yHtEty701pc2
xtGi55PS39XXdsZ7IGAbk5LQxZKmYHnmutJ+KIc55pwMm/T1jlXxscBTMezsru46Qx83JPQ1AELD
urwoiuBBZoJMEga1CTy76B9CxYgqd6StMpmf7g1RywVKUumY6R537PYnwGOBoqo3Alp/o8C+VljR
/nZclDngq/eTc4fa6Wqqv8jZB5cNZZ1Y1NlX9VlOTTTdKo7zDOwQ7Beutm69P2O6ae8soSL9jqDW
Nd8kIlNlq8u1enhV9nytXCQ6CbWaqf/zun9FJUafidMuzpZqjQfSCNwDIhqm3W3wcvZR4QPbMyzm
q648+CFUJC5YJnqeqt5VgJUVimOztQFJjLTYqp62Yr8+JjSe3sWQd1Tjl7IIshcSejqwbRLL3Q8s
hZEik8ep79GRR+UP1V/eoyMbIyYxgEo9QjtXg5sG47dhmk/Myxzr0zarqnCYw9fyG/uhCk+C/T6x
BW5XkmuzorMOAsRK1dOyFBHW3cXSQN+/uIwlgYtZsHTbM0n3d0/BSgOKyk0z+8CuErj2uGNGe7lE
9+EzAl0vQwHCxYVSAkBuMxBtPzgPZDFrXBvJjODFobhlwWt76ros7Dzxr5UTMnXDDsnKQG7ErNfF
yrorhKQm+LqfsrZZke8MgkFGNrXms/VFKlY60Bfh8AHwZz1riyrr8L8smTDRz3BbjgJHQQO2YxWY
QOUQQPlzin2lOWLIEHmWmSdThMK69b3xZJNH9Mayw7jRaUvVf1Wi8zmc0jCesJM0Z1WmAq1x0mKe
YiBLKuOUe3RouRvFz2o4U6ggFrlyZ8BmozVemVq+50BqGs8UdUOtQoSi+q4+QO6e4x6tAuSngk3t
VFMnm0wN71Uzs4m7dIEnlC6ZMUTTmBN/1Fbxn6Snc0O5dvmDLqRqKXvyw3YzgBfqXzyN2Usvu191
k2s7dDpNFROHwPgI7VxjzQSBPBSZ+SMRzJBqry0uOB8aFjZpk87vi9B7mfxSB86cPeRlktVmen0V
nSEzN+RjPxWKEC/Y6d/Ic1tRokV1mWFXQvNcR5OgmgZc8+ccjzqcHjG5DJC/AjW/llTiXw//UNr4
fYAbl+A0hKU5ldIuPDeLmzbvEMjtvXvSDsYNErJ1EfJgnkQJKUSGm3sCstqfJgz07QcP2jgF/KeX
FslIQzQ1vZgRJty0I0ZudMDlCP2cUX4w8rXbQMFNZDmxcslgC7OsImLU7KcGYVPXycIqvpIQ+Kuj
y7GLKGYyvTPMApx8KzHh7HtNCJAgWCD840CT7HpCnuLwqmRKTOaRx0q/ky40s+sZId4Q2SbGG0Y8
H5aU+g2bWPRGx3ylcCyMYtYMgVKhNlgdV+wqBaAx/d8U1emVSjA7m2tjIMcq8r8/4xXOEtLhu9Qy
11c95dDR7XGCSMNCZWPhGIHV3kmCZk+Sc2FBMKwayZgqjD69/KN/+AEBd19oaHIidt2hK1EBNAIm
6wuDTeQIp/V2CYzw1a19vQZkxIIMl2hbE3nONeT9T4hzVBWtjYp4p4FnmG/zmUKo4i3S4dQzTIi2
I2WX+iFMCxOKvfDpWfljZVE+8olyPzMxRBSMVJTlIbQt05GKDWM4tUHguO8kSZIyzRg2BXmzNFkD
nlb31WtDr1CD63Wj5luVNggSjYSulUrm0FTe/zZtwUMxvmPl1JSRZRTyLoxjeiapT4sifc0P6JiL
VHX7tH6fpNkLixC1spvTIKl+m/rU/MENFmhYc9wu5LgIsXRhx43M8DnEEZg9iUlSbVBogMbiHb/9
4U1Ct01pAlk6kiOgyjR/e8NzJXPpFZSNWeq+EXzsDB2FrVoQaR/M9LrUPggiIFpMZjtn++KXaCsD
GGTjxzJQ7qVP1dmEnCztw2yM1N2teWqs+k47MRn53LIkJrNJ+aSBCS08sVwDtVsc7NwP18y1rH+D
kF7IFIQ1obE5ud+BDxFRUcWPuMan5LEvhdf91V3iRKfOR17niAG1r2LgT6FkRplujH7qQmmA0rJD
LaaTa89+NxqCI4hf8T2yFPq52onADXvTQ1vAg/crggTnBqA2VH8Jwp5+REcPmqkWJ967hhfg0Y+M
ccZaEBj8H8Cnsx3wPic8LZEStMK3Q0nqr/7HHTmUkaa9fhvFqfNIY/eNzW82Gy3LRz2ipDcf8166
THTsu0zNEyTt8fDvsGdfhULUSTn5w0jlIWk4K5JYWzNyeW3N1z0+NpCW9sn4ABTHesln0nD06NEm
ZBj1BowkyOcpe3PGq3rRshYiIPKfIY8wAQDHeegRjxPHSenofKAXu96nnUYhsIE+VmLeR/WHGKXV
jEQRqESknd5tOfVKzFXvvGRUWtrNztVxZFg2IFpo5Z17kNUYRo1CNZqKQu1p8afoFYrbh9hsLDEf
zRtoCvt+dEw0rnQ/5IGqoPCd7q/rf1ytnNvKhm/V66hp87759UlS2dk9qxgI9pFixHOaZyW9GS+m
4LHG9YyhSQ+unNFDBGNfPq3jpMn7l3alUrPUhGxwXEcICl/BAKTdruAg830sWMLtbrbC9NiSz637
Pah99ae9RCMXrObqQPEJCuOhPv132GuEEzJ0gs9mtT2gfuaSbeVNHLhcGUpoBcRikrxCIWK5SQa0
GboULQtIS99gMG0KXUbQfMldTiQAoBYThvC2t7jS5g3et56vvJcqQCRyv3jb2azYR1OFb8CdUQfc
H+O7RMvGy5aM7mnEkvotwjHehyraYZO0PlzaVcLVAdeRgIeED4dZJnuqUax5YZwlAtHW2DMUmDHx
BH6zPE2lmFxVHLJ6fHqsIuYVz0eW6Yo3Qcl8LTy7e0ckniNNebrz9Rvlr6D802XmMsGciOThdhF+
EHKcLG4KxbSxwvqiIKbjoqfOuRHfR5ViA4T9zEPs3wuRzY0smBKDK7Iy/QBkOM/UQHQaG6S9IAVB
SLS8giEHnmzhGWljPafsx09UBVjBdgclaN2QIfc0BbUf1iRhPJADSBBVU0gS8oCHqaJE5yIGdA1G
yaNE1pkFBEZvRwMY4xFsGa7U1LloZAXpD8M8onUhE3y8Bm4Zu80d/JudUlsrR7uYuETtMP0TLB5g
qYm/QC/phZjLZbHbcNtXJi13or2nPHOSCEfofAJhkTf0PLmJz1IMv3Mtz23mn/JlDILOKfqQAW0p
+BfUmLvGUSGvj3R5xCL6sciR4Xx+qDaDTM2r0K1Wl/XrrOFHIt0e6kQWtzHrT0nOj+HNumSRxxc8
qGOJFz/F/47GYIKVGrI5BfdAj+Zalc00mMpWOmJv1Nf78B1Or5IZj/ZMYmPxiJ/0pKhwbmnYfUEQ
W+mf1BUk7ENxl84ongrbAhwEvatCPucSrZysGKLqumWtZs5J3o1Gp5eFx/vGyEphUtx17WZbwu3i
zo6KtdAcHsgepV+WMf5zbjC2gU+09TPa9Rx5wgjBw3fuquD8HLso/+u/pE4rWGcnmGyjhk4b5o10
ZMZ2P0oP7f/kf0WqPieX4Y1d0yeeqURByVYtRHuO61LoB9Ev7e4F0a0X5/RKH060zX1ge15PnjaC
qk/FP4Hc/9hr72yB2fpBEaGdLvCBVwkCWbSYsq6xxLhey+iymyE2+xA/XQIC0oRrGWx7o6wRHaLr
pcE44GWDoxoOUqc3+89AZoSUGvlINyQdYFemkUEICs86p3gFu0HUP2X8mK824Ihv9ckxqb58u548
MaNjhy0BJy6QkB2fzcieqeIY6UC269gACIrp+8pZEEo7ygH7X9/lpo30Ujvs9DE9q0UJpvkCX6pt
TuxMkCkv5ihR3542SPjn54Kldbew9N3SYAwEsIMvXIuLHT0DQ4rJXlZZZO56uPpAhZy8NOlTq/eX
9W59CI0YXCW5ta84vdgBZmkgzimTb/FTpksv/Ro/Ee0CpJMVy1AWN8jdrrlDNCZ3QFSI9IHDZ6vC
/FEPywd7mACPBg2B+0hvwOTN2kcwTDqhkETfc1pL9RDdrhWZ0zw4wL48buIPeLj+2kas8duCQqi1
cwJPrqh9UsOmM9l+EQRdKkQrXZj50dI1ZGoj5vOxWICwJS0oeSUFpi1wxSZkXX5vs3YBwTrp8TTR
TtqBrjwniK3D/mV22Pvncg5RhFJ+ICGEPs1eHDdawTSfOJp+ORSuSeWZI2gOWKL+qLCKsyG6wFhV
KmcXG8a82szRgNYJ9hqj4N+MZt7/KAwOIjnQFAkR38L558U3K4Q6A5syyIk6xUUmeqQL8w/pNUsj
8kTh1NvTE12wCVUNjPG/4OGIPe9KBlLO3kcdNvYCevNhh3pvfpi1dtlDkhEtoc9mvWVAlxNrwZbP
9LHyw336BziOoeC7iJv/fJTt0gULmR7CXYdgZQ7IfrdOR5p0abkLRHEiXqNydkezecyJuVE7OdiS
X+yyw7koMybELZX+UrNr9bJKvv0fWTBOmWXLj7wC3RP46uLmY1f7PNNRsa9+xJySzW4jPeJxZpAW
cFPCDivCE0TOoRMV2v9eljo+zuyQfIxNEsFgqGW7QEiUJDGrgG3POzhO5ciyLxz+q+x4m+rwmMau
zGXOoyddlrYvOGuOz+Fg1YJAwwQTUp1yIcYC2PbyADusv5PZDvbEnYWYk+lZ7Q79Jm8VKl2HwubX
8zFvLeIUjvlzH+8pOCvBS5ZFLP7biAFqhXIy1W9IMIEu9jS4B556dxTFVfJf7hHiEB8EII7qIMaJ
V0FaG8qI3HajewjKE4kGHiPjKbkHdUAT07peYaX+VZrPze2ByqJ5/5eiLC4f+R/n4yF0DOu5/7H4
lLe7CenJe/2HOnR8C5O4HYvSw/LbUcWykKzUwOjvXaLCtliAUYkMbsA2CAqCmXI0FggfU+o2wGfF
nsZBIaJRtk8L4j1Wv9pa85ZpIT5G4Ap9a1xzD70GqsaybEhICRXLmLY2lVdNXG1iI7DW0Vg6gk0m
7KOmX37XR5Qd7UKC8UbbIn9UO9tnBTCeYZWvjqVI3Q9oHaO0kiy7xnlXkmP0HiJNIBYw1pFITmh0
JR1a+pFJNVsq2ja/BLB3VnRJtBRhRkZDZMuM4aXM5Jw2DXeEHg24fk4yDlJh/Tx3ubbuShDixmSy
D/1oahBpXSGXWmbB8TeuehqqSxGJuZvkgBCOU67nQusVV4DFTvhp3u0HS+Zwvvd3WxXQ6TIqigN3
ereBcNEaZE/yzg0qknXkyeCIv2uPDmfTsS3ziWkixYd5CMm5TU+pRUQNVGPf6ATOTrmPDNaUnTPU
9+I43l45Z8+s7Pwt4UcQ+E/75zCqdQOaCHGmEz8Tq3TNGEEAvSdbLuoUbuRyAj0orS3HKuHsWdRL
1x0Qovpq7v/wP6lFE3SvvSaiZN6U/SDh1dwTrsU40yFKIP0a45ywWxY1K8Rlu3pcQN/CuDL4cjyT
sX5qbQPisQCjZydCipCi8ihTQCoX2jqtz9bRIJIorazTorFw8/5cU3rjAxDMDgxXV7bU3Hq8ltEJ
oIfr4QiFFyYspUDqN2ya9O4zr2eQVZuX2EIgnF2ZG5tcP7H0wTu5fB3n5oYycEtCDVPSLfOkeOnq
Pfmn0DfGfO6YOGLfxohSuChDqveYoIt7wP6HBjnB5LsCbtTCNJc6V+SmzdvOiRcXoZKV0Z4Q4pN0
Dm1kHdsay5oNx9U/oUDW7ykFmuJOscpQGjo1ZfbZEe/CdBvJyvYemPvwzhBecwjJuu5iRIEwGPVN
0CB8EAR7Gz6TnGjin9JGa71OO190NNWwKceKqZLnePnv6/5/7xSSJ45hICdzZGB3z+BbJUlGuwmw
aRbpWbqCBklhkKCQmS0pEx28r55jgtQEIr724yJ/j0u5QcX74+OPH6Ebc7pfhMJg4TWXJM9mJWnQ
poQ2CuxozHEA3VoPDMqSqY7CZJHOtLXj+qVMI9pnRFQ+TsJZHs7nZtcXem8CRZcyptlFZL8MizY8
lXXCqhhqPVu+LNZf8BvZ5MiBhIk8/ZEYN3fiJ0dX+wwM0q/stCPJwjgovUU8dzrPcDoiK9JSpTG3
9AVPMSPfrIdppquBbOxnZitBJelygaLyRuRr2iEajTecQO4B3i/T8bmGK7z5ZMuA9hLKcZClPGtO
Z5SMV5eSDVrqnMDE2NjNLhXKjPLKNga/EZTtIbmLJoPjSD4gftgYngxNAJxkgHxdabG3aRj29nYF
i0dTKFPwOevtZODXIKsVONrApBxRMCcf1GHcbC6CCLxnKaG2wIbixUPwQ4haqOHrTPpF5BxV5XMz
zh8kEt+PkqfMxB9Y78qtzi7z9+PFJR/hxz6bbu5EgfMUX6FGMWlIESIppEDnEGEMMvrFJwGSmuyA
JnpVYmMkfNhOMIv/68s2wtsl9NwiOXLC/t2LCY2svVyYrSKqR/8/CV27UzxSuV1dgZR7b2DsX9aB
EVmC8Dw46xhHKTq7Nz79XfgTzPS16KzOd2hxg4yiVXDdA0uWuyEBsLweMhaDDYheqIi81RypZbPR
UiRCEussLVbuaRPhnvwwyrymwe2eJ8039IGWt2/LvRzcU2v+OKTdrPrFNqjAt0VXn04JMpTN2Sz7
LgxhPNvCdT8ZnXKRexamkZh0QDmFV9m0Hc6ckJCTfB7CRZrCuFs8VGtGESX2amkTxiTu2H3HXv0G
aSd7UoNcXdzW6c+hQiVohP94t1xhP9YMg6FEYxqH7OyxGjBdZVcRcA/8P/uODE5lXpQwDSqFfybK
gFL5Nxd7aRM48hJHRJTKZuVLdlrq/orsqJxwyz3CMySraw3hhojCJ3V05xQMsA9D4qeFeDU4X1OU
aN/w5oJ4vIhblqUB0ak8blKg71NDzc4GVyH/EoewBjCmeaQoSUB/67yBcXWZ9pSfbSplVEHMTBjD
qFxOJndjTFkCF21RH+kwTBS/qTK08pl+owbd7LQ8/h1Nzpe7rdA9S15AUK/0fXPJe7qo/T6xvw51
gQ8zzh0aC43w+HMHEPbj7LDGDhn9Sn/YrBFz0ljbQje6f+zoZRTRJ1Z0eMO5SeW1pnAxH0UaOyq3
F1MfsO4L3VPBTJdvMFbDto3CmZvbOpAzD8RRx8NFhp8GONrxOrbFM6Nb5tdCSRDxLuuzXNDCkWRz
/bmQiXjTaYVUrQ2YVWEE0AazZuCqeTCYbbMm3TuqegseMHnNLyAob7KL20NXy7G9It+vXngk0v/5
VtoJjIwe/lDAFXs4KmBIrxbGHK5xuNslSzWd7eCgvVpeFhLwFewwbXqmL05soPVLcKtBW3OwZOWD
uK04GkjTsbGF6wdGh3e0Yp7P+8OqExbVl+LZS6fPl8Sb5ucxf7aBD5tFkXTeRrRzAx/7t4I7tJxj
pxoFvXkUDvO2jF0DYog4tONFZC4fATzZFeWDRkjFHwsDiTImL5PhJ7To6VWZ14wlX7L7g5l5WAvU
zEUaitCcCmK3cZ+/QENuwQqD4KXKBF2Kib/zV7ZD0lNTHFOGFT3CvNc2wjv5GOFrOeMkXUE+FtnF
25qeB/kZ9IVZxFb2glVmNeVYua6BurDNeISa0+9OogY+ZC7IuMcfVdu1KBv6GE7xqZsW/5ReB3Vi
hW8dYyQE5RnwQCtxsQ9dDWFqTdDq6oT0dQOq5MmHOCgXc6jzA0c/7cNgA0WrZXrd/IEXdN6KZrh4
vpSWE2+Z+tbg+o0xAlvzoGQVVJvArndrBU7Lg096Zbqrj+zqdeUx99CRKTiy8eoktZ2MS4LTupFx
axmc869Q+zJR0L7yxu3ggkEr/Fx4c21Rv7QkawY1FM/vddCqb81LGkf5NWVvJxScuUBNYy59lbdQ
tNvznoK7NPqV1Pmb5CmLinRhANmr6MGC1JH5bgnfjIKwqkY27BgQ1RZU/LqUw3Dpqy9ioIgu+ASK
bAZ0fmUaFhFso9PrBsMwslKFu7vGJpShoHZQb77TyLaU77YlbhDYQpe3FQzESYvUq+o0zJatZpbR
88D3n0gX+t83j1gWmmjdsHT456fu8KcbS0sVkovcXp0OchfZqmqHj/PlRuo3XiNBvjcEW7aH/aaw
/furkffycVmtRySKoQbiJKAxwqNG2ijAVu/UuNY4j9dG18ewvEWsbqGyvFOm4RXeama7PCIHQalu
SWkhieSG2AuXx+i5a4QCst/DIwhXOg/mTGZawze6k3rqTmpYQOtR6oZuoZdhI8IPm6HMY5Z1LEt0
QJQ/15FdpjfG10wSny7vEMjchzz1IxxaB5LzyhueO2+N3ma4sJQpHL+MITO3VSRs+Y39x9u3tab/
Z8zWpeN3bFmFrCFcsuqSZ52y+Vh59a733tMr9HSWzi7Br3jd3Fwz2VzNk60sc4Dk3TOg3uRZr1fw
vvlHg2h4bGBpUavVulexVlMhXEbSdPsUZ6B5aQgRSooDj4zqFnErDwzT3dF5/7rzpRYIDEXmiosy
I/huHzGdmqMZTUo6eNwm7bFwbqROI6ELYjLcG/i0r4j71eOvGL93OW/+9f9IQCpxhx+OULhV9O4R
ZSY7TE3Z2xw8LZ9QHhzfWck7RyzI0xcMoHQqnlGYG6AhTrj7uzgeVLM/39v9YscjjSDZMWEHeIUm
hkWpR27kP7Kz1TKRbnrmH8cNK+ghGqEs5+WQMJo+1KvjnzYCr2AlOnmMM2+SDhIM8Mzyzq5W1ota
2nxXgiN1x6BeG8OZW1bb4UH4NgfmsowfcmPoC+z2JUwIXiHChkOPpE1UekD+j2I/zeF20zhJDiGc
13pWr3jaRZ2atTelhQmka4CiIakYBxrL8PrO1AGVEKVdZfpdDjg4hrsI/pHsZh9VV46Jwp4yQnUj
cImwYyXDiY9l5VDfoXvDPz5EFPE5A+y+qck6Vv+/nB99sQux8+wuyVnebxJWGl69obR+8fQcgbdM
m5LhgDd0HBDGX/kkghWEdLSgc4rXHNfrWPmrao+xHvjAjCNrmhLXjO7ZvLIujghq+lpEI8Ft25cM
HH8XZ3jK+41avJNJ0kssPdCxkXGEDDuRk/Yi/S/W3q39F8UtrIqayqXYpew35qr2A1f0tdxjRctp
54dSpRamkNqixXE3kk8g+xonZ4vNBKNMqG9/eJVYmDfQBV+lPRPP8wHbszWUPK42EAdRjg6X8j41
Jnc96TSfMBO/GxaVEMRQeh11HUow76AKsWrsC+opGwmQeFZ4PNZJqCKMWrxP6W81iWD1lG1KkJ9f
N2YeZgJdTlG4epH1tQ/LbXt2DQOs0pQ66UIB4d+v/9YoAaZDI7JSnR759uvVFz+85w9c26kdiAjn
/ewsxsMdGFn/lGeHbOZzSjnhDACcnNwpIEb1+fONPI6MLDJ7jOYdSb1CGeAze14mus/Ls65WfU+2
N8Its6Xg5Of+PuQj/ljKx+ttuw3bCxdZCXGM0DpYd2TALZRCgK/sklRYZDLX8t3Pk9lQN9YKd482
l2aS1jHa0QTYsjIG0s4Jbpvz87s4Nh+WJ/F32LNzlRSqq0BNk9rWdZCO9+/XVbM7ZFaIM/ox3q+S
M5/WHfuOPMzjSDEBWO2F1YvqqRjv0rZT0PrVoxmnMIYiiFHa8JpYb/MaHxQDRB5Lb2FluPKOdoe1
2UiOzFR12DGa/oSnmnhpv1B35ExGFFpGS0cYMYunUwU/rtoikp8Wu3zAHF4fu9wW6MxTTxVbl3Ol
fYlU0vnds5IrE8lnYesm9+x4D8ADUNQV825xt6Y+g5cbHXreci3Yv7c7bKcL3nYV54SNrqlIVX/g
4BE71ithJFhWB9wRIYEadufZvefBKNdoyuPh35QcsbeXX+T+Gxpb2p2Nf2aik2cnT4AEqeo/ihXv
ez7/R4k5ENVzxg8uggc1+dAfcitUN5/NbZAanXT1glgn1mM5gRy9mkcY7mJ1YqYSrQuZRo/deA1b
R37R6sXTu9lfuw1e227Bn6sb8f13Nt3+M2fB0uCuc8oA6MDZuVuyL2QvzSxvvV6/MDoVGcUNOKhN
foQ9kz6gQ4wF1LGLn+fJt5Xxee2gglh94eJKcOsK37bOfhy3hArqMSPzP5QV3LAR6E8rYozRuhxv
Oxt8Th+BvQK1RKq+O8keCkfrdCUqgFAmnfvbs8tBfWm3qN6tGlfX6qGA2jjpdWIKnnFifqGGFyn4
ASEyAk3++NuxADhECf/rAc3lGtqQLXYUPKec/EHyrK1F56OBrVoGzdxORmagV9dsDqSkrxYWQp0j
MyOZ81j8aj+iuU7dBtKjZ2u62fQnSxAedjJh5poCe1lCELfna+Y43kc00AEKw9L5x9iZkHWTebC8
6OaNzlPwVZXFHl2c/hPmRHZ/qv2CnP+xLs4FoqNE+oBbkcgXtY+efnlw/uGrC+gfwUp5jLQjZx6d
/MHDS4YdkWF0cXSt/2n0yrACvYDR6ykLbDwYRfpDkdF/Jj9NmEUI8BdCJeQIp692f1Vl82UTtSyE
pGtgW+WAJImdPoNCWhIjM9tCXyyQqnQpNRW3Ko/4U5tO6+63NEr9phF8IYtMkkXKeh3KWOj7iZg6
3wxjELO0ASW1slLGakzRvxQQY9zVm6DARwlnFN2fVBGbcO78xbccmnljq1IF0S8yHPeSQDwdX6U4
7Nk5gGaVBoKUboez9nDxMvFRkEJ5+j0R8kh7vnTmSwh0LyWbGwbG2qX/Web0OUGO6Bt30oT/JpUM
iKKdA+R7jq3F6HceScehRkuLNY02Q8g35FLwPEb3c7lEuzTm5DNs/asjjNOWoo8Er+2/8JnzlS9z
weBIzIDHlSbYNqJ/EHzwvcSUZeChDzLU6pqJGxMP2u0Fyyv4u43+qNR8CE+B5HOqKsH44N4fjpLU
mVhD5nlUFC7EHG4SSCaz+mepkYNdPPs4R0nqVzTgeO6ePxcn6UyKG9yztW7XeCr0C8sator+M2Xi
jEnP0D+MDO4Sf/XVUVYsSpsFV2i08vwbvYhFGq9afEZDrbi4W4nKcKIgmZ0MH4cm4eDM7tCGI14y
9wlAMOZk0enmprYgjYSHT9JnwXbLQ+oYWcBuurwwQQtz1gqFYUhXVKidfjZQ8HnZUiTqJKQ2wwaV
iB67fOzdDjM5V+hPvQJkuX/VrN5zYBRUIpGm6ScDyZsnom0UOBpPTWo6FM3oT1Foyqu8Fzwm91vN
40l5J8e64qd5pj5q4x+zB63mrSHD87cTo+pcvg0rPjG9x0EKZUGZovaYUGeUg7ZAqUutNvfkso3/
RjoB5CuttSCIpp1lVpGU5X5r4XySPEEo3n1uXqm3pNT5w5SWC+ujOgU2kEajFHo6HpUCf93Q9xFg
BOBD4fId/Q6sa7Efg1IJ776oCTrgV98zZUkKvzZpzHjpcpq9b5vpUH5kDXU2erVb+jGlhOXcLmsA
LiLDdNEtt2beEHzmL3oqxgoBJq4iBHa5Q+THg8nBKMIuISjX2Z/wSQchzdn5kdghdtxuNhukPvcK
IHeUSipuPwlDbtCgu+mZ9O87YZ+xe2dCaGtmVlOZcDIeWJaOMAe3b0itT6+kLTfxw8KbSBRImyaP
NuzauqQyAZ5pqVCmfrEp9L85RTmwO/Xbp7SjjpuEnCQV7fLqDvlXubGSSmTWAkmBPFAbWe81LhZm
1LZbUAdOV51CVIum6gaTi747b1WhwHSgmsqGJBm5HhTKP8ic7j7MFYWs2oMh/zl1JM0oyjM7fIho
sQtuUbqnVtlt5yPRf6SkfG3rptFt9v15X21wMVk+lwK4s5LsBZiAawnV/1G80jgKjg/T4shu3R1e
LETR4Vhh7y/7AaH8qAkey4HbyV+n9bw57zeAMl60s4jQ5V5dHCPAn/qTgqjVMtVig3ErNXB98MK9
73Fm33xUkTzIIy3rvGbEG1jt/CN36qfRBtvqN1dRhjI3YGXH1fb+kQ25ORZY5Lzp/UgYmlbAt5SF
3/P2IY6nnuqXvr2g8rJjAebHxSwwMSTEDAhlh29xVf+YUYWQpbWCcm1Fvg8vT1Y0j4/IW03X9iIC
Eks0dzcrRoQaHGK995MCbSBDcHkNQvZym0V7k4wGOMmmP6ozipOc8uowFfn9DH7yh5pneA1u6kD/
PWQp29Jb6RangDmQ7dl4SH63mrm/kycwF4ytzFXUDKO4HIRqstQVgdxIOn2qfEltW+pO9MeXhy/4
Rsau6Vi52FsAelAGJcEBL6W7QIo+14SuidGE9D3i3yV2Bm+Fyq16tf6rbrdE/y0g9QEjSZqTtCPf
NjCwG39qSdlK9PzKB5p1s82dOZUT5/dg8ngCS98OcRnxUgyR192EnPeRXRII3HLV84WkzK864CEO
WsdkaNNkI2s4nmoSSihfwQWunjL1QiA/xHVdXXlEJX+qdigRpQT/Bqf5sh5KXlw5b3suFhV8HkE1
jRrqg9322wvfF6tkdmL6c5DP3G4jmAzxDeJm4gVFMcST4xNm7eE6Od7Itzj/BP/fHjnmSduLIsEU
2bQiJv0Y9X16jWfcLHqWGnCG8PwukGdoQrtNHFODXNAXszfH6zYz9vuja+4LvDv85s2+rqSsjTia
XpzA97pR9s21qNqJYGjlnlc4P3vp7WXcLx7FsiZb5+bEZ6owVhgbO0P9VTJwgWvEzl1rum22hMYY
HI0YDiic3oBrIsJUruLk2KGf7T/siGkoVfEgUKEQ3SC5KeM/fzU5mYOUCVsVw1wBA/qZ8Hs9hJjo
kPQWLrYilTHs/g2VZX59Vc+w/gJ56FoRjBd9GhLJO6y3tUbRJGzssooyPdHXJXUv40mWmAH7SdQ9
d71K3Mmfp4uxES70BHTVu3xAA0LmbCm3t3pAq2Iw/qnGaOCR8Q5X98ku8meh93RN1c8jSZI2pHcP
+0oB1Bzxjxj5p7zFy4ibCfadSKo5Xz4mlfcp0MSc/l9fDlUB1F/nyhRRrq3pcecz5UTMLAJoY4vY
DcAOOcH+4ssEkxNjzGXzFWmqfcMmKJYQXtsuVK1NMZ5DzUuDGyNHbBnU04DxkWywrirTO4oLYeFY
O9Q8xT5YkCM/B1ho5KL/wkcyBG6jZpHDTNsgt3W0QXuie2PSDkBwL1zxmvw+h+FUFWBQ/2O7KYPh
PXf2z2UeL9VCEHvPsU18gR679GIloXvZcrXLDP4qtxTT5YuCU4itiK4joXFK48BfRAvMudVpX7qG
bbxefR1hbJIcG1NvI/9/PGX5E5GDTb9FQdGV6O6Sjjilu+JHJqvWIIXG7d5fVUicdUNUB0wPLj50
yw8/r+3TGPpMQ9jDgr3R7tdOTVan5/3vMsAZsv2d4IryDaO7+HRt8KK9e7aLJcoIHFSOMwHbd45a
W12QJ8hsEtoQdlnfv4oyLkQOfaZ7B0isfOnl/GduS6IrEIyHpOnSDaqXefn7jvRqpiS3lUJI+eVW
9wBMpNpkuSDV4IM2FpkqW31wArejEGiKAHCW7/Njz5nQHNX5TQkwkiN505pK42JoBNWNDiVg+L/5
bd3MY7SLh2iybC1lzvcoapasLOO8HQsUXdytwOw3WLEskz/9xJwAb6n2EzcV6NN9ZYtY2byrEdD7
cjmpEvNxOzaYFSAmfcuIgD/NE6KP2YhElxvx8zvkMSzZy+hqc8lYpRalxcyD3X+86z1E41DhVa88
XXChPyTgyyut+/R0QJid7VXtDB7U/Nv2veeZMqPAJBCEC7WOcz+K4h5PmofVdff2JxSKXVp729ZE
80HVg2g69zuwtM/ZusRwuWyDPYVndkbTiKy1owib1jLTjQVhVVdXzMSDrUICdwGju/4Vu6bHRDGz
wrlU7tlOepngO8ISPypM4NqbwXpBqrqAm9ZweyZ7KwWbQZyOUXbnEsADiMMdLZw2nxBmFr0wqw8D
FinZt+/vA4UUn0Dg4MgN0JA/DYlWGCkonWRAYGrs/+HFfmAJ8UA4fiEEFj+/wEfzakeOUeL0lTwz
bl0XqHaJo9OOS6F6YaZ3/kBqtiDfr7gzakgNCt3/zM1ZLjCSDx5HPZhZpkIKx0kQ5L5kI9+4gsfm
Hh8q6MgQ/Udt7MDL+mD5AePlXMtpv3Zc9D+dNKhqI8yEk8NJMbzqQ6Z44EDDYYx/HbfgAfuI5484
FtrpcO6e+Y/85sJ6up0U5Bzte9RPrcfwJde4eSsfZEbLiZBCoNXmVRd6vQ5oVzlqWpgu5p+zttge
0JDe1hqZ7cTeNqyY1w5oWh89kwiqAEaGcvm86Aw05t1DI0ezQeQ4rc9W+RhIUtZ2ZH4PQgWpfVJv
wwIKCdacoDhOSJACsOKgaiWvlkz9nNHloItwgVJIaEXwMJgsuKqccKq6puvWRpwLte7Yw1I+iw/V
hSlQV4aiZswYhpbOxNIK5YqyJKaxFnjufsxPqC248QC+i1kFG+rp/3VeHYs16qTTmWZ5kzgB7NM8
cgSYuKHz+DB0jgEaahHaxBh5cRUWFF6fBVYYUST8wxy1dI27IxzACczVNloQPwhVzxtN9cF8Ofcd
0ID0wjieZ1oV+T0D46aPeDn58hj5ToXdw8Y/urlNbYWLyMO8Up59TFf8QE3ZZ5BIxrPAzxZLNdCW
OmVkuRDXxFhrOfmNWSkKx5vWZxNVXDH1/hKOt2rGlbU0gko35lQ7coGdz5NppW/oqn7cBPFJrgdO
Dzo2l7irHrWQJzhhxHh+fDg5n0yTnWPAti6Sb7iveJHqYw+VLXloV1sKkRJ7bsFtjsrJ7J3/j4Jp
IGDHSrB/Bibg6HJ71Md3jbk94NT5bea/xUdx1KX2VxSTH+27QH9HKfuNddB5JNi/IXUC/uWsB8NH
kwvIZ8KY+XEQHOqoE9UE9z+KlVFpXDC/ppV8R3uyB4YkgP7BAO46AI2M8W3leewGWcL16xFn9ft4
TyBoTiVUcHLH6kmoiP0ug4Bt5pD/eUQKRtahyHH9uRIWMoGKeMXDICzH/IYX7feoofslzR88eBJp
GnfrlnMcQxdoKfemIVbvGE7I8xoJIBpQocFA5r4AO+J1fv0cI9GGCXjsg+/eB6FlJcFxvjrUcO8R
rrM//wV0xYi2e/vBKfNYPUJhozqHuzx/xkk3jj4KK9wGZSYGPSYmXi3IjFxja0p4vVXAc0VVs08q
bQqzUiIJ7SkGR8HfKh69PlM/hewcKgi2vllrV7VFO4baqQhdBz8S1SmnTTvHdlCtO9mSa94Egska
XQouT5XFZM+ydEf8i6OK+c/t46uW9n+U6aEDsrApkiAkXycDYRWUAKubCh6bkj+lwdGNCICTXIs5
BuA0QbWMVMNdpJ+RVVvBWqFOwKpjfp20aNDGwM6EQ8acaOn93do5vRul9rM6GUzadiD4a0WlSRD8
GhDsJlbsrgOD+wcOXQ4UM2GbxilmksWLEr/sz9J6bf4hlAxga1dSbeOPYiwnDKPGvbyZrbI3t3P2
fjpSckw8TOdncTtMDoV3JyiGg+v+052JaIiAfrCVzRwQzQJfQlHsx+QzYA0MvHYbEuuMZ5s1N4HY
0hqs3vGIoV3/LQTpRgkOIF4ARPMV7rJ+TP24fFQJaQzYXSQXie+/8pg8kmoBRuxPBup1f7rk1oB+
MQuooebLiMH3rani5QyiOiWoalukEJu6c/2NWBm3MR5mzVwv1/PHxj9p8HpEwGVEZ3G3dD8yiGVW
020tdCxLYRcbBkZljDxgCIwnInL0wpnP3Gc3dd3AGrtu7vlky3DbhLi61gPxlHQXNCe42uLzB6xT
s/z5PzoARYmSJEfDtzd1IkD+ZWQMMh5nvDkLwLHn3iLvIVBEf+fjD3OMs20wal+IisGBHYhTQR3f
Hq0ws7iSezFsTLiMM40es7IJj2N0Dt27AK7CqZL6cwh3NUt0FZDTjIfqPccXjGuIzJUzWyetH1Nl
Ciw2rZ5zho4Iyb/hkVbx9Bft5GR9BJpOScbhGXMiVDwlTchxMXOnlFz/G5dFhN62xPjEvhgKw7P1
JFYyB4+VQx6yWdmwGIK26Jf1NHuZ2OuHS+aPUW9ogg4T1g10zzOC5KcmN2aZna+AyNbZzQnpPsJA
APcKAFgILr0Df4rcXxIsIAIaClNxH6tykQd30fZhguBCoTXmdYVrdK/Pp7vJVrMjg7crn3cOEeGw
X1Cu6GIQkGyKxQlJDJPVKYrzg2sdoaCHlXn2PYgd3wdHK7U39zPuQrvxU0qTc6Vnd6e79tiMaVrw
OKwqatZQmqV34taZTh81jhkUC0GrxBGEeT4uhLwLxSKPDBkOUgGs0avH9y4LQARzNktVDQRd2ZrW
OFN8cExmgyIrHzojLMYp8j2mgs4w2l5SngoAyoO1Mp8cLDomERAirzg15s4JK6m/Hblu+Nwo9mVK
KEi+/YcWFbQ5QqER1xwTKoPCd1JlAO1MadZ+JUT71s/3KuLSoJnGBpocHO0gyn2LWGSiERhCmVP0
bFICEfZ33TZRyTPZ84MPDTme7dlY5vw38MvSpm9g7K7a6ptZ967WqO9mvRHylO1zLuhCKdlgV2YC
tLdPoNjAvrRDnuRsF/tIvhvQ8oolP0L1TZOULaFKXe6IjCvfvRnpE9MneUyV6hWBLKMO9GDwe5pj
bfa/TFHILX2xhgzo6HzwAMUmbaHAC+S/QDuQJrlL6fZCFUE8MsaQ/yGwLO0Me9JdyeKWFrqYqvDk
rux6hFiCvhL9BMGRwDPG61rypJ1P13rZynfKSXh1Bkp/QCJbCVQKAUGObi6lsCeAS5bHC4c0xlog
q4EN0XJx+msmOBTDUO64qOJQwJWux3xY1w4ZDJ+c7scFP5xIR47UoaVm8ygv6w6XYq/MZMmMFH/X
l6Syksgl5CPArrxI6PmP/CDvi5cf0wMb+fJbh51mNYkuQVBoOvp9RWkF2j8WXT//pUucOEpUdr9z
yHXxcECNKRpa89PPW44uZrbC0mt6QkTnZGrRTDuDvcL1FygBqcjO9sAPtdWAFZCBuoDlmcEWuc6d
ZqRapdhNZ+PsYycbU2gE2O9tf28sAE+aBVz7ex+ayaVJ5OcMs6HNxTTnjKWVYE4SWidSs9t+X++U
C1WnpZq5fDD6fLdFiHyOw8xYF3fTzqrKK0P0rL2zxlhWiH5CVc9IBeB3Ti15y3Nqz9d2CxgyF8Gz
dd4qG6KGm53HAy0xalZB6syCfcsRomua6nVNz1SSFCyZCAJ+z+eM+GSqjZubjIJxA/cFOF/rbUcx
XA715rYJgTgi60zUlWl2uhNJWt5THgErUIlSqvSJ0rpBeuUz7ebVmyn6u6d6pQJuLCiOpFEbZaQo
gbLdOiS4wd/iXk6o2szwrb73p3EWkRMgFXlCL2nuDfxUqAMyJL9WNt4RHwylHt0x0qobJl9KI7Mn
IUcbJk8VIj0J0aRYT5HrZBZCbemnEn8iTSBJM05zPI4HMFaX1LSOaDBHSdkfdnGCf+2sFwoNLWOH
mGlqbnPTpgYbqzjINiXEa40RNP2KjwKKVQZWtKzCAY9DQnzdT7qSFTtIdr+5CMHCt2IKQKJS/+UQ
xvuzqgYZz1n+cMFJVTZxH1XOJnIbuVCHxfFPC8z5bN/lHi7xe35WymMcK6fDE8dp0BfLGaoWyAbE
B+GvDxdXF/Wc3iCqoKAe+/a/Ps13tATnvsNWvgDbfq1u71aV1rC67AU/qaB9bKpoXZj2uVOCt6EN
hlAh0jTIUWU6s+ltjhozRxpi7rbbvisofsA3cVtPaV9n9N3a5hgRh2/lEIcfgysHqx1zd9bQJugp
jleGZIIwcBFDOJZM4Rtu8WROqSfa7A+h2zYq2tJ6QeZKebt/MBqzN3T4NhZzP/qjvLF4eOt2rqQw
H6kF/9bUkWQ6qMaDnwYMcfIgRRld50vndc173xtPpSgKcBAIAQIEplaFyFbJRN8dVnhiyt3/+5Bc
GLJPgW6t12m8Jees1VYv50hrvhDr54DuikoR6774tkpT6Denx/4ClSe5kdRY7Ex2PB9zQQzQquGa
q4SyoErfEzyW7Gu6xT5U0bJHlFlubbvtEGQZxS7Xs+9XlfI4gwfXXXoXwo+aG55oq1xaDHkH/9F4
AnYdkEbAliv+Uah9Ay7WzTFGL1Dk6lNIGcvtt0HzlWbpi8LwE1u6IQ9XABdSnwekHdwag9JDF146
MVIjX09cBILlbK6wfUPglI4EEkYyPplAzRTB7a+e/50grbLs9sCUFnqKKgT1btvb9IMbRb4fFnUI
IzNxS1cY0Xqh95UADzgLoFuUNSBzit1ThsauKlQz5KRnkY/SCDH/JK7K/GoPKBG+Eg10Q5wqK0Zw
+atfhhvHubwLFuL4LrbY6pK+FDQ0vwZTT0Df2qAcY7vv5TtjG8SLGd/OyzeHTb9nsZmNR0l1sr3S
VyTT655xD+wvk01kxWKlt+s4r2FMivpqlfmCkTU70T00p1lSqx1zOR3HgrqT5p7tbMHb3SNoCgtG
plXT73kPZy0nCXiQUIVRxKRJDCbWOP3LCBgqBNuSW7R1vD2WBI1Is+XqWA+BFSLnv8dH4bv866ec
aOW3tcXEjdQw1MRghFl1bpat5qDAe0S7e+yrvVhUdPV4KdFvkHju3RZ3iPUQHhi4SPf+PVpWOviU
vQRCTagILX73JGxTE+lOoW9huxwa8lLpboorWcLS5NG5N7qDuhDjmSfThd7krVykT199L4ASi4Zx
45sJZCXJ0XHmjFRXUluHf7ngQpdRokmrYDgiosc+QLbC5hBjZePPDhA6y4E37UJn1dJIgp/dNOxQ
mvP6SykMarNslqPzbrnkPgfeFFCY8CBMVxqX5n8XnrygnN+laimvZ049sPTGTeF1SWGhGsZhBZk/
CWRcu4ADAzaKqFiYvdq0sj/OfKdeFo+JhBHhiOap/gLCoHFuLVivVRN6dCS2CVt1CLeXdOJczmux
5brsDJoHFwY4G4hndrNONqhARIuU3s6zJDGbcuujrJO4i4r/p2Rbn7t1TOCwOJS3ZE7w6VWrakkq
eQ31U484tJriovsVTtK4MsLbctss11Thoi0Whr23uev6lUb16NprykdkhWQDP4iYtIhnYIrZ/cDn
SQpy2Vg9pAINanBjL21z1HFnEp9DP+LghjuYQDudUmpWNX2O3Uzb53jfraSD34Zjr+U5fOUUuGhF
jTOsStfOgMZLZ010klD+vWzh76ljjIDAYAPxS+UaTaoWtgxqhvMJNijQ36QhWG8Ot5Z9P6++eHih
F7Ws08qbY29qYIZwHgpnfT4xrhMldT5gTqHh2tUQT8UUo+dXhSbsGGSDWU/LNTVSmm4r3MAyHpyu
u+urYThP2uULcYvjAkWzTRVUoD1/KWoZ20LcTa6UBn2+gujgK0obWD1oSCI6dWcvKaD0RcsrRkJ4
8D42aAw+gJM1tGjmUVeq06mLFcMbPaZa/0p72BznXspYCY4kim5szEfPC786y6BZcSqgebRQuXn8
9SfrniBIzOF9DsSmJKXcRA2Wr6mj1FMIYZ3t/i/JaWsRg7whMPjDiU6/Lq3L6QL4sl70lXugiZWx
TEHC7/BivgBDFp4wqviN56OTyjY9dqf7XSaMwAXMoZVra8rrvq/aWndIjH3XIcSwa0pBGkdyvGyi
OPFZ4ftfbSN2q+l2MIyocJCqziKvAah5qPF1PTMy1s677xkcpfNcGvhkAHcqioS3bkbhq+xeqnMX
u3dLA1fVEgEhRED96WBnRygCfWM3wdmP2MoAkjJRh2DjUlTEDrjeA1P98MVJq/4bSOCJd3EQ1qsh
R1LKrH2eQ8DZEFKnfq99RZk7uoGrZyBpHHfFTC+EIoKhSCtVwfsgybkkpVvaxVCEddnXQojzDRMx
rvbjxvLc5FEex+LhmWOo5rbT3w7UObtyRQJI5t3e3IpAiKuCDC3H0D+O50nPB02FjATtypB3Fxky
MGf6Dm4//PimkhKLwCNuF0TuRwGDPfMi3mJnw20yGuKOR5djrSwLJ9YTG9oX9929xPm0EWXUsJbS
99hr5v1yEnn/a4RODvwtv8+HAJNRHyDLdM7RxvZggSZVc30JbX83HDcZ4qHZFiARw8kzcpePSVBi
l2UeFSQfPJETu1jfLkzz7y1v0X0DHo3RUgEjMfZ62SHcQbLbbDknmqfF38T6HV0A/qfj6Gi+QomS
Zv8djRPXTZn6rvJTef8j0CBLuaClXbL4HJY4A1T3WjURMnexad7/nRzOcAoxVE2KW/W3beRozV1s
6csa1QjjQRjNdqd/X68nIkXS2VarkEoiSAH4CrLVE24sH0jsIYKy1eyrS4DOtxrw+kQpPooakNqD
I775aKYsmKzkNfVIH3boBobOl+mbiYpkA/io9BcVW+iCafwhtNIdvgO1i4EUs8a+/xgw5fAKQRYC
NrfHFqL4Q6RyPFGKpLV0YBKfPvuMth4sShCUBib4ualfaImXYnR0rg75gVuehoIgOsQGVOBPPHgZ
9YzrsxMiH9wKcysp/VmSQZSheyMPuRGlW9E4Esi2pxey0fI/hGzcLeWMc/3v8w+a0+rhfbU0uV1a
BhsyRNoHedtUcnY92p1V87K2LA7CTFFEgLOwe+yFi2LiGLLkvH1ZUN3x+/jKzDIqM4z3FYb0EjSD
IlfgxGDdeJUWu3HkI3upVjAYrs52rbhkYl3gE3+BQVMuz6i5n0jR1EmwaWRIqgNXxynW22lP8AZk
z07omcTBYGxFhG0fz5sNFaMzsqUzLULT8y9mnqcMvJ0NwYl/Wt32banCJlY+pFYcF7w+E+nM7tBs
ZmUIUDjGvVU3A47mqdncEQeG9+XX2q5ncLKcPQsa546fBPLFW2JyGjL14YCaXzPbCNyFn1abZ/IC
h/pthwINIFqpnIqhYEJD8Iwz9tfe1qasXMtep6nbIRMXzxUywJRZEeR9JRqVkOKzVaBVfOMPy1hk
dQzTbjp8IBbeMWimZqyKXS6Qve/4dXZFtmZokYyVdY8kMDPiI18KnowZIy8FRXG/u8wqIQvDaCcT
lXBO+vnMpGQSfstrvgaaWj+ORnQuVceSqllerzGm5YqvHTkBPOftNDU72i0U0hbptQ0myGkn3vjk
CRFzn6MQgBtRp9gggaccQ9JO4F2TzMz+tpH/25OOq2s2pkLjE1l/bqtMdHbaxSLz5bkjRtyQHSrZ
Z7jFQngbASgH5jtGzda7RFTcRjZ9d7xTRMIfdQX6nQvcQgffesLetrV0KfisvTMEDDFxmk6S0MXS
NG0DabIxYoY73TzwEq3raK9aBTGGGoriORuXtBtP5yu5n9HDJ84baFm149kRmmIJv0yMMYuNl2lc
nlRIXuRvnORNzCUF5zuDUdd2gqU+N2EG1FcVvuhzoZNMXpe0SVkuqDLlR3FVnFEsdj/HX/avvV2R
XkUmoCu2yFt2i9rKIzXVPiB0zwzTM9/wjSqcq+945CdLtJk+vbtnk9oxnxAxoQkxlB9Cy5HuCUkj
WrRWul9KWh45rzS59/fUPntzMOcqY1PnM2RgX78HKsceEmoeADU1g0oYKIFaLIKGFVGdgkrBNag4
1xX89VvM16RsTo4Szp3+CvIZIbntQjfqktYUrvjavUsPVe75M4VyxUJTITHJu0xxJxswJFurOBDm
rr3mX1S1Qje48580J2N9o58z2fdG2Y6BQZ90vv+qEFrIX7A3ObDIY3Q50I2P6lNpjX/bpmQgs1T9
ZbHRSyye0ErUvVIh5Zd5X2uvHlGUmwbNIdCajP7QUkEpCEM6MRMHufiztRSwSqVH7t0FZ2WcirfX
0USqlHMA+EAYujtEOHsCc6Gdf06X6wcgMB1sAuxl6nwiwhORr/WE4OYrwKArWNaQyTwVJhfSQDTV
6VOQA8fyFTvfTiEvfCrrPeB8dS35z6GoU2wIlCJ7DUtI1y4DgIOZ8mc14jv8p5UJ4qXpXCEpFk6Y
nwTtY2SQxtySdZtCua4g89uJTGxfHYt/5koVrj+q8yXY990GB/Wyy7iFgYu2zW2EhtIRZmRYAIwp
8doXCphU62eab4slnm74OmH6xV2R9YpQIDFrcdNry3OaGK3X6wRIevYKgn4bljulujI13Gl3GwOF
9uKaRJjAOXckMpeyYQH8nC8EyWJ/k2w2ngTtFmEm6tmOWCMczieF685Hm1G6kEGJLZhFWruXYuof
oHIvS7TGoG/mzB8eJ20+Zbjzf2+tM5ivZFCzWgHdeLWv6/VoBOGGUBk8S2om28k3J4OQtWw4VnOc
Ad1xtrpS/VBzQoMvffuG8CC1ITJJZl0ENhQu+cc1bTQwzJqaYsr/jmrZdRO9Qoq29OW9rbdiFnoC
U5U+MYxEwd8D8aSskM6vcCaYDfFW9CoRL56nCeBbZRUsBHOwVw/bOPDkQkTFSsHk5oHtXjQ6s2m0
cRgu2BTTO0yq6/9zIQYq4k/ru4EBJnC2VxXaADtaHHoQAyBw4UXVGVvdJoFjQ3y4H3e06IQR4pF1
6OBgp7t+jxLydabnd0WZRmzDpu48UyDLOy5vf3tcgNqqfSVmwFkHT1yJCe1FxWs7ZRhXVpuCryFS
jZWBtnYTRGHt0LNI6sjN9NWU8DlkU4Yk8FEuZB32haXn+RIDJt7YTBepSELBHMCMB00vPK8bV18H
Tyt3Egny4z8ssB9yvbAVezm/Av0XdjI6R7GQXYZuS+sJydc9p33aFwmJ9Y/7RAlom3OZhgBjq69Z
I23vfUbsCgN9czrnDMt1bjJoDlMDoMs1OkK227DCq4UqrMbQ9ldj1AvHq1djfZYt6Pb8c6ecTa/T
L3Xfk8hk5aTnO6vYsdGu1bOdcUVnHDytrAASmly7XZA9wEynuiU2EGqOu4gVC3xyO72DKr5SCZ0p
oavmBWnAkyLvM2vAnUfCwiO4cet+ndcweJnETFKTH55iX7HcVpzNqpelAQojHk3r1it4rqurOiS9
QQ20KI2LcVjQgVfJfEqlU1+dOfY0vyQ34L9gS7Bs+UKKnUWm9lD/n6SFEQb0G/bzveGVmYcj8mYr
1hBsPMuIxd6Xc4AqYJo0Yg9VRr3/0Yv7Dme88iHzwEpcgmzANuRJ/miGBb9Ug7c5pR/HCRh40Fyo
4t0/rJgj4co7AVUE772ClDz25eWgnvZkmldel2s0XKv8ijlGjjzJe2Il38NPswQO6RNw/n8eWau4
9uvSu2Tc78xzCg98uBBvaBbnX/hnpOsoBebdry95Dt9SRZYhDVyqHQzoP3MPMS/TsqGYbZBEI0Tc
jmcD+6KGCcJC/S6C2uKUKzknC6zbYA15uyb7syHXYVFDNT0BftwgF0ggIcJ/dABrDAzEfrLOJ9H6
grqnhitlgA8dj46hVXNRjQXycFj5q+pTPD1BSLM36JOSDrO5WvXsx6o1E1f/cq+DmKYCVUa2b8kc
JVuUt4gruLDxaKCpCxncf+bnSUXkx4tedZ+Re58AlpdCBTqG3Rf9r09g5O6gR/vitvIeRkj4WW1Z
Spj87z3fbzglcP9bQQRy4hCVleEsOIoTeV8B+7ZInyqwDM88FCk8VA2D5sKoWIqPOLkMO+0yfrEo
/AglQ4rkuE7Dq8uXR8WnzFk2jjZIHSLFtG/S3WstOTcarIIQY/KGRNGTzVyIjrklQ21nrM0Il5o7
jMBW8/qeMljhVoegfX/KWsAfROv7/599W9mYWu6I8wlkG5ErIgJDZS/nPSNgB65PmLxDimdXGl3f
vbuOHMlQhg8bu1lu4M9/png+bUQRe2XMfSWunaIAQ4cmUMkhUv1RmuiAtjwmJk1lqgTUXdLsapKP
gLXD5M65n+8d60m6uNRuY0oZCheke33v7tedj1hDh0DPY1RiVfI51qMd8Zx26dS7Ki/987WiMjGH
9SgusE2on+R2JNHvnUsrqogWpjjAnyyVkcCoWyQQLtsaMJVCAFCG/s2511CTxvECOX1ON7BCa31u
LUYSfLV1OLzmtAeqR8wzrbBnoiGt1ywi6GvRJOQGxb2eCq8Q451dPJDC2/Zwf1NNci9dkOtj2xLX
Z3Q86DyL0vRXctykW1q2tswndghqULWcpCcAOgZr7rO0/fMIH0foU0x2SsXIQCirrpCOLxRDbJrO
2JY1IXVZomRdFW8vQGibaElIY8+643DrJp6vWqb4leAzAMv5HUR0hhrRfqiGwvG31p/7Ewhwp/bC
s+lCrVIvFA9j+zkWKO9ticfuDlfH/1c595iCpfPnI97BztX3JRtPyyA+JMqGjfPvSnw7p3js6vlV
CDb0GJsLzK3ceJGKj3aBIiy+hgvIMKbRueE45BT/v6Pq1I6bg4VJdEyg5YugGbHGnys1UIRP1Sgu
s+47+OySUDTtiNejCoILUpNsbUCTHIf8dHoJbbVRCvqVmXY6h9nT5uC4keGSiyBgxtZe85wvpy4o
qD7Oxn5RTiXUocz6SIP/nJNKlKNS9fE0/JLsB7Xzaa1rIsBPVgCRr3mb9LYXqTgfpyZDLm8XPq3a
85HsQiTwxwiTSY6PPaIKpFznAW2lQgxls1g3kCH1SqMxFlCGBL+1v4Gx8XYtDvZCw3P4Mpdo7UgZ
Jt3qyoGwp80UJHQtsrmOHBgCMiViF2jQKZYlNghp1X8mrmSalP1kEb5feGbYTjgZuIvk3nsjUPwy
qkwJXxdECHuABuWxfilj3c8OGYLJvvW4FEt5EKYzWyQQi1VMV72KcR9Bcf/186Mba5dsRTcJ1x9z
4UpMNjUmqGR10t9MNacFw2QZXst7wVRvzJ71K9KK6+iikKVee+WlN3xuvFrAkuvTCEHpZkSTlNEZ
Sev97wzQrvJ+pUgUWkltZq/j8fuftQl8tzYXT8HSNazW+Nj2O8q3Qdz2+wY7iQhB+3fGkjWhP3nB
WnCojhNG/TeJ2lF4ah7DvVO6OiTVnkXVkYDdjwFfW/Al0i0SM0d8vSJCI+86LjTlWeXdgr70J82x
1SLcIzYaNyaY2fyWkE5wsmjKN8GpUyQJKi/gbGmtY9cgcYHWx1FDko/4r5w5sQPqkR6qDtbPovzB
jijv30EXYz0bzzQb4dDceglykjimP2w5S7BnSuqm2maiguVuKZlZv2yLppLgKkchY7Qnel47EXlu
HMuJ3Jel8OG1ZEwhvXXGt/yYZCFYPNDc24Cu+33yf62cIsXjvFjPF4T6mbrY4XEdJDyv+xwD9Z1+
vJ4cdvl1leh3YdpmUJjiBXa7JdWevDIb7yS4C34ziXvJrdV2HJNf8XTV8sjy18nvVmFRH+DbhIY4
kjATV8i4n6i5ZiAZv+AUg1VxVtCfJiaU1jw2pUoLwSauFgEOotxdQjKdKEeQUIMWxAZtkyo1sB3v
o7e80dthHLKTD84fOaNNAfbkXZTxR2IDAvBTcXUToso6kSMkoKTDevXaPXeYM31M7Jur8/It08vE
zZ2gj6LQho2UvpO5bGpGG8SgL2JEGcooERP4LEXq9T0fwDiLJU1Wr1xtdjQmQBJRzF0b2BtVxNFP
Kv2Nu183y0chGoWB4JdIukg2HkjsEUALiuS1NwsO8u+HenHDQQ6JPuLhmKT1i6gfdgYiEmW+mdZ3
2QPC6NRV0epEJvV3OGH5J4Ucsmwb72HWqBRZMoVerEbRTPPPyAbnyqO0VHepi/nuowAHNPefXSgN
AwZIOYfwx0ZneTKuwID6loo9Lm4QV2t2SXILDTLTpOLg6XjMxCr52t1UN1LZfh/b9C7TGj7M8TQd
cXFUobHfXY9dUiVvAplV0UfReYn+aMQCYljv0hTP6bS12J9qB5jkX3ybToezsurXpM9PmRQrFICp
cLRie5KLUlwTgAXWc7+h0B26VnucubtGFGPic5fhDt3t8/NZID7L7l6emkV3lYHmmKbZ3LVqZlUc
NEsEi86PR0IGauhQfuXckPgMcO8lg0xH7rXSIllbmiwKIz38b+bQy34VOw+9oQUcoZaqJUtHqHlz
eoscqClge40iKzd+pwA6WcrqszCKw8JKY4Rdi3gDEx+35PlUIt2ZJIjzcTEvxjvO0JiuvARJiXeL
FDdHZ9SdQG2OaQA7GvlNQ4jvtyA19C6sPlW3uUoz29a+tghBzBbVs4jOIBSo7qk9LWw13rz7QBiR
7vb4xKLVyxYxsACWXEEu1weUiH+uAXN9Ubo6tcoLbbzWigHLgTVi9pEA+tRRTS/ZjkXZ30bW/okV
+2TCcjuCgPj3tmcF4Zjc6GWm5iR1Y9Xr7M04Onvgaht7esSlMh+qi/BfaKJ6KMOceCjUCnZACTB0
I3VnocBrXbu0+na9Q14DmIPTdqi31knw0CemI3p+4AoQe2opH8ytaW0QvRSRFDCDS9Xcvb3TezUf
BxAOolQBJOySz3q8A/8fbYPG//CLRl5BWsj6RR/ICsSx9FxOrq0hspE2k5RNPY2hbt2DlZWBvlnl
MRI0y5YGfZ3+hZ5hCgSdmAp0+3Rbi2EZ64lyPOVfXhBPz2KLl4tQb79IOj+t0KLv0tJZ8zbMuR4r
mqv4LMqQgnUZRLNMP63uYyRoQ06Tk4Ki6XpWqqaur4vkqNB3OrHIxvJ8WFADzRkbT06WAfpCAiU+
8MW8gmy1pEn7wUCaI+VT1hTDl9Ef51LPB//GT+lUR406rYt2E7y9lA0NLMYQN/Lf84WO5u8UGUHA
4brs/8lujkSVdM1QVTdoG0uWe/0x/0GHPg2QjSRRNTuPieko0S62M40/3CUFuk+emF5sRRLgjj5D
gwf0SnQs0gamXFfFUgOuHmxaoVT5jQ8xbcagWQhufLJDRskBMCzEwpS0n3xetyPMjryP0LxLjasr
MCPOC3qZHdNwsul9wgG6DJjOFVYptamnkYsE0lU/tB6C6Nt/uN7ZvFIyLtIdPgBAGVCWK2kHdEwr
2NTs/2/ZYDItZrnRMnqC5TaLCIIOGiyhLIZLMrFLISD2/vVQiC6p2d2PpDK81I3A/We5bw4sWfN/
nFSBQ1JBo1KB7Exk4pxRdfF95qRqXWOSnP6wxaiXJux8VlfHLX3MJTqnxEkg157vQ85CgeMtXH4l
ctYi8Y6e9WYMqBDns7uahs+O8fzNr94lZB39rA5h/sRNr2XPEwfIWORoSZAsvQg21XScHIBAG26V
eJnSHtx4AM2khhP19LknVcPSa1cv1J3MG57ZRHCpoI6a6EwCFkueLGPv5Am8B5a+IU2m4+UQuVVm
tMIKdS353gtAGVy1j2J8OsPG7a5N16QnSLu2Ow3Lg6rpWUh3fRruszG2O1/60HipWvclLspeOxSI
ffYtPBS4wk+eqgl96fAYBoTFhd5X2kunVZ8Pk9AfdRFqd0F6/BYgfp3DRFPAaVV5VvIXpkF6Ivwq
pLHDriZRRQQWC6NrdHwKu2hVRXVKS4vEA5LcS6JNmXvInTW+h0BDOrg8n9bXCvCeTkvsIZ0mZJQ2
EiZIhW+sscd68BNywWiJekLZZtA9RgWABj6p1haY5lVPz88oPwYoi/a++nkFU/mJtaoI7HUnd7vl
sHSyh7snv3IyYuQtwFVEurTIZ+7rjeOIh104Awo8/eF5IYV7Vw8TUv5cRJSdMl4IJspHqFwlkCJu
lEfHMAzqlae8X2QyMKT7BleTvydsW+Or1YsdEwaRPrQWh1AqSOn8S7krkeyg8D4jhqB+dDyr7lKo
/swF4mT9F0Kd6ipwB7jbH6/sm/qadeeB1zCgUa/inqQWUb1Szd2T9lt6G9bsXzz2euFTK1V0Lr/v
J8G7OqcXUV3CNwE9hbNXVMBHrA7vEoxpBIPSxf57ArQHTQ7rahEzpCDjSaJBp65qZkRMraVXvkFG
ArNNaAsxGlDR6DOllg1CnmmBittsmftRc5Y6MqxpjVXYyMlEf2GNQXrDc8c75MY33opyngAaoAG7
wcweRuGMZ7oa2xIYyz7jTxZ/vu4wRsbmNUjHFYUpaLseR3dq6ndj58Q46YPBVwtazUfGeZ3H5wlZ
F0vG4+iVqS9H5pXptDoBLTauXOCjw4qrgs74VsLDZ5FaxdDuPZ+cAUUYE8j1hgAl9F2p+P4s2MTX
wK57k6WPSx0dCW8W5zLdf9ebLkZxBlqmyB5JW/ey27bMPJnFAglisHKbItG7N7JPmQaieTZR27zP
2iZG91/LiU/UP6QPBuyTB3G0MpTsWSdI7jtq/MR++aY1SZeiR0e7NNCNUl5A/yClFyE+sAwMubmL
RdI3SeeX7PrSHs8saFhfF6MtKAvsuihGJtx1XS7hcXJuIa+NQ+XnTqM07bjh72YRT4G3jcA6ZuQK
l0zXXzLl+zmX7uDYb+AJIRmlY0niQFeQdJ1zKITkGdwWfaPkFiRiKXgIE+z0jYfKYgfg1zt6GeyL
MILzDCw4uejDTpfUo681EqPtxRrRaykzbmOE3zfZnWr3pmYiSNsdI+cu4jwhBVfTrMUR+DQwKk55
siccGK0H0KWloKqgiJymt5tPoAeee2oBYUH+XCSEnSuyyu/WXJczsm9unc4ORWjfb/6ZyiJaHrXu
M3OAEBLk9JSgrMsOWj3ydUSrVJOrVsNpD5vqKSblQMgRVeX2jxdIeJegY5EHB7IyFj5ekl9ksulk
rlHasZwf1tW93uJs1ona20335+uf/GXccNxp5uKdcSz36fPDnK72Y0vpFDt4/JGyWbB4OkOWtZU1
y0wZVLgWUXghWWFTIpY3MDBMKEV93eBgGoRxoX20Pf1RRSRaOH1Nx+rW1nlLcAz/4CaxZYH54gie
cyCFmgf6VJGvvHBEiQDKWl7L8KB8AdfVEyOFCsrD9Uiampml46LEgnv/RdXIFSapoclQpCE3XoCr
vgJi70+EY9Q4plWqM34hjyFLt51xHvWCSiWqQb4qlvxoXPZ4JWV61sU7+FWZu5vhCCpwXjK/ZK7B
/sYcum88/IOaWkubgEWWjHyPgSFjwbsF56JOxphlpQrQbN18V/cZB70Y7VvH4//RusOSQud3xcr3
FzeUIkbH77AZbriG/OQkA8OrCflKKyv3ddTq8AKzKRfoq/jP8EWuqUL0r+ywNj7XjWuE7dZKRwYb
jHivPmG8Aw+Zy9cVyN5E16BRxAco4x66za+wR7fCTnzan0aZnthmydERtsQUSI1yr3Mjw0cicxcD
hRR1ygtTrOlplb50XEYGQdyMwp7bqztJxuNnDXnNQaMVTEcB5LqU0eSvATNQYPT5AE9rNuCt9xHG
EcIj6Nx4G0XFQmYkaT7Oz3gDt/I1aPwQHKKrPp128+3DcAyFpouIvpyBrWxskOyLdcEstALoe0ba
wyWttoE6MtW/BfXee/SgMQ9PFgTTqnm8aHM3gkemFK0g0IjkHcVPo8tMn/IApGEfXAcdt1agbPZZ
zoGJJJGNUeBUGw72CXge8/5SEwpywkiDCVsmyQc9ruWEpCREPxSb2hxZakoLouXkEC0QBY3mv2ET
y31CuXXburuPsYHSv2IvkvlGcfb+pUMe3vCYMjC9Q6TKeWXcKUWSu4+mf8Q6hUH1L9VvMsmeztYA
RWLDTQGIsjAKqRgChQGyWurqSC6tU6xL5tuhPajhOKWYs6v4e3765TiS+05gz7Km3SPDJ16yAlNd
Gg/vuV6rv4m83OiUuw151ExjOTbymVSb25F0FsFUtPyfax+98tW4QsucynKrxDkRdM3PxV7YPgCk
SpYoiLAIsPTNo7tacWTXDmKhdDFLULyyijMppWvaygSbJbOiazqIA2UccTwDOOTAIHVJrTG9GaD3
CMxdCuU/i5R9xWB8EgRFtF/L6jJxt11g89qLPHWedjkcbQxf38S0ddyeDxf04yuhvF9oh005nLds
uyRE2jGW5tJT7SBDvm2pDApkuCOP5NILkczrMKBu7j2YiIx8vnKqNY8F/f3tVQOcN9+cKDduO3HH
BP7TvOlgCNtFDufCkrI+U1yDXaRPbPRj/Zk3qHrwWTHqvozH8SmOhqBRuecMtgRlD+Mzw1wDUi1i
GGx/Zy8in5/Bsydg7QhPKreiMSpQoQiyNbRWf9y5wLnma+ThOiMO+oMLe/iX9/NcXoP7dDD7Xeul
8tWF1PMs57Nyour2/uJGtJGtzgdOt4Hl6Dvu7BLo/EbCUj6rRMZqojfJbSch9iB7noKnssvVtWY7
OzHHIzdkEpGm50AZTkwOut1SZ5SHS+ZPwa8h68sV+PAfXDuKwFImOt8hd2CRY2+uM9GVBuJ0kOvU
IvpKhsnBKAtYVfMZSIav1Fr3SyyGLVD21Uzyx/D8KUvBuZW5zc3cvwZK+zt/gZe7Fo0sUBjjlsP5
XwcvZgDPa059YKBVutV90UmBfpfP/YJpG9wvC1Q0Zd4SHiqs36sLBoxt7dxzLcywmkTOIZXRJxTP
ZakzgC3epvGPp9FbGNnUvjwsnr8nG1MOzP3hjB4o7AOCMtkIJ+qGd3fG8tThSH4WiCwT3EfleAMK
3/h+RfPi7zj9q1GbepofELz8E/T9J73aJQ7eIH1kMMSRodz207pDTv1W7oYj5vHsGHiVjKvjwwB8
ZjGNyElmoEhLtX/xPVT4Y0nhXfI6l/6lCgofM9L2o8R9uBvslg5+wTt+QW4BH9tpw6NDn8V/0wAa
FAht7UgxR3bkpGIlCE1gb5szN4KyGwIxgQFlk9GgAurMK5nZnM/crU6EbTzzDV61Z48eO44u4nIQ
sI3cjJE/oX/enHiD2z6R/ddTGI8hjXTgPTLMbGIaw1e8g5UgjTB6wZZUbUfs7s6gtglZ9DJS9G1D
PomRPLmZmKzSnsAMzOi3RglFxPEVSfcWuDo811ExSBEJar4w1XldOnZJh2uh4EJ6c6e0yCWgwR6c
2bL6kaL/9+kSOe5fqOfyPDPtvc9CIvBU2uxaoX0JcdHOvlKQDrmgtDlcC/NhGNCVNP+Lb9CBzF/R
HDyyuy8/g3lnf0MDbLOc99hbODUiudNkqnvoChyTlS8JIku71wpFWYtAc7H8HBDGlThw/GbacQ8i
WVaoT4PgPThzR8/xT0XRX/PHm9MnoUe8xXiBMBjMRXqHc3pUQk2GM7ECv1V7LJazy4J+qoUtxL3Y
Ei3/j+mdvfzdqTrA7gcEFE+XVwxN7VSX6uLVOwr1jBjbfeRj8o+n1JhGBmh0hI2y26nbPjPzdxHX
tnSEibeaxRsdWc+Wu7uPf6tEcx2dYACWAsrtCnQ7gudfFQPUz5GrZkoxGHs3Fdu7KBS8PnWOuCUF
IEEAYybhu1C+yHxtblIOATseDqr0vkpLsfD4djNGAexwGGfoH7oLdCA9jsmdovqoC7VCgjks4cry
Ez/1eqBsCsH+FnQrxfXewbes3qKEKf3pHleo4uej5T8yPG5os2Cm7WRw1XLIJ75j+/OhJaVALe5K
dP4edXE0rwLPV3YlW0KgywDJyNrdi077yiq7vE6uJwfoYp0XjxjcVc+KD8Rb46nhMSAG7vQqRbvM
XEaDI0l6XILg8BRBKo0qSq1XiFh424aNZECTEPUuMzibOhhb11qP/dyTZxLYxomJCHd/oAOsfC16
vMzb0rXaEn9ojbtcYSrTix3cOLfnqZ2icg5jg/VO2GNR3BPsUmqctuE2lITpv8Gh27rPugKkMZMd
ZjO4dEKmqv1vD6TlBm1CYpiA0BGESuwSUkv1qWiy7C7zHw3c1QSca1USruYZAox7JP+ULGuoJYr8
KfnX3rSe77Fngx5kXITn7jcU8WjT/3U3MC/rWbUPB6doY+AEvxBgsVHOBuPKCQ50gkhMgjWLLfxl
B2p7eFFj/RYqY1iP44W7jLv/RstX3vXr0cKot02m+M05fyvVEjubArIx2uIZHglhE6jUqDw3ksr9
oGcfNW1dhMBDqpBDTf9q3VbO2XUzHJr8mlrRPb/s3NDRaeFaJhR8bEBYRQntpDsBqX3LuFnDGiV2
W9plyLKZ0vUIFjZ2tILPl0MnZ1SXpoW0bsKWN/mEkcSYC95lJ4weqMml0HgsjyUcK4sbsZZEXvSP
M/UOveHRuqeMOCST82c32s3XFkgrzkVqQBVaYcgJgPtc6IzjFBl/1NNEL46IMYpYA/zOr54Xj9IF
zSCERFY1febyuOp6rjQRRg9Imni8WW+2hCJNVQUC+PeFAIT3P6IUTEOnkA1+oo7irUOtkzgxhSmy
BgkUI/YZc6B92cSScUL+04hJtERr3b+eH44kko/R1uyAZsOdpmoT2DQF+EpqUIZTGolToL5oenIc
71l5H0H7ogiedSnjdD5k9ANZUN2A2bcVm5+3ufIesZgen3gR3wTxYVM2ffcXsfj0gbGyDL6sgFGt
hTubJdlyiycfzU+gtsNmyIt6y61Vk3apH/fyI/KwlqTIsrt7GufvY8gMkHSUnM80gbZfOgZ7F62X
j9dik7oQXmPROO/hT/cG03M5Kxm/7gwBIKhqDpQouQqETJ6PZ0BlOsnhAgoIzKTzQ6phZrUP8Bgw
37XvXAuDCNPMmnd5/YBKJw9s0LOtrErMd4T23O4zuCtyNgA0hCr68eSQgVOQq2kv6LIipJ3wFOsr
a75SHFFaCogrR7ZTJuEcG/aWb2+dc2hHhOGzz+mWV/NUbjnPCI29rk120mxvgun/Aayv/fsOsda5
kpcAcndzXmQ7XpEpT0/rmNiNrXfg1L1fMZyYciqJ1hMP7nMsqkGpp294clhIMqG0QbzCVl2RD+4v
EYmMLgVH6sgQyciJ3A+u7nEYcmGzgvw3TRNfi/+5VizTGaN7tjKVPd7QFL3XMmahzqopHw6V2iFw
ftNNmUmbiNsOef1vYTcassZoj4XG9u3w1V91xOXJov1xqkud6uFubLD/tWdDQtzgb7qjarw5dIW4
mb8MuPA8LL1wUHZvLS2lN1jThNI8S8GphRdxuLvt2hhemGh8B6XRTXQKfYXn5PLypnLfoldajkfM
vyiI4p8NehhEf8+ESM0TwAvky03GHC7LQCuNh7P2xzvT8TM6+fy9ubvEf/KHOCOS3I6wC4pWuDWL
T3gKL5aZWBfPd7IjDHbrgJ6OQgaX3wa58dWdoLe8QIENe/b5wkngydmSZ03rTpObpgpllaLNDvJN
3ODS+gDA0daY4cV3B3D8lueLM52TzVqN7eDyu2+f0xlw6GpuGcE5Ewsxdf2ijCcUWALnBO++HEUc
10vMVWRHSyUAE2o2oR1HArRj/ptny03bYPzozlBOvPK0aMu34vp6pCpmTOOKPwko4zuvi67S+H3K
kAshMqwmZujt6sOjpvjoTDCrwA3/t59LgQEEcLQbOX9KqS3KY8N8cDiKiaF0I7zMcQFMOours+Me
9BxuxwGi/qflLXAw4zTO8iPhvf6BchxXtvz6x0vbQH+E6hOomaFeS9+9OsdWrHiYtO56hmPcqcQu
Y4CF/qv/sHJqMxWQMOA0vJzNi3VM1YfItvA95yZTlviTZ9PExKVZu34BDCbA5NvuFV5y/3rykems
LzWoHChj5STtT/oeABmYhUhP+s05i3nd7QqoHDZ4Rcr5PRWXfJYAX0q7exx/EMzQkzqQXztaUCsT
l2ZZGBnTcW6hG+cwNMBhrnp80DQEHvGqmrlZS68mAUAOtHmX7diQoWtgAsvwTb2sm7qKYK9XUkQa
fRTFrSHcI9UTm6IGrHgYoasInSZCdLEzN32I/ckS4lPXirYBrblpZ3/phirCnoiguvOYdqj+9LxE
j3mjZlyR6a8lsUIR4AWwSRyp9zSTqdCQCZtSvhC0Vc1x2f91wuitZteHrksGWK4IBqT2SLlEU35p
FqJ/111kFujWI+1DK26cN9/DQZH78JDNn96GymaL7RGgHPZ92JzgEFR6unNQvvUAO9nI2T56Y2/d
tqNtnQJI11mAEdYvX84hD5sPF/kGBYmDmewPC/kxN0zJQ3NQAGmsXCD8kiCPKXB+U7DBYdHMLcZg
/ML46T+Eo9iErh0ktZ3odemFK26OIgXL9VQZxJe7RMDT/dluNDJ027VkD450hNpxFX46ikso+vXN
HUTQmDtvbPrOhNPOdNU7hVrNITkZyBsdUe//FuISgpROxc5mmmnSl2ndNS+jdQafJAspwIUSuN9p
oh9diWeP4P2N6DG+peTHFW5iBbMOHvmtcn7NsxDFrj3dUjF/iFoJ+rqz3itv3ans8V9Ao2qpsdew
6YOc6+0IGM4J0OZwh443cNervsvK31K4CpAvCrR66oLYuTL3tQUcn4SiDLWZnOLKWD8+noVt/0ud
ORKSyGdUzIii9sHfX4J1nmRDKB/UaytN9FtQf8qkjUtFHzUw05lidYsqeo5Wh/s5W/f3AK5WVP9T
XN6uTtvL10PDNIidLzbms1ozA4z4B7w6kcKVkbvPXbm9UOh87NMHPV5td9k2pN7bGIhAyI5WVAet
nsxcbdjh9R7828o+ZSnLkRC1Y50N6RbiEvCoY2tYUGDpzw+DkZ9t8XYIrOH1lgI5q6dsSkWc5IrW
nDkJerW/ETTppkzgSswWr/EZo+6G4YF5nmkbPgnIbmx2p6yupZe6NopiFxe0LSsZ8799n/bQU+QH
WNKhWGECvIWg2oU7vNYz6TsQKhVzFzk3Uvo934RmCiLBKzaleIEGinYhxRi2A2N+OnUe4fvae6Op
h9TJSvz5eIa/TuVLbP0zoRiclCdcoVglmAGnIZ92xRhqB39Gf/KLbRaMBNZE+cdQtxAAxE7gDeKE
RMoo1m2RGLuOwUia1xqoRBPHvGJIhi3VpwdQRJYayLNxim0pthofKlKav+eWa98kKe3qQEfgnOcG
pAuQzf+a18WHpsvig9maW36J6l01fjtyMnfebkYcaiJNyDSt7S33s6prtmaKTDXwIzh7iQrEdSgk
wOzdocTaX16Xhp79uROUE4FEYaLaezTtjec09pNBDboHVREN2b+Qf44hmPc6pcvwa27gCxmhrkCG
R/R01wI0Xvnyci+2rGUfWWSyWjYpczzZcDrLKCZlIia+8nMPE5IjEV2MnWTVGT6dVWi4gO7tNhg7
qUBwtA2XrZAoFBMajocT8YDMkxMifyZrRNJubFaMLmldsyVyKoUyquigB7RsrVA8fTQlEiPrBG6y
mBrzL9yGL6ZC4l/CSo9o02Wzq29b8IGqIzn6pH1R8qFRCRcM42l/pfIb+tTb+ZuUq8gkuDyxWvs/
+O/Up7enpu1EjmRfhpE/y7vCwOkX7IuNplhEQ8SEM/LquiG1dzTpCl+6v6mN6A39w7SdME4S4U+U
Gg81gWA39f7O2fnxGKVxe8x4qJsM+wkKKTN+fmc+0EBwsuTgoQQLoCrG0Yu2SV/JE4iTp13WZqmu
nIdoaQ9Qkj/Dtu91bNpn/GWTf7cWKl/dp+IhLcjwh7RX1bPlZG8068OKMVKA6i28qWEm65sdbQcM
jdd0KtfOz0MtdhW0B8J98q3RkrAr/Mgen8o02VE3cf8H22kllOZbcErHymK7VRv8WakE/znQxoVw
/k2ZnvxUf2lpcb6KU9Svu6Ghr0DmLl+YSsTKuqyTl+cTH/MK760mn/Q8XGTFeZZhfiPqEV0J3xOd
+nRZyYx/wpjlr80JrtBnjD56NOJCnv87kdCOYwRsKB5wM5OIxrDimqgfzvHNY3FHK1PsMsvt4Hut
m5JvSJubfrtEZMILyu8ZOn+jtuWLsmNr2prd/zM+SKT9RinstTL+OWwir8b5BEFuNyIKkJhchZgm
RbdJGJATJ5ymVEy15HciiMeElueD74N41YL5UZGOjvBezxdi8gRQWZZteFMDQwt2lsZFj2HA2cUX
nZ7U+jXxcYli0du8sLQSOkheR97mFKNqo+vo6ogpawRcHfkmaEd4xhBvjyLCF0BhQ2/jvbr8QCcH
yCUx15BrhAu0iyKoXRPHvALhC+DeoG5GuE25v3YvEf3I9Z9hIduXOQlW/FWq7zGBiCAkoGvpfIme
IIrQ3KGWbw9oTA2Avix8uMau4pdd+aSiFwZZOetVVvc65ktq0caxEOa8ZFNcU9Ri/SAGhbCrhzOm
i9o7XyYB01A2x1nF3zDEpqZz6aaC4BtZzYZEKyAMHNBU4qWOmQIppIJgDibiNHpRAcQKKuNszLef
3gVghEmmrpmiHKn9R6Flp73fBjxuLVAmglBttn+LYZfeQWMTdXo1P/T5AbEdoD5YD8wDXPFmv7nb
DJetAS5gRvxtXJXRr0OKeJ4nOcBirn+bfaq12m4XYRwlk0TjiRwaKDMFYYj70g9TymWDcjJ0YSsG
dtj4liyDvoTZ2HNNn7s8RYXLlyfOmtRZ3vhYh91VwLNS7tuFuavFyQeBDiTwsDemMThjBraur0CS
9/nb56teT/t2L5HDb8dz1w9QT1scMPwFBA+dbrgR5DWURmZps5SvWG9/5m/kp3l8d6qRijABsMOs
PthO2BWmFJpt89wPvMwuAK1f0ixOR4YOyTkaO1a5Cbg/vqJg91ZC+eLSQyVUUk3YabzyU4eqA48Q
DvBq6xlhKCJ4YfZgC7aEy6EwCFYh+1HYHJTgi/RspQearS0RilXh52y8IAVhEHKnLXuYbd/PklzF
jlljZNEJzzVdElkDbilqxrKMcx9WGssOPRz5NvUMjZ858moBRJkh+HJaPa/BrC5ZRGtzK9iPNN6P
5cOtsWmi9P9OrFaJFWfJ+J8/kQQ5XP3iziboYXCaDLOKL1Mmu+NcSB+sE3hWOiaUs2p433j1LXDT
tWsJAhAdsxEvmNAlWqPfKPM55EbgsFhJnMJuxng3NZoqmC3/FoYOD1poTuU8I7ehAHLgteUaOCOO
azWHfCnOErJ9fNuL4LBJefUHnSWmj19Qk+4qGRnkNODWwSHOgZ/p5KPVmFWDyrHFs+cfO+iDVwny
ThL60ynxYhwesVYljGnUL/wgmwkS+xEwN1xlrj8JhMgadLojYARWr9KlRmMioOpWeYzfin3QsBdQ
KuGCTqUu8QKoyfEnDsZdXwM7DqQoZ1w7u5CBeA2+xtyY1Fh1p4nrw78+quJSCOVyui7LAu6V8+ir
jaZFw0yYA8fGYcMlm0IBSBaZrF/8JZQ+MlCEZYv3tGAnoX6091Rend/qIsn5Z3oSXN4W264OVHE9
eqAAAeGcECJl93wK1Nakw7ZHtvNtrlsivWcHIzVLXPj6fqNgpmXV2PgNqbyYu5VP6Y/RZPConvyl
fXYDwndnQbMrdTGwctuZHiNp9sM9ywTvd+4PTRiwocWa5wF8lfboxq+SoP3hfXkF9xjtmZXdKqOv
xbBv2JEdF0QXRW4VFih0d/PYAdlJmh4/kIXVn/CgcJ/mQiqHehoYdOLldmFZxNvrH/Pe4EPu2New
67Vc6vsD3ZOTd3cIHZToaaOXnGiAjkRn8zJrIBQBDXim6a6QfXccTJMz1ndXhoO1e4wANoxqRwfi
IL5NfyIsDrC/skoIIEUGNveCOPf1vT8H0RuxPcaEe1hhkrUfqEFANxqDWGr1MWzCXclE9D/LT1rG
q9DT2DVvQPMJmi1ix/8BMs+qtCnJ+bqAtuuGaZnu3sneOf7AFrWHCDG04MtJ3B72eKh1BrjxgDN0
UY5PciBxEFf7ECV2ZFlsJbMruE9HG6GX0jmPJsx7dbSx6w3VISTwvd3ojOpeMmwE4F7gskzn7xrZ
hCM3TIG5M6YY+u15OLrAt3hK89hDfUJrvq76oxYLqQIfgvKd382eCNz/Zr6400/dVsxTAuTrfnFo
CNzE3POjMeM3UQoB5tdoPXVq5wPS/8hqScxbgrGLeJsUqlvDDh0amf+YlG9V6bW38MG5E/sRs5pA
XAakPGoQu6qZ6ftci5cNvztfzZ8IZYdp2TU1D6ukD2F2/6sdA1fAxzZ97wBSsxRbSTiTMfxL/OMO
i8TSHR4SRUgObXCYZ2/N3bpfXf4rptvEUD5DOBjFzCZqB1ZaPO+OHjHjtVyKn6YGb5ykt6lbRGEC
nyfMr+LPqgInDWYdI87bPuvsKozIV2py9yhkbUygObe5g63GV4Dz7QzQkeyw/f70CCGcTxlBtJiS
FQWBMFzWEnBLubAM6YMI8jwJOtMZkym8Hq2HC/L5rz2/zQ8e9uXwjKhXkaGhe6I5SeApBbLpJjm0
F4tbD170/ElqsxEKbb5wqrvfZEKudgiz9srPAsI81ohJn6gdQLrRg9Nowhj61XxXQTvb6f45mZLx
pBROjQiNXLcgI4jUw04QXXiliTZ7O1/AhjOIG0P2ulDylQmYpCMh0m+H0sw0rdzSn9hkt8P7PL+S
h0gAMA5z8vMBJ8cBR9GC0FALuJI/TAJK6IKCwmdNo7xPvqMBjtDnRA0+rzBoM/StZBEWAI4Yc1Yj
Br8d4c8MDWt6NlE4fIeExwW7vNCrXeIBzPRHEfBAD0NvEsh2uVDrgAKE4PNYa/8W2Vn2C2UxSnCd
6xl9WAEmPPE/5vocnCkBqIrA0lbCpNygofJKoUxKEIFGAuIEsQrOnlSQ3cy9Nw+6RgGrBPDnZXvY
+ZBT77drlAil2BilDpcfrch/Vj2LNqJz/qesMNREamQ6vHTgMdDaiwgQEgfXWzSLl9LS5kZQ8SaD
+8BywHZ68HT7ynbZkK2tv/ArZKV73+QRFZiXUUngUH4iihQaRIzCYApotEriDFEt1wtJSn52pO4l
d8eJlXFVWsUFga5AGowXmLY7H1mNzNvpGXGQFwXLcR/dlXQY9xbEMBfqlKzej/ISYDPfR12FVdYw
KxT7uPsOP9w6PpGbvX7oOrnoB5SCEqZ7Sg3aSn1ad+wyCb+ABeVXCy8B48Zxkftu2rlYNfMCa5S0
FTu+rmIgy1w1y7panJSWcWJMZS1Ex9VyJDLbVyR0q1/6A6J4iUGHq6JJlqfT2LbHDeLnOhCN1Sow
JD59eEs+4hx7zF4tMu1ss0FHF5cxRmR0UKfiAKv2ZKJLAqgnE1W7Efcp+TY/v7EGz5uT77JnIT7c
DcUxGIqdLzlT7EEIGrCSRV9ByBcklkR3TIc8DHdAPwDLiYbRwy2kwW+6DjDjT8L/crtQ10AhZr9C
5SkHDsMkZ/AeK6t1HWEXSsfSFvy2NAIYoZxgix+SlBeypmuC9U3acvW7EvnOFQxw2K6cIbpf/lxy
u3Dnyb4NBACMh+oYnByRV5cSzic4rIHhxwI38NJfNdfS8BRwKOtsCi49y/X3r/REIFja4jMQhP7z
S3EH9nwx+0O/2xggPH9gfSltun0i76aXM6fDorcm+uo8CnXsElHLOD0dCRi6At+jY4ddOxVFiQr3
TPcx8oCLE8w+5X3/EcuC6j5msaB0ak8pQg2h7hxVqZYH4FRSd+q2KcFcTVio0FGGMV4EJeQP2teA
Td91rJ8Aj25rUUC/scaFVR3W+kxNRIrwJ2NWgfUqhzjxiLfel+7ZsKqeKTBb/F5LEb3E+mCEtC9z
7ReQdfmcoNsgQDJobOMV+X9ty6IWvym76LOqGXTx4FT/2n4c2hTL2opo6YJ3PH9PBtBNw0RsWGck
vzYs1fcO4Pdw5POdkUEQmvVpjTXc43XrQOVsZpXagiqkr74TuC9sW+NCCFFma7Se7qc7Hr3Ym22X
7D5nXAptRQBVxBdnHwLqnAZNwQ3bVz4py6UeGDx/FwJiSyE7LLuahJngfX49h7XHFx3vABGgu/ht
o4rgUGXir2VFxkKq31TWv2w6+4mUjeDbAJZMLmPm/sQfFWkkczZ5m1w6Z+24Dwm1yEqt7n77iLj3
3MfUGGiozcNJY5nSTtmXpSyUknO3QSeuyZKQvAfDTMwjW2pcxkkYvru0aK85zPfFDz7T19pqBUKf
LkmTW8Ra+AmNAKeU2A9hYQOouLLhcn6+f8/vmV/dnBnii6DI4dc9jCiRQSu4PHrEjCsUncSeGDzm
fmFhRGpuKj6qHkp9vWA3OAnd7URM5+bo6rCw/FE5ORN9dHMLfKezncJFMjE80Pd2ztZo/ZxdhTXJ
zXUcerM24/Q6qipuG3xvHZgF5TXYgc1bfNLKke3guKHL0g/gqSBlVQmwjyWj+mCJL+w2tEuh4HP+
NzkRmQs5ZRqTdgrlnC0XCfvxuls7SzAs132PsrH2QMVENyUF+DfX5P4IPWaLeR3z9v/tDcefTnT6
rVmM0RPU5pmxXmH9mJzn7WBPW0IydJJW9y040fUmWDeQmBR/2hk/S3Dxm0Fw0fCAvRjQIW5ppjPG
ZUKbD9l6zbkhlrCGp0a92vof6QulX48AQofQtrob7QOP4lDV519ITMi035ZUiyVUfaM42fj1tZEX
sKQ5or4M9rKIVGkdJQUQhdN0TTIkJsaX9Nm1avnxjD7np8Wbhd1V3+AYL+uX2M1f5Ls0R4aOGK3L
3o+L37qJ1QCzF0mG1m8CIVX1JSiO/luLGiSsGwJg6Ck8dWLWRFZh1QGU/lfI8MrbTuEaJaQ7dxIv
dpLkoZQGkbI+qCClqbla/yZVU8ZkuiW9N7pm/Is89zrGkes7qHIrwxfH+m7S7YTE6PwsXZ/sZa2N
GjdpJ/fVZZiFB54ECZa+0j8CbmTknmHtnTH6vf8CYaIuk+CP13LKc8Y7WNfNrgcnJVsVhxaW9zQD
l3vUUnBcTz1aQ3MrRKv18+i5PcsfsnYAEPHjkGlxs1wUAowDuuwdii7XR6xYaqul+jb7KEx/id53
Gj7udN6fyZemDQ+AeimIkyMzmV2gfYahNnUDK17ZfdHOtTQwhl9RJB3tCSJ3VfEMYjniJL9kqcx+
8DRmhweTAv6JcGS3WZ46+4DdU4gK6BK/Br9DoOlGEgrlroUpvDdbZFvI7s42rTLQO30zJ6TO3YcB
qP84YyxEjFriFNSZeL9HN9C6+VaPgZvsbM7MZCwh5QtwMY8qKR7t8KgS1pTs2I9P/EqCe1KdqIZP
IDRlA0DGvMcQ4JlYqj9jaVS2AJZSNRep6bCX5HcuIDo/Yvu7Jkjl1BsxlO3gSsmR9gPogN6JB8cx
G9iZAW2TfL8Tlqg/L5uTEGlxVKf1OQ+Frng9nNnHyjeDiGZbBgy45+6pifOTItQ3i99CYlLOKkiG
f0G+nt3fSqbMtTWPlJS4JWaM//GYy1acv0YQjpdUY5bn+5a3FQJVQn+QugzRHYYp4xykPXuejSiK
MQOmW0jVApX3j+g/mv3hHjls1cuvH8Ft67Rw7VJxPmj14InpWaFtk+XWo+pq19PbWv4kHGJ3eVZt
VOaD37mEBrF0ClXvTj0xLqfMPEinw7x/ts0yzM+oZ1RFcPabl1iQG1CoDtjROtioq5XZcaLI0fKa
CFnh72VyXgSzzT8VYFCf3ZXskpPH6CITMhOJLHiMfH41ydVJas0Nb+gJ2ro2B8EQvmIEvM96JGKJ
VHRv8mBeRks3c3bk4nvliUoOKVrxyNIvTsJjPFTaPfMPge27pBMlhMZbKh/iSeGiA8J9QiS4qTfz
/gAruQcBFE8HSpbmxlZ+labQbSFhrxS83ODO5MhOYP1rTo7va6Wo29tzXquhO1k1os49rsW82KO9
+2b/eeI3VCM8J3oK8B8EplqT9lVX6v7TJiC+qdNTWRJVZ4TS5UGfmyBIpv8hjLZ3hZ9rKIjyRszt
3KvNckfw0fzpY8O4y6wWjhGhp5WqZjn1Lngkha0DStaESNOgGaosiPH9bwmUOW2ygR5OgdGEhwRE
2FWAH7tGJiTViLB2xenmSasSyVVFeS4GbJh98xr96Mww+oqUt6VKTmryk1YpWrnNs8ual9HIQMx9
5h569hFUuez+eynH4hZi2QaGmiUabX6kDo9p+XRiyt4Byxs0OEJsIJRyx0M7qcym/RNSvPDY+/ap
lC5Fd87FqqtOmA79UV0yNgf8WjuqwTTCbGpk/kIk/Fe88kUENwxiBIt5EfkHw1UQyS+ZWW4AzOMI
Wz9XhIa8cmW8G2KrpFVQWlwKBgUrmkmYYRmbTWZLxZ4vftAxJyJriX5Rga7EfJE6xLfpZ7udDaRj
mjdtEwlfAaXW6dahkUZpL//MeZwuMncEQN2HQKDogeM2/BvHGag65sHeq+LVReol3FSO0HZVGmNf
kCVR24/RaPXG7dZac2s4HVvIIq4j6A44ZP6wawwFSJGzoCkK5H4Bg43FoR9pLYNGaNUwncsjwCvA
y3XYH2JI/u6y7CHm7J3rrVIgB1Ol2v7No03W0kUNubo7aJ9l87DrNqonIWyz2b3ePmsvG8NOeE+9
xlxtFssg7I96pivhu/Enm88vCoSE/vPv++VuQgzntt7Di2/+1TufeE+y8RXY3Dcm0vgtonYotRGX
pB7D/xBOPkaHJs5PCM7Q8g8N860YVybnQHdf6gAe/jrVvdImrfX2hwZ+F2Tx3JMsYFwg9D7Sk641
xO1A5CnTMGNOxGpUT1vKzPhQA7IchGWsjvrClwJD9BdTqhN/4+8+AJq11ei3l/ryflISRD9+TfLV
QSOPYj1D3amxNVuQhyjOlCnRfHTDnd3p/p99e7wjivbnE82L4QBAKgW03q05YDkRH5GgrRwOI918
NYO5U3NQLa0nuQEQUtNrgD+jkB9jzsEXpZXMGA3KiGkHM4zXYtBq8p9wRGYv2RkrZcim1EqVgFYC
cV51u11YHmuRl/9LlvtYyO9PupexdFZmaa81mVzXqi4lo6FxJ0zQgy2pSTCdo4DxgmAszQ0dTDXe
SSfFdJwoQUTJymBn9/3ueh1QkwUs0/LcysRctyMOT9QCM1TpzlpWbp7FveeoeOMx3P2fczBnavGh
nI0qI34LtW4NqMln98mrD/xxG8bc47WfvuC5SVpoXLeIs0AQwwU9n6Ho9kZ2b2CIcPBJQ452D6PR
TN18RKLQLrCW07f1aqn4C9fsVUCkPwtIUPELQde35IwBlZZA6oD+XQDZ+hx+6uExe7z61SnI5Hp0
e98q71dDytXgIr21B3kQMBsAxK9p7GovxFMoeBinlo9p92F1iNFI/Uyx5alwM37po94j3MFy/46l
lcUCR1pqFVDFvjEuBpXrN4nBB9L7eNGw7ZV27AQ2GNyT6H7Q0XfC6xR+dElDFtBgu5iHZbW3fyHn
Mjxa8esuW56RIKJtKh2P8HPJi2LGw7xQfbQnSPVvTeAk6/6+JydnIyHX0pWV2SuE19WIfOZd/J5U
uxpvVM79z94AAMa8Su2WiJj1HJHGAGsa/60164Is+/WfxnuhUMMTFZrKmC8flcEcJ3bRwyCJu5ab
/Ve7R1tMiWffLCMmwAZsxMXYozOP4g+tKThGJFEsS/yg7gnCX7PnHb78f4AO/h4mU+yZe7UhXgvS
zK/dphdAgnDIab2N33/0hiCTGe4Jb36tDcraS8VJ7UdkaEXThpVS6f6GavvWP737sGZwSt8BVi4w
4Krn5sWq1ukXDZQpyUL98M0HgfMF8l6xgbEECHVry9SM6AQ/9jRJyt/ET1HB6ndn4ZQj1ZuME4TI
V7q7Ibb8jQCvwNIKmF6jNUx46WMdaYTz44zXoUhiJwq40qn2JCTJpV+FTd0PgYqJ6H6YugXTu2iI
kJrxKziy8kg0r+eR5oQWdEMxzLx7U4XbxxZUYLJDADy4rm3m5Tq0NJA0KhZqwH/2ZgABemH2GcOO
uLtnMFNoY7Ks4/wZphTVawhL2piru+lfUXB/p4oMkHlYDkFt4RsyhZlBOrXxrre8Hw3rfdaHCDNd
79++1EiaAAR+Rew/1eqpDLw1Enaf7F+tMjc9AL70OTe5KYOntmJA3IZWmu6FsgwItLS3ZOXUcm9P
2qYdQ/ROCFwtcbx5/elIOp+5/zwzwVUiUsFuxMidQw3I00BSsycUomV9PY4pCAvUhl7FymiHaiZy
uXfFll16u41GlnOPji1a50QSFh6UcdR2Y5DuP7/bbV20QRSkw9Puswv/EriBd4ku3x2qrACRxX7z
w28gDY6qqcKxQmwDdIX0soA56zsIzDIyYFC9uUilq1eTSgSNIq4dzUPs7706hPVnZRFwX8hqkDn6
bxRFPpcBsXQH7ZUvS7JAatUWMZ5+kKpPyOO+LR0cg1vHl5myzPbW14Z8OAdI88qPa03B0/nrQVYj
f65QYvxLbANwJbtuGg02d0gntfOUV2HR3eiSdN4Jji5RStigKHnpRCA8dY7XMTvOYii6XQPMkqA2
bW2Ty0AxPSB7+49vreeMZz1aSyLcp71iqPvpnBRanwFSFCAEE7MU+Fs+UilumjHuPAQ/gP8RMxDD
sf8GGpHu/w2PwH244g/bvyJ2ihAuz/stCpAbtZh2YK7UN3HIWRqJzhVpyMBhdzs+/+yF4oAPmj1B
dXrJlvNsyw/oyJHBnFwJM39AeYuuDAXxavGjQGJe/dns4UMLhJZp+iDX1CPo6+MFyedAbCZXaOKi
6a6UwfhtdajqdtfgeHVQ1Bjkw5QAohPIxUHjk5B9hrsHkxvpt0EtmiaMhH/aqs1373F0cEIO4Auo
Y56wMOnSYJfOC14LpzuqlAmQB1tXjRVCmSBQ2ORAqgu5sxy/X+VDNyDXgXzDe6mDWL9Lg+r61EXX
54UAWmIqrDxf1BE3r9GH5UfKAD+C1Yx1gsaryBrf27NG6mM6IVBn2L7cLe/n4iaME2fHbTo+HGir
sWGRPeQTqeae7i8jt365KACguP5TcWS52TLUCAyKYZ0IBaOHGCUrjB6xzSz5p5sIO0jv7kwuGPHV
DZ0EbWJXtzdWuHbTOkFjh2+NA7tpdCpqqNI5CblzZFYl5IBcEbUMH6u1bbZ+ASK8odps7XChriXK
fLUODf1P4BEzkQ4cBrgtMzCGrOyTjVmveWJtY/lfAnWUC3J+P/bskwXQKIvwDKdSrHITLsMKKIX6
F/AsUZ8syso2v2jkL60tDkmQpgJ0oP9lLfNCR5QdnMDfjhP24jfwXHe414P0gHfN9tDBPD4YoRjK
aRi5a2cdK5Q2Ot10csHRs/Qyb6oOWt5CZFTuj6YubblocbiIAvuh1GqI4L2bmlZk29uUDA7nsVHC
5BVDnWwG2fUG9HyC3f4nXI7P3cXS6jKXVQK47Nl7vVLKtAklNwKw3QmJnt7ZfRT7WZfwH4Ha+sdI
TsWu9hbUjQ/e5zha7qEL7205Kxb7hmWGGZfvQzKq7XiLJybTiQ/wtyN79XmsiHnaAwXizxNlEmFM
fiEmocg8C3Vrfto6gjwCeiIyc4X1SBpCSgsJ4gf61bFNqA0AWvceWoFcBkmXuNWX03xVAwK7CsRw
6cT01Pf8tSlitZ+gT/kaTSPdrC3qwkAFdA+H5sy5W5lLkaybYsMtPvfOCKuOTGlEXKKNrEutwV/I
YceY+gnld9JUBMHZgMMRbQza2UCikHLswti5EkYPY0rgExrCK3Tk7AKnkXG/wRMURoy2pDd1aTzf
Qm3cYrEbwLxeRtbQuk0kTqiZmCOSt0l73hJ3MXKy+RACQt8OgSH6bblRQ/KUi1KTBih0uneR5UBn
sSVjySD4wx7D3sVstyDAg12ZN1x3SlIFlwcEfcqEDnw88InzJSFXQ+icxC78A73zuDsR8UogYQHv
x9z7t9rxVbHGsKLRvuks9m46r2b/U7aVb6K+XgL4m9zv8jMpfZkmxQWfj8p5fUO0aUFivnn3FJbU
tPsWF8BYieFgVlpo54IsKiEY41eBjjBc1cQMLdr3UZEIPLS9grBCbyjHK/IYwbPybQDC7dvQtLK4
D9veWNAxCRYXsIS4Wi7EPul4oOrpq7SRRH9NIgbciXCUJ6VuyqUVkcjpmWPN/qzOPu0f6QvvLbbb
iU9lLM6Ma5zbzhaEUwLdh/dRmTH5s6MMBfEm25NyO7tU9mPsKbJXPPMKedntda5P6issl0uFEbBw
uvvTwg5kBnz7TjF3ELiewfM1Y5OyqGXV2k0kGxbgTN82d8nOnDZ89bfWW2+hlJstC2Fn2TEwYJhL
DLjKHpGwF/SZT+CUivKBIKd4QkDxmmM2NUHS89QJBP5a8I/GcuSetNeUu73lrvudBoybxt/Yq1K7
/iP2XZMnnbX5MC1R23PH418vG5CrDEVYZHkvuUQsrGSi5KXQKhTdO4lf774zRmrikjXfeM6n4Q7Q
F1JcohQ5pzPE/IUWw4mpBvEWhJp9WW6qcsmxOgzY2hFmdqR1BSFk2bfZ9I9L6Ba1yxLr+/JQjNQV
E89HW2fON2KTq5uUr0PdEoD8/msu/tQtBswcZ2ux6f8PqGYHASysTZNqgujb9oDG1ph8vlGRoZme
xFnCrtAfo8ExPo43EhfO7sgN/xwt8/cuiccoYC/XPH37zX6HL0fmaDo3vygyPcpLHaLEpDegkW5o
6+kJP1QNAtcggc8P5pwqyb+EmkLvd4vlKro0IaiJsh2pBzdF2fyhRytKc+pPdUU3wg2eyZOQ5K2r
28R9JX2SK9CF9wzzG3UUnFqfKjFN4I9oH22tXlsobs7uEAnaQaSnWLe2sphglZWnFwwLoKYK7123
X/2JihuTWJJjKNgqdYFTNlgf8+2BOtuyhHR0NCz/F2rLCWGZuf8rrc0rDPELqcMISUapBchxe2Wc
Q04IKrSkSOMp1eiY8aJM7kI4f2tltDXnNs9fp17Ux3CIXWMFIHZkvQkWv/6vHv1aPYB53TTg1URZ
pwlacsSpmKWLopAccUjVJAYl7W96S9yfS3GDMv2xcIEWPKKuB/Jv0H7QpEZWaBb3N36tHfoWQLNt
kDPrlQI3X+wVFiikf8l9zHOhMEBB30v8rjdt2UqXcCXZKP1DHL/OaW8fxZJ6ZP8dwNZ61pB98KUW
+LYlW1SelkdksFdad97/mhkHPZC8mFXOWpqc8urOPFRfsYzbkTri+bFeAN/a9sA1dAhfw5NG0gTJ
18qLa/UrAdaKY1jKKSFDC4cI5HgHjGvtuEICZ/lv86Eq1AjeCgLhrm0uvzCqZbSNsN0fh+nrnbYj
k3VUbVIxWXqzNZhr3gI14g1Xp8RyUJboWqx/wQ4dqZ5EVWh77ab36JTv1KOX2j23UpojxJUdM7aN
F7fLUTClEq8Pp6S/+uy9d9V0QBedvn+CnwFqzXHmgyWwiPkVBw4IL2z9TXhoRnlHBt4OvMMiQBR8
w4GVRWJSagj0DFg0JGSq+8edrVzjmMJACl4v7QcqG3CXshrjfzlgdmmfeypx1vZDaeU01KAN4WRq
wZxQid2/B65YQ/7gT1E4Rk4PbuD3k++jHHhckuAVmu/uCwYK3FGzyWXqg7v2nfKBxxseR79Iq/Cb
PhoxBWINAtzOBfcne6tPmL6JiZ0zuX2e4eHuFyQdN1KdoGdB7bVUw2Z3dvgGGlhLod6atWFu7obN
tuccOP3myTTSVaAgVhJbCFveA60E9pYX5Iqrx/PVyevKNLpyXfgnmr60OOp5grrsQSz7fURoi0jq
JLOLrC0/dxccJZGpIt1iKoefaBxZ/Us2altQ7HEBvXHx64IpwdG5j00Vi2ind4/p6F5Rd58hr06B
MPW6KwxvXqjsVbo+Sgstr6ffHBNF4RSGkUjLhb6BKHdAU4R3RtMjpAZ0h4s8OtVrbD6uRgbm8HNK
Fl+AkO/d5dm1GWE1fSt6CkGvEw8jXqUS5c12EVxfdlmRw64hMiehyauRliH1ov2j/5Pdj3C1Lkx+
LAngQVMY7H8yeVQG34dYkySUuAqbR5eXFv1Kddsp0l2lTpWU2PN4GGezL5wFBO8eoqA2yFoE0Try
T/ypTtrRrG9dBzm1qOpVLdwRNBa4oJiu+F+MMCXApgO7fGo6aw/tT1fOI5nMxhYojlHClqeg2QgB
+S4ljDhZWbM1ZY0CzIWakEdCw9stTYdCCqM6UqyDBBgQ3vKqkISUFNlkc8V8A/ALo1nAtFNSBA3p
A8gV4NDcgZSedyGbEo2M6yKtLeZO68W/+8nPHvtRURBrBBe2k9mXVWa8n3x1U7KKOJ6+ARz9J8Pw
A8EWztwSBeI1hqBy6I4X0KxrGpJJZgmF8/FvioLEoF3lHEoMQV+sJWCJWwnpJW8RK91W4R21UIip
l3znSuygAOBlxymvfxYLSgc/zajBK/Ok5gHnyQD4Msx8ts2CULC0DviE8zi0Zmnt4y1GM9EAQlpe
WQz7VU+qU+G0NgneP+xhRpZuo2YbVt6l+/2+KwTpBYZN39ICDWCX5WMh7HUNQ1Dhy6iYAomGJYHj
jPCd/u9TmMt9sgdBLj6K8w699eXKTpBiiHrontJ8h88ozEgwFSlPl4WLQ69cjQvDnrtcCF47C6bA
SOmX7hgBZMLOngZy6uui0xZEXx1xA0j+kOJ33QOBk63+gBqE2C2Q8uveDXD5JU2af+JsZ/fEeOFs
mAjgo1ugtw3ILG4aXtMYss5g4CfnMJhOUMKs48EJttwIMfleoGFHbyFbmn5k7u8KxzQBBouSenMg
2N/096KPzTy9FgZwxE11kwSewrVH1wUnZiBOayUuJ9IQocmUyoLjE4j1Vo49FbAjq1IrcQ4ptGhf
32mVoNGWG/uBlNZOCYabITdXoXDX/N/LfE7nMUDrBT/o0TEpvv/IfMS7x06dHkHsPGNgh04J1sCt
y8m+7gS8g2Sop1JSg2EtZ4Q+2G1Ug8BA+22hjyralAASdSuGO9iQuInyV9eVEzrGxRJah8dsPNlf
fY9EWR3L/s/jYILGc4JBmHEYljCa6jNYVLfEvEXCSyqFJhJ0ISnRPpC2cM6QIIFKZLDBWyYOoSDP
ErTN+52YHoGAqTAGL6XfspL/Qcc1laSqxcqiUOR/e+PXpReLpoPVWzSHFdQjq4aLHTMgaVYgJBhJ
IXfVOXeiYV6EZOKoA+zZCdmHO42jrE9duuf179LzDdqZchbjjvZvGWgnjMb1o/FPLF1frzdrCz3q
DU6EFQIGcE27bTe+UlY3rp+hQKpYzr9qt6SSxgTVhBOw3s0Hz9Rb+N7QPZv+gpMH6uvqzCDjXVpH
FYtvS5vUloaItDHz26aAwth9NALS0057IuHJAFcaucnuKEm6WdQlUMwHtJlcuRVAgbxzyG4YrL9X
APo+GhdoCcpzUlwjdQW1avUL4TYr11ZvNVoh5IFaI9nT7eYbrm0jIEN+SOnCYZ3p3zcRuHX5R+FV
Trz9mx0opVvPndIniPj+96LQjc4ID9uyWT8k+zIx20If2xmWC55hYsCeo8TioLhjsy8HyCzgL+HV
t90BH/xGPI486gzMysv5qeEYbySAlyzlQ5VU512/Rm9IbWpgYs4IFZDD4mME1QmSKrSsE6M3OEpH
JoT/CWo/Qa7X351qzcoWs0sC7eJYKTJBoScwe2V03hjQCMi+To5CktKn0iGv4gO0Dpeq3CWHjXZq
39mb0TeERyJ0ToxBSjgnNM4W0jTTVA33B8SZLPNwCyIIRdwROjkFyS7qbpzS5b4Im9QVIPyFifrv
N8xUzEl+S317R5IqAmgWvW59eSw4i2tLyiw5O5JCUrMdEg4fbWHWGrmVVdhaH42WKMmSja+4vUzf
1VHvDAdvzDh+uN/1ZDWgPc/i8GzYoAoYzHKDjVRLMx8A7OKMG4ufD0cDNncibk3dUUafzIeYDxlA
7GrJekN3UnDmyxbnB3335hd6ZdI6/y2dnUhWZ2DIjlybg3KBFVsQeONpC7htdfifOK4jv+9zCsyT
DHHaDzbnsfrZfG1p12kfRDf1QQ5xCMcGfknA6pIm66hO3YZJM/fEL+ZKRy8yV5oVJDn2n9cptWP3
At7fWWKCsQwxNrlSw/wFU8mPnMX68OEU5DLf/ZV3DMc8lrk9x8wFjbQ9aRU7S+ZP4Nq5ReEjADkO
uF5dieCvV4q0rwkA6MNA8pHvTSQrUlyQ4/MTQfW7Rup9enY2KVMt5egKeMuEYAO6sxcycOMgx9CL
r2U0RtL/ySC3WsB97+ug8xQ1s2Z3XmTxx8qbN60npsWp4MGVPSRj30MbD1RYzpwwbz+P4MplpnrX
fj3DJR+z0icF+Ad0/T9T7LTnkvCy1UIpaE02Q9ABynEiU5aVRCKGQNeeEXARBH0w4lM3tl+Cd2Jo
FM1qYBSSztAaNPzusVfjG9RgozNJNckyCTWz/euoDFUism9OPtnLLphv1ZBft3Gp10skn/8zPEQM
F3KaIinG4wmll1CD6qfekZBcOMLNe4o96b0jUxGW51Is3fPYrTRYOBDHxWksA4xHYwfnpCz9zlse
J5D0wss1qnLx6OLBr66npYxFK7EwhitT/lIGiYWB8V51S/Hq1/9CpLZC487+cAZhiQuJwdqbek9I
2fehi3xPzyAh1Oy/YdZsvIOfctbHO/3+66p2EHdA5epiIQ7FwMhPyzkouM3zQQbOJw+XKZVRi28t
iv5VvVEDb/55Yxza5jG6rQfUDHppr+FqFKSYlTnKpDWbZrvOwHXBxrlwAc5XYdSrvXq8/kxuKVre
ZdzVXxkDpyL6kGyGDG4Y/DUwpimcrpB32qfiHh652T/cNcqp5yZ3PAGcDVASUy0yM971a6kGVX7c
0pNG71ueNEJOcDEEzXRK9SyTp0+CtUobZOexjAE0aLB/CUN2kuLtBV4XmY4z9nIVJajkm9RTupnL
5NVOiUZs86PcNwYYmeu6SfRY4lPbOp4QvmUbM8L+f1T1M2ZDb9PAU7JeU5wr5oYsBKq5cVIrBrwW
PLzuxYfWbLscnDnijhI5IaQ4JhvCx369qRxyUzEARRggorIKxe6V+12BMG5d3wawDTcOrD/deJ+t
CuZC2Zl6wtyroNYU2BZbzmZRjPX/IsxcgwCYJQoJHvDJtykuRKvN6Q5cUK9ln+F3ItuIHy8N7/EY
Ei81FEWMDCTaeMK+V/52Qij7qe9za9vNYJ/Rx6wGxceKjK1aXi4ve6xbA2aDyGP0ep0R+nrVw9iW
Kr8fL68liIrhZqCXVd1DzI9gBVDp8ZLEfi/NWjTx5noq6qS4NN4H+04fOuiGn45uDmczMWjobrGk
/VkIU/vsPqyexK9o7hiEiPwVg/7E1YzCTLXDW5cIpFyqVSqhDelgIvMhYeWcWAQ1fZAF7z9KWpGE
gSHBso9VQvfzLTArsuyKgxiT+XVjpp9rTxt9PspgDyhBgkoHaGXJYybG4BCbdrsMuTSa1Q8QulvW
b6A69Qgtezuyt1GfF3bkcT8UfCPmLpJgqWQRvnkN8DCOfGFXm0JBcUSqXFONHgEiK5mjBA1q/kIK
0FPhPmJAvhtJWPCUav7RWCcrrpWSVm5eZnUg9CY46Gaq+P4mvqFrTTr9qeIPh9U9jq+X3TCFF7ne
8rjZyv1j0ZMYBorBRLjeOWxs2FiiOZeKwA7eyeGad6XVBBgAkY2yrEryb1AhEhy8Dn4dvbgW2THR
bxVlTtFeu1HEZNf1X6hCzMW0oYUsVX/6MsSEuYH+QWUnBywtSLkSZgOBNCrtSJWJ5O8NJbIZj9TC
2QQD334VoLKqIwMBrdprPdjRj4VHbC260BO4SzViOxlh3XlRBoD/9cm902jJ+mul5vM5i1k9755w
Zwx9W/RrAS9rv9n9Zthwv0HLPJDTPGXIwNRNtdGLhiyfVlduWVaEqRIgrUrK/b/IZs32LHbTSIU8
ius7tFjH+D4F86J7eFBbHT1nhsamCKeSa8a3AU6v3SFNQ7vQUgK76tzwhbSzi9ZlxCmKqAA/SmXd
wIwSAkPlk2ZazeYDo8ydYmHMvw5/pxBzuSaEsDJXlx8SGdJYgfm5yPRQSfxetGXiNR5VTNQ89Wu2
MGbyHLUT5qJBCzrjEsLLboB5MlTrK31D6k+9DLdhlvc/8gvG0uZWeb538EEdui13yuwdw/BlNfsn
+SobZ0KqOLssWtZ5Oq7F4i3QnHj7TUKbuLMHcAV48mMCdV1/FYLbsKk3eZ07URhApHGpyJ9z/m4f
x32t1xa+dy0p7PXWTAC3hStP7kwpB538zRj5tGnrcg6arrXUnERSaath+pPzB/GkPhYKIprVsmp7
NGtTgQ0XduND5z2nryxlg0joIgOBztjhM2h0ObQtlNMMIaDOvnh/DMh/ggWV0nlo+Pp8AujyZ+0c
i0Ap8YjBWpb+32a5V7qwCpgSFN6pcEbuDDU2UTU/FZJlNGgBJhEb9cCXQCiCBn/beWbyBudiPneH
kYOfaBcn8LwlZM1c94dP8C7iSOLxIlq2ccHSHkfXGg91SHEV+BVP25BxrYVIDkv1eaBRBNJSaMa6
o1vIjnrMsuOF9JVTxB3o+MHimNl0+HP1w0T0MecngpyuU+rVFEtrKyMFE8CcHbAziSW7qqvy+zur
9MtngSQ6KBFSn3/6BT6des/2Ywtu6rV2LWgU2CCmK4w81edad7jGMlrdJdlU3wm2S5UKlyqpp0/E
/n8GbWCSaAaPw27323XYAerVwCqqSEGJ+LnohnhUzgEG+XjzUl4rokHIgSWnqpKLWUa1gBxs/PVS
pSUhSz21ge3eTLurR5AwJmlw2KTAGfc9COh8dBQd+4lr0MfYP40z6+Tefi2ywHB9i+Y6BxJKO+md
A71vm8gjMSV4ULeetwCz7tJi6HBEMSvSQ/x4SQHUtaFhJrOt0z78wWxxMhdiKrb9b+yFw+2HoC0d
L0QE9QHMky3b6RFKUE3X2gnPkFf5QfWoT8V7KQabIyqTMltfvl1QkTrYSGl7qXBIMacAx+iDTtHA
/92W+Mysfp4e3y/2/wamzy+4PNbW4iWRVj2SFyxJpY9dryJwmELR2qLZQTHN7DFFXvWfIiGAWCaI
61aghRR7PUHZ6+mISU+ND8D2T2vsgP28e6EblDh27dBfJW/bNuaJaXGBzYqb2qWPjhUPicTeaSnt
Oml4+0ZpJLEbGBy4ci/p38+PoH3sTG3u/cnJgxV3yEriYt/iGHOsRTFb2V2zbXBUsMc3aav29IoW
mSs8mTz6fIpPvOtdKPrX5f1896WzVESBqsCy9W5ij8DYq20ANMrPMC31Nke5Fuw+2rhnJRFqBNNA
WAtakDERB7tPho9AohWOYPpKjc/eHB7QIv/av0sDIGtWqAroPO7QEovpbDv8bPddmF0buaarVnCc
KPg/okcd0xGpToibFyC3TdO9n5Q/R6go31+l2zdBHTunHPPD5zf42ztQIsbGaayVFxHv+jcUFesb
36LSK9CEBkJ1O+ENSVBc0tf/dVHe5KOQRSKkpXxCXWAfgg4hk1Nk7QqU0JbqD8xYjcvOwXSGn6tq
F0VikG8Z3s7DcCVk9veqgP7jSB/cn9p368+3C4tE15gEPKFUyo6jF4CHaSgJSiXWHYhMTYucBScG
nJ2WTR3TbcdOyU6CqSbjFQDaMO0ZwHeT26nYsu4t89Ok5xDf704AUCAY/Zy3PHDOL7wmBvt8C6Jr
F61HoIyMUGdv/ZRwte81FbdGlTdyVIcu07+1Q98bipxhhh963bj0vj7kKfAKe2zfgcLWf0taz+SY
id3+FiB1ioqcJ9/JEEXylroUIY3mQZ2BpYu3an+kDlV9bZhWGJFCpxyLF5e9fOL4Q0VK9kflwBzx
d8u8GMZ+sBghtLmm07YiZn9TvlV5aZVtJbzb9lVFQrjSk0Zcsbw5Ro4wdq8026J241FJ3bRvhZLJ
wcgakkmM/WsXbrYjjX8ywk835xCMCr2jjgJfQOP8rBJ7B0KEUja2mAuAj0vNy3seIx2cY5XFscdw
U/B4HSeTLHdF+JcYs+cBWwkXQTpZxgQCEYYdrCXMOpIdHMVBAZwE4zHAx5FrwxizO9mKT2Ca0vEF
J/4e8nCqxow9H0f1CGOW0XfzFMnybMbgDEuBNNyFCrn6IdFqa8KdsAn18fHafuXTAXESzbBkl11A
OKUC6PA3p82a44nVTXfUYcKhWHUjK8dnVTBC9zEs5hvpITUVX3dExfOdfrxrRH9suQ8viQL9HHvk
VUsfWBEaYRYCigwH7jtey0CN2f4fh0iQjRpms2fWmF9AAIUvv3zdEFLu1VVkZjIaUcJSpT9C20Z5
H/XuBTWXs7Ks4y+cHCe7VfOuwkuES73uMRg4JbYxziKy6ARQWAuNgwKT96Bbr7ac1yj3r4Nb33g+
olhxonH18CXEbZin0ThWX8aheSe73dNFMwaQOABEX/6Gj0fBkf54n99t2a7iLknSqQk68UatBVsv
sAMYwmrGmZ8B2CtxcuQTxQWDfTYA4RtaUFG/Eeh4Hv5xYBqiZ2tdc+40OxgtOK8mSqNpHSiCWUti
Md1KrWHFQ/sj4vu76Zyv74KapKUVkHBwAO9omIH7spT9ANV+cocE/MkHULVDOlPBEhkgLEA4pggR
HzXTekHKmfOBkbFq2ZnlDJwkAwQciErjgsg5bZ/ZHg/p81MUZT902BVFxp7emAXkUZ2011U9JC+I
FXFA4QpjOfBElpqjpOEsjd9KTklyo45ikkSNNk5Fta9HkqVBEc06SSdOYL2t+wgok7HphMiJI2C8
Mj/FykM/y/7P5cfTzjRdUXBsJK04I/XeOShwHftm7zn1vvPA02pCqUet6lVtfwWOvf0x9O28Fi1C
sYwsNnrT8KrBTtOHO43HMQ+z2BMPmGn/k37abiHtQDcYspuAQgUR1krrWfOL32KvbSrCq8xN8Wya
yH2wt1Itf5cHf6IGwb4+EdxpoX5a2HqoxG2tef1moiZ6dnS6Izsv88ye7QYBSPEPpqeAiICKWWNO
zrRaTMTNO2Xbh1O9ajGlqy09U8G4etE2GGreu+71MO9u2vMd6w6AcelXEDJn+Nx7ShWQprZsxDsj
lFFIZnOOepsAu2tZxfzr35rWn4TpRT2JH9BlIXTinj3HPnPyN6oNMuOCiLQhJRXTB/FPlO+QBHWJ
NCEAI4s2cyiGJQpLlB5ATAnwr0CvdMFOwA+zeF0tMhX6P3PCHvKUwLugbJ/GPUTKufnoIwmvZdo4
o/NO+oEAO5vPCxiHxRHTrO69sN/xRtgpgmQCIM9rFzjxIdRh2YZh0OeKCOD7o9rupsGpMldigmuv
aXKNxgwnQvwoO+afxhRPrTEbs9NJ4Qz5/diwcquriHGAJn9T/pXlCtr2byt1o4aLd1z0mddlQ5rF
nam34d9oPefuEc9tOixmW//epZ6xRPHXI4H9XVXbnqVviMgQTmUt3FCtSLOiUh2DTNhN6KS1RrmJ
dZ0uoAGM7YwRySSMbdtbU4ZmM0mj7OFH+yOm0QodqPTGrsa4pP9uuBl5Kp2SKPgDTHYSTn0zCjgY
QTCSGyIbRYPYB17AusasC2hEkDrreFh9hZpWoZISJp6LJO9c2uLAfIXLQXyeiEwmRJORntBhKVIu
S3FvtTGLScCEk8d9/Ptm08wZX4yrJvFeGANlmpcywxU5xseYX26ekIuW7wATc0ebe9hzefgij0Z2
nYZAkLccf1Q4/SD1TvDT7htyPPmgDbdG5Hh2iHB5FyJdo0711VqmoZQKG5f+4NTDL3c3qAnvxZq3
Lub+hYoOhcXiIA9eSsM3tgdWJTN/fWYJ+FGPrQtsisPUMeE638UwybqBPhxHcB2AIjAr07uhCo2O
6VrEqV9MRmS3r9REFLv6QiiGfqJJQzNi7weLBKb91c532v25wnF3/Gh86qB79SG8r66w6IuUyVqv
mJ2nj9a7l0ZBys4D4VDZyAjXzXFiAdh/IbO0teBLAixejVXH1UwDB/Ue5QY6tBtIAO0HOlt1ElO9
w9RZMfuGMpfkaN2rkfb6khKBg/4/SDMNcAOP3OKKK5N1EzSBhWMyPcdYHxyCX9SjL929Uj/qFPCA
me9d7YGa/4FVI8dwKzZNdKziM/4g1rhxCu94k+Mo8vbWEqr7O0TgwLjdlLG2uygEo93ZsQbm7nNV
DtWT9UHcY5s3jX25zn4t36rjbPpF+acGcLLAzJ4UTHFWTrgm69NcQym5/AdPWTc6IMaXa7KByt3e
/fc/+NGwgYoblusqqiNR3h7qZ1kRwqm34L08z72cQXBDUe7soN0E4OJVwaACr0RaQtcTlLUBYo4x
g7YyjUjVP1HqC1eMEgdiDVdckehGPDK4VFFuf3I2aOLLXmf+Q8i9z9cK8C2uRyahbYx8t53802cA
IC0FIPvpZUevZCkdLvEQZx/8ADGnVDIcZ1MvuVXBFSeCWwFcZ4vAxZs8dfkFDEO9pScs+/HdjKlE
GaTw0mOep23fYI5zukV2AaAoDL/zfltlIez4+sd4ku/fXYg0foiHri5/oosU1o+6yuLm+/k/gdvZ
xdbErTy2fV+o0JXXLyOASNBJzRYoVkdYcElHGlAY/c+FN5U7HCo1lssSZJoBkueqQspP5fCtR/u7
qBLCda1oPK5HZkEqUIU72KkeB8P4N+feMoJ3lAm1z+VjwMvljFIEtJ5B/0iXILkpIg8SVwAb6JLY
TZvMtTjTYKJvN5jDa11pesXwmzfiUIyUwmWkAH6+cpMtEUBzZn5jPQbfserlnztid+A4Wf2Jm3ut
MgKlK+zdPvZC6TlQNYCqb/Wf2uhabUvLQ/Ris2I9g/i/R6oUWcM+ejl4T4vm4QmE9IHLIJ+lhC2V
KS352XNYG5rm7xF5JcUg6s1ZRzrOe8ln8TB7bFPfJ1ktOz8i71jhI6s71eMi1A+D/wCPltgnB0fj
t7s9JZ5ccdb+HibNl6oS3fdyxI+PN1EmEc1xL60xhaCel9h2xFh1Hj20IuXL1PJXjF5Qq22cVdGX
tJX2ZmG9pm5FlUIeV/L8pLzo54qaGw51i/8sRd14xHt9rvi88bCjxJlCgmfR2RsI6nK8zIftHo7r
2RPcAttlybSTHA3yppzF0lwcc9EAfJx0QozVJ+I8MoPPadk0XUnORdCYGdBj0Ew0awA6b0HypuU0
j+qbKRBnjV73Q+qjirgaJivbyuTLeLkdDCUfbiA329h65J82Sh/rO9FQBiIAITzeZOaCd2Epvgr5
ltRnMojjp5psAJaPchc8M5O0SXRSjunkaSFf6weO4yBRTPvjvr87hdi5izTFBUJfpIgbB4cHlN4b
h0a4LstX9nkmNM6FnsI5PU9XPxlee/9lx1yn2c1puGrfPNjy00c+CUVNR0GD1+vLzJW8tl5bpPYE
Awx50mGwcMx9jwGq9WIuKc3QcrC5tS0mN/7Kpg53s0FfJdE9Bjfbc7ljrrQhQbgLJ02/mG4guzJx
G1b1GvfNAeXYLqIoJTz7lYyh6aI6ZhEKzc4AdWTqEXdQlG6bHFvDP1tIjqDd6wVyYX6RHNYUEgCg
689DQO1iRxEb3hfKd/JIGUhGkNj8bSZOKHOmJ+hlnXc2G/dB+tEKe4h40QC2wIITxjFyhpPDwkkX
SN7j9oR9dfIFDuxyUmvSn2WBlSLXWQe1vCcEcPDbag+96xvr6FLR1V/0FbX4PteHyb3Z7ZXfzH+C
XRBp69zc8dIHOBOnY327d5W6c0s96o50b8/6ZJim1BG/QPiFENmpisjlDfyYOlS3ZecfBuY6hcxL
s+JdwloAcmnhwD7AohvBK0LmnQSOJ9rUAsS9Hx0BrQvTDpSekGaU3T4XhTRKK1rt2ARUGjvixrwR
lUqvuJaKdnUaltQTSv7koC+proKS5+nZB+rGTmpuHJOdtrR9FGld9DFKkRhRIfysnm5TaPMLfKKT
tTbsWA3JwPwEMhqJ+y813955Ywbh7GKBIJO8VWOmpHpif5TT7g+xsVqVr5PbOjz7eaM51nxPfH/I
z8M71vXPzKEeEVq1vkyqVWdd2//bISXa6bGMi6nSLEF9deck5gtN1gSgD4IC8ilAZSSsGuIwyS+p
iJz2/uNxv+qcCeb9JMIwwi4GblbqqkMJy66gJJYiL6Jx/WAraxX/w/SEi3eq3y3LNte1vugsMeet
g+X88oVSTOxMUWYGakNLyychaeWdYMwFILQEB50r4BeSLUvDPRvvjTb8+GDw+/VdSDNj/kS07p0u
ypQNT5Btr2i1thj0A7jhzZwGY8lQ1tjyX1UkD3dQYywZUGq/lxRSiODivSNZzumCGRnec7+X+QqU
DCCJHfaNzT/LO6BXmVRGCcoXE8m3847Txw+KabVphMy0Db+1bzKYsiRP0c92YrRAq2FUrBTw7SIr
7I5pdaAiX0kSMzhfxZozUPvvg2LB8zPYyYZzMQgJ56HJVTx6aqWDchsu5hckcXk/al4m1z5lH1E5
IiC0El0tAlwaIO7s+edCgeaGnYKvRIXtN3CNxLz6/FuwnC9CSG1JETVlVYoKr1nBUpl22WnXz3Tf
E5oSqzHOdObu1ishUhTTPp1DNwPqbf7u6cIdYL1xIN75LBWYMXSNWwzydjV9F99YsGhH/MEZP79f
HyyPrXfKmeOEA4bwlQUx0we+wqEX2vCiZsoeg7sYnuVG6RTORMoewZm4smmNAfzHxX/D5P56Bfaz
RkXGbaKRhfZN9rpywm4ENlXhZ5X/o/pNZnAPrlgFqEZ0BQn4teQ3UjTC89QVF0yGx8UtV6Hwml3L
9lMYZrwIvta7rcFfjWAMqTUm/0BTcGUlWZvnE4ZcK0lqkkOrnilbbiGMCVZjRxEIXOnDgCgPkJPO
T3VfUnXbPCwRzLAkOcp+5qqDRDvXKEF0f8fr5FHJh6ZNUwMsSPTwThflkFyseQHQueJKQV+n9ZDC
1JYl9w0E8coHt7bpU/gcIYf+Bou/01KPS6o8kxiPisZVS6XpZusp1ucHO4TEPRM97thBKqYanEPk
Ja4iyqvb7NlbLF4mPwm2cC2YnFiW7RwyQA/wH8TU/TSrdIAUDt7r6kgYc6gTeCXQaTLsfffd+Ls8
DHMMNfeGEUm/Q0JZq/V3gN4Hn6ryOXNkWhuKXBCQiZEJvaLn9DYDdL8qAkUZaFLnX2tqr84pxIS7
HUAP+tEHwH71SL+ZVIcvx1SRRmpbDF2OwHnqcU0sp4jy7y79OB1My6uSuI9t1ke9fSScRq8MPkWr
twk38tWiGSCNcBxmqIOLFhK38C2kEzrl1b8ljmmPcGts+HaU3jdmJimn0N+1v1OG+4RUsz8TIoPh
qwpIb2+nWX8cpBK9moVYequFGSldVQn9pAOpCy3XGHqn0Bc29JOGQLOmd3eY41y+IGSf4YKZo214
Ic8Ueo+l0e56hdzSZ1sQaKPBZSxlQUxsto2fKA8AZW0zJq7iKdRz2V9QjwAJCvBzOZ/JIaxOmXxf
k5NKImLZoDCOOUn7qVthD5PyTXCy1Y10Rc4x/eriTftBELw0ZG8/jft12UliTrDDMgz82GbVABgx
DllPN9uIBJCiQjV0LyxOEf8cWvhG9eH+S+6TgUNUJnFA8tN0Avb5+3QS4eWVbIk97iJ1afKuS7lz
HSKBTbOuN3hvr1nA3A+nBIOI3rLgTArsBqQBooMgYnI87CoqDiXihp2LP+5vNcOAoz032+anHsF9
Y8NnWnE8hYopo2fsp1QRupfFEzunG18LxurSxI05QvYQBTIRFyJb0KxX9Z8+19BMq29NU9Lv6rfS
YJzxhgWuUOYHqG5bPphZEE5oFPlkCVzi4r1ARkR7dN/6ZDiyeDusirBguRkwucaZlqZ5U6PJaMN0
J1V7Wy1/7BYzMlKaTsDK1PJ+Dz1BIFNeno8YbV4yTerSYXhmrvPEYKRx1OyRgxfUcHSbzTDoINio
lYdlndGkvHAIeTywLlEnGXXYJy8FHLQAAbC0lWqO/OSUSroLTaCGA23SD8fQTow3hYzWU7GuCwBp
X3kkRN7eN2AoYXNFd2HmSifZcmhOKfRU/qC6mKUw4ZrCyZzs+I8tnH0xEjJMD5TTYZel/+z1XOwT
EEWAcuyiYGDW3A+HneKt9smo2tPPPT3xbmq74YI7Fif+68vuIxSvB3PRSjseg9i21Nic1tpj/fR0
MZaV55J/P+88MEC6D/6ha066yHO+D2Dz7tHsP8CKDompePIU/qmPOVeKWQ52dOws1Wkd3D+lWAJT
CS2GX5pDWmdrz9DCE60GUYb5y6BOtZhZn68ezaZrESqwEIdE3yAnkYPlSN0OmVWw9anhA4N/wlCW
hp4OHHboMIQLQ/ekmHIF1QLBEdGt1JzjcmFhfW13lFx303APZKIuTNSyCg0P0+RY6LlZSfTeTXYh
+MtXsJaoSNT6fwDtaXCIYMZ1cHk1as8FkFStoUQ4tV16fioRm6JFb/Ns1BgmmXfxtNDWdOg1W1G3
/T3FUzESmr47YHciPVXU1s39lVambukngHKZUGa42sAEK6uidb/53oAfhcre6SCfI47Ra8vsBiyQ
dlGpQG6oZ7gIkvZ7n5r9lYg+Q5XVhqdACwMr9/EEHKmJabcs9lcS2nigj910mkuoUjBG73GByr5G
6mfTIapyWmKdXq7Dx3drfOL5xY/MptBoMqWdLrPps/JsUM3VKmAWxXrqiI3E1zdcYFE241V38xgp
lRMdMYBNZqklfMweKR/c9vvGl2LHiWsvwrQMErnnwtgYvcf8MVdqcec1j75Ni2eKj/TmWvvy0Yej
hGQR1jd2gNPTOqz6bTQIgVbz6NjP1hyCFmLBrm5AuncdsGv45FGETFtHvC7CqAUNjA0BfLTiTju1
u2HRzYwXJDQWwonXabdZuDO5Lza5Hu4+TyFHtg/OWZG6ameSHGxJ+n0/dkP3KcHqsPTb10e3jTcp
gZ32zLvlngM6/reJCLUcTIBTjPmGfs1t2LT2Ep2uWieKeA1WeSZJMTVPuDHhv/NQEKSmfIZHi6PX
Or7MbrtV9l98LBeNTPXTKsApRKUz0cVLPQnGoGvCtOEm7lEHs1uZjBq6JRmxVAqA1Ogje6PsFlWj
B0aZ+SGr4mL0ov7VPb+OhKXq5va81ar3rGeGViMuI3wmTh8hcHsNxbClGCKczWr8UOGs36pLSSJ6
YtFO+0vOcQR5BspkYw8uuY2fKS7jNVEzQmuM11VEezwmeGxOkBhcQh4pbOmxTTZEc0JIvxFsk/a6
ucZ0hmS8m7VAvESY3r9eBD2ziHOVUDLSpHTWUVoo0XW3wZyHmsrpVcemYx2fKyyzdl6Tpd/DULhX
1UZo8B9xh6LY4Cz0tpBWGW51XWpe9S6j9V6BFHRecetQ3aGxQ06l0e9bzV8Lokj8kc81ocR1QTJl
hoR4uL4t9NpC2tpdflTLOepBFuq0oETR3woCM8dMgTkjQA0rSq37pKQJIY03ZT/0L8JTYzd1sT2y
Prg01594RFNqYYD4UKh4+0LDiXZAdYnIypuiIiWWxzHa51FhMI1N0LyE0W8rsQ1oL+WkbefCILb2
KlKHa4Mbc2wgV/hjBwELO8/Bu6DlekYmjKVIdAylGV945LMnugFFmKXLPiH3RuZaPd4aIOu0PZQM
hNMKzQUris3jdbRZJlpdMEO5ZLjJiXYqpDNEIwi3BDfEGxYuhhslyOpozG8epfw8P9N+aujgbSLV
77FHQ961CuJDeJjXIvF181tF375wV8+gLyPbDOqqpNVTMP3Mq9hq8MspNlbb8YBLkWxSguKNfspP
RZelkDCSppzq4ovHtjsDlfikJ7gUXVwTeOoj3rOpcSfrndGCLhPsAAAea8FS0HRAHAyaIALvdgry
dZmQceaGK8mi9c9YZ44uIsqBml3QstFHuWOp4Kwg+HSAGNVif3iNl2plJUkt2r/UerUIUxYYueOz
an0e4mEDxsnmIHbZgCeRYjC29WI2Adm30F/xzKws0v5feEb2ynrMxMx78yZ/LBJb9gU0yxfkN2N7
CDtgCrRdOACCRNrH+vVlvcRs0VkhT66ZWssuqGp4n8LHpEy+0E4X7Qf5ltDIF+tWRrkiX3LwykV1
XX/F6ceYgi2Lk09V6WbEKufe75tIVuZEWc7e/fsSqjc38CHvAsFFMjsil0le+tjAY6BJXyG5ofDQ
uWDKhAciY8aeJjuUH+FWE3MbJikf2eBgAsg8xn2vcuUjYu52ejeCe8GR09WWyaOfDwgojsPHpqGn
uFe/5iWOIUamapQzMQ0kbw/lQ8XpuFshSDt+RcYraJIIaap8uyxPnYFPVysqwPWFo/LNXMftRczv
pAtTRWQXd4/yoyBDk4T/dCYHUXPIovCAm9XDfGGRIquUzIKJ+ZenZcWUX9gTx4yebx10tT1frSAY
FAa1F+AlEnbABE2/oiPco6RZFKP2Wv7MVWTb5iW5c3srtApcQ11cdMGcf7qPoeUY/WqiC86juubu
vDrFdp/nmb7qwSeECZDmFaBCEfh9fSNXUlcgxu2FAH/iSYWjI7fBrYWMA/GgOXC+FU4E1Ghpdmw5
kfo5RhySq2B8rPioy9Gc8bOtrlQJMJw9ggkHe2eZRoJjSBbvLCecYBVDiSifQrcpZ1aNuFHpo7EU
SVSoSfFuftqDDzusHF+h6QlUTlfwkNXQ1nSMYUbdujijKzmR+uaSYme4JGb3nrARzJOXj5oov8A6
vNY9AGmJnq7Hs28H55yTe/3pQfwITU5ISZfNrol//UaqH9n+Kt9bdQ9EPmF8UAMpb8SUfjJk4Ku5
RA2BvZrduJ9393zXzJiNF1eWHp/CcH4eQQoTZ/+xn2hrjDOSAXEqAYL7ewGhj4pObQmzePjnabUF
EAhlU1VvGPV1r7kOjwk5BHHTCBwR1qSQ5KGuwLN0pLpY8Fon2uQJjaO/5Y3+VmPSMyspB75SeX68
fAps+/1umLPqWQQO0f0xhQZZCES1iTCrfyMd3PDUVIVNQk/oHYUT1oQ7j9Nulmk0mt9+GUpiB/Q4
URe9+mRgm6IPpoS/HGkl2jSf7iuwJs01/f8oeZTV0rr00WEWKBdMPR4K6gFpCqb3936jMtSc6Gji
bY4Z75EUrw/8plvuO1smW+BfAMWlTp6CErnoR4tt9ODphLbOHRfohgnbi79gh+fhCe5RenHoZ5h1
Pb0Wradl/3g0CAZ73nOMRfJ0clHfnFM60Kg7Q3I88bq5wMlbUU5uGFdOjdauWvCqSkVudPgk4ZcN
tVsFXlP4ARNNlyquRlPYAeIkg1eD8hErv8CYNYxYRW6GIWo70T5Zc8lXymBE6MbRtgQmt32JXhnk
r8IgSTEaURJ/39GXB2O/o7xCF8K+ijMBsf7ITz9n3pGfkRxAWdtBYTFjj33T6FWGUo6ip6yK5/gZ
dgIS9jA1gQJcFWWkUiyhHbiJKxgXk5eNcNydy3HapxCJtLv4wZ6nUTA39dHaWXsm0twFBVyTgbnu
TTayMyHNMYf8XxTvzPBJ8r8/KJuGdTEwZg79Ihp5SdAFNPLpgQwFTla3Iwf39P3WmBzaJcjNiQrS
uFW6GRKOeCRs5QYjnF4Qn/MalFyfaCvbScm6ehbmmIuJL5bJodkJKsjp1HG7cPmubLxLnwntDsAm
xE+x2/VOMVbAuqmExO89P9KImk1vNPDD6kXmxbUZisywwvTWO6Q/ZdQjBDgDrbAOVwAfLebNzC59
im3S+BlgJ3UlMoa+zcH01MEtVY4VyHRho75rjei24kDRrXw8I+0NIWBPOlPLZW7Flo1WTMOl/hFB
8kMU9qu+QfrhVVLjTwD7tfcCjN80JuYVdHmL/tHCXh5kb7yXR66x1PwRNufVvvaVekqYuTuq5wwc
rC9fX/LRTi/KkMgWlfVbarhKAhX/8+xnPQqk6ENBZ6jTI9JHzQR0kAKK0+hmg5wv8e6VTN93wGZy
rIc9NwGuFMwuPGUwqeHiHQ/PDjK6IpyF7/MsOvxRf0RbEyeQeSNcdHW+gZxazBD4FlHVK5ARU3l2
O6aSCw64vwjsUwOKMo1nVzusXM72ley/pcTLghJp0tU2gLA/yTUnw7v56iLQp/PW3lj9kjnXCuIm
o62/NRvmEeCJ7rdBW2dhQ8T/wmhABId8H8FWV+zlovUXI2sBeBcJVcXfDiv6nHcf/QLqxCnn2G1T
JgO4maNs2o9N8eI+OHP71zbO0x0EVEu11fjKZz3XjBJkdTKDCjOrpQ7S7C/T5XdHqBDCalyCn1Nk
JNXbBlyPrAezPze3ZubGKIEr4qZTDkWAbNhKpXGRZcsInsjCuC87TiRabPqXuYPDKabLUpm7y4fR
VQzp2DUf77/yIZ+CViUptbaSNuHQLQBsgSRxUInGkE/0suAHlzJ7I3PC0990VCO1pLfzUfaFPMts
3TY0z7EVHoECCKmmaKb7PdDkU4R4bd4X9Ri/YayHIyp8njgB7ewJ0Et/Mk4nsqpTiNp5rL0AMNtw
ZhrDnjSVa4XEyRuSRC5MY5wSOGawBsOcfi/CRxuNWJDESukvuE2LMDDbTll1kj/rkbKzKLh5ISvZ
nxslQAT/D3bwP/1RbQIZFAPnw4SSMM8FPAvHLoQy+pSF45z68Ye3XmW88WhH5/asj/KWubGuFaaH
I9KgtKFerISupEflCwf2rYqocj7OPH8E6ERkm0U39wUTbbcNweEveU1ACoHYjaamR8KEgACGI/ma
of6gUwlWC+YHib9MLbKHJjishOPcq++bMK3ynRXbIRU8AzuoPebsFzKnJlIQaZ2q/9hJmqDB4Imj
JJH8N9GczrlatS4osIC+6agVKAfjkUMoE/6HyKTxCZVFwBk6uivbD1hxRaAPii8VjLLW4ZCcztBp
Nzx5TeYguj3R+WOMGG6rplbl/GsDor9RLGDcAKyhcdKWSTrkvV9+jFxfFygpRFEAN/3Xv/NyBbBR
CZIyGVEScZa/ryzUUauin0GL+AVq/ulWZdBkYBFL03xR1LoxSFrz5UAYerj1eqcfFthtnDAHO4ss
IVCLJeycJ1P/ZqI63GUElE2Vz8G3MmT6voFsRXv1+JnPrrMY0uvamJfHcsU/KPL1ccYpk+MDGO2n
F/yDlt0fHOvjpNjrjRXFmnP6X6RNRZNH9NtSIi6XVyxcdTjz5M1CV4ruXEa+5SC8nkfkYocfK3C3
aVYnuUDsFqVAK34i5cYiyY32eeLUl4vfOvliyQa9o3qEk5/w0ZHv6Mbnj1naTR4+Y8kMGc0xLqX4
FJ8dvwy7C/nch0zZJ1Yakb7gqMDeUDUtzsJtKqNGOXswFGYfFUVByoofR2o9gSkmfZZkrh966bRe
Vxua7PfjsWUTQst9ZscajpQf2jhXrHCkvB1O8FaMin3pQ4e/nVBPZrrDR+cRSmgU9ufw3vdifPe8
tpbksTJuybB+XfqvoQLIw9PX9ruxA1dLEZGR2NZo94zELY0OwBn1aC9qa+DIC/LzXaY4J3zQ469p
V9xAwaMAQMtb65hbrJ6Pyju9TAEIFgjx6aSqa8Nu6agMNK0CUP/0a/LKfxshkuDTEv83WT0N7GOL
GgfMWXke0mVLbp8H1JvB2KyPMW3NMCgXA86llmkxeRcCK8Bg1iWUQv6skdP60VywtW8XlaWLu20d
QwJQaaj8FBUdLpYIEsISf2vTexX6eJJMuDKKfz7RGvZqCYl+ZT63DKNc5bo/nzyMAQ4w/HgVk0MZ
gxkWyRqw8wl9cgUAdy+wgKxzteDY/upcC/XciLxdJQUIheh2Izzlhm0MDGFzOPO5HKE2S8zGcN1T
RJWN7CGoGSThFrhKsXpkQBb49/tqAt2e64Yf9jM+VmH0gtzkywu1BpbnLNMk01Ehn/Vmvcb06DFC
j4QYiUYH5xnIUy+Mi4jBM/U9icvMcuScVSZw7QhDLsYH2FhFyuRSq4Z4bK+tN4s96CAGWAzb66f4
9DZMVZqGkGav2xKJskimSZYeYy/niavCoctgdSJFMqj380CjXYYsVU55RgQAWPRcP9ylBfz3RxFJ
wl0IwvZv5/tdmCjRZEPejt11L7MCeUA/lFT/uA1YjfBYk8CfJ4MXahS8Lo/hPdxbA9m+LSdInm/p
3PPVD/MmKLmYBudg7IRv7ruFP21t+QcF6LuBXBBK/3Y8zsjqgNn2SonogrbDx980SQipB1/O3RGr
fyfhCXqvn0a82U2LYv9cV6GqvH4yKSS6Giyl/Oo3V/AGl718fOJVfWBempcab3dwDtcpzqe9fXQA
rS/nM4yfsTTPDgbab8IF00ovfKf3H6q6GpJzklqHpWBWuO0fRmFoPqfUH8mMyfSp0SmqxHy2KjI0
Q+NK0/2+oNhpryTeDicw39xewczu/Nen7GbFEMIvHdLm9XPzVsu5VEcwA42Ac/AO34DWRFfpl55d
sI1IxMCmzg8LOBRboccqvY4TIZA6XHOWq1hUiirbizUxeRphWiYgo/gao6i7Gi8uKWAR/WlU7IX4
14n7Ytg3lI/o7SKpGH6lJDePzvNjUBwTPrj0ylfrNlYNKKfgA5K781VGYdD7YlYG6ysjT8P6D5yB
pQecCR8snRwZSmFwLOhAY4dv+08Dd8VKYDNiETcPA7R9AeyendgbhJATSRLrzCgpq/iYMJXpdf+s
CfAxs/cuscd/DG6BgediW5GAZGyPgbrZjqHnB88mhED7IS/QywFuF2fg/UxoUS4/TeyhtcWudFLa
84E79OUYCnY3NMtpLBUOPFgipa8SYHP7Gs+L7N6QfnEQOMORD876FlykFzQQ6FHpjFxyippW57cX
CPC/XyZ3+WRu+vKZlMIxQMt84jIvfK6LNbUbPOKeKIKQL1lpSWepqdif9XwkxcukL14jWrSt3hgr
7YCe3YdvWH35sEKxWYXYDODFN4zDX7+WLny+ppOEi3lN9TQSmX2v1usJNJ5ARWAQJq3MCw89YDan
DtHFLGhyn8tofv4wosyflYyRm/u9nksAf10PXX+Atj2nqeCFkp8fPWVkaQoWMbjO1dIof6lwgsKK
okbSwL3p6nqAvF5Wk2TJTZPmGteAAx0HMI10/kFcFFvxNpUMT0bt+tvqd5HqoA3GZjZ3+t5Osk5X
MJTwVPA5WDYRPuTM/nlR6apOmLx3/NszQyaUgyNuwfUSYgzLZR/06VafKyK0tzqB1dI5klPWlCzc
pGCJ1HLQj2IY00Xl+7tsG6QGXUrz/aplmH5/LIBmSfrjaBsvxXJsVxh7ZXnuycM2rd9CEhy2aV6d
uDaqw7boJtdBbdOH4WRV8bvmAlaEgM7BmWtw7G16qUyIe+QYbl9XyNTQsLQcAY06X2HeGMqdGJYy
PsgXQPQ6VX1b82IIh27G0jZyGlMZ0r87393lnfpsVSoMEwv8r0vYa16EkAh6WAXZ5X76gdOBqE9o
+ABW7TAiexBb4iHK+7EYd0hfDcGZ1bNdhKIMIBIvdjoouRk0fCcvD3wFihuadJFQaONjfxFe3VHz
5uKnj2M1yUTWZw/tEbgty+nHrMxtpf92F5iyqJZnQW/Cx/gw2a8XfLvJgcmNTnYO3+wI8harTDUk
iuitI/gWWwa9z4YHSEy8PoZkGr7zOrKlrM1+jv7sYKatyhQPlAUdF07RrytwebJS3UliCZOZ2m42
ep3dz8ZPczHeXWLF5lJP9bt49EIeFfAoWX8eEZ0UR/6ekqlk8wiuRvmqpkfDMZSblJzGyhlP2jjN
r5yfWI5h/BgddP6SAZ1FT+huQsV1p2553ArP7EuAAm1iKIu8DNCMzN2NA1kZNWsFpt60QKl7HUCb
c169xLKg/wxfdFOsIMMrPZDVhwveLQLaaBiOjydFV1VBdouAgANEG9smSEUQb1PjUWmo3VP/YvD0
2P0rQcfG1RNRJfTv04VPmPy67E84jTLOM0Ay+lplHxPYINADVHwfeg3CrkAvz4aLQ8M5hzAoOTZ4
2waEh6GogZ2CAQLYUrkYLUDuJi50EHZYL2kzXeMUCfHwhY+3oak6Pqc1UiAcppkE8cA0Ce/kaOmc
Bg8jigxFbHHMW+USyoEn9nwoFsbVtk7DtS7ilfZNFD9me1CUxRPdE0XmyM7qmMvce+dFtELG7lOm
gXeVNt4E5ee3KQEzuHG5+5kgIa8mKcQshIgCvUjEX39psnmJDRIhOrgP0VRUqVQXftT650KcXv11
3yKW3X6+URR6FEasW/HNT0CofvGIziVos2gMPkPo/T6GeCyF0N2b/jGJn+SQ7Ttb/n8Tfuf0ROPm
EFGueT7HI/Iia3MlH/mJAShV/PvuLbLIs1+1DtnTI8JHzWoxpWNNRu2H4ZUUIRZgz406LN3Jmczk
ZKejAfArjwSz9UqsKlEVQADLfUDEB8QiSGZl26TSYie/7gXvE3g2515huHH6gQ1aGxLtoFj/+naI
LwupnWKlVLN0iIQlyFkFVnhBEcxG+T9jMenqyra5lV5UP7kqz8N6nUW1esV7ngzyU54CwHCy9HRn
4/t8Wzd4mzkirWna+9IAAdaBmW7SaMbQ+qJtTOuvsLkWV1kP987MnlLMRIAZXzRNG0xYA8NkBiD2
ojTfFLK/63n/1S2zPH9yIHxk40uWQ2Iw3UrzQDdrXgiPLaQ0tOdCiFIBMSpRh9yHs5wZVWC2Xw0N
Muswvtuqfr403YyZ4/K57w0VLckBmq3UNgtpqJ+u9ng/8icrSvf4YGN0P08dHaYYPvfnZ3ROhzts
xPkGWLIR6LTmUsKyhICGRuCmQCsU7LQ8ttTgnPK5OyItB8mh6QghezzjwmZ5cU1M+0SobQbsyE3c
4XiyIYkh14b/Jgo8J4bANiSnTvoLBtJ2ia1Ea5Irjbf33EDb2GGhP3s21z75VmyZXuiZbmU9AQa3
tRvLFF0D5sZ7065HKtN/2TeIppc8mn6rXu2pqAzkCEHEypUdkTq050JkR8MMIkFSbYtSOushZuWq
P4XQ5opUIXF2v2kCdfqBA1WDItW3JljXz+qpkmJVhwBa0X4fG+chNHwM2q4umWiLEbWeiWhRIMwj
hZO2Tyf0RwjyCsmw/c2Ps4EdLR/kb/tlsDe2PTz3bdBlFcRR8o6Nm676RSuW4aIAC9xH5zXAQGkX
bMV5SSNjr+143A0oKjcJCiYajW6HnMV8Dd+CwszycCgmkUcuGMMaQfA1AztVHakfUQ7Ua0Fpt0S5
3gYu9T3MLEHsWruLOpEmmECIsbQ3ENhqdUd0QOhpky7kdDzsZLaSHLib5ZaU4cM07Uf566GiePuA
7ZF1/obB15YZMFT4gN7Rtnc1uzDDmMNW44BspuYt8UMCw3BCkh6xFwqmFdoRBJfZucvxigmbseo/
tEw/0rH+ncgtHUPd2gCnXp2Dm04a1UEx33T2vphSxzeMtR7WLwsbNMlpSNGd3InIK6Xq/0sLN5m3
XoR3e5gmneBqaZ8l5N21vtix0LbInwob2p1ksPWHzil/M6dzF1pkHF30i2oFW52VH8Ra0GzQF/dV
yGIwxGqf9dvNENyaTHQtK+Za2IKnWNhnw6mRsRYaIMNNsaRn8ffiOEnTOpy//pEiqzcm/AK+hBBF
vRjw7tWsakLzaA7CKFvjaWw68ik5f0WnNLHWMvfzvsneDbt7T+jcKnvBhVQyEbdPG5qI+pYpbxfX
1PXwOWJL/jsCKDuN1d/lv3IVI1x7s2o7Vavh7Ml6yamkKCAO4Qomwgrln6I62vHdOS0ElWf2ZvW/
seaxPtShhk5bmezJaFIvdo7UhfY6kPJhqDzh8sTH/b0HX4BjFBa+vxVFCYw3GqN9YO5dfM36hKqu
tVk+94YsLX9SU9RBlaSRQG0Je5jB5RmtgiNZk5xO0BrEh7KUdaacPcuOJ6EJM9TT5guFOtJnKHDK
qUOen8wJRh/3eYED5CSGszWQWJc3XwdCEIg6hGllms3oTXkOn2vb2sVbFX+s8Uri41l0j9gBtbtU
VyFWLUtGC9s2BnQHHqxo8QWMBq2CQP4oiUT1X4EE1zdqYeobWW9fR5YHayC10Tkp7FKONCN1FFV/
pcN/DE8Xa3J8R0kmbZ7VXg6tepbalD0wKWWM/xosFN9k2opyYeS9maak7KjXIAipFsrrXvkc+55S
rnDLiqBDxk0qzFLpkxlZt8PjJtkrX2LrFBZBcPmOSqrc/RRdIHwf3lgTr5qpVLr4Ua5N+ORRcTm2
y0aMdEIowMDcQJkMZA1O1yA78siq1o/l/mHfQ+5pRmCaKiPzOlQmWyhrIlmMP+2lFnTrvxmHcARh
HlQccIf1onvq3iuNCQrWfYE9b/Hw4kVdtH1B4gGSFdC2zz8Tgf5LxQbZzhKwwTz6YO/O9W1le35H
VNAA2Snw7E37IOCmtMeDIRgFybQzX90/JViW+iyTz4/CHbgnSTkE35kyal5f0n0XvA92AxMNb4lA
KDtJzTclgnOKivaM4FPgGzKKDeNeSgBINfwlh0bPtdpv0xvVoq5Fqfln1hWjwGXcM8jqy7GH/oXa
b3ToEYD9gJuYbcT5gb7mXT4UMT4Z7ZnusxncXQiYf3mlpk7cWVyEE/hrSgvkluYXdASPiwXplrTg
PS3vBartsaUHUz7EVmqKuGvLIHKHZSHx/lHWzdE+v9roG1ZDO1oiN6GCXNi1rGLMxjVJevuLPrTO
PUK4ie5z0GDhvMdpdjXfeuW+exV+rxvwLH7gPdVEWyGK6zhHK3qej3DspGkeN4N2HKgE5R8EDNFe
pSQOCT3lZ0haEkxSWtmw3k0Y2vn68YFMI08ve0dveVZi11filqozcdYykQ9/t6Q6LjteWvuC9C7e
xCtxGttsHnMeLgZtDfOQtMvUzeTrnDg2uGBoAFzrK/uk6xl1t5CZKVLIvRYiR6nCug4YEv18cDui
EEr8gK0SQt85+uqsSAXWgNlciyYiZaBMnVnirU+ojUQUGbQHNZHlBNWEer7WUxA+2cN7cvihp+5s
gQTGfDfH4wmTU1BoeQdlg/NFEc9ZPAT2nGMNHxY5ysYHmPW0nXUs34Lj6jRgBMNB5UAKvD0N4XjV
U3Vb1B4z78Snc3QLjWDiW0VSXh08gUSkt4GGfYzpV6QDtKR7yO2rh/89o/xByhQhs4hom4bwUcKj
SSYhzILzemaYD6oer36OXzd1nm2FMtv90jMjK8D7oMVjpAAaMb2InVcxkx0UbS2YGmylyC7ktkgz
Aj0w7aVsNZkaj+l6drNUsMfS7JkULVL76vsGTX+sNwPebyM8CJwjpR0B0NTqtKTpd7is6boan3Qs
a1VjmApxiEUzrcptfAGyObb3EilXxQIlTxJlwPkKYQZ2rMU25s835PU4DcjS17ons9DYcJPUojYc
mNXkvXjnC+6jpSCP10qMmsi59gaKZU0sO7w0JKaHM+wMmn8EO2X01v/BLUsim+9ktNfO8YSjG6La
QqBW6eA/SCbMKi8nOBvs9M9+Xrhii3Y7Bhi3JkPNlFOo9JhSr5r1uSxVE6izwYVhi7P1e8ROuySM
SGs+XFWm2s3KwpMIZOZhNVYqW10RuTaC4ndq5PwzSUy6XBTvpJmpdeOUd2L/tFhNoieR4kpJCw90
MEySNHR9X5lkbwtQDVfbyllUx3M3cZjY3GqZE4mqq2siSgW/9pAKv/vXq4LjmAJcc13eP1RSbBQ6
HCI624ynp/FOXmR3/aVTqB8JZhkvvFS5QpGz00m4e+l4fLCT3BmcfEu22i/5Y64nvfaAMHqAnYoB
wGQ9C8h0bb7xGFlkoqTe/AVePXgZz3Y7cwCbhreVYziInO0FXyKCzfeSRZZI6oIecS8ogSWZuIGn
bVz8rCSZKsXQxt1HAOpukyh1PjTnxjl/gHLyXBa69FTntSUOWKkh1RNncFYtWP3F26/+HCrRwZiR
F5TZSHK5R/fIliavDntg/8vUTkHIjCitpJYaakI0TgcrzNWaLwZOMpoOcQSgVr2mxsit6xocVxvW
eDzNlPBjzbmavRsSy34lS7QYzKR4ppWjCgYKeoPg44cBbVz+hFZFFTGGVralLbSqjaYi0qxPNNed
gKugUVsiqAHtT5eWznFmIcU9dz4GmOgWhwg8tR1DWCMUMxXwpw3snOH+NJISyB8KfD0jPUVgJGKO
4CgxRAlbSIP0yqlU/xzrngqKr6ThTWVt97Yf/bNU1VCoawfERTZarWx3DgOxNoZnNfErNAHPR+Ua
75gS+DuAsM9Yc8FErANzbDxJuQJHlTyOuTb3zFmWmHKnQP0alITnAYAjNNxHMZNMJ72SvvGLAhYV
eYSWkIjj/aO3tS8YN6BH/uPhGnAP2pfUs6rB6TV9D7WkTXMiuvp+zomQiRPO413YwHBLN+T+vqRI
z1PN+Vl8g3N1df9tTSxKv6h8N8OE7QFhICLsK1qCxT4b/ao1jz2NmYtmiHJzwou+Phq5OFGgJF/R
xrgzRT4SvgdBAUZuKWbT5uqkYiFPGjhSoghOarw6ahBaedYHZf2BzU0+iN7xdONweRK7i6fqWCCi
IvZzQoBt3gSQ9d1zw890e0zxOk/Dj3QAQnzXo2XWIKzYiLjszJ2gsEZXtDNiAB3LA/FrDzPTAjiP
VePpM7jovO22lSlzUQ7d+bqbo3JS8toXm+06Q9evWgfAD8b9rG5aknHe9xd9c0or1TBjqpz6XvuS
7wQnHdveVOQaX5/fKIud5J2NXGXE/txA6KztepC7RybwsiRJTn7SyrDDonZ2+1LE9BR6PVaCPash
tU2snU4V5W0b6KPs4ILm6/d5o+cfvMxgQTCyAS6pZnWoDknekby+v6GnfsAToW//BvNYC1LXhl6Q
mvCr2Rd9GTYNcyB8iaKyMj3heD4qipF6jX3KVAwRktsZpDnJcXtSky2gIcG3geQHUX5oZ00jRHqv
bmrG9uVgtY024MhX4ECTcIalw8o0T8DJjUfurUZ9f3zhAKjKlp7vHYheVP0360+H12TIY6zk+2Rr
01vlJ2yIgI+jtQOBNu4sX1rHG2JlCmZnUZC9e2dz0vUFT1c4PRUu+/ROZkLOqc8kICXWgPOcS7fq
JE8UmzAoZAKu8W2CcRTXMoXZ4ttGt4lqDPEOCcaeRpm81DWyiwxbZ9WW402IYzYYQz2UzAaA8sk9
0kgEfplzUjriK2nFcDxXRQIAvSoqtYyexVhWDuRNjofJOF5WsRJb8BD+el3nBKgELoG5nVF28dSC
JFyUqtES4MfXHC7l9C+cnWNktWGgE9nLkzGaHw3cbMtFfmcnCmPoaBiC63V7MsOnlSbw0K5mGZ+p
x+K3bVg3Q9ZDNO+Ikep94mKNU+ZQVs6Ow1RmS4wsoUXmE6++/po6Oe7VRX+/cu6btvyLpFmGVjf6
YpM26NhSqNkRSwPDCGnMzonDDYu+f56kSzhAbAZO53P1sAQJk+fmCsqmg0kAbWYm5kCRfR6/9ItH
wOpb0Joy6/6MR0IhfSP+iy20Em1kAAu7qjXdZJy6I75/TZ/hMK/cq3+bPDNZwgUrigiUK282gBpk
5WuajFhEcF65FcAMm5kRmYVkK6Ba/xeYew9+CWHPLt+DRkul3lzSL3bz8ViqsgpDEKFGh3VH5/Go
tMoeLgAuD+igXrmfBbchF2hcd8PWwTBRbRYqqPRbspQ++x6yNTYC5bpMHlsLh8xBIOQ/AdNeW3dM
nP5OWXkeFkf4xRloWQwsBeiy3Fm3RyEY4wfAacIvtb8Bah8eP/D40GJYY3eC3udj7z1fCIX2rPDu
AQlIruTX7o8WagDqJwdKjMccUliHdZTVGBvVh3DyTQifEglfe1BS3MKlA2+TmFh+ISelG5EWXxVM
nsF2MS4yaVbCSRwoOijv+8RBjJ12y8QRTRcMbI89Cue1L/z66h8UN9Fkjr0cjXzxGTwcNcLX5Qlx
BaDhoiS2bMBvzkVem7tKJdOI4FT0gUEAxVat8AGZBuU4IEkYQ3Ea3D+BNJ4CwAHC6e8jNRoUvyYc
JGLuN/TINkVXEWB3gIxmyXDjfBLBgsRr+pIU4PJaFclxVTq05J4XjmyzmgXMhuaPFQ1uttiYmzKT
MylaOt55uAbzsULDCNUwsmb/pFuGVckjjqwbSbGp75vE0gb6Ku9/EgipwCCUZOWArMqU/q9UutEl
yTS5CT41rE0Yk51YYyrKrKwR8w4N38h2/32jongsKMjVW/tAfL8Q5RX9wpFi54HpvnWWqmvxr+hv
UWrAw0w2+BEREmQquxQHeoY0AF5gIZ2R/FZp12moHsI0UIkIeTPiNOKBBQwH31lOlybS9dHLT1mw
UV4yZa0juXNgRIX2cgt2xg5oInXQ8HlaDEgbWNH2QJtlrvrqO39r3UuUnYlxauyyTLOe7jRnOcBh
jTh2eIE723SVl09q1hOjSMeWhwB25qcy8fmeyQlhj4C3DA6A7frEBN4i1GRKSB+SOkGtP1Pd/dez
g4sYoacWJm8BWXhcS/IEGS8+NfV8l0BPov1ssWdNWifdt6rWp/W2kMQHbx6Q7sXg1Z0Z66cTmNpA
9KxJEA1LHq/xkZEbBuuMnf+JgQZuaPbMZeDLkQzA7+nRrUPdfoEZBmZbvP+Yai6aB/4dy4erd2cL
ztc+ctY6TGHBerMoZR1AXgpSxB3nQqIhU9KptOI2wXJwvBJlgDCiys0f5qV/qy/jFp9agfGhknMA
le59ggZuuJWGe2qiZ/k6aML45IrfNitPKODfSMziTJrSY0h6bJmvDEB+4EBhqDRjkFS7v2vlu78Z
J1EfiSUC3MAv1V8I+eP6/lxxtATKoRXngi2bTTOpy8VE37O77rPnYFs5/cDnQJcIUsmZY58H2R8o
lSiYhFPK6X+CQQUmFcDOtSK1fdQ1ANZn+vMq8Uf5pM4bL6USkjA4MQhdpTLcOTn1EddOgyrq2r6d
mhSzwqtCpgiZPW011XG9797Zre+AgJQpYo6VrboCL7a9KzjafxdIio3AiOfpu/ZQcoth8kZOj019
tvLnKcZ9YGaY0FVeg0UnNd64JoS7tlydgUk/LllYpVPWRlb8nfWbMRxl4YZUwwd205gvWcLWdR/e
QLyKUH2KFJ3BJ9gmPiYdDD7iw7gVBJLCtI7z7wcJl8y7SD9zwujTdaodxgYYT6UpjV/wRH5ZILoM
QoELlm/WqdFnHwOh5LoqUyVaAS+U2W7WHQ4Cts3oAyUPZV8HlVYKx5NM4FVA7S/jYJGGxRFfBLGi
Yrtv8BUnJNCMmt+AYenQGB6xrWc6adw7/XyiE3SLKNg08O1YkrVzUlrc3OW79dyLtvhS0hnp680T
x4oQ+9O9kTn+9uIBXKYanEci77zC/Jr+FdtC9OKNm6pRTetrtTQinAw9CJX1TwyO/cPXzDCqFCVg
iMwr+pzvQuEjisYdWNjdNBUrTmGdx6PM2Zl3ylkWpZz4duoaoDSA/VTBpuSqJC+Gl2ZzN7BHBWmI
LaheVAd1L9OxPEooIbQJ/xLWFlhVafSGKywWdG1K2fCZHnRL+lSy3TVpt5hBPWTFeRuakPjpxz0S
mt3zq/aMe+lbr6Tc4AffSEKEXBkRLS2RazT+Jpo4D9oRJqzLIPUGJtQbNtNZ5EcPqn5Pe+K38Cj9
5aUFrzaMUB7FkJ24S+1BtT16C4WNj7qcXpvYmATY/JDtlQ8oJxeM/u3pbJUlbiFaW0R/kDfHmtP2
kG5lXvzKYgBWJWv7YQKWVsuk1IGJjyARWHEj6GqTJ+RUSdoaEcXD2QSQPnlwb4mxiYgD7elpATRL
ZpM8GuEngxuhorXKolQWwTIUnb5KAtPZNa0DTFE1FmCoXJ79q7guuLfobaH73k/xKg+9QaminO0y
P3PvF0R3RR0I1niS3y2IeuJPc+0bJED86senLpCXk48R9kF1gY0ifKVTcfuABMJBjywZtThQ4QDG
eXl0XR2nW5rDO+vn3ch7ZTk0i9guO+KJzq9KzSRgsiK9uyVG0qUojRB2LucWpVTazCM/CjlQLGqt
Uyw7XUSndnMF/FE3P+858X8yLQdSNA6XkV0hmMfYX1HKuHwFJb9XuJ+BHbh2bm+S5/nrMwfqPZ20
vMvxeNERWoqVAZbwYCSJWGv2NytFGBdMaDomhqXn25zJTtcTlzyuPGQhLRAWbTtHMSo7VN6+xfiH
6kv0jfa787pPIf5lAVWtGh8N09jU1Twib5T89Hb+jYcOoYm5vC9tkgeOX4uKJOMnF5Qqg+YdiJmR
k1csOhuRvFE0EUdZLjJT//3eZb1/NI2slE9RRAP49AFcZoxRNJaiLbig5fROD03AC3q+C8zwzec6
gKcDymZpr74NJGpH4EwrgGEsgA67PeD4uftw5oCQjEhdwtmJLD3wh6iH3LsJmC0oO6VIjK9Or27m
zaEKKjAXYuP/pp9BTHNTtiTSCYHkQUznv1wHqrpl8pNtn+UwvJkvIsEAK1CQK6LgS5IdBhwruFmk
FeCMmB/Cv8Y7jqsI+GlY1q7JFNUmvj+Rc/+B4Xdm2j5vBUYkPZORkumjBdSdpnMOIZgoBoBu2ugq
/4yFQon3bf2tghJVzw48337Jj9/5gPTBxO2fBJtxxWDvxlUIxjbldBKLUq3++qzXoZKu1eJGdldS
Kmqw6B9/EOqPdcLV86Hqf3oOFCOMYIAxu6mnlBS/SWVGHcmEpfaiGGw0M7eFyG2ieA6yC/HE9ydN
XZYt3t3q2YoZB9aN/6RlU/+Gz/IDgIebMc3wgjXIwsER2lNdKQ0XvkCFiU3AKOYdsGv+wtzyTKMd
xevZUHJ02T4hnP706FOOrvOvmREqSenijk1fUM0k8CJHXDtS0vaqRVebG+IwnEbKYKLECeWfcXL8
L0v4CJaoKJI6M0diGKUi+CAGtry8bRIQYOkXblUyjcLd8Jn5QUYizkX32a5osstlSp3kqacOEhPR
h3RWThkj1GfmTNWge4IAovfAOeYUVs8MRpHEqz7XGx6/yaH7Ew02vdTZuEyJjL/za9FBnsvK1wy/
KDcs5BflDweHEZzAzKXBeG419GDXXyBKqWbEYckan5hbuAjUwwz78m4KczcIh/rdW9S30OIPe4fN
Rh/0VAsSHE/J7vUGGCqykI5uH01mObzvQfEHJk+EFRuGcn4wU5V3n0xcRKs5gBe4EV9r5ZkfZDLy
dWGGyQTdv2K1DL8MB44bljPb3YLiU2z8D5oqGeR5rGMqfCmhhn5sX1WSBL/jMFx+vWGu0ZEWJ7TD
DEt67LzLP+xB59pjTNMYbj0oE373MNnUjN3xppRVrfjHKL1naFep03FpBRc9s+wCAJpyOuX3A7M0
m/q7rbo0JSAiadIk9icYqBBssZP35uKaxaRnoZ7HT06wbUIRAQZE6C0fa12AYyaFNKR9WjOE59sE
/0IF4KVRF9kp2UW/sOWnuIJMU9vf6o2N4M4aouvPjzd66LRnxYJnJgKq4nwTxKCrn58iCOWZJSL3
dzBFl91Baawp8Triw9lbShiejNy7ghUFFRPVSFi+dHI1SA9THqyERtbiCqNX8n/+7Mbp+2d0NaWQ
DP3b03Lw6iuQPsNALR+ZipWyyzrr4DQ71YVV/dQmRPJe2mEt1kSg593jtckNvABld7DvjleRwL4y
/gcN7mTJHedpXtEfgRPY9b+urxfobO1QbJVzK4t8md9nnZXeCChi4F6ULwKUqTIMrFYTCNQKBgNk
ct3e3He73/RWTAZkVWcaQkrGbtnxjNLVlSTzlG8zo6IrEIUvPqupnD7AcfNJgVleBfOlz0F7hntg
2TNC7ShvO1ClMM8Lc69B+Lflo3LZE5aQHbKw8DGk4AukbmBMzFWWZg0xOgFpVy0T9yt41DUCSqXG
mm5BlV9QUvVxNoN3vq4kHDPDdtjxC7qw+eJPV6WeVaSxlxqEf6aVgmfZsdSlW8vNK9XDE5RC0J+H
g9Cv2c1GeBjEeN8NOWc0muVVM7MeAczkVHbl5D83U67FyEG3d2AlfRoHfXUpvUqrW0XAd/OfFClP
Zcse6/oO3YA/yb1f9L1xe8aAhgLHOBh04ELZg0hidzEZa5Q8PeGmkzntoxLsKcrU+wTN2t1N2oB9
y6sa3annaeE9/xWcucUXpTEjknT2mYpFDO039aEcvDqNCG8KLJ2dk2bHcyFomgatpFLPIOWEDlLL
Q51RMyNMTUCAlfsVIHX9fPmlZm7/GDX3QNc80cm589Hrvn/l/wsv+doBVQ2bpoLclE+gJlak+/cE
bg36sFoBEvPyy5Axx3fXrup/Yq+8o95wJfv4RpNt4OrKNrcFTFueIf1Z8S4f12TIZNJ0gyVIgdH2
29ngbKk3NtPanW8UK2GXkqUCwRL1Rf0b2XByni0prr2SXa6ThCpQhTTJuYKz64ck5uxEfg3ze473
Qmzi/zMCcmXPFFBMzndwNnVUtpHY44m6MDg1AbfjU/pB+wUhhVg/2tkwSHURwyJjNp0WFwFWcmDb
GUdRZw/fHA0P3hQvJs0WKWm6467FbM+OYF80DQ5r32w3H86US6Wp4DSFlCyOmesD9A0DQPrq0t8I
GswuLUXv4qRpsTsSm7Nv2gKJaBWhq8t1o1RyF1cxw6rismGSy2QFJCtnaGidjuhcUkDJKSFlW9bM
5vlfY18sw2HQ02kkWhXtY3Cgv1Ef2CMXx46tJDzIKfpIYIwE5i7Vwj7CaXo3AqAS0w4b5L2gAlQL
OeHUlNsIvfpdCeoEWmN7zgrjUcVFqp8RCDzOPjCoFubMfMegmbOL9CaiPGJ3LbU5VLgKf8dcPrvj
Q9DOx/TVycyuCVRVp1pxCOwnTrcyBcG4pMVkvRYfKZTlhgH0AGcADY0ZeVHnAqZAhZiwmZEkx47q
N3xRNn0BhrdtLa3U3UoY9twEAX6a1YlRyk+g3bWEclPusbDqc3zSVybjlrfi7tgNv1QnJTc4bkFE
vZbwOS1L8nDS0mcpbbLd5ZTQJWopPp446LlVnj6y1isg4q4732jOt1HWdDibE3n0+9fhMNsGn38U
VQQqO8f/xBFpv1AVAIPYQP/yWUu4d6KSI2Mzwkyn4froFwp5NoNW0DmX0Eb3V60bOR6ktm5YO/pQ
1eT+dfiaqWMS0SDFcS5e/UrdwkK3werRFoMfTw9aoLOvWXgFwiFn5lWY6aeFYY85B6xR2rTAKFPM
dOG4+ypo2RFsnKmzjF/hUF1nI4gIrazuz1ppyZq1OWrBIsVveEAmHgt7iwUWl10JkJZiKSFNKmfe
dOJZ9ehsU0n/L25yjs+mwP8s7MLO8oFzVmUfa7h8+M8Qh85O8e8ZZDb6sv3FnawT5Ity7GpBSNT/
vqJfK51MGaU84CNQFaYxG5Mk8l8Hmeo8GkQY6U3z1PDWouinLDc2WU30CVw4XDxiC5HeMKxOoyvO
tp/lHUX0orEvNCZSyVUOP4QgWfaxgnPIvnpoNYSGXKDpDKEEQAuJOMexlbDXJGhUlTbztS7tkGTW
3uAKsnIUADYqw7GHTJTC+OsByMIBxgln3itr0cY2h3teIUZbIrTlD+LnyVz4mjEypZNqposdzP/R
se1Ay8Ksbx/5nuBCGHVAp5G5mPmHYZoFEVQWTv5J/0ibEfq7CrzSrsK45Cx0NKZrXHrVMzoBShFw
cSvAGLYLSIMlPk2OFprYPedtsiB75yPdIjKES827Nh6jIv4KaGYd9sLPChOteK5ItRQ043rFJ050
ztONw16wU9L09rdhhQmLEKVNkBpTw72D9ZRJibTE1i9fbJd4/1zbkrN0Dx+E33wtcbJ/0eAtzkxu
GbWhj+7R1ZV3DvHz4OcMbm9WkXG9UM9uwAHKlwpF5RzCkRQr29XnYPgsHZaeAiuPileW7+uXdBK4
bzgt1D8XIMXskKkia+zcCSUn03ZoGxlOpe5QiLfK4bkfS2wcD4i8oLxVN8KHNhxH+rveRsuNUg+0
FJm9s1DUvpplSTxEFu3ql1VbnUpGk9C/oyLsG2ZmUB0Atqa9Eg4FpFt8MbYx4SiifDsDrGhSlMkH
6siqaNShx5/8MHdBfsA20DAr3nTNEQHAWRtixJs0RKuXxspPPWLazQ9r6fXHpHWOBpyh9uiYoLWl
1VI4wFoFPePH7u/SYbQ5eITPP1M5buSIsD6zhvDT1hmYp03Vcg/T7042B3PBdaiyvOGEH15OjcJ7
bGmZ1NFrNL60saXUTcBwLrfZ2rZ+5c+Fitk++5NAXYnQ9EOeR2zCyljYmXuhjm5GYu9IiavXMb9Y
gFRRK5/Wiw/aUwcLrKgOP38f5S20OqnxB0CsufyoHMtpFUI4ZQodpW9R/wQ8k15d2jUGkb0hSNnO
X7jMHIHwYzO5FZAdiEhg37rrFUsmrmAagmaVo0EdgU2roKrSQGK9bH3vtRbeGBqM4L+A5odLkz4K
YR6iSJ73m6qNuH8HrAdJ/qRkpFIHrBCBHzsS9yGqXrgFYAC4A+VoBbWP56EP5vlgmdtUkk5/cEGa
j8OavMr9Tr3LspYeP6iYQ+DUzmW8HG9hwy4ApX8KHIirsXwVoHZguprykEtLigy3H7IWPfnjC7gS
yE0ASPzzEy8p//WPpF9XjC6vSswMABTOmxogHObP/613750P6o2u6Ib66N1LwWyJ/B0qjZC2ME0G
bHWV/A5VEvNUfmiwXwvVqcJA5lTMb/m58tSBEOY4P3FEUexQZ1d5b07lhGcPZ9ECT0jHfTo4U1Ux
JqdAJtUNvgPuJafh+dJPgXiOQlPMga1t0Ew0j2FULudp1EadrXYrEkxUE404C16awmjx0lL1kC15
WLAb0T/EsCeg5uWYWdKIzvHIic0cfecmmz9Zg0inqoJMB+YXNQsW3ZKWzyRS4rn4zgm7qxbTDB2t
nHjOD+qyN9dVfnpwaMkURkif/5F17SIgLaz0xkkMfBLB3GzaWr8fGnWkQqQs8hKqQeQ6UIoaI5lW
xORqAv+r/1TJCVsSe3ZB1cwB1/0WR9802KmEl+8mARA0CMF+Oi2HFgCcyKH96Igz0RiZh+GSwPFm
kD/1wstRGCzg+wC8FuczR4YDyy0fkA8p8OvLijnv6eA5PyPUwjqPvCpHk/778c15DzFJ3dpNBrSS
q523dplB0XoqN8eVk/VY+CPB+UDzNUnvx+2G2GnVWrnJwhRTpPIBWcg72xkw3bdRanLuqPm0Vnsi
cVz87R6O+bL5NfwBhIIDfMMpKBA+QDYMfAMRVPLAZmY5ZE52M4CDRqu59G65P9Dqb8MLFrcLUDYo
HMBqAJLb6X7/WDw7ssIwQcCi8Qvg6YqW8JxOkP77LLMfLtbPHTEk4+MT0OAJ4KaFC5PIk+hbyeUl
M5XqK82/q0OXi5cOuLjcOiHFeMCyqpYD5S2cRiqNhfIrvGdIlzDJ9o6BJjI42G5+WLVMCJvT837n
5iWY9u115hW0kuvQfR8bRy50t71ju5bTVqEa0InllOsu0R8dewfeCsXrgpx5O+MdSqLd6+GP0D3d
Czko3rlVvz3O/rskbgLiwjlzv3zYmnQAyzoHvOfu3bPHztVPVy1MjZMkFxn9HtxGhTskYGBLN0d9
EHYDjwoH7jgqSNAjR4QLeRDePXpuXOctsUn/Nm0HQuVCKcn7Hffn1DRIBKFb8rdNGfYDThrALgoX
tDiFdgaJQbY0EBFKM2bTKrrxR6+I9wsk/O2tsUnIjpmr+rNMQfj3DbExtTm/1Fq9tgKxq2UFCECP
r5abpDo6yUfkFEwTsnHjmTxNiqy8CVVEiP4M98QaLIutt9Cw+NG90SeV99ej70+dzWFs6d33JXbU
m/DoOgRICOP5MNToV4gYkil3/GVmmzw+tBqKzttONZg0GklTm6nnRcJ+kVqfPkdHzeqqQOhLQdZA
8dT0bFhglKWMDnof80lN77Q3HaPtqxqo9jAZYTo4fHzDqFWLw3L2hrikNTjKS3gRJ67gBm7GVpla
2VCAgvBC3P5yqDBjX4bhWfZuQxLrABzzsqgY2pdWAS6IGgJ/Dh7jDKXstGGZm6TQt9pY/7L75t4+
EghGHDvSEC035Z3zLf0qQDj6bSnN/RCpX5Ucy0aA3knMsmXJWQpZKmRMIlPd1aiCANjGmv8bOwfT
fAd0zxJ8W7BeEkRiykaEMlajlvvEZd8njyUPtcQLDs459cUjPIMt/qXCfOp64Fr/eklHQJBeecI1
FV3++stp65o8ZhHszl+Gifm7oOIQdSba3GCkr842M95DmkEPR17wcefGxk78qYlfRiAvG9ySP5U9
Z8Nlsajjg/EWSBAUs0IlmBwkN0WoHuL81Qb2JS9LXeP/9kgXGv0vPFhVInL2ilyVMZK/qzDh3w4h
CNahzYesQPIvuYvGwGZ8/jQNbQX19RH+RGJAcRAHhSG2VVxdWtNm/GvCaGTfMPA1U3L+5//4Xnul
OnqTBF2mk9MFeOpRc+0eX/o2MIqUyWdDbeKdVRTiQOQtz1GnnI+wYUsOBUhCtu2NnciLfmu3+AkZ
KgTbahVG4x3rDc7vUyY+mRr8lYs62EH0MGInq45bengO2L2IEAoJNLXtF3boADDSL1NvVZ8VQUfd
wh4iQQyHK2OO6ZAMIvYXL0YYRXmqOhtLEd3PHmnmUsi30KP4hFKKXMOrMTMNvKH73alxg1//AQQP
Ro0HqVDs6FQGdZL3tr8y1Al6UmDShzDmYITpHe4XlwAOvQaTaoYCt7EZLZOxXSET30YUNinXjeXh
YjLnSA9z7Cco7NrOHPigisCSX8VrBA1W+RWVcILd2bhN9X9EooutQhTMmnXRr/qSg3WktV3ZoMg/
Wayuiwx8ekKRkQzVuHxwmCyF+BxHP2fWpI6tIJVbUMMgXrbRG6YHaXNtYPLhVYY4DdLeCgo9Tskg
Ne9vJRXhXdC0gpe+YC9HLM+1IQojhOTvIe4nvog176aDqTfpyveX5VXi+8Pkhkp6E3TAbvvw6YZx
3Fmze6vkZNxNGETpYKJp6qI0bJK6Jb8IcLQchtc4NO3GNY2GgrVlwj5Eft7NWdCXx4310MkdMRS6
ZA92we4gxZ8pgqavWG+YflvA9WYciMx+LS8ctBjjpYoFYfe457ikGL4fj5qHDFU6lmbz8MQQPumw
X6DLl/CwgL+p6B57T+L7wmgDiGH5heXghJMZQ3h7LgVzxYUHtKIYQZdKZibsdGnDtOpXpj8I4SJP
Tpbf15OAWQNm7U5eaLWWguytNsqc0Ju3LfvfE3A4ihZjxP/nae7hHP4lmiywnJs7A4Db7EejBS/G
zQT7OjmdLQ0WExfdqH8SFCAQXzs7DLFFxAcb8IY3ZggnvWTrjzfM+4RI6Mt1EE+pfdGwHOzi+tl8
8j3p3S96Wp0wkUn73aqcYLGZjHSBvf4OobvBkQwq/XP95ba0AI/T4t2K7fPMCA98PqPfwqa1YRrg
zB3Bo2ktf3uFgU9lGHLnHxL0fHrBbgfX+jvbbCkaypZbeU1q4N7xPonbkE82lj8wquSamoKRnGdk
AaajhTbi2sT2ymnmb7smJusMdznuPgtkP9iA+V/AfCh/Pjx3mKyzDJMPoxfSRabvI9ii1fjZzqH9
OyGLu2gZNLuuGwOwHyzLyx6b5kQzJ98XKGUff4x6oMbYyDIPkolc+BIwRWe0qsFORj/M0uYdMRhC
N1Eai28YPXlaC8dQDEkW9ehAF0A6SzxjBwx9U1WvUv33jxEk89gvI4Venv6l8w8/93El9kKGzdwG
PeB+Etg3kq5k9P7WY6E5QXhkz3Jh2xE7wm1PQbsVqhsLPb3HbFCZw69ARiuGSqIFioYPP35zKMr9
TvhHnzEqsg8TIjpWCxbhYsP80Nij3n4jC9e+U9esI6dd2LApBGEP0PvdYDCCB2+N2+QdlixP0AXi
DzU2ag3kuj/NARLhMPUDVtYG87C5LnGfzlqTmYD3PT+NDfrJRAFKHwMAKcf1NPaGp9rOa6xMNmD5
pwzFQfEXuQ1XhJabpZoG/nJ0SETeMznG74KYbyYYWoortMP/QFhtbBvJ0SuFhiQZEPwkVC/c1CaH
03/EcfzXR4tHhH3QgwnPnQbb0XOer7NuVWmcodMOzqChHbQJyKXhnRKf6Frk0snKq1iyuh037tCK
iW0arDgBRapwVXAqTyjuVwf4O1Tz37c/IMTyMnXX8a/fTSf6TYsJdXjV4NFuIXxBFnR9U7tXCy4s
AgfSn4BglQ3YwqYY8PqiXcu/QXxcIPO5hlt6ANFFy6MATiwydh1G4W0IGYpK0aaV87mlasi4VBiW
61LBd06gubFPCNcdgYAS/2/eBd/CTgJQlCWLDcoO9HUhlxAj8/d4NPfD9XeSuHl22oWPt+4Gb3cT
l66PDOYHQX2Sn+E5kV02H/nvN87CFUuIzILmB8oWt4R/Ta0oTii098m3uvnNPjqFP+EXHzJFQf0A
CO4gfNP/yowG9FItJG2+pKe9H4Um3nFj0pdO3aG+iCRhQCeJr4e4NIcYqY2n2i5z08FIKn9hxMSv
ZKw7XNn3ugbhBlEj9gqliHN5/47NSR+iQXjHNfPTJxWYMN4AewuNdHVwL63UH20Arxui1PK5XoXv
BQQExZrf3JTJxtdFs1eExq/eS4VanVNqUkXmwtYeASpMKRSi3g4Gq4mGB0q2WAvydKJYzlTI9K9I
V1/axixag5Uy0oOE2rCwvfVq8OjlqBwxam30sFsZHHkzSeS50ItknD4FaxWM0CZy7VoV6e+Lawii
IzhtCSyZjGiul56v/F641FBn0p6cOBjDnywgctqXs5VQtB/KtqXcdG/sZC6MnWHTYMBHDkSpydoI
7/o7VsdUzFA3kisNHgSDHpumxQhwaw9sTpg3pBWtjFtVbJfglQWnN+9yCDgwGsh7ehp/mAaM7Evf
midCJGDk0CPdrP4MEzxu9wsYuSFNWynC9ckQjwmllnzE3IL/G7dtaFW9a+pLjsYkyz/Glf7aZomP
Js+ZyjWZgJj/H48AGzVHP04df3TsvrFJ75snBCGyUGAJwEM3aKvQtd/coyMS3Qe6lmzIOsMAM7Rd
9TSfkAjnc9Kj/lt59H9L2NIFw64caLgRMiaYEbDUV4T5Atw4Vlpi3t0vmVrsfkvJzleYmF88uwzH
c2kZUJaThLbABoqeEwHfq4ZRVHfbyrTo3cpgBpGSRmWqgm5kaNOwQnDXaNrcTJhzk3fzs0+NQf6R
zmMjcIV6kCiRMijbWmhZICuXxaAZdvBdVWiRFYRqDH567m/sTvv1kfaKB4wooMwbFJwnuFtzaHnS
ITPEFtS8Lr2GA1d4EMzfy2qrpzQzmlnK9zI6PofRDnne5MUg3tx52uMvjCuW/NxrAlYmJwbJWxhY
UgqcNzb5qy2Rq+fl/Iyu43EXWLXoaW/XgpExKv72jDVfQIGh85EZdmK99ZuivsET3XdYsR11mR4V
6REhLQTyPPvTlWoVKpB+m4/uOkxL4Klryepe9Oi9NsU7/nv6gIcXSK0CA+CwshU5ocsJuE9cta/M
7E+lpo8SOI/Nd8i0ZGg/gPVOOjs28ickfIp9F4sA6vgoVeO8qOPqj/3z3wtegYDeuBd5lIZICLgJ
jqLzhLrP4BmVhN3KRrQ3YPVOb13+U8805w0bUgVBBS/qvH3sxm1VKVvhGkrzIaON/817Qrv+izd5
A728FZ3MvMnNjoyTxtniPBpPK4FSURvAa6TU8vbzKt/vlsdipdqF3pfIFnLQ/gO11MdLNRNsPTro
o5adyEKUdZe3QcrVVY7fuBsaQKmmyF/vilri2RNX+NAWjlK9Fstv9B6JaJXK4ccRpG8AGz0gdoRg
qPo+IMEDWNL6QvklEEneLYgXWrefU53nOJwI0UzZntJ/DYoe2yZ4rtQezuC/f8F8T3/hNy9JrAZV
/NHOoKae2pAW8aZBo/LQrHTITup8j4UtXOj3Jp3t1eI8432G8MJh4r58ri6A9tss7hx830xfmjoW
9q2lOIEl/d/oIiRsKj0+Sh+4+nRtPtVxpTt4aQn544CEAC4/GN711cpaIEYN2qeHtLL/tk6IOMtr
xcQp+ELVBT9q1aTXgRHIXn5DreTUeJ4mzBkjFPVf1pIc/6SNA3DmkwBkRb5EHS4HdtORnRJ3694H
VTwNv9C0B2W/G6DHfW3PyRhFtY4yluqRww0o/hsq0KwCoQ7vrX/QquEQboeiNXBFkrraot6Gj41n
rQ5vxDOpEVO1mepJH1ftcYpyU15x43ABvuBaysXfjMz77cmiXUW55X2iIzKlt9ja4Epo0x9I3Puu
ZjMPVwk3vjEz4adbv0Q7rCu1B2mVQ+DUgUoGmDak7BisstH27DRzEqavYIc6wV24rCHxMuuwQg5G
iYAActTTqTmTEetqjD74WJC+2jT77ak0gV+447i1YDuptHSh+4V2H2xtJ2hnzgElhfdJHVlCvLRI
MLOf+za99xAYVyYpeccvxCx5nK7+6SFzaWPBRb4JUkpgRuNXoXkqGnBkPbvKJB4ZZF9HwuitD0fN
PNrWao1eTncJHei0p6SE/vfgy99N6HY4EyrFVdtd7cyHjFT/5YJEFW7cq6LuEa30PnGh/6wjS/0Y
8IQd3TLeiiSkjTaTMupMryVuAB5GB1WkmiZDYs2IHiCaSJnqchJtr6U3p7raNEG9FopHdf0d5n7W
KkEUKVtM5oT43qIPUpNJpbqs78PhqZ+jXPiB4uGQ7BBx7yLH87e1po9g9CWHqY9R5N/8w/xV30Tx
9cxHtw2zBwzhESDTuCfzyoVCwVwhM/JVQfqghAT+jlNGDOy5lsS1LK+QTEWblyf8ujknOH6d81Es
T6FKjhRx+S1sml5dQsvO7cP321+mSVbMKe8Z1dwS+Afq86kOfj7plzcQ7rhhM80IzRasE2wiZMh6
JB+cCOR71zhaZR06PWlehj0YfyFHiP1yAY6unLEXAIUSu6OKK5skEn0r62syqmLcYX+GfmEvqxMu
iK+dcH5QZSqQQPoKXr/asL9OZPDkJOeLJspD9G6WoA48+MZZ/RqTafcjN9ODmHtlgGA3WMnrJafm
Zw8Q8K0u/IrwqVOO+dJlsz7gMsGtbinpbtToTEgr0Lw7Mw732ui2OnXhSstdODqqIjugJ1rQSaAh
CKpTsPyflf2+PGCPs+kgKPm7lXpIiu6XT31FW/VxsYFM4SZuBRB8bIfX9HNRHzwUMASHkmsPLYrk
ZFygeKNW56wx2cpsHUJEAunPmqf6u68HRA8mXHnw81yYQQ/66Cjw6OWZkXMYHtoWPvn/JKDwFXaI
L5+oIdkzLHNE0wZKyIW6Zwd2rqRMQPcbjMeqYwnJjGo3LKPP0IoPx5mHTTbaguNCD8iRWsrPfg7O
qllpYEK09PQpoCD4sZRWAhhUTbsz9rPDntvX7XpUY7alDKALQ3PULgSevZodlcrP6Ia9A9gQJHn1
UhYack4wx74paZkXPPmjc7bkelrIA9mzKq+oeu5NcM/JBlG/TZd0Cc7W3Mq0mCx/lvg0gbzXHwqQ
xZ9QCzPRKKRA3QtcQTUtvjjTSKkXEg2UqQ+gmbUckTPm6AO02QH31LcxmPUB8GNTkLxdZ9BMOpxD
7Ttj2SQT2W0Y+BMqhR5CGnZRSO5onlPDZbd8mqfRrW7nexuPnN5eV2WWjBJL9by9m9gZx0Kt1KF4
IJnaeJt/3LWGYfsU5dpC4IROVNl54Plr/QrIbgnD1usDTBOXo9BFflwWK/rTq60vHtJbMykW3Wah
z6sLflLJrJDOTtPeRrkr5H6E2J1F9WPNXSed0Pf8DohuGtKZqctA0XiPD3roGPTlVYWHRdkCHYet
DlBDs6cizHkOKO6V06arXoyCdHVUeTh9aXz/UVPAJvLQdMgSbSjrSQBcJQNi8f6UR4jx5Dj3lxLK
Moi2Urp18q0BaboXj+zBJU2x3RU5nCFkhAoftuiaMtEPTn0lPbL77wXHF9WZhIfw7MOpBh1lTaml
JmGVu9x/fJKAebh1HbrdC7I9ylCO/HiXLT2zV9aVGvS/p37rY4xiZ1rvz+AI/9HHJSO0YpLKo7Na
QVbeXIeiVbNpNyurhPy/1mqfk38HUne+178X3vx6Uo7Yej6JHc6TkTwne3BBfJBuRxF8l8JmebCr
oY/njaioesTYSWZzu6CcgAiKzIEbI8kQS8lYuJgtTvuR+rIwkwcqOmR7f3mN7gJt9d9lZkbTjKNV
dLmq0dbhVYfCvaqUN/J6g9xC9HhE1AP2zX9jxbArL0QdNpD/a69U62fYe1+7pnWojzhlujdX2aGa
wbQlmJLOD4dEVk1c5JIEIw+uyyXzfgzic4D2WL6l3LnUtMQic89awJ54vspHiwyVoftopUxap15L
L72K0urCXmcRI4HGemT/94bg++2HqtLcVCmb2a9GwH60y9kgm/D9d31+Gf9uoiV8l8naOIOZwCqt
KLF40VddL1YfgEIqpKsCJoi4Dvi7k836O3Ru6q3TraeX1PE3+toCFzs5wrPzh3rYVGCtz3LBp7qU
FITZqdOzJykQVMQQTt7YytXNo9tTHshVkFR0JecPW4LKivIrAlLMq9w6FGJfWOunzC5BrWX6UTMY
WlBOKPlhxg9+X8i9MCZhtFnCOnCwJYaddPbqpyMBnVab6jz5C6G4R+LhaFqNCJMcwkjRBw7i/v3h
3k3QLakVP2S1Y6JIYYwL0kbpJqfnBOuAbw6WcTRgmKunUSMRhaGwG+kAesKk5sKiHKAiCKYtqwTF
Pd0uqnUFhfqCEnrh/dZzKMut4MdFd+gAP/LjT0/nKckrldlrOBMFMm1k12YnQU5z0FpTrUpUvLkG
zTZntBAUyDR624QNLUr8YalBvwCX9ISLUM7x7CerWNP9tsnHSg+udLqIxCbciIrR2xf4teLnmqV0
hwpDdxG78xUatdC/67Wu+7hBVRdCRJvNmLAWA1kUQ109pVjdX2j1jemWHAZZ4vWZ0Qv77iyTEvav
6C+VjUrd0C74EYnHl1AadbAQwzDd4+RfnktKqt6giw6jb5QiMHs+J3TCRr2NZ/qKU0yoj/kPG96i
wx4u83n0tBEeyw72Gm+AScuZRYW/NLDDDQ14ThC2IBBzXD/revxx3i3NrWcSECPDMyF1tRI6Blk+
72mhMdff/JM3HfRk2H4NPEnYt2+kRR5ZDXtnkitR6gIHydYZxAA0X3BOqMK8beldIZQ0OF9iVstD
uOSKCVU6xeVYCKnV3U4euvYo7RHXrKert8hxLvd/Eudt7wKTiZyF0QZ8LTLKa5QzhshvrLQRYadb
PXgtmXRXuSIiMaqotHs4oFQOn3RByLxj/XvYhvi753RgaBDWcjB/B49pbGt1oMSMIFyNRFf8Uxv1
7VYehuEUaQZ8ObiDdcY4mN56i1fHCHs5qGoZu5T+6Cfn0203U3GiPJUCmO4dbYlc8pAkRof7lMWh
Oqnn7lQ7ZgDmmMQahksAHE9lZWKQlJpbvgsuSyjEtL+Al5K4awxPaXTgdie3ULHoCIeWsINbHcIg
6pezq2y3k8g/NKDsCCTOQx8ZGvopRtPTi1+2gozD+efs/kIrH0p6vVLrLuKX3qQvfF6CKADEgm0Y
uB1ly7qoTcrykbLuxsf/GnaKf6IfL8FhcCFWbS3Y8c1jCOy/sJzMhDG8nLeS5JLNUpafmnI28rMT
ydqd5yvOTeZr58nJIattQwboj/8zzvvDtZUCbw0DvvvmiSZvrSQbtPVA530Rt8cyUwoMY4bi/u3i
weSHDZhGg+qg0Gss/HwOcjbCOnf7IYatVRlwkXev2A7W2UiETwCWQapjHgVfD0Un/vpJ3wW0rhkv
SphJKutCYbekJt95HQuVxYVnTcV/Zj1g8m6iZ+J2Z076jhyiXe9KEqKk8g1MXyeBpFSI1iNdZTIU
PjjMx4C6n4QFmQVGVOovGcmGh26ehxoZunRzBHC8EFwBemawY69/rXhiN6hlxsJTakRHX8osPhNm
CQNc2/09XgzkR6nZH8H08EeJGoDmCEWFkqb/R+VNCnT0EmQxKuVIED2V0jjN+uC8Su1YPZ3308at
c7L0mLkqvkd+aA6/9pHNwkX5ZSWY/jOzSpR6vd5X+Fs3mtxq6m9l8uprHSxHGMZ3x2qhTxMXOnTW
L5O6Yc5ybzj4jhYuvNX16bpiu0XYXLtlMV/JYPKKouPjIDaxmZDs7kkwEWogWU0LYGMkduT6WnGB
/N6nKkd06ZNdBhe1Nu7x3y5T+z/LgUFV8H8oyPAAIGjEKbcSb82/2qIp0a5tmuCPzjBI1/+OjvOl
qYvrGjsGSXSk4ma0sBr3emaiQYVlBnwAKzi/ESBa4qIq66V+O8UtVdfYOwUigpYTai14EMqj3Ijv
fIFveT4uOX2JfaT0FqcvdKceHiDjel9q3r/8WLO6l9CYkOCKBxxV28uN1vRwSb1o8/rF4f9ikYON
+rGtlTeCBEdyMo9mkY+GS9G/PM7rTg8UyqlbjlYapzbapTg+VT18hJzbInAZa4Nrh08+yCs4ZQF/
CFpuhclY96rl5tUD3eJhRwjxh5A0U3TG1083iVBLwd3eK//g1r8TxRUfCWL96PN86c0CDnCrGL31
4ZrZcBUFJ03frHY3RAXKgPL/hShYAlKI2UeBcUYvxwgKlhzgrYgUc8owo3LKgAskBNSsCiAyu1kC
HodMvOFuv+c4QMuXv32LVkhCWPbj8AGnJ5hsPq0IothFlbO5A4fkYN+tYWGdwDvWAZbZycSfcTlx
UgnPt4QJvlnQmV4S0UriR5EWltM93P6Yrz3G6y1mWY75WSoqbloQW3VMd8bHphLBscB3bRi6RgZh
Kt/KyBTBRflvZozyXlbBQkwkrrdY5o8dtfI0Yel+FukNVWCzHeU0aEeYP0dvTfC9QaqZwIFxL1g7
lJmABMSNneoEmbVR3+Goh8qfpGq9dWrqi+KKYOPSBGzt+beUM+WbZ1NAFAdTLIDmMUNdGDw/lXfU
sjwrRhU+OeQChxa4LaJOprKLwInwdOMVTwxC9nHPONh3YuiyX4Btl3NDtvLiQdCwNamE/GQJFBm3
JzAA5WsfitLE3IhXD2gRRCIqjktM0JlLGillAT8Yk2EYpR/CPWgvMiGLyZNg2HqbhRASiDSFdK2a
QmwdySpUy10R2puwndPcjSAj20J1zjhO06mQO0nGAd6limVlyB5iz0hVhewF7fKovbY37Rk1oW1u
SOCmiVbsDEXJkQo9NTEOu1HRBh0hCwVnW4dey2dIvQkvbRsfGGXRh6bzX72dFEIwMZoxvfKDi0bT
UBd+APSa/JeVCAfrecSfyDFGZShjlK2xiphhj8z2cP0X4ClBczZyZ25xAKnrBPiua7F3uNrXY3RB
V0zaVp5RRvaDyRTChVxYT77Jv/O7MBlDAPoytGsfonSj16DzaH+9El5drfefmsnqOm56Pg/+H2gY
I9HUogv3e9VD9bbR/bTOwbdnTX2jlz4XVJR2+w+7ak/TJM0QZz6XNq0SC14UEl//MOHZUR5HKqvY
SvBTpj+zIPQr6JVQoiCXIbU4LOBz1/E2gsdhHOp+lYcWDJSVJoyaAy+riBNq9Nn42d3v5KYKU/Wz
LCXfo+Z53YvGnlI0pF0jqYudvMiOhmn3qiRBMCBu1Jj0k1LLI3GrDEeLIU0zNFoYoFkzyCWkGnSd
fCpkE75g596d9MjAk4OOO0xFAmyMjvWjJL+MuzkDw/e+AfDkMdGJ2/XZX/ScFbmTuzC7MWdPTsuX
+dWgOYTTan4Mfu9f4L4cOHwp8Qlb6O72L4so0zyVxgK8oMBtM656pkX4oBPGWiO+30nAZJw9tfr9
y87T9D2x+mzEMCdfO9QizFUinAu3IP6H66C/YM397gRUU0dKTw89oabvJmq2ozEj+/mPiKh6d8Ko
Xb3Rq2ixmsDPCgbsy/1Gmm9a+Ey0+5dduoloGyAzPL3TypI2RE4Lxg/1izMeM/fSTb3Nh2NR9x87
36PULgiQeJaUnNu63mKiW1YZQWIUYCWLKc62ZwejAnV2xRi+Z0zY+nwQvOawMgeS9n9Sdxbd5WP7
oWCMybxBgnI97W0CBfhKBnEgM4jTSQcUgyWPG02Q5ZmwPTjtkjwjsnEpK9IJ6y6XZZ3oRQlNwUnS
hB51e2xzMcG82aQRpJfPpZ1lRF+pWngRR2VtXGirKOq3DyhYtOKeZYTe5Z4uaMaFv70GTnIy6h1X
wkFTODqZ+VO7sYpmBHLpT9tledlZS06o1id/iX61ny0tVmCe2H/vcBOz4UvQmOEnbghJMm+JafEQ
suFX5dsc8xZWzbJVuiTe0Y3eZemulVTOSqDUvkr+5N8YnccbVgz74DFY7E4+VGNFOFR6BgJajEZr
uuOP5aUu0z2ZmgN16ycw2Uz46hW8tZBFKxhVqXa6d9LGl0JQMAaMy0QvfBwvutj4MK4I1iGtSudu
mNuQPivBlV/0w8UWjXAARRPfmwcS8DJZvFUcSXLawvE9Rz0Jje1175LNGpCyvCgF6QgGGwCi1MXu
wYqZv4NM5FPBlz6vd28hPvBrXGQ1Peo3FRTsM/Jt+MGI+Lzq4OCq5UcU1gjiOV3JV9gm+7alfuaV
kaaLACKmfk68iSd3Uz/+TsluyEB8BmgzTtokLF50ml0+wrblct+UoJlvssLd+tLnoOrD4+roCJGL
0F9PaJlowbrCtQI51tdbVjGnIHfsV27k8179TZ0pNjy4a5KDFJbu4LApTPay52xAy2e4EYzKS2DD
JJJOOf54hk5urZXdwXMerHxWzIH8Q5WYET+yGFHwxLTEIJH01qg93hyo6ypIfyxUaDey+Wx0xCd8
wlK0n0Z2s77qdTQieD+bSQBHmTycPhD5Vsa1GyZJh/0gSvXT93Pqgs2YZxi+D/z49HLPpQ3CGAid
fYhE4L4Q2m7UkgA7BZBcmoAE+qBAA4ByC+Pb/o1S2oijLOe098jLuWSExW+Q5gOFPrsb6tcx7mjd
7cxoFaYAczBSxZOWVDCfCN+wvLydkwcymcEhjkJ7MyIk/ajCsNXU9AZjxPSnxmSsH0LrsQb0E4WS
IjZAIsrMM7HTRXixW4tHJGbknlWEP3A89LJaZSGZDJLIKcCUIXEh/ddAhVUJDjXZpDk90VmP9Nuu
V6lF1TVpcglPd0s/eIG6Ts2FX2Op8Srd2w19sCO0WCgjlNmr5EC5PKXdMmV2n7eBn/nG+aTJZHm9
UQt6gOcUeUeAis8Q4myyQYHQAmbFpBiaCXeOSjb75W3PBdL4hytjQxwa3GU72i90fDWQyG77rq0A
Lpa8lbCWpxCrNHpJ/OumsihfIb9VYpT4RDifQ+sFTJIE1r3/odWMWjcIhAX3nQNu80XITxDRKZjw
1F6It/eGYP6xVy2WX6dHB7/27ImhmCuxsH7DXqWrBEjjbwltgSaQ1Q6yje93qy6bQC9YXPSi9QWf
/wIUgpnr+/7TgwjeSMY7HrUSwdCA2RkklVvlq+c5Mc1Ah/BzdDMGe6+oFPWcaO1MlLZGKzGkUrHs
8CUa2pej4Hf5C4QlRbMZFveCN4hGb7plinhHHoFp1yZ0R0+ZjC5jYvBhuWqf1xYMAIn0NNJYI21A
rZq674JScfTpO9V3OtDgsv+RBhGP0g0W5045xZLtpVOe8WAgHcETG2EoAWgqFXIwdVkyQNrWk/G3
8jnXPz3547uavVhINb/YhNBqsGQ7qux6Oa0SovtVNREW9j+KDrL4q6jrv94QIRcr67dqqOXPVLz7
LI6ndt6h71+bH5hCPiZFPgWenqnOWyeyaS+qmJUHrVeVi7Dp7D65lXPxNq09sqHpBWxq/d0Lvlw4
8ZMOr49iWX4IPELv423zwv0Wwks6pfcwfNq1k+cYhmDrfO+II8MEgvUqwOPLqZgTKc+CN+7acjbN
s/fpqYJVdOFCPHTOFrOJ1V26Il8JD4fB41T7Ytsi2izX7ljY9YhzW4R4SGo+gNEzsdWW/c5SnHtm
sTsqmKJfN3mXrqDgeUYc9ns1v2SbEZsyRRA5Ba6Nrna+vKN/B7yyssu+xbLV9j5PyCtwwFHpcfe+
+guRA9CZGaZzIFCUPvWzz3bib6luF9yjsQQZydhsR4ZUzXyl22L7aD7nGgHBv6Yy/Cavq7G5xqPW
M1FopFRj6I8d7aFyo961+Hi4jTa6PyBDzEnDzrcEV7kGf/oQTeZPlCcJ28I00hzW17fh5ehIWoDu
kDHO07cFUXTfwLvaqO7QOz7MfQa2ISJlhFyI5enaKjZLy1moFVchA6Q4j4TtfFY/wczZMn9F4VUj
6HclmNE/ocNakQybsPTNGSV9PijqZna77SXmEtSXEKgFN1CdP4u+c0UbYuyGaMbIJmcC85wbWoSX
2pMXMJZhc+uf5laNlJseP2Dxmy+N/vE/wHa3936bzoIxERsfjDksmFDnoFTKMTWRjsxaJjHULF9F
1nBtN9Lm1SknYYlY1TU5jKnhvKVhjHZKJqAgKYo2IVgfTkjmyRK6Pva4zE7dMP3nrDp6KBx9N6dE
PhvZsme2WTsMGB9f5xqI+pPFinXP9mjaa2wnVaon+AM+H260h9zwgbEhTtnSfZnJVy72ge21ONJ8
sAjWv0IhCHdzesnux8lYhfLkB6H80FcolF6SfqJ/WYgbUTZt1S+TzXE/9+5rcpFm+mMjONHBR6pJ
PdSMX85h/407reLlZTebx0ylXbmr7cytpVUO4p36L8tYW8TDQ9yWE4FlhaS4oxcBe7IFk2s/ttgz
HYDigdJim0ylfZetKD+bQG+5rtwsbzG91GhY0JaQ+ivIUzXtEu2Y7ZSqzADBJje1DicrR5lHDMR/
lnusAi0J7DUUm7Gx10BOliJwXINnDaDbhVdK+PSMG3NKgVEtHBxZOw0G3nlAzKAQG1X5BqBZUTXg
F01mzE2D3rCGTVtc0BxWtxdVLmRCX2TQX4OhwkOAU6R4F0HHKeVHrO40d5wcA39fyEFc/dXRKww1
7EMjWhIT9SlSata2C7N/w08354eUuEYk2dYvNed9Q+brGLscOQREB1INAah28JjSpjmw7kxf0nrl
H4NxIkKAh1TPjD1cV7riKKOv3IPxrMk+XQenMJV6CDlRiMlwynaLvHpjQ8/3W1P72pqphEoBCn2Q
Wu+OQVlKOY5RGjjTuDz4swU93EPgyAA7rSda713Hex/uIlvZI7M3gJZiVrIEiH1KgCV18+lwfbN6
vv2m6Bd9XgW5rFye+Njel1dBtjsDmKyP+/JRjvQOeoByFGaSJIkYj4ITI1RjH9sAfrvK9ttEyz5G
9tWJz2MkQozdzehUN5m9rIUd/1vEp9kn6mZ3BamUI1AIFonbpyo5idqMzmv1oGuvlAy24+4i5LQc
Q0NFRYkv2AADmbxoRT2dENUW5RTRr58rHedNxdyqDc5/sUdheTlnpXfRExlkLC8PwSXYBxQosDqS
HETQomq8W1PEMyOrqnAwbCswe76bviXrf6mAdUjiH/mN3c5w0EabpYDGaPfZiiFRROWR+SeUaUDY
FxPRd9U+SUHxRcOfJAtJwAho+cuj8gP47kSVbXEjmWZA++VvXLlNv5cnBKkodSrBS12HzU5zxgPw
qZXNrg7Vjj1XM9PCkFLHNCy4zApv84ajv0pUgF16jBdZff5OwOkvd602eQAaWSl2nIfWYIr0zuvb
sWgr8J86Mu7CORx27vHxFMbPWwtnhV9HeRfHzpO5KCApzsfRatZ1DZzR761j/sZFvwY63911Gnki
+L5+hKXyxpao2ceCNbrq/NLIzlt9v7rJeCc9FVp9VSxOVzXaFcAnIJnHozLwBBAqtaRrHGc5956e
Ab9VPxqHPeRqfYV3yQh8m0cT+PVExJBaKrDj/W42B27EzEkCHIe876lNDxybsoIYu11RloUjT7+9
IU5affKGCVeRVm5jjd8jqtV2SOB8VbPn8tO/dOcO31Vkx2jXdjLBGdcTEhCYhBtA9EUR+gs/VExA
MWJOg7/M6x+ng+slmYEn6Uz1Xvso7OJwuuQfK+pNrUy8O0NzVbMHrJHc0iWfsIwVg4xcvUDjsYA9
npMUgPB/GPFfs6tGRkuQazu9Ar15QoSAvoBaa34J/McLXNMnBQ2nVlUyNFnPTBrRZ/JyjQgzt1Wa
imWBVAtgEm+3kkpMoeEWa8CQDBck5SDfSg4oySffryPGQnho5A9zeBec4MLhXmuY95zSbqPCDj/q
oml9Qd9OtCer1Ry3ESESZvm1jLhbpynWvAETcRwxEeZXAU/fpyTyinLp0U98quC1jnhMphyV+Pmq
wPc5+ezhJlDP+Ms52Y8n3/sZbhUrEHj9Dmv9ZGSLNS5RJyuryEt7RB+16Zguk2aDGvN5g+9faWga
PwoGmErhDBm6dD0qsl/UKpgDfS2qhBSDMPd9Qqr8vth348PuthRMU0u0Jsw6SOM/xK5Q42U7tWfE
fazbBhcvQ/lDPf8JMGfxhbGSqi13+CreZDuNJApzze8ObVpuE7VKqhw3PCQja5GQooHS3BeN4CKp
MYbbgkFZByANyonEP19EdPuWDOrfOEc03qnZ+SAqE1pcPdSb+3wo7JKtZOXYZCH2c9Q2Dx49lIWJ
PbhQIjUAzsI/dUxVt/sFecZtGSemEI4s7YoAxehjCxBMFyW+WRfz8RsyGxEc1MP5WM41D6Hr7vY2
VMGJRw+lCraAC06KqdAmrXHcgqgsNeZ36VuzTWeEOHBQU8dDRwfcjtDvEb6HQ4nBUeJlT3N7JLhY
WYKfSdq58dCaIH/m3SHQLT79gZeDCORsirKF+GVfkRWi05bipVmS6M0dbC3MzkbiMolZSAgtIaRq
NNFxPSHJQplKrAnPslo6EEnAXV8hblAn3awFOYvbmERYFXKDLGLTB7YujL6lagmWtYQneSdb1aAa
UJ+EseGNYCuBlS2AYB/OXIdoQC5F+GQXHps2YTJZ84BpW1l6Ahu36bNynqczCQc5Sq8NZoR/Gy4y
GGvizKemBJFURGri6Mvg+idfxEdOcU6VZNcFYGaN9xGt+NL9KmdW5pEW/puXBKYaE0ttplIdHAk5
230ZJEfJFmc5pJw26fjs7xkR3tqiPqUO5sZEWghk9QTSWr0i5C0JMGrD0MVlVWehpwwfD03/z4h1
SnBmr0GpKdEABRMokFv6x6AyfN/lbbxatC0zRjAk7JFrnEWlepAZXbYVl1pLdlUzIeg+/sbe8reN
/R77LI3zvHg1M071ccd/r1ZQSfXBmEeE20tlljbW4FN8HEodTfQbJiUjObDT64XJyAGGwdTzkCdj
v4tEMXxjlg3ohHeMZzKK3Sk2g0PQlDOop9LpDlenEmhl+7pSzf9oAy0WWiH4umDPAgNbhYohmQV2
Qq23TD+IuquNXCgnXjOlHwDFTIDHZ2egY3PnSKOB4XU2UBdq60Tg48DUPVYbirse45gGn8FNqQGV
9CJSAbRrMUiKkG6UmQKNFo4gX6nkboc2cZoZsC+1W1ObzGYRzKGNfl/c1buRZD8JSizzasHOe9Eh
gUHFgXOiJaV4fgygsi6Xllb99xDF6x69DSl32FMbScbkMBM5218nWGeBIJZAII26KQSk+TO6zjGz
+kwXtCp4RPepVDIwse6Y/VRNj7LynP3om96g8OBBb+70HDlHmmNrAqlTrYONbaRQ/uNEnFrtyFwc
DEAtj+w+voumRA4Qg5az4/toDiFaXoD8HwrnrfA3kjquK16WZfy5lVjn0DgFR0ksLz8KTdGJ30uP
clbwdO1ngeKGcyhibSrHnfg1QK3UMAptenq2abSqwysizUn/oPaH/xBTZmUCNSZUS8I5IEWJ/br0
k3SrX42YQ4pLgd6Op6oLbWmMH2679nVjz5WGKoM0EOeyUZd9INZyyYKszlCMZtQCRHXMCCQWLOc8
mxWiz6l2dGCK/nYWVJYGz92KxYuEJAKUIaimjjsyXKcqJy1y0qd3xT93wLW+eigItQpoCSM7tyRB
TONtxiX3MxjTjVX4MeUhObe/+nczubAA18KuQnr0Znm0mxfg7OwIgVaHyF1Ee9GqERPaOlpAmPOw
fqElQPH9UrjKTkfcH9zkO1BeHeByezvCDQKjuf6j9lRfzGHsIz6yFdUtsqxI6R2pC3pnlNtEVNJC
obhDEnq0kb93RpseaoP5EV6wEb7h4O2nGV5qrBNQuP3fgn/BJN+c5+hKAYThdZG+D22yTDQAJ7EK
EOCquXd3lBv1EiNzl0E4bPNc1/0D+KlD2tMG5/sakVhQvMTJePElTucruehUfl0OraTuXaO0qSnw
Clt8KaK0hWt66uTZiJrwWiVd1OPvJofCu+E39x5eEKRmZEm9lZC8uhN9hJx+HmTQ9g7sRK5Z202Z
njRAsu9Dnv+g6hyEhhrfqg2JFq2J1AixgPbAtqIdIRsf6pvCQxoPDhz/gAwt/4Rbsj9Yp4LMgd92
Zx6TKnvdX5cJBXmI7dpi+c2YFvwD1QnCoq77d1UEIjIfW5GD0feeOpT4JwCI0bBmGrgc2848TJd3
bqrfj5mw16Uyy4VyHxaKZfx4sukzTowT4w35byfG7y71SYGFSGQrnuTCHzdm0Ko99vw8J/3hfST+
133BeOWMr0YsgyFZaLvm0660KRIy5fuhIww2bzECJWJebLXlJZL/yRwcB9ehXWo0jKwoZnNc4lV5
Z2HfAhI83hkYDlqj8cmcWzfSozM+fcOnwWKDGnC05J4apK9Samkb71LxPNeOBtrumQY95Q17xNJ9
dWhuE+mTz+od8vBg2xxF2myL9tWQ15AXQvCOfJ8AT6N4VDkgHwsurPvcrY4EiCvWZDXsCg/m3f9m
tGHdUDfiIXfhTTdENeKZdHkCMAC6LSlwFK85uECdwUqETzRF1YIFON50RUWPcQiQZP1WoX4Qcc6N
OSiBYi6RvD9CU4p7F38yMofwb3cPz1s2OAjtorxMuhNl1qZRglfgW/4/D/e4kAQju87gSR2xMpZy
NB00ZeNqQYOAz/mchPWdx1XF9WvmcWxD4QtXMTy7qMz5kkk27MChTsbzfnVd7gi9d6HNpD4jyCeg
YmX3dUUYrQRLO2GQD90ABx3AL08QMTa0PNgSvl1SzajrRziLXgSbXf9StWZlm/P+SDIBBSk7emRH
bdyFwYz9M26PypbNM5zR+1pJTcdX9OyBfmtSQFk8zVoLG45N+VIpdi2FdjeXuQMefbmy9x8pemkF
hmXr9aMXzj+d3belW2rlBuzYv4ERQBp0UV9yE4yZtEYGWuKAFHOZAg0SNPcB7GhPLTwCQbpkRMe9
2zrDpHKja9Ewcnj8DBN6NC3pQ5hoe+rziSVNDtN2XbuD6tJYU8iDdRrenuDQ4D+kOaMZaPz3Fe8Y
tSZsBYQifb9YNabvy2wr9OkwwdDD42/6zDyGmYqj8U3YB2P3FsecBz4z/psR7ZYv1FedkvidhQg/
hm10FOsZdyNO7i8EPAwxSthrdMABZppZfOHmkQrnE63MgmMx1RI6nAxFBobcM3LkQ8o6ZoBx07wz
EWEervx5dlZK2Jdw+9bkvf024uwP8lc+ugV5mnG0HnX5vKefadwllkamJmjggnY3Bd7qOkAzXP22
W5jlJDT2EOiyNxDQY1XEX3PV73H3AHIhzI6e/HAqs9BHlJlSsbjFMQf8GqZXgJ2rl9KySyJ62DkB
FMBbQxNFkPH42XbxhfJLh9p+bbgx/G9G+AaocjheVwBNl6QuLAv8u4w2Wt1DJAGkVPgGBUrVPYOO
pmuW1+EzebAEAlZ4nrL2Z3EfaCRqSTekOgZKarYo4G/8PE/0oe7hleiBKoIwuQxpE5vfGd1QrL4S
VvghY8L/DzBY7rIKXdbts/zuuKRrWQ7TLlqHCla6QGOAkT3HTbtbhZrGy/yjEm0E9i1j21Tr6Olt
T3y8bUx68523fHYnrTnU7Du59M2Adl4c47lRiq5g7ZD8LeYlBMQ2HQkd4zFT/IziaibGI2sz/5vV
jxXo2NBuiWSHkUNln7Nn1veJJ3/M8iCafmJKiCeArYWsgqwa/0/vvdrqLsM4J7JAH1mOHHArohV4
DUEXb6BrdmA6tPTJtd48qBJuyqjQb5wimNRWySJGHr4ghk5qvgQasw6FbJlbybwNGKzUfdmpNBKP
zSc1synaHYHvQJAIEBhjIKGTPcQq0hpKE0J2oaxw9AYUeBbKNKeF9MJN0q18Nr1JygRgrg/xlrDZ
asjS2r6s/6sEe5JoNDMI2e3KG9R12WDi5CKCU5COamTQp5ecpx0WdQ6Ht1DtEtXRgBgw0H3cd/oV
dtUwwP7VeFGYEaPiIViyoxq241L4ewmID3eQQqboPRQjn5bMsVLb0z/aCFUMgNJrefXddxhIBIF3
DV5HhgC7htNZFiiCBfJ0Qft65A/WS1RyGgjgoETWd2L+PB3FR+zqMkVpbJGIg6S2YPsa1BncpVEG
ERqXYqO1/1Mpwkjga1suLnqlqDmYYvr1HPKvFFs8puAcpYK+qffElV78xS9MDUMclJNbiVjfWIVV
hUueFdeGYKU3wV0PcMOIYtl96jWa1VjQ0sFvZ0FuwzKwENLW+02DsyiC0w1Y7p7HnmLDfEqomTXR
WpXPeLoWToPmrR9F3lDX0EqbUNgCZuE1EUTwyI1TNpr2absGV+rMxUVJcjm2ralvqMiW6MMVMFJl
a/4V4Od41Z/F/iBFJU6fh5qVFWcq+SLGE14R1KS9ovs5sPTBdiPng93UnXBTXkzaCwcQzgw5YKAB
CxJbmn790bzJXmsHyG2Fj2jR7xSP2nwGqEol/7jsxot+Mt2IqWb0T90dZxnDRdzMw3ApyjEWyJ7O
t8CASk3PJF7s4nbyzQxeWlbWFc6PP/BrxMXuNMEXqNilgINZvTlU1cep6xoOZ3nbLHDdsNZsrifM
56cZFvKvNpB9CsoFNuWSJFpdMIXK7s3pLUimRfRP46gQsRDinFzGlce0xxcO0fRT7gT0lKKCPlHl
AQZH4E53mf5D0yDcp3ZjbH+zK40XBM5F1512nxn6x75Yp9Fs/ooGGBkLjh89gEa6ojDHsY50ZMUE
zY754x9lXZtGRUm9f2N6SD3vtGwKqbktDdCX2d8VzAA19F511sxG6xraQSHg5zcUvMPPVF70gLXB
z5XE9DM0f1GQW/hvOkzJIKvy0TqcQbBHvtHg9hdEr2zu7H5LaEbRZj93QnDVXVeI1cOcwzvOW37g
C8IZNG86D9H8qft9jlA9wVu+1psKb/oWRW/an+6BYD177WFVznr+hCatwLgLoJHaDh/9ul8vAlC4
ukn4JN7pjBQMSVVtK0UWlQL7/qqZgIZt3BKP/uoLJOi1WGxVYNXYca+I/CUhJKpd7oynvajbJJ7g
YOiOMQUcD2te7UM0Pt8CJL2V/MRuAX6fRsg6MnEeQ1sLqqzhFAk1+8hqmcbgaaRDYHU+a1U6Qk3T
PB05zSkmMqpzTGXWWOqKMDL/6nmq+5HubAab0kVzCMVfGJ4LJLRDk04PLccKLf8NXtp0VsY3DhA6
qi0i+VyN0VbJ5RsFoBUiVt87EDumS8w+H/mJ1IQoY/F7tfq0MZvG/KYSEwr4QX7Al74zjRnbTQb+
XQokESDsZFVAakcNet+CVZeeMEv34tdMrsDPrQDSAC6azelibQcEafhr6uEALi7lzitqwlzmbqbm
pjvqzESBl96GIAFk0t7L+Ui6lJwBBCuIGrqCDkfNDvBQ/iaOtyGmhxzyrWHtJRECPNkn1+kuWY8M
L3/I0ePOo/MTmNv2CXR01U8PIT4WdcGcqPLPTf8GB5YmGA9y3S0JceUo8U7X4C1RPBJ1ZSiTTX38
5ahZrpL4ZKu4RdyH/ehXPjbYZroonySQgfh7AbgUa9cCYlNNvsVQRUTvEDkMzX6D7WYwzXBESXK0
wMiudW3oEQu2rtiVeqm9e8LEe9G86Sr4peu7r3K6UoRIgjZHlTdPqGFCTY0u9uYGOEjfL6hWTet9
OvtaZfDiaBPJ37kPCzBzT08gpOji/L/V/xNoPuYZ7akLHV/r1VCizMRGF4/o2YVeZ/FcFNZnI6Qu
5W2o+pK7ib+k5glZbhbF12G7Tze6lTHp1Vysc488wAe8B/lGATOBVdPlBT04/DosoF/U0KSpRf2j
slc25xTpr8dxsC/j3+2UYtMpxsSrhdz9B0s3Aer8pPuuVAMhrZ1nY3NyRnbf/aZIf647g88jSzdK
LYMtPtv6ixlUQfiFsV9GrCZsOMNJkMA9JwhEmob4gwHYvQ1HbbFlXUsGzA/jbtLeMrSFrFgZtbnB
0y1glgkUdAg5oMiKrPmHImbZWGOghiWhyeZV+yK1kbDFhCwH6ltECtgGKbgSt36wGe9es7UKHOJw
xAUf66RyAVpOpvGUU/pWZ9OFIF8fOUoOs6Tl3Ol09rkn6q3SIbWnmKP5WZ5FEDROsaVmcWEOethR
YO81qXUrWcJ32jmZ4Hf7aECZHz/BSyzYv27JiaMbb3gJNulx1xps9NTgCH4akQ/STFuPXyNxo8Ww
qVSKV/ig6DEyNsXWCDLRl4Mn+JUECTOCuHuoqRGMj8slAgfUGbs3j1apa60Qx4ONbgj2/9y0cjso
+/cNJOleo/IYP9H1b9ThBofot0BJSeL/OAkvyRtPHFzjNFehBtdV5dX+GuA8bvmL76DOQnGi9SVR
cmYLHAa52D4KMGVOgBsEh5CekY81I+qexrCzF5j6rB1zknwrufkhpKH5ae35aHdGPCfuODsO7gQI
+nYQJA/mMpqet29ueo3YrfC2TjS/9VyVcqMezDPl2ArBfEc2/1crxCH0wPMTg4gx5D7xSmlk8K6n
5AfAD0vcHF/cxA2genDkc98zkarAvZDHsLMMHJTpS+ailyHFJZ5XRzQK+RV5O6WTgvB7ag7/froC
tRuWyKhOZ1Ogflvl+nTaHCbu/4AsG9SkMjS19ybWaCpA/uLkeDdP+nEUuEdtWe+d0nFCPaGGKkgc
mNhoMFFTh8Plypa1/iUPQY6UFzuzC/dmEQKCosy7fuxW6NVhsn77DIqfYQkY64pPWjM5/SFYL8Ej
+Ao3Do8JRDGd2pPMXJzLBZ6uy2BYzHmVO/Y5bQNCt4sqtg7lx1FD9dpgPoxQTN6kkBpY3F0Fqq84
yxlIiVt1S1kCB61TsJ/JNZYjdvF2DEMgeHegt1SwCxYloMfJESDJzSTnmm9kxUpNKB96ARfgbO61
pjidHm75fY9b0NAaleUXttwP94mAaGdKRXj44Q+ewsv9K0aXq+OvB3QDpf26nprmN//wCf9tNFVU
anzplvU5EhsGNDgtwKDQid5qQqjcvNC1LCo6cAwtbkg40z7iyRwo6mQ8bx5g9rk4PBoqlNKLy7+T
JWx9MLTqK8JJUBVE1bb8YxpiFMEPqDgb1zztiY0AqWjZD4wfWT3CJDXx55O1IoIdaB1H+rL85k8P
KFY5YbKLzCZ+Fff9zHogTLuYRJ7lhEIOKd5n7i4U45WWclqKZUHdKFQx2KSXuEmACkUoRenV6/vk
K8Y1uXPFtPad3zNbFeqkoKjoC8m9bTZ2jglv3Knq+F8XrikCa9yEllMZcHuaaPzPl2WXPgbyrOah
24U4SXwT5r1sR97z9pNEbKkMcYnW7UFmBvrYrh0EORcFKfkiD0QJCGJ7ysbAEANULP+2W9Bo3sK5
5r9qyPhyM1bYtQpGQrhpyQyydAWOK6vTezDQLYmErH3p/22zWhYH4qcn3XixFZMRAa55PLYQM4AO
bSJRhEWndgDcnafZ22Y92nESIVqUe8ZA3bFcsb9Bu1sUIxcAc9OsOcg9L7/PDrPISeY8EoZ8Ox0v
gpq2WMQpjaw3xdqRr4E++OTdu7GuMtaNMUX3jw+m2ALK5LUZ4pzWWgt+eQymWs8rlFvQFK8fsr1f
9e0ekeVgsQP9ECCoctEQqH1CgSsVjFGsi6hyAFag81FizXwy583n2NDH3Bv3y+LhIpk9cStkBScf
f7Tvrz/RXmOZJkxbK0ZXr3Uygia03zGZU2n88gg5EJdUdVOge5+OJDR8lZqzO85046gjmoS3lbYv
tTLygHD/sTBZSnSno9kbq4xGT1fRpoJ0zsgfeyRS434OZ43G2lMUXe4yY5+wF+9QRUm/i2mWLkD/
aX9YeT0ZDuIs4ssXv54mI9C5REnxmH7jbrdVO8ps1CduCczHFt341+lCwwTQM28iUWwtU0yyQwZl
znEpvyfUEDRFbGOzLa/+LP5uNpqaMIYYhHGUgevgZ8hODf6xZadr2D8ZznHDxlfnEnHtVXxLLbug
qlz2YZtn6x5dFNPRa9kiGDENZZXtFNYLYigDTO9jH2F4yOz2Pi6JuQI3WV7hhY9AM+nKcW40nAcW
VjqusNx8r6kTi1UYgoEj7w9PbiJz491FJMG4abqQFrGVdCwM+jv2zbSwaQH3b8NCh3tiqim8gMhj
9SBCA14Uqt0UN5cYthmSLBGhaYZ/Vl/tHTsQY2TaFJhOvJA2j3L2uCcTFBs0jKDF0PfEEJuSIBTv
PG1rLVnZfJJbV+mtmva5bHl/rW6hhQ2ufjBGFpul2BUC0pM9U1xDhqt03r/VvX49Sx2tk08k5Br7
VfSvYdAr4AuwYwvkv3mC9/0Fd8qP6IFSjtTaithFiHCyzPiq2Er03ImQMulcm314bNE9iHvSqBuw
+Nj7W1tu2LBbKFzebC3wx7OmKrS8xAPOuPT4mfirkDnlyaYDXRtjTSO6Y3ACBTaD+ud/pOCSAzvC
nUEeRdRjFMQlgjXsZObeFJrHT8yoRDtqfauyTcG6uSXPGXuNg594xmBnOtM6p2UJ5ipAp8G+4YzU
zS1BrH0BwhRyp9glzzpeaQviVi4+WmASaEkW2khT2Bt+qyGESaf1H9b1VLPUEsX0lJJvkyv7M5mM
+xikHEDfKN9i502+TgXGTobW2gG9SoukeZRjK0XPDPZ+PvWScBqohCZspNBMmPlXmlNrosjuIKl4
ETacJyEal0FSP1YoHfcx1IVS5VYgD0qH9TsjP4tHeSsALNaQsDC7oH3d7eeGWk9N6a7rUvs0khj2
befIe/06hPyPZZS+V1mmf3Za72chuxodIK7TaHCgYEW9j0jDsND4FfAw3bdbawvapVsw3fyY3hL+
CG1x1va+rAGLnJnU5UPjRXYW1iCP/UfIFKyztDzxnTWNKFsMRkNNPcAr+c29xDEz1IA90sRO4QZI
gygbT/HC5Uc/M3+aUw5QxDYLW9L+Wlcw83jdrSs8vq8eTIgFFMzvb/aIQhsfpgxGgV3Wgi3++GV8
VqUv/wujxcexjF68tRq/pYhGOHt/gnL/ASEzz3PKBFLHmES7NgBdlnwA28iF3+sIY59nZGq7DSYA
v3LuYFlrzPtnVjeHT6KTHhx7c63Q0GVK1WT15z3OF5vkSSe5UrOX+0Z1tbZCyJK6UTzqf/vbdTT/
GXvuX2NyN8rU7s9/elW/vrgmFOkjXZuAQtscy/nHt/88q6s2h3BFw1uw9Fy2ki83ySulAt2B2oOk
0SnqC5nzIf7dx1UKya9JMf2B57N8OMurgsNWkP4a6HlaChuB/Z2k2S8FrfNkc2LoILIbeGR6BX1W
4e0XsI985JBcWgL24tqlKDCH7gJjv4ilSdrneVofsJdZUwduIM81ew9iaCsJixLn/OhlGqsymPBm
BTbuNUz56zPuR8Q7bxnMgYII35Syop6YVkN9ZoiDW8IwJOfbpOdo1dTSjI5ZhihzTXhEAhofsIso
HflqL66d7ksAj/m8+m2P9RQ68U3RavWM0u4F3VLGB42+dg+r/uZYjpJwXRir/y9fgvP2hgHk2EZc
lHWVH2WOwvD3aZETZvNQeP6M4ImNU8qaZKWkXMt7U/hyD4IZZdp8kaATtn2NfIs89tPYmKMhPK1P
yOHNyx+yP4zQkK1QMiAykR6jhD/bPVuMf3YJSoX4XPDkfjvojgq3hTLf1cv7dkSbUKvCybVMP1c0
aGG9o7tecEEA/SFI2iN3BSGbzfdWqBuPTcU/081RlbLKtzicRfGwzWXRioexBbKmYWY+cIh8Vyxl
O1Qi1e/BkPN09XZ7FjJ4VcSIF/pZalk7nIkkgqkioQ/HeY6949zYoT6uoO10RfrpuG4vLf3obGdn
ZlYVLnHs2X5hW8Fcf9B1jmEyjiAvhpXPm9uy+fGIvlbHGVrQcUCc+0W5ykVHE6emQuOD1uML6sTD
9mNNw2ff6qSIARoxZ2qoxRqf0GQsAUL3qeU3QlAf5OxpE8vYPG3u3JloRKkB+QQ9DCcXUf22mMJS
o72v4PlvXxckfJOz19LzBae93A2huNeGMUI9V0d8p1uNlRuTRE/lkxeDfI0LB8AhlXImhl4L9rj/
DTHAqYiygfHi80IvAhh/DyUGZMriYCkoLHq2AG9gRlS2UU5kQ19MI7h2yA6+IUFBRnEAllMG6slW
g/A1Bd0qvmKmndrbnqvDTLbRnabk6nxfOy5vSNY16+DlS7kaukx9x/3hiUtUW0mi1WlHX+zskKBg
eMSugu4+cY76aabgJ3vPTm4uNBNWot2CsDTjerPBrhu8oENa9OVMYmHPz+7DyjrkQklUN1SyyzSV
6bYuC0XFtr5zmrFX4HKl8ZandwYtBPyWrkdLtQ1xcxOorZ1as58UtET18oe4pKYWU6DmDWAjwtZs
65jiDBOyoGvMMYGkZo7Af5HeXAByHsux64HhLeJLqfu4EWwWrwm1ezt/FOZdWUSEJbBxfQqQ7UQl
uMyc174NYwgt6j3q+XQe4Jsolwk9yPH62OhPieDtisn7jGfl14bxU7OyCzNdlIzqbF9lYBHQz5eF
Y9+/dUyDVYW9h6XVW740nj86EVNwkDl0RvwUt4xR72HWRGo+u+tdZmRmNu+0jup+6CZqJMYDYjFy
LNKl6nTIEJaeVvhKMy8ns4prgP7PW2WI4B1r9L8pAW7weWwxXdt3Q+e1c3x6g5ePruAvPzzHSRME
25vOhHTTvX+IwFOa9rmeTGxjnigs5im+e07AZ80WguiMQ6eEUXyWAgVvWS+qEK+f0nLyGeElajQp
zpqJfDgc81/6rPE+bP+sqT2FPhNFygKMIiT4BxftGonD+I0mM5vR13D9qFRHX3Z5nNQcnrPVgC/V
v8vpeijusmBKlIesP7z20elJoV2O1J8nkbTahToQtlck4xBH1ksjCmv8764tx+59De1Cryeo1LgN
0vyxUt3niWQ9Eh7md2TtkzcpNPKkW5qb62OSeXigZ59M6nJKf4wBoRxKIa7B5FXt5YKgq15AEpJh
qTTx7rc91xN6mWMeSHcC397sgg6tcTISqFWq5F6aggCMnbWCB+eAH2MsIcO7gFtnsONKyjDCpsAr
f624IpCtIYXaTUM0sV9dWKqUlb2+GYpcTR0qzyhYzpkV2C63az8tGpL9eaKK+pfuwBOxJbP475K8
pRgWh6DyIZMWgs8uOG0gblw3Ak5oWQehJDznMIcnDCI+xwQXYQ2+1ufE/ZpeCnlzVGF2wNK3RLN0
wF5G8+tdm8H7aOfTZFXaHqMVSEGeW1mUSX/ABlxS+W/dTBUvkFSgBgmjljnUaOvEQGWmSb5feBzv
FQf4HJz2npLLsv+vU7r+S8YHM5ysaPHFioDA1ldwoq23ozQ7bzoDmKXSUZMODecsXTtIsh8+mAOd
cwZ6L/smHnp5hwair+a8y0mmW39ga91OwO2TYBsKZ399qJBW5erS7MX5kD3jROcNPaHNvAHn8ypT
occd+xl4TsL1zeZgk2QDyi24Q5fXFvM6kc+G9Tri+2EK7ltNgOD7bgzQ2pcSbbv+mCNhFnHo2G3u
+Lf194sjW25cZJfYofv2tMT18oUZnAH3OQKjIRzbDN6jTtUvEoO7yl5DzvVKl3hUao55XIjlrOnJ
YRrkJLywGVqEoDJC21r6pm/CxHz/wapVP9DjwSEPsDztvCtb1aMhHVqbm5xH0STRmhtYRnixvECq
Aev78ic0zZ1gflgQ9kq9WLg1SSahcZJiyxjuKjvJP3Ka2M2FXw20dVYBBlwOGT6BJc6IxQt+IpN/
poTowuqVi1iK4sAmD76YrkYUq273Cnb1U0xnmDYNxn7Bd0jus86ychbHQDCVRddmG1+BBKpet7IN
ybqesDB6YpARzzrDs3OKg704xWs1TRKBB0671Oaxbc45eT0S1hSdnnbH9552anfxST2hy399XZ9A
nGXfoZOK5L+RoixK6nhRHvgHh2wkcoQ2JaIVWDGyhMCDxZKtpYzmUPu1V7OZmnEDy+oRxRiTW8Ni
ckRjvo19BexLmjgJXVWxMC1QCZav24Cz2id1KL58H6NLkRmv+eq2V3IuknnewLMJF6Vy4HktpY5S
kEqcMdVILaAIVx9rM0VwkePlXfUzQEB454tipauMt++159Ubxw3J8fWAwQupD3ggkdQ6DLpFZarW
m7qYVdVsge0ZENzIau+cNVFhDzhzKLGwp4KX0rQ/YMbah8Nj3MnPaV4ej1ZyTD5pP+UZKrfqPPog
jX8W/6OTNP/joUZJZxOe74YLD74S3W3uRWChIttY92NWSNJ//Hs5Gj0oKriXWPB3vBUvGxUPx1et
6YMDEYdIKXHC9rCfHOo68hKO0CKQcTqcp2kByK2cHJdmrbGeFrat284AWOVM0CvHavyVCjNyu7zl
YI9Pmmp6uv1qUmq4x7pL/to/OCZxBS+6ngvKZp053lrV6hz1N91LvQL8uIzVw2brydcHTltpJF87
Od51mucdC7oT4l0GUQjpfMSKS4/7q/vuTmVZRQrBauUixa2cjlZ/E5orLP2mzJg/gKOmXPyxSUh9
tHiCsxKgcEnf+MQJXxNeeMvBkhdAo5usGfvGGrCkWANE6tbysVsmz0vP3vbw6tWw2EmV74Ma8A1p
3MbrTB4Jui8VyRssVdA2IOC7MXmkCtxj8VkgTl4cLQX7JKUJDY0RwVvv9K/jhKGKw+KOopaf0d7O
uzzN+9kPkkIltkRvQutaNzyVmvNtbepCFfuM6LYggbWBSyn4E6kGbjJapLvy76rlbIrlkwI/FCkT
FUz2j0QEK+8N3D/kcpy/ZOxyRMIJSlyMtV/6djE/m8BNLpU+qtBynI8B2RR13cfJF4MxkCQaB94Z
iKzggtqozt/Cz6OKrVo4bak5twuS+eZE3fQ1g48ZQEZr8RMoKtA+wWf1s6lDZq6XZ2IpPdVJxzU7
i4EZrOLYTu5zY9ZSvXD/0jX28Wq5mz2r7xP8pkGKG6cXqS/VOLiasfvFJlHFx51mfERUfaLOEzog
tTFwiFxc96Sjpt7R0scsxsYC8zmShk1PbL1HcZZwmsmVUIbXwmCut8bZQz5PG9bwOL3vXLQUTRVd
xNzKCUMs4/hHbf5ETuuWI0+9EDOsY8I8na37jz7cC4o7CfFzGsqatweaiPWu5qRyGXipPA0ZYESm
1f5s+lOCs2ttxbA8YluUt+vrVdW08x42xMb9fXgYqLOMyQ1fbC2Xy/KOF7z/Vk7cNpX1DMGKvLev
EMpJleNKUQKdt+Eo+mvfYE1/RiBz2iCV4b4X+8x5W27J+3oNiS2ND7BugKwPOPrBdDgnQoPVZSMj
xx4kGDAAmonRI2Pe64Vm/04Ln0z0ZmZGGnCmQcQPllyPobVXV71MftTzV+KruvUyx/bth2EL1ZGq
0s7P7P8lBeoc0/GsFVjZFJbQOJaTSfjZgve1gn1Sxna1fbj9LlHcI690bQ57n1I223GAFi+3F6oX
WdDJiGJRynKlOSOUnid1idY/jxvN8JVvBvtsfZ4egaAn+PHOamXZBGA2wVMfias96cTc4vhJ1HTu
SP4j7cwJNmgqQmxZoljF1Rw/sH8LUC45+dlIbXRNuaLZf4OFOYzqLuNAN85HJIH0fyq3AFm56+sx
0r0R0P8+VLZRl4dJlXVwQhrdMTMhVgDrflxqizTh40fej2ddlh3hCpWura7lBFKqzEsDNSJ4TJGH
U/a7OwKXIcOx4HKE1Yc15VS+sGERKm5QrRAvA9apk0RGUOrWpqJ0YXK3R4f3z93V4yorioGoWRck
h80dfdGUKq06CEo1eu95WBKmPxrun6CofpnvT5+sVv9zxllVc22VWIveDtwZXzYUFSkcdaU7PULW
4VfQ2uMoI9Q1IcT9RlGgIdR59Qwf/3hJkCsnG6tvrJM6FKM7DhUQdKev1P6O++80My3VCBA7md1H
17pEJJzHOpmpmjc5IZW8+RHXLo/OL4C7vtEy5CRWHgtowHgHsabtM4jDsAoDWU6P006KNuueHcaY
IJuV3ji2JySjI35I/RxbFoJZbKqa5UqQ+c330pYp7NiwaQwm8qNcJeyn3qXaPBrcqSF3zxLzPNqn
ZPV6+lWhN3VRqwroYg+hYqLlc9DMU0uXDjEklD4Kl0FH4/HGg7FjJzpDeErhpoJ1fMYchxy7jZot
DPkfGlzpTC9O44/0oCUugze/eN74X6ZgWStAjdo4l+ZJ1E0ahrxLQ5DHPqIZZkmmuN+clY5N1YYp
qp6z3ZqIeOnlf7G7IYifK9lH1ZUBxyHz5EAs9TuNJsqvnmXUehvzNp6y4/11uiPMAxblEwqAypw7
aNT+8aPoJocuieQSk5Ii0GcKNlJnW0qOxvDX/PFdRP+JY+fOEtCIJAFP/6Iye1dD6kzmlfEf6DWq
MIqmhlgMM3tw0Ri46+N0SJwCEGteHIX9NJ/47Bqy7u8qzIlkzKxBeMh+lAqpnrljWJLlkb3FOcaY
tGRYlYM+ELEY0glPG7aPq4Zj/RyhD6wIcPkkob3e7vE3CpcWmjP5FEJo2CBV2UVF6wGpIpIGLPu2
BB0AGmIGQIt1WdG2Wws4ach2kHb8RtAYHOloRw+Psk7PWkcATyOEDQ75VyscQtMYRjwnRafJo2Rf
JlSEgSSWX6iHtCxA8P7pzljpHulKOdxV7WYK2lsR+/OnZ6/SABItb2vpRf65X78UUI8K/awmGKK8
19w4d5iuDBhnx6gcXKa92iqcnslSvGs6SUSAHUAe/Isz6PA59/3wFkMdJs0DJJWQIRQszMWLN67q
Y8Nn0WjOICZJh6iu2fTnqeS8hXHcU+J8B2tK5neVFWW4M/1N3o+Pz/QqOEwB2nylrMtoCnZFfTzN
PMq6Vn6gB7mlSPslWjYMylyFxu1zPrnGj+Ek2GrWXVefHXER8gDkeY/h/elKdyp14wlVaUnAMWOV
NFeL01p6ivG0TYOZjjZ+rasgO4xIjbq1I64bH6W9Mlw19ke5IWeU5Xd0ACt8jsxABGb55Ufy9TNM
IBdPSlm/vxDOMWwfuO/X9JuRaaecYueVSqugg6FO05hnDoE1f34JIdxGjFmZMKGkxoORLs/XwNFq
gkiYlWq9cZAhiURR8yopgKHMB5Km7/Gv8BMzUrGFWVVWKxMuUazbb6csxvnS5Q/NGpGu5kX0SHhd
Mydow/uLVP3DcRpjzFvftdAWRmRAL1x6B/Fc9AVErx6okcuyRLy0nLkqQzfIPgjMImlyI3UUb/1x
bEYTDdPD3198wfw3LVNdci43REEbMxyStXTPAH581Cv7IHemcmN8JFesxIBzowTiPKTlNgXRCbCr
l2HtB06kXuDn2F/DuNpF0BbT6hlLeykfjqn3BsX2IabZJd5ucQUBGQjU4y1GllT3aWmV7HeLCeZv
mBQnnn2CYyGvEE8CTctbUlhWNqWUIojuxcB3cC9LI34w7q+0+nLQxlewDkMiEmVRpgQZZcCLpkgd
lFiv980s0A/H8C8QJZjzl0VFXLHyf7INj5pljkdthyUCSPmYwz3McnlMxLLRmuiBp6flQ/akBOLT
mDVZKndOiIHQFOAnsquFKtJiuv30gt5CaUEtDcgcaVj9QPwggLVvlcbY0cthwZACMLhk4086TLbK
OC5rK+BzUY7PIM94DwMi9mcB6q3cc80p0fqM1hnjECkEoET+Zt9kEEw0T7zjc90JsHxjg8FfkCPz
ts5VB4sAlKSVc4JunT2KVL/6UJLwlDmdkZDI0MxrroswSz+3zm9sP5CR48yAr4+1iwrmAPLbsIjM
DRBXyzhbkQI/ucTtZh2fs4/vNM2gb/X8wJe1AUJf4XmsNqaeiaU/rHJ6vTi1j0SvM3CLrZyyvQbA
46pPUur40OHlJWSwQirM/to0jzXT/akGHCzXwLEfQWVALA7p2yNEvZVzRpQyobc2gwIYa930OxhK
UvREtJuFbn3GnJEsRrqFR+UniJgs5UIKhsVkNdm9VHHoI7DoMnbRiO7ap9KYczNEoo/BoK6STaui
tcNEGFojYDc5AXisrCUfjVO3K+cEHYhJtB03q+uqsH8EEmVwtTT6IYpA5hfp6oGB+dQaWHATkm/h
IUNkq4PFbywzVMo6lWdr9CB3Qil/JVFEC12UC5E2fc2hwTpGvTgL874SVd+McSaQGuiIu41E7Jh0
R1wL/saalbjygve6oYRYX/VZQl6Ms99jzor8jxYaCjVg76EKNgRf9BhbJlaYhPMqYRTV78z+UDLx
IEBDWVfx0it/QPXAlNdqPgcE5p4cffYx/1XQqLA0W58nH6FAb7i31Uz0LphmFqCWMGvRtrYOwftN
WMxi0zBXeiFpxV42+I7AcuU4yDDnYqXUsDAhDYSLwdsP1saYYUSizDaVLv5ZQJ4sg00yPQCatxil
bfa+GPYr+2FB64Y1/BTjYXzTkwbipHdkE65hXIBJHOW2Q9MUlZBNDkr2F5ehU9V6iORA11ybp747
41NVHNN+wOHfbTcXVJ8YClHfLEV/yKEjvk5Aa51bqMCWo+IQhX+CHJtVR0oNPC9eSZzlcF+LMKPj
bRjdvjozc18wpdwpbNZn7vNXIntEw+6q5yokkCEXok5PzaQ7lGAIJFnmxajrHyNbpI2xelvM6+Jm
y0aH3U4wYrHUuSMgR8oz321sBIxWASpaSe0m4LKeiVMHzo9OYh6fMi7lLlCmb5F8edlYFnmub1Hw
yJEHMHQEJvrY3HGCbqTauVlbnRDy3AxAWcYvRcdkne2iSQ7IuTDBgEibft/nPkCWIBUhsyo/vizi
wHmn9+JFyReH0Gdo/jaTwGjtw6W/LN2eSJtOvX7KqoAdf1IfN4hPet/zUvO3oApLTffoqeOlajwe
KldqSFp7dOyOqBY54ywRR9nbjFcHx9NbVr/1yPXG6iYVbbs21+i4O1Af/e/v7neWa3F3gYWaaX8O
di+QdaoqDcTEKbmH0ACPXtxfHxNIdnWXxfE4wC5Fa2P1YtdFDItANgYgbTo/R8OMX1AWHwB62Oxc
Laz+DEX9EDyfOpnRKEmh4T6o0TttNVXjZEtJRfFYfibVYDOrK5eAP6+vAQ4rfbs7C2AolKc0I1Ns
xU6EEhHeazMZakphXI1RmWa8RY9EHc2bKVaF7/h4dHISTZqSiY1ibHmhMOSA/2IP2hxOv1tWI6NJ
p2R+MmD78++JXxjlRasArtlR4gZ8RWM6qnLImNdxiJ5DBj+hnKjoo1sGI5NsjnDUYPtN9XBAa3OA
7aau46ntDblleUdQNgNfnfX3Bc0na1w6EngBwOoMtVzdRofc7HrlYPJnDZBBL6eeFUE6HmwNPBvU
mVXD/x3m5rnVn96S6X74Wqzew+dhrS3gksG7apT2u/Hs3ln6Ke3YgDS7RrBYA5/5VEKCrwFFjn6Y
A+DIheU3BkJskGWyxBSwYWHaNT3SFLyDdo+zzVdybqJa1I7rdv3HSxnB33tDUiekWQuYWDyxYSUQ
N4vKI8alO/BAYU7d0O3icqKkdxgwR7oyqM+2lQVta/nx4ibIAgy9J9UbuGP8ch00hxrJ0N8VZfG8
Wi3HPL6I3MyfOJ5bllqHQISbpOi9xLyPZX9O3UApHt9aDzGJjoRbDcfAaOS8QWffWTsD15eMitQ1
wzLBchJltOfYkhJXhuJJpNeKKy456JnrHFNpDz+9DzscmIDuujILZO/YdpGiAZ9N4l+ph6soJaOp
yC2XMFiD3C78s+B/0Oed80Ln79pQcS5DgeHEZQu4WHmZARtfsDypzQ/R5qZBfklQdUNy93bHoVjk
TAPHNwJfYJXMSwABzIM4EQpXqGEV7QsrKYmRaxv55Uxqq0MQqizfLDKX29sHjC+lEAF1Qj6rnvsd
TITHrBNwZ+Yoh+6YUGHABQhn3rFNledmu3gMyA/EUhi6I6R4s0AOQk0zTlxGCbqKZHyC2sJuJHhW
t6lsUGUoo9PHZxZ0jitakE3r5BrxfenasSQbBBBmOHG7CqJGhY0F/FmpwJrFtame34Rro9FXhcHy
MHy8Rug/wIR0+rEQ5p4zFEk672nftgv1UN12P+mhxIskE3tldR6kAEHu0bi0sCEKEytkgpnXQKMh
20gKqXzwRSJKzPq5PuyLGnxl7hzbxXp9XDl3Ny/G9qWsBFLJkj0TG2wBFWxRtHB7kVgdsaYmViPr
a+oLXIrWHgBXryoKLzwQB+ScfdGb1gwUdHk7OfITDiIRkTbum82I3y7LOAE6y3fNM/x8+MO147yg
BvKBuSD4xxuvX5v70OeGR3Gvv99ODnw5U8snNNQUuzDihGBh/rV+QJRmj3lNCeyD9Nvj2tjTSgVn
UGW7TNq+zZJuQ6In3OSsnMg2y8o+iNhh7Du+oEGh5I/dbeQGhmi0mG8XwjCInCskY6PKqdVD7obQ
0Gm6eExkN7bbRnsP6/W9GteS0tmpLD57CzS88GeuzStTWmuHdbUkJxn67YaHGBw4h7X09vOB5psS
332OLn80biqICTKAFpSa+0aytRo3zz25ajXsSIOPuWvJVl02YB7uG6lLZUsVatVbjto3B1Celezq
FqrkGJxS0t4PWzJQkOjt9m6B19lDVkIChAckbT3VtH8aoDIj6DFjugLhHW6i+gMYe4QGV9UUafCs
4INMypf9WSss+LkGW6Ws/OpjtpkrWB2L00YXy8LNhA72cfyd7Wk/GK7c+0Khb6TpSqhDVhGUzGmW
5VnMCyNv5afDflOhi3eEv8mxDEaZqpbn55te9RH967ljehyJXHWs4cMSrLv2bAS778ti9TNnKigS
fRT9Et2La4CqfKQFKH9yCuYjqhteingvbx8VPHmxl5PEP/OnB1UV2HxWGseQ/KG6+znkyyyPps1T
UB344ljbDwR/oiIqfkfCFYwIXF1XR4P0cTVcaaRy+sTUbNTatdx3XZ7ffmmtggVFRTIdvGHP7wHc
zS5oVncaNKRKhOgv36UTkp+8deQBDolurFAbBJarhQ6LRhTwfE494xcn6ibkigex/ewialG+Nsp1
AUcJd2udhdGf+YVI6GAK/oG5BrceyXCDLjGCBwFCyUlBYoJZX+cZfPbtjUD7lzxUE99h/wmercSi
KoWu2yAnyaTjNbTi+ugdAvgahzAF4vuYtsj4VUxwBR6EsUJyoGIlWM3YGlNdTGnTx8/V8sGQe+LU
2E9QMqQPoo9clF0D7KtabfdmfLJY8pW2v6TMX3poQ6KE4hsKH54VDNHwfwrnoB3+/Wg4NnAZ80CO
q/OT5wQJy8xqD18EDWpAgWqXGRzmxfGO7uPj+Y0fcLwzCtCuNrJtSjXcPn50A5slWWXqm+JozIvj
rOy7jymFndSLJ1/+8KIzLdl7L19W8tmKeu06ZUp+Yid6ZTv6vNevAHbat/jWSOSXWYL8W1bKxbI5
/nDJ3NLiD5Zhancj78QPCQF1vbadpWhnS33KKN8sfUKQtxT7KzbAhSNw7KyHBULcXnwwUmcWHDxR
h5Fh6+inyNFyPdAkTY4h5dcwYTBY42doY8OE0HC1Jv2MWhskp72/qIFjnYhzfsV0ZTLdyPdS1jCa
g/awG/oRHI4/SxckYUY+qNOpFLGDFKJmkKYbqTtacriQVqkd86nAAE5E9JwnSOEDI7fcp66HEcx7
uHz7GG7xeeu/Xmg4+Yotu9borLHq1cD8+/QmDPr3qg0DvySpLCiDCXfEVIXJRB2KKRJJ+XpRZYLh
aFeeHBwPmfkbnn/MW/DYIYgCfWdATv0JyGbkqT1elyFvI52fNu6p7kNBdmzS0xED02yuEvJUGjjd
6cgkx9aTRavV89Jeuqcc9MRKwj/9Rl5jj3fIKsSOUI6ZDCKwNayWcsyO0LHq03BG0fL/Emj6zmec
uURw94Ra0yaM5d7+sesMub5349JrOJ5wQgbKs4/pOAjofdUKNbkieRGxfjojBx+cnpQWtkGWpdks
7hy/bPlCZCpX5ZJzes6hSiK7jLyIQrwvmGeEG6p4auelRI9En+NJ5KyfGCbWi2f5meOuvsK6sJpx
p35uGr5FXUkxr33LRUUM6zAKT3DQ3T3+lHeDNj5oJJGpJiRXkKqoUs05Bgr+CD81YrGZ8OommsW4
IAvXPkM+wNDtfpqh8g19HDkHrAA6RetY2bC/aBKF4IJZ/Rkj8TDqbWsj7Qv3ZfUNU+IWnh4clx7K
eF4xjqdrKBWgRsm5iYfvIz3CVxshRntbt2T/IXA8pJM/0ktcnNpYUXsrFDtH/VXbf/A0lEhwKWas
y4A9yIJjWcyASnsqa94FGiXT6vhcw1QprWQk48sv2ZI27PxIZYMZcs83J417OH/7fdQVeOr4iaPN
HdocS/z//2q+EIGO/KfN0kycpJfaP//q8XdWdfqRDkFFFR6vGJE4Lxob0skMRdAYJ3SCrGkqlJLM
R6up2GkcbuhrOhvV5tt6hJn+bF8d1y8bP5SJqWz6d8Z3ifBbb2Exoc9jjMfrvhTBx2neTV7tcXzB
6+S5QnltxbWuHrD6sv4boJd1+T78qJH7yyz4N1+Pbs+tehQnmAA6X1+/04bHxWlkxlKBgSahh2eN
ja4jLFVyvhmS0DvCXBE5vyyG4qALGhS1fqYcDPnts0fcNJE6wB5AlHG9fuF+qhYLfJ9luxZKnJW0
7EGyYfdbKs4XdrOJiH3FmVMciLbRgyzwnyf0oc9W+/mKJF88mxkqppRpD7Ye6lmTXpX9IQdFFWKC
b05VNuvdQ5IVQpqmzS5ofX+2RcMHvawZcnZyEbKCUE+yaOIzK1iHTvvLTD1xhXWTOnzsLBl4RQDu
AV6gE3/CBb6TmFQCuA419JTE9pgKJLiARiF9bVRA+BXPnwbGakyGPpinO6EpI2/c/dd4/STClgkW
kEzVo3GUARLc5Bd2GwlNhasrh5HrP45xNgQzahWXxM99gdc9ejHtWirO+dZOcawXsLLjcnqixdfH
ARZWosjJ5nFDVuqXQUvjy9EUTID4I6dCAKWtnXxn849EtfFSUwBPXUKooQHfDnYk2y6vj2IeTTF4
F0tYHvpOhx5Xwt13PX9WgWZXv5x9xiQAcP9uNbqqe1VGT58aYRzXwnVLYi5HEsCcMsT/osapl2c4
aBx51+IRRC9JZVyAWf7qgAdNj4EM7hJBOpq7lhlCDYYPY/UMjgQ2WoWm9hk+ZtgkNLIPhlHokggU
zAC+Oj7k57aRz8psSZL+MZdxfbUgvoRi8g089xP+EmV2v4ClJcHkSb/XQ/gF7No0//b1DuqtyeN5
olpyPCZS3D4BWUlk4TJxC4+e6//V6uEofFbsudpuZL57+9w3tNA+v2sQoRjuFb6Xk27JlpeUVyUT
wOYKe6gkUDhDO5jnZLIv3IVGioghJCr7CDfNQ0AeZizjorFVApLlJjMOPiAT5GdJQD9xbewTpIOH
hQLTwl2reM211wuzG+DVeALa/Uh3yMZzcBrVAvAqrXdLzoJTs1wUTybobmyclB8yoWYuKG+x2H8o
nHReNpCpP9wB73c6qT4p8C2Am5puDY+V58LsZ/P1/TvAG1zf+bsYRj0UnpAAGDYMXe6xSIniC4Zi
oTHwQK52ymWZ3QxJEw2jt1qFomEmzB7j8/hQv7zvAPyhNIY5elzsvlJ8UUlhp7euwVEMF78llzd+
+m01Gcw13LIyGa9U4fWFvs51JtYSpIZpoHN09uJ3ZeurPrtnvCinWOHLUTnYlSba1NDlW+K8OASy
RxOnFpUWZMcBs9aIxI2lLoj6X6dss9uz5llsUbYqeXo+U4/5gRtRKTPotpXjeJ2HnzwdwCJgggvS
dRkGxlk0FY5nSlkzg6VRfASsn2sXu7NEtaX79LHJOdoFSEVGYIIgswuvChxuz7uXbPy+LW4VmcSf
BDXhXeql0WdDGM33dpRuPhRPwxVAkz7W71l6KxUGUPKK7jfJ3qPCNRDQX+JBQvZxPpmC23H9y+fE
vv3Vu8AsIxO0SyF0g5HgQEsZH329v9JHDrCsErKmeBUU/W2CnUBE/SftiXTTUDkJQZyMHvexMUOt
6jn1LHa/1pdME0t3MbR6WF44WEMUiZipwcCpKkqnwW6KaZxGn82ntL0a8LMU4+3y9DMOBPtXNgif
FTnEvnId19tFNEAUk2+ilD7jv+jCi/v74QWSVnQc4s6IZoZedVA4K3VlrnZetqsNmyJ4VuMfl1Ch
5aLR3JAo8BH/Ii8QQeg3K3A5aB5NiAJw4YZpQmqfvtmN6OuvkILBHNTxaI1N7TJ+45RZQqAfSCt3
dxpfIAydZyJDb6MVI35+d9Zt9PiGvTL7vAmM0r4ATV1F+Wn+iWfM4hsU0ghWOWf5ZmfmuJTsM931
bbOb6iD/mnN8SIFfu9g79ntTCGdF+EAZT/pVOA4l4mdIz0wNTKy+t5ChjMKY48xhFWc6c9dmwdtN
cOT6icKoX+lUxsUkmbuSDcqP4UqZO7wBXe8lcOud5CwskJTqKQxWtv9KnZPJLmvpLQzFlZ1HXU5V
tqeyp6rHcaemKVWmrngVDKgoP/Y645O9Q0wrDLnfpJ8HWASY8XH9+u617LVcGGhXptM+ZjhKBs+2
z1ZwsL1hUB4JlZXaSw6QM17ETuRRt9Pi4zrVLWGDaYlU7a01uPLS4F89CHgDFOXQO8OTY0NlFsPT
d/3gqiKRlXba6pIQ1keJ93jITPyv9hUBxZ9gDYAEeFLFOlXin11+4k8nf8fcUjMBJjp8LikabyzR
hKHEnSUP16XkkIH7KhoIRbMWre9EU5ByBOtP2PszFIP+i+gSJuypvh5K9UbG5SYLQxOqDd+2Ue7x
sB2tGutnvVhsL1C9UkPq6T9NMsiRLdEqdqgecxEgRmqdOiMpRQzEE4R//prnJ++ozPi+7l8gjOsS
ZsW/Bs3qwpSmHSDpEYeSs0uBCTFEihB7FvpgSqnMwSIqNsPxFasHzijorGAd10C3x5xFQc5EF87a
TgzBmRdHJaGu9LL7zweRBHnhhMqSYewc7jLsvXPCh1cnoXtPB7gB/fgGsOUMMtjOP5Dq9o8wdp76
1WTsBHq0uiq1kW4HVaGjvfQIIF0yIwq+B6MiaGXYqje1D+AycQmbuZ1KOmMRdRjaV6SoV8LSEXGe
9r+uc4PMnKYw1ADuMpqD3rv+7ayEB1QbMipcp40UJFWoUOVZngm/1xiU7so8xvcSGk1wa7y1E538
QqRr2B9hR5PyemDnYhec0pq1fZhLabx59OVBrvuVV4SKt1/Cgj/hjsvfylipPnYNhAdptCDvMq3x
GWzmmmzZsNguu2PQsGmPvQ2yeQqC+8HVqyYrL6WbkSlTXGWLGJMDxRHES1NtNXsDQquKwa03LcPN
hXw4LUVU3paKW1vic+C4iiTS/ITwLmfiWA1iQeKHw9uOLe15WFifzLSgYE0v3llaZ2J8wwKs3MNF
79CB781+VInCWOdubHt5S8K4bifWVK+4J/O+6DlOPBE1zQLkLmLGs10qxMPK16FkCSYMogf5F+kw
mOiY6NHtQJ9CDT9rd12HXikuALfbSuDOZtUpaWqp5KLj/albapggDXa8jZ01g3ieHAvtBF96aeru
Brry1sPUiGUmZoTCFwP0aEhcZeW9EddteLBN0TUPAH7eV+/4c0y3D2B1LFtHzFjCaebM/j8tqVBC
mm07feWgD/OX+Wr/UmwrPjPt92piRyuha2lx99L0niqMM12z+R1mZsXJ6HTAFfMYcZ27NB4gwZ+R
yQ0SibTcLSqZbILTJhO+Vp5F0j9BjilWL4gpkZPafDRz3937vSLmi8/HdwRXKdUkKegXnLTpUwWB
N/xE2bfJCthV6v9WjrBEtJGxRrhM4sJ3WSXsTbk3/bUe2YpS6rCxymRdyj2Dnt9VvVYd/tvqWy6w
ydBBq0vUSKXGRuI4gk899swKMBsEVKr4kS8fwSg5w5gTfqN3NFnkDCzAU8y5n0/PeVtFAFgtr6xb
u2P07JqAMmeu55kXe50diSHCmIBbJtxgstwy58odTRz9lYF/QCGrFh82tWWJMuJquP7NJGi7YmBo
2c8ypyK+oLqv5o70QOE0C85qNO9e8OHXIF1jo9p3wmhk3sUjuDi6l9KlOpcIOUpYHuVw+BEe7sam
mhqWYyeSeRFcP8mKwDyvFzY7dPivy1QQnseWsMB7hYnKK2OewbhWdEqHdFbluwfufrMmPa63d9jT
86iKFuueylkrgPOv8wAf1bJPA2WsV+WJkhmJAL7oY+UMPXLNuY+oP/5V2CmkjWMEudmd5+ZIvJFY
4osr6v7cotOKXpjBv8/bxcrAOZkbqi8iRiMA1wwqV0C7+DhoVqrKJdX8szZl7iNn5PavLiuIlRBu
9Pa96T8vgTkNJSln9QB2iVVxp9kyb0xwqDd/ofgbegkQ0xAFD6tv767VFeSFP6JgnCdzfBYqCubM
VkgWMVD3IdVD2tZnORtZGbuKTIAKZXqr2kcAbQy91NhH7mUDl/szmKImJ+v9Ca8GNaIscmgy1CLB
6S6GKadDbhN+xOP2VGA8FbUTyhLeIn4hdUBqi3AXFeVPN6i7ifbxmheQeJHj258TosJpZsUEiEz2
bQIoyuRGfHua+YlCXqAuSmVstkBLW6AN1sm007BTwiHu3aQ9tFKvN46kOS3CfiJY97ln2Rm8WHdS
GG/F6jgI5OsOjerVYU4QYxWovP3jTSRLjaBwHfVPMxorLPoIcVi2CcY9ERj3syGprNQlB5XHP7Ob
Tq2XvlsW9/YPLEqIz3gOHH8dIW3KZ4wfQCLehQMPiaaUZtdjYNA2x5Qbwexd0OGbLdDdtyju+DXQ
TkXOsNCZmVyL0crZvVlZIYZbJAONIXL7X0Vp4Q7pIBqF17SqExcef8RqXFQScNKBOuCSD2WWrq+d
3FACoXzeDNLg3YnGmmIZXEvdeWFNtroTiVRDteM/AosK9rgZLWOE6gv+g77bENMA/DqfaNjSw24e
I90UK/ftfrzz/KCREvQPT6tP3jb8KKKzbttEQkdHQuVwmqJu2ihhDmsuSyZ9ujAkZuuxg1iWtGoN
N9IdY0wsbw2uJIMr3zJqNRx1jGZEtLeiPcLHghdu7Rf0xJ0hfq7WP8GKJwrrk6beezu5vKrejUFb
lzzDYjcvy8j5p8Xs8HzZfrf12CIfDLmoJ1yaUpr5Xs3Eie5wuQmPKX3Ck+eTXzBzr/HdxbMHd1lV
m8vvw6m+9vWTfrbUtukR+iTd1vbdx/eNB9aSAokFu7yAjQerrIBxlTj5/EJ4agCuS00ffLWAShrc
iJTTtJBLAUYnDyd06GKex59zjHB8gNXEzNpyasoacHN+gn+WWKgc1/iqDbXjN9vT8XFbE8UPZgt8
k+lQmywiF8C7kbJuFu9+oW6ec8UWFAGrTEKudNH2w1BxqLuuEh69NSYM6Df0Gnfxm9qQ9qxbd9r/
17zb9wf7FjDPFqYM/bTi+yNqVBxKzbAjKk7C1TritoRAZDO1UdDO286edSjfBltfMoSxuOTwg8b3
HxO4jg1BQPPIrFg8KKy/M1d0xJih1FcrPMTK1PBX/MDLtHwEkQ/vQPbDETx4wNgoEtZyv4/do+aC
8kKJ829dTMKoDXN4NvIfrzF129yZGUYfLMJy/q4cyUqm+/nQn/Bf3EMVFR8/hBwZ/X0n50WlUcG4
KfvNpHAHfZgFDpx9O0Nx5hmaK7YIeJ30eup1q4/vdql7/cMIAc1nIHRCt90fc551wtQLysvddCRf
d2Fj9NqbrUrM9xoeT7YxK7oTQHwq+Co+8cutMxpHOgozA7qWjJxO8zq6YKSU3HBG3tNSdstlAr37
pMTXL0J66kryW36YUMD5WsEKqnpkY2GkZP3s/K2wK3fKpRk83dQT1WfETrK+itfFfEalNMFeqDjT
yfxERmNHqO5p4mIsvoNMi2AgmhAMxpEKhPLqXHZY/2wra22Um1hNSFVodQfo/IMqdw/w8SVVfTrp
gX1O694r+rM73ftFE0M0oRNYDKfUZv8emmEaxsuxQGp3UoVMOKSOztJMxgdAFokT3l2TF89vCWb1
UK0/mn7wigUt7W27fZ/pm+k/sH6gyAFiqbEfNbRM5ZTPDAF9e3WACFX1MhR77m22rImX6f7g+Hq4
STvk2qmEIQA9Q9X4q/YyxI8/N4Bjg4cuXgYEMBf3+sWFbUSQLTkqzQ/HegI2LtDR1B3Wo/y0YKQp
6ylJe2EJKfSNA03oBCr4pjVObch7YwhGsdF8x3ce8Odov9ps8ntDh05upwZRIq4XmXHg7L7es71S
RVrnw3R0vfOkAE1mXuhZPD28zMrIYzzsz8S+4M6e60j8Hnfli/0ACnvfvgN1pBaHC8gGhRwEuKDZ
55ClnOINldzSb385pqR474W8IpS6ETf/5l16PZD55mlRtzPANeSbe7mRHAjhK7a5SncMGA+unpMp
eeiEe8v70CpnEAJgDRWQp4MeKykhmSwSnrN8H8izg1D16m3hrLOWmrMAKi/B94CoZP89BUp95sfw
bEkh3u6ZOnyVmk0vxLybx9j+E3g7KB7NOaDJfzvZG8SNrkUSK/SyZX8sP/66xc2Tbp68sesJyuiy
2tk3RsOmaSuT9sUAcMLwAPJuoP8ttpYdeAr8htQA7WXQSm3B7QsTKW7+gBUHCBGMdUSlOtrQee5z
31yk1+GkEendTWQ/Phamo5LRuuTbloQxnIuWAwLERNU+FlYhuMEcq99GIPEB2/H/Yw81Qx9Wii5o
k85ss/Ayhqr+DGTQCBdECw+n1Ha3C0uxpJmWni9oE/+Vq9agqLQys2KkHrcYrKSA+C+iWYbtBA2d
Wckcz/LOG0qJ5Nn46GWbOFTbK+iMXJGUbgVExHvLtSIVa11HCpHUQvTj+NrDyvG78IKpYFOMTSww
K9HFpg8UNIX7oHw6vLr0Xeqk7JF/hTpELAZJdyTLp2GnNFn1xI9VRJG/8cT8oRIokrG/rdsDKg5s
Djz+fBkf7H1qvVcBWvOP2nb9S3/CO/v+qxjyuaE2vyf6Ho6HQIyZ2IwysGG9m97K5GHwHGQ9HLG4
B5Uf90ChAqfB5LUoGrS2UTDGnIoeXZ0822yVV56pRu7vvmiTglfSFM7/wPfdHKBbOKYVkHjC9XC7
wtZmONEGGkbFX/imBuyupoemdHHjvpihGBragoinNYnZ1VKCk6lBXgswun8llaK8y3TRf8yiQipm
Ha138Rv8k+Gty/4ScDdEm3vq0sa/LRbqwhHAM7HWOJ5aJMo+aC6nnV7ZI7/NfErtxc/Ro698TXig
R18p/CPvvajoyvkZc0KbvfftumbFnOJXuIcIJyYE5+wYKdjirtsTxNvpnzxcx7CME1RprYff5enE
XiQ1LXAC3b9ZsBSGvuXkkCr4Ujpr3KKM+EjHoacXxkKXIKSRlSJGnWrsmVgsFNRrwmMrG+KymZsG
HE9lm2tD/JHIM8IAiI8TkcDPkJXCcB5TwaMETf8KbiAhsPHATbiA2re/wf/cYTnWIBvViqGL8f/6
AAt2aojawbr+2xwFUsl57J2uxDP+Mg4S6sG1UuqXcBmWryqCphNNJTHU2dcSxi2lKJEF3tjbGyuI
ejZRGXHL2iHuFz9SweZ1tqRNm59nbm97QSAf2GbbeNbjjFnN1BpSzVe1oWqyH2ebY3OGf79uhpqc
mbbD2TRcejPjKGvIAaYD1M2EZGjV/U11BMNtP1YgyIbqP5oHJ3JtFYElXGVv5q52kkxlNXc4chur
Djeuy5YpDbmkqgdCfzHxFWj7Af6AvCRN1gXjGYnU4qkTkP32LgzvOVDSGf0yFPPj0AqcA2vsR+Ik
uySG4VWrVD2JqokPio2bDPL8FTtNQq1gdyOQtjSLuUTKlfimpQdW1HZSW00ZqMtPj/vtQk2UgPHz
prcnz2NFrmlgdBduul6WKMgl4u1TiP9cpCrRriK71M4sS1Jl/kAxdHerlTqn6xAyC5ooK5d9vwB7
jn3LigA5X5ZSo6zHZPa2x3obJL/o8MCh8XQr2qRAPuQXPfk9spwhNcZp7O0LGHx2yimkzhtVE0Xu
5SjDZqobtYdPzIZzjd4cibL3u2yENRdyOA8e5GK8pm4IV14JLJ1kqQoZgjXFO3Jngniu7NabdltR
LaeaATZkxBTrFnhmtbtXLw4joDKdNUMWhg/pVmnl+XH0BoM5VAmG0eijwQGcOR7R5r1+ssJIKD1h
L5SS8UFeQVwVeBuVOsztKfvD2GIVbUqNq0r1/l1WFBFrlJMr4hYD8SkJYmMsADqJVbv1KJuCGc0+
3qsuwBu03iP5Oc4nAe0MdumT473RmLNu9eqBhcZQwHadEutfh9Ln+bM3xRucZl2BeyJRWkc2rCgF
oKMMHUUEVCWrANcQ8axDhrB30GY1eTmL24IHKybnlT7E3/LoL/Nr7oZwhxhyloTYQxO2j48NBgK5
5Lt0b/9WN48zZePozEzpHybI13qNYWq2yL+OwTI5poJ9HjY2gofiY/84qdhweMizSFbYFNB3oVPB
3+MwnCgkSh7PILX1Ek2e3kDl6WRqj3zM2U8u1dK+UOMd4/3CKDOyOXZrRpg7h48SkGWCqbbHL/gb
7LlYZfttqfz+iRKHVqR4fy3GZW+xdoxHYXf1/YBa+HXpDWK99PTMHaUJ3dKyDlI8EE9U7ASSQdj+
U+f2zuxMEQHVI3joE/vacZZ/Kb+GwHduU10fWkIXaMzl4RdetuAc9bCrGeY4WG+H6NNCfuf6qoZh
im3GEnS7MEaOqBSjqNARHd/LEcJc4OV1lyYmSqeKxNS4PPzYh0E3jKsi5NgVBRV7HAdQZvZkVnte
rJYNtlrusrgsUSy7JY47fMZbMKXWkdO0UB/F/qWmuaH2mkxokY1fyqYrhI3PPGGwtz+3MGOx2CoF
9ZixiDge44CY+ivHc+uDfdBjpPwvWOjXWSn/U6+WggNSumH/POtZbZzP2rlx0kFKpyKQSbMErHnf
O/P/2t1rtAU+4iHz3gBOHxuSqenR/L7N9BrWjrIO4T+GWjMck6iId12nynXAvxc1ZaLgrS5mRY+y
dfqXrl9ka2iLeUfT49SHvp7ehFzqT7R0AQNOQN4k37JhWpCY/ZkXOrqdmlkBm7CDB8pF3vnDC4Pd
VprSQhze6JHOG3DaJaHEvbH9upedLAsTeCjjnYmh+l8OI0NixY5SgNGD5sZ0+C04/U5KAqLJHiEx
JMM0c2rfY0Wnd7FisbNeJanINgqBnSKCYdOG9B5B0ZqfnAevBdBgNxxDWlCMIvRSAuu0ysJq2CE7
fO7ilxtLhmFlQJakXjN4YBzck4N4A+R5TyomaGq7oBGbNSENbndKDbjttvYXkhPdMRayKRe+gtHS
Cf8nysBiXDHrfZ/93UPsa+eTDLWFJvcF1yLbWPZAnYO20cLWD1YUBW7dHHQLzu9WLQOtb7HRHb2c
Rqu2jEXKEVpT6StV0itDwZ+nBaoN2diVX8Kd8Nuch+0kPSIHnKCj1FbmLgQI0nPOe9p31YnS5H77
EiYENlSy7q+MYkqlzYjCfkFFCqSXVQDMOSlbwelmz1wAsAVZQP7RnJ0HjCx61YdchkpW5kQ1Ad4S
Pghjqy0ggH1fc5/ywOOPv6abS6WA5igdBUPykAvmAyJgLuldOzkWbkHX1+V9KeKoeHc2RMkWSx8Z
0Jgg60bR4my405XhZ7sOAN9ub+qdWH1Aw0JjSvVva9FnIcge9mB7JpzUQLf/SLxJitUr9ID2hccq
KAk3QDzgeIxj3tUVVQvDW2srNeqvUZ3tzGsB3teZXDfBPtMcIX+MsoNt13AUIDHx5LqZLLx4HYu0
OWQ6LptsL2ScA7c4MeQDGJjlnnzia/EuVJkmNdObhrfrIOhAhKoxV+YS0x1s8btKlaVW3saSHxKL
RoEcMUO4/Eu0k5TWVzTjaGH7LaSeEBlhtDm7vSkkSN12qFANi9frc5Ap8x+OBNmMFgoPrKxxYdUk
W720vOx3Lb4TPqmBxrb3aSIQ67cuGv/PabtrdWiwPOG8YjUSOMTuaosxnGribAXLhW5I+X6D/ze3
FRQdPUG99m4XFrVMSQK4Iv93JhZCg0E6+odQ5EhGZMUNP66YjlR6cz51CrYqRcdyUEqcy+qRKNBC
7jN255luGcIlD5C/iHI+x14d5GR4mOH4m0BFDWW26n/2nWcS4OBNRF3QEjmWpIwbfjhWlZrjng/f
wRicDrjtZTqa9gyfNET8gTEqGu3VlH1X3H1z3UkVaxIpsJKqScTgV0yiz8I3rzA9hSRg1DV+LiN1
wNTuqhHT+Bkk7BQG8bTJrV5RWPAQEZuuipEy51GzVB0RWkK9A++N6ODdolkNQLIKAA6EzReJvy9Z
mm7OYEr1zI1TKbnqD4KBNyihxBrLyBFnfjuQONn05usqvoVkQCwCmZ6rr5aqu8+q9AedYyvSYpAS
O1OpJMWcIgW1EfjW5ndGEmLwFpBU3qNO/O8PRO6CE2W8KrdCJPWepQcvMa4kckgyVPV5jHDPEN74
TYpLGd/+WazUf+zwGYR4a+VPbGOtzA3sEUzGsOUshCn9wznIB9x4LcdT3ymgazwc9gGddGWFoTdo
rHEvQm9q1CzoSLd/jfBIi3l01BTov74mRmTsey3fFfotwEpR3tz8mnwoAvK86Qf/I396vW7PsRkO
7Y5kBM9I2SMKId9wRTbn/U+IbEOo8EuxyRwEj0jsqg9LBkv4JP4I1Cvo4Vtjb6mPlN6EbbCpe1ke
pqp6PKtncgQb9+UabwVEwn6aLc81G7iAyDop2YBBPVbloGeIGAFgWS1B1S1Bs1Rt3HCxjDIDaNHL
oFcNZ+7AexXt8xzkUbnlFmQJmWvjiMoZUnJX3G8x9p5TVxak+1HJ42IaqeIg59KBrZHFiXFkTRXO
loQGHStJNa6adrx/kllF6QVc2vlDQn4KlCKf3mUxptnUHjCJi8I12iosB/sCOpziDamiYJIuy0vO
bWkNHVYoMqMAnAy5WgsfJHS1SMa7Pb4fQXW+lbZUmGmoc/Nhw8ld9TQRNxzmWIGXHZ7AtlYGDrEs
/46uPnz2hTSu31PzhSOIz+NOfLWihmptlK9cH+T+lc7hj97gZm+263xkgI7/5FCB7PHl/eC3R5+l
sq+/nDbsLuSjQ0p0HH6uZ/MDTEv56t4yvGCzGH7Owfmfpm9lz3QsfiuyuYByaeiufoEoQ0fAn5Xe
Vuj8JQjYXJ2fzAToTBXQ9/2Xs+90RkGJ2wQDHhninkuEmA6CyPDpMAZhbjlUHnRjE5b/1SUXW4N4
u2kadCdBZPf1Q3BJZe3frmrMntXesARXDM3RTClS7ln/hAPHYuyOAebPC7wAXt0RUT4x9Dwq/W5f
IyyLSa5JBxKATP11pMO7Goc8/KEiNLNBFSx5C6sLJrQujgMhWP74IwSJsxxW4EmasjPg+RtcaBMP
wF2Y2hEMDNgXtNRpfb79B/lslMU7/kYzw6LDbwLZkkedbIsfJ7nYgM8msIvtluM5mcBJgpu38tGk
Fwr91gC02VheDHgsC2Aala4TpDr+cdLrfQf/AUBj9sAHzyGDY6Xi7W9PinR4sRVX6WeYA8PpUBzJ
eaXWK6ulmjaQSIB+CM96EipfmnRonqeIiFScKhU/XTEArhF3XXx8dUM1e3FPbTUSpjnyCwDYHs7k
ZrFB7Vw5YFm4xCqqdb94p1y/JO1H9VdcAY2LtMBiI89SWqssxbYRzfdA1MWAvz+Om0bwyZv5alyn
UgWFD0klTpWcIp8SLPs8hpALoC3fI+8QbiRoy6rh1czIBrMnLfgYPuJX8EW14YXXdmjgrAjnP6RB
pbZ56cwR5Ke9H4foAAuZwRI1Mine8y4/ht7SndoiHyzMh7mYqsu9iTeQARa+53GPXrUHdb7mGNLa
bMQSX1AEgJZ4IoYlFbuA4hb7KGXSfocEoIJN8qUe6DxSmUgmwPolOfK1bbhm0zXrYcxbNsBn8mSW
eFXDvlx4/WsBJu+evQN/bLJRiFnuJLY46oUMupkf2h8AWRL3FKCFqB0WqizCjguHgKgSLROOhXJ9
POHmGyciBC5WRR6kI1iOcZv4P862mNaalNJTnYMk8hIb5vvFdeC5MlLXoJVA7t9FawE7Ao4hDiKv
ucHaqrk2azRHiHk8LNExdafANWItBrsggy54kEo/cVyZJk2z05N7zVeYbLietBF9fiSzn641nWwy
fM1CITeMXzMaQ45Labzctjmvu2GB4nEgP7/wxweDfY3mR5O5qsWHxzz/On3gSj/FiKJvOUvnmJKW
UTnJAoOB5zhaTkVP7+tU7QM67EmL9upYcG4RfH4c2MO4nWNS0wJPM8DnRXRmEaiT4YZ/+9lFew+z
+ikqRnRvnlUGlByqNPKfMJCkhjWF8DxrOgfjLzw+9Peh9PErkXnYMoe75JV//ujHqjuBPLHxCqju
safSRZiort25ypF7V4bhQsTo/8J6tCvObjrGf5GaAeRi9NVVTKNnEi9/4w/px0CUrIWXZZq8mFvo
5StkRz+ZpEJZCJZWkNEBKPgwbf4vjscFCcJl3o9nWwr0saDnPXyiQdehnx+Biiy7hae1E+wWAw4g
6aJwqmmQ8qThPEWWY3xt6o9m/g0os/23H6Zf9wbE/D04ictE9+6i5w0EBzuIME2gRAVT0rUcV3Mx
ah+9XVQTj/sPcgpXStwxVV9oJL3qmX4++r8+Jboeog1/LJ0yWu8eJza0gMm2VnYxGOWZblRe+hH2
7A6/+AX7IhUaIi5ayaP5W/VvN0y2wmgBfBeBRijS+F5mresSHf6Z696Zv6rKnkd1zsHi6hQ3+eoQ
ChG0zRbp3bnQJQHw5H0GS/Ia8j5utvxYPN0YysFxCqCajqbhjP3IbKKW+GEvOvgcLA74Ri8h4GXc
lEwBO9FEGU7cN2UhobVVVG8mBn3/4HQ171H2KbJHRh0OZWDLzK6AX8AxkjNNGjfoaKfLErd4CMJo
1CmHkvZiCy9HwNpuKAdWXDfArPmS0U5d0E/Pts1OMDEdAyPpgE3sBobFMFT/chz8VbGmZcZRrka7
dv+t6sVLE+QTfL1bW2kFqak8afn55gGtRCXfVsj71iE9fMQkMC6fGPzzx03k1Au1rQKvP+ZAvHV/
ATXM/8jNRUPoiyVomufmEBmwGV/fxoGDVsx1TLi8lZbGDCzlL+L9zMKIHuT18Hf1vcAtUv9eHBW2
fl65PjQDNoKvynwAP0YITu/MgaSdOCMEXGHc/fa7zU7u1JNMcxhC30gMPRvrkkJKDs7YhN9AZ88f
yGNlAtqZCZMJctIfurUEgozMAvfr24RTlgxIVd2sb2Gzvs7B1PIttRQi5P3+0vWrEJNwT4d7tn9P
RnxejQiCLmzKhenu9Dh+/BhJNm1OBahQo0HDPOrEd2stH6rLaf8Kq5i9DOWmI1IdVgKYsI8fD1jX
zsqpzevshsSpQIj5+Vt5rjj/MhDX/7QocOncjsRwHxuobfUMR8Hhx/cFV7spkOfkfdfDTdLP9dCa
ZPyJvBHPcD3C0jVUp+nNz9qyUsrr5gPckEgKS8/IiNhjK6B+2mJzurWduIIZYVGfhEsn1KOceelc
dfcQZgiQ4QoT5VNw3c5exlmhzoMTLKtnUU9J5xdzZ+8MBxVBUOJ7G9k9y6nbIoSSrr+xfb/6ZWob
PmkkXkDcFl6f4G1XIF0bf8PU/hP9E7VuQe86yzmpzOoCaVr/zozMSiV9zZovAz0EvP1+o/fSygTQ
yQqu8LnQgJafhRgC5HUdMW/sevHsoViFLv2mSWi/JU4mZJPRfTACzLtIMzlzXxzOyeNakUuGkdi3
oJLst2y1uD1CmSu7DcXSnXZoXXrz4phOQShaTQ17jCvvVMtVzRbf4jm5zRdvEdqqdp7L3TxqMjJV
M1VhAaAvBYp/850Yg9dBCamUcfq7WWnB7CMBsna2gU8dX55Tb3XsPZIUYIFMbENGS3EMyA+3O1M2
3iTXtuvxQ155b3bEzbEh+KxGsbZcTRKjZ3PFtzXq50do7ZTkLAwb69+HDN8rGBXm+WyYJYw6qjb5
2pRyGhqTKnJ4j84jwD1SswU3PkBHNV4EZ9bgo1RUODhu6N74dj7F5mj7Mb6hBo0cKQFC4wYWxPoU
SdCEmtGpVpnJ/MjuTr5OhOjBy1ZPRiI986xmIfEntZeRjaM1AA3wURNjweu/k8s/1mi3EvWQvGMN
7lw4SWdibEm0OmyC4AojZembLl0vEn87qS3Vwd4hIOq6wti6qARG3+VG8XHDSIu65UOKfy522TS6
fphixadDwZDgul3kmO1XhW1i0pqla/bEkgvi4CWVZ7TVyCzql3ixgUpprR+t8smCHb7AIFCyRw0T
EhqkiwTQk4guyyRbNakY8++GqiHHmZxbdJaeD/g/QwYLbXLWJqQfgOmPYc6fTM8KQ8eFPFalkUej
ogkzlRkowphOHh8wd4SuJQtt/S31v57ia4QLtzQd9UyswadVSqbCGoAQeZMLOrldFFzueW/2cZpJ
aif0/8OYwnA+hxroHLAjcI/EvhF172xhAhBZsOPRmaCL/5Grnx0p4WXIWt8BJnRuLNDVvpHdA+C4
FxTtvV//5Ig0h6MZB4KZl0fW/wwXkP7F3/kJw7Ng/IzrdIJmDof7NUjkHcCHTYbpwtKF6Ey0u2Pe
H3TPK/em+9pwYeD73ot+qTHipXbd0g9X8DrcgH7M89zHK4akW2Gw16i0vjk+c/Twfv0M5cRbEruX
F7Y3dBMDE4NmZSlpZnTlkxwkguoiz10BhTU5WpJGK6wELLMR29/nm198KszYwq+ZSkqmK5ek7ZWf
G/KYj5aqp1+5Qm48Qux0p4Vzm3AYMxOO3LrRjcYOz25hCIMM7TO75UZ20zX+/z7RMuWCyeqjx49r
0kkBIYPdtnPUrB7VBQFtzOft+Tsr2MB7GMdkfPkLEbnrQrSnXCfPk8jupvlh5JUsix2+7u+TJZoi
xAOFXuORaJPL9Y8DPVEPriSfdIkyw+OCx4x3IFjctmXm8isdZln+/eJGhOF49pa/ag0ChkCCjgJP
OyRc/GzATgBKupi5kLgjPkNe3wyfYu0N8Pome3KXaRU5h/C1nyar706Aw3MEVCEJcj1DafOraByh
s774EE96wmAXrRFsfmubuJSfmKel32DqT6I5jCfvQ9iZfdIynhEigHsz9iNu6rBK+sOLb6Gjf8uT
E6PrLjx+Eob7bYYxbTqxfJN4gyak/Ld0w4vZtYeeLsUHQCmCN8FNxnD88pRaZ7lw3tWvq8KAG9n7
CXtcmCsPdQNHsZOin/i8wYEPPpdtsmsvoe9vG7YlPX17/+WbfnnbzC+ZQdqAIY/wIxRiHLJeX5c9
98ZDTULl65L5KtGvCE4ldhDD0z/zcC80Qv1ncEiMrrDSpcsnGF4Y7/HyraY0TwtaEENdNGDwF2W7
0rhk62oI1z0H35bz6frWNpa+LLxN8uPaegc5iGYdSUnfSntDZ5zNXj8n49vI7E0GPc7HtruHmqdC
Fz28SheuX3untg23HoxjRbtOsjghWefhriwxV1EZJgfwJclw2ZvzCCIQLLbzk5FMsfpkQxtIFJI/
0ZlRhyX1geieoTcYgTU+NlnX2Z7U+whtd40C7tN5MLwkQOkCL9WtsAsvl8NJViMEEEZn218FjiYB
hvbsbcoscO9FBFInKTdXAuGjFySJB3HfnZrd5q5faotA4xqYC/LudBHTBKbZhm2nVRK4Myxg+f1m
/aKN29g8NkemDP5/AAlH0Vw83kczzMBvdLCXWbcPTn34vUhYeCAjm7FWbd7Z5oDIsqxOAz+Xjy6F
16wA55hkQCAM6Vjx8Ib42OoSBFv/bqKrqygsMx0X4+aAEUT7Ir9R9yOcFQ5hw4qwBRIW21ejTgqe
gT+xgY+PIPdCLR6Pd6VrekUz9UaFYjY3J/81eNRNGRyVQfsZh7+u+lWUWLpmPC+x3gCmhev10gtS
b03HZXuXQRq742CpoMcKfbBLCJbbhJqgGZ+ePD3mcufmdbWNGiWau0fDq6yZV50xDFIzz5Y7pe75
AV8MNNFg7djkFlo9tcO76N9n7PA+uuc3lmfWuW29l5vRLdCcBgVKjrVxahBtVcgiWGCFXVwwYF8X
OF427t44OE8pBlSVqwMQQk3G2VDE23vT+HAo43RDFUC0XrQScB62Bypcc7ZB5juG/RpfXJ1yjlIQ
ebkoZk6s2NpC7DF/egz/U4ISIdHWxhXTnjaQ3SEijp9Bv8hwRlZlbxOfVuMaJS3GOduAYShFpw2a
p68OITxDmrmpyITHQ7SZPCevSFXcnPqLEweUxj7HR4h7eYLOadBdpk4G2FpXQdT5PCD2OGxZCXRO
AxKIbRdgV3oOJnwWIn1p1jReXQy2V3hhvz0JGUzpbDn5rvHufNShDKXy2WJjQVMJbtxSsF/quaWb
PcoCqkycOiL5XW+XYi5nIbspdrcmy9lE4sY/ZFiheLkt2+43zusJLsc183Po9dYdZOhiqYjZOf7x
VL+jq26GfXl1JwjP5bP5g4dFxpUPFBRqhqrPFlAd4JOxiViK6v8AFwo6DfAZwB48BlMqTyuWbjj6
N04jInT8p/7wzOJ8NoqtAa9R7aG2wdzhnojCiD0anvPRsyrs5tho6UjZdsYaNpilljqmM918fiYa
8+50dMQKv7CH03YqkRcO1fOduzRlDb+srZx7KoMFnkwG6Nhjqvc0DDXKOzgGlV4tCwVqzX6nZd8o
6MhIGqazWbRDOrz2KAVnnPmpIO0joVh/R3LnJ1KyRuGkB+IODOPPOfUQRWeewnW3jtDq2ZUdPduK
KimWpFn0WtGyMOW/73Xvlud+itOpGreMDPk1cktYwWcXxPz462mVG9BeU7g3g3MqoVl83n7wYxWA
Rhn29fzqir6s09DJ138JIbcK8DURhAcGAa0wmkynGj8O6DyQ5A74A0l8WaE/7ca1rScNRssTnddE
VV3c9TUOsqovt5X6M0STzbxeIBGNW7enZgs2q7F0GlaPY3n9lPpjj/MV2hnbxiwbaCkPXb5mkQS0
/KXyHL1Nr0RrMgEJoYMpsZ5fx6xqWKWRx6flD5yLiiFhl3VpJaz1LsTHJMyV6g3P4zOOvQ3dXuI3
QXF3MOHL2ztOn62drzbRsOW6y3Y5u77CTd7el3qu5OXjIYpGMFgcETrVrfaOx9EAZmZTH62Z/DuL
v1xEcwDk963OeZtPhQY3ufXHE+KL+kqk8hxNiKCWSOjAisRUKFGPiWhfWbqPyUFxTi6691q40gYG
Mdz8DuiaF8bd16XJjwBNsy8SuN8d8RACB0JKblDcBgJiaUXh29MZan8KAjy+OOgqe09dn20wjIbQ
lTxfnLHaKZUP0a6kTzxUFZC6RI6G392pDSFNQru0v7Y1eeb6zbhlYsy2Mb1bK0VIXvEQbuxSPJwh
jCNx0M3wP37ckdgDkA/TNQFDkCzcSEZx8jFV2KKnKNzLxczrWe7hiXkxUf93xyZYsvjJBpn0Y6n+
IEhTbX/TKIiYtD2if6S4SJKzKQroMhLDwTK9U2z+TCQpl1OxvB25KURt78PZ9minjvRN/cDN/8ZI
ui2rj4zgL5G02dnRbKifTfZVvutCEuu+xd+oWW0ctepJ8uYKAVpox3qFdNU6LeP67PihkPzZ/DS+
XQYe6gdvAEYEw1HNcPdN/NatxsDnSZJN81bMaKUZP7s82E4KzmF2cT6gtHG9dKx8RkFr6lqAAhi+
FhVnzy4oSGXdtdcJ3bWYKGv+k2dq1uBPNLPaDO55CAgQYQ0bZR8CEV4St6gyPXJ02Dsxgqtqr6t+
bYdw+Hy5rRQ3OS1//wpjjg/0zKm6+US2wXeFCyq42ItmvUr1Gzs6PjS862IWMk2xe0SvTYXbDkpF
9V+GADMWwCBlwPxlW9vAYyxn/tLYp5+QO49mdbS1stimVArs/6lrwiA0TI3EScohkjo3uFywFgUy
EYo0SWm7WlVRGlsBl+Jfcw/CS8pdWGM70tOK7H27wo278hgTtnJsi/pkmAvfH477AsLGQYNYbc3l
WHF/T6lD+0UiUIWIPxmT8Kxnu2T5gi0fjVpLH05YlnWW07Agbh3krnVUg9yKc+3bTq6Fdw5WvC+6
lmi9I0kKBZD3e4stUmFOlGrcFQnHSbapQDc4Ad+tKl5+27888H/IHIrbqSoBdxtVt7nJW9e4iaZX
Cu/57AJ+0jjrTmge2VtLOqjlWqnywtJwagkj9nnAys4BFOHMIFWl9smzkoQXPFZBTKrlPwFLGx+4
pV8T45qkoo5ECJQuRDsy+qLun0jDGMYTWltCPrDmilQoN7DbxaGfy3zn8mhYgXhYBYLdnFLYBpy/
0U0QN074mTPG7iS/OssJsFKp7E3FwyE+K83+LvPAHmgLOZGvD5N5J90R3/zD6bMziT8H7IDC+TP8
jH4KDVpBwTzaRMPBq3+6DahUuqhIn2BiTuiaHJ7M06R3gGAsfmb/0L9YxDb7DzqvDNDTFsPGsgcT
xqqdNTGkk26/38a499VuL9yHFan0A+Y/f0HkkHOKHj+xLMRv6cB4Kl4UqPZwLUcqu1aIWbZ7YpSx
oRBHXvNtTnTR5b/SoY3aAFjyH0rqP/NqvXGyrOXz0vguHIyJLE2NVZYAgrROUH6PjV/bWZuxWfFo
H+UR0GFZq75soYrCZLO/ThRRR3O5e3XFfctuf9W0Jc/otO+ezAK5nBZ3jsgvCCmNCxq0778nh8ON
0rXKsNUYPxlFWUpN0KWHzuhMDU7t/EmDsL7j806qUGhYPTySYEVNNul7amwce89HUQPQJ9JZ/9Gn
NJ968eSZx+aKUj+ryozatMWNadId7W7eqVZZDz1/JYSecTQskR6dQ/3o9zKkaSGrj5QFH1t3k52n
ahulfxMCaIm3ikykk6PEztWZrZe+GcYxb+7RfloKsZLtvOmthfAT1L9U4iS3m/+654rVQt8/lGH2
WPfur8lFjPbH5eV63xoxfY9lXKwMj7TBabNF1mNI+ebpYqT6wpFBPlw8Ny80fkJZ0FZZH/e8OdmY
rPQSmMaapiCK1EXksmitSz43rvjOYAXY+0GWj7Vy37blSNbpHe12ms6GfpdWQR0w9c6MM6zJwaQK
SK3ZfB6/a8axGBUzbn82YfS0P5Wm/CkHMGRZm+WcdEz+jv8Sdn2PIpC+FGyhwa4FpYRZ8fvoTGLV
Ye2w2/taH6U7TGJSMIyQDyucmuvu8RrJvtf9uIBJ6Dbo+KYc0bxti3WQSaevW5SIEGG7N01eLBzM
OheHU+vXIlsIZmp+IbGnDEbVRCW/oucp1nSsYnxC5yyeGXqq3GJqQutLGXcGfMUS3wzf2V9sF7l+
2LSoW1nqI1gVkiP3Hq+q5jTl2vstTF1VEM4oV48uCsOSOMIX/0srScOJK6mZQMfVB38YeabIyOQs
fCKnzIlA130FiRDkEI4onqTretuRDcOOb2HQxOZWefzqdoSBHob2wpfP+jKHdnaUpul597xIoIbV
gWOX8sBPcvTQVGvw2lfFNcKqjA+PRKWJqm53yvoab6N8lYkf7rn30dsd5wchXawl1xBfzg5fE3AF
G3TlEJatjfdOgjT+0hnseg1lle8e/Z0YpjJtVjqNwdQxq1R630cMvc0C7ph/opKUn0wQrnY1+Plm
lsn9Q3zW7b9ynapSHIHgvcZCR+jbbA3SC2VPwyHeKNc7TI/yOlrFJblS0Ho8jlV5u13B/KY2fcAu
xpTFG0nQx8L21+yXNevPT/NeM/IQj60kJbq63oiEA/hSL8zt36jlWtVngLJAzxSpqn7pTkETg30Q
Q8esEguKY5gDKbe2a70NsE9+t55lRDt8+CukRG9+d3XpRam2upa5+OjtDMA+lVGaCm0xYBQfTfNB
Kg2MkQLbXnc9o9cSIVfciIthoqVm2GcOBcvdjKOZJkVCljZoayv87zHsMOWgmiag9nquT8SIOX+m
sqA68zxkKNKELdzFXwHGC+YbOtaSGGXhS3eOzHSOHGu/clYPaZPP7AddrzW6zM+mKULXLq8Uv37Q
bCH1A0anOf+QpYo23BKj29pQoSVJjPkkgiMfggU+d0l6FrUFUJvPJyWyB0yh571jxaTvOmcehie6
fl7j70jdYwrlp2I/AJnjp0j219HQLJ0e1q2sEU6heW48NLnp/Y2Q3qoA9R5lzNpPVLuhsdFPUohE
vjQ2KbADoISgFQ6gl41Ij8x6Lx9eouyEZu3onGPdW1PvCZNaqkNiZZhtdZDt9RWeW5oXuDSk9Wmu
2f6eswCHzN8LJEgI9AdB0D32bxV4m83qbLBYUcfym7xZ+yQdewPnsoRlo3QlmHgO4HC4ywfRqG69
RRB2EGmyETg2rVxF/nanMeC+KYg152PozUq8GD1cxSZxfoU/pEU3mJpr+jZbJNd5CzS9uKEd9f50
xssgvWEV6421hu5wJRm3HnF19o4NkcUA6y58AfzPvclBM0SE+L6R5VZLX1Y60l4zS4AvnBsc4Laa
/WIlmaFxIV71aMAzk1OdAETKe05/gHNukHdP0fXyWx/faZ36iTOAA8wDDdbE9ATK3WGjAqarnTpZ
q0wJVLCW5C9ZkAeSfPPzATN34IHLqF+ONDnFjQMXhShyMoqpHmaxCg5ulK6Cgmn5TntKICIYrh1H
zjlj6dlHvDet7lxtfhmcivgNWCi2Mrfs2OaaTqpro032a5OkflBRlWZn1N8RpjjMA9UG4eRCn7e1
m6TXWTeJmxvjCbpo/XsC6Hq7k+pRVjnrV3CasQ36HEB9hjtjH9evScmnrjz0uzHcWkCCDhnWmuuA
qIbS8q5MV/yAZrJ2axIReaDteYYgMScIp+8o48E7F+xwZuKbyNdYWjNIuKedUqptVh4EN2Kd6vaL
pAQj42Fax8t03acgau5g0oD4H+4j3ePsNYXYTCizbT1aF+E/5wNvmCZu1v29v9rtfDFn1vd0HSXF
AF0bYxrbxII6TMZVbG7tAwlFGUMBrkrSZLAnzU/hav0FKFgobLn0AKS/3e4zKouJGC5aH5oVPAhq
kafPAM/eMWl6Ni/3a8XV3OpRXIlKQX2aRBu/3w1tIZotKHkfj4jGlmUA4QMXGd1SgaYU7C1DIno5
nEONuA3JpYVR30F3+04y31oKmHXy9awSGfhisYJwOfqB2JwcpQicjH3Z+SIlgF92vREhvUmv0t9d
GURZM/zrECIZV0cSSq8zgoJW2e+sjza8mcFxWAQdAJA7fvJvJ/dXx9Si8hSYZOVgt99jbpCNn0Av
YsFwQm7BOaVyTHX4ddYMNpxQ9Nu/s1KtpQEyymujZ4Q3jkaGv3Nq+aCWsTc/ttMjo0IQJZsq+rA2
UnRIeqJvOB7wCdOfnpKsPoJA2nDfLS6z7Jd4jo50YwVkFuxbqRv7UD1uMzhzQqODF+Y0SjWoKhx3
oa6aba51ZHz8hOXia9fG1Q0Hz6m7MXYKMZZ1QvKAhnkvmiZf65VdxXW8HbgS4PwGCMGBPDLjKKN4
l3kAKKCFFF/DTNXLfsN2yx+e6bxArWPoMJgIQnmpp6FRrD6wLG4+tQPs8FTrLBkzNsKDD6tCB/XC
cNqBJVIKD4ILjqCX6Ng3DkMf4wwCSCtHFleFko1OMwRPI0rXGlhFlAPxmtohHB/8iUrK5vFFHL84
sFS/OZer7V1oreGg3OoaEuqSryeopo8UTXGqgGGZyVP9a1gpgSQiC2htqA9uEgcU1BmL5vCHMN0n
a+cKtinfNGji4IfqauAHwDY0hdlRzobl3ePHT8yOScZpTvwC7wzyJDjKu9CeMpbMFuXd2ni1Mxlu
lYn41S8ykUpwE7BIzcQ/5ZB+bIfj6ENQND68iqi91rbxL5anCLSVLsOD86DdXRr7Q0b9JAS/r1Rm
p8uN5CGXRieCfSKM2Iu1cSypKqiHP0kqkdBUn2TVyPjkKdHJBn97q82PWfLla/J2aj6JKv6yQF3P
sVFcvf/cH10Mk4cQcZfzMqekSw/69KVhgG2kEBVjO4uRAei1HeXs+Tc+4irEKwsPUF1HMOgADCaq
yU74wbIS+pNJmtgG/jDbfu5G7BCITdYVpIcKJEbbRPIKk31iwSLdY+1OvSSG94sxWfKcLcSutg+7
9DjFBSMhjopk/pESlAQAxBfI0B4EARmgBnaMVmKMIjZMWYfPKU8gk9XQYjvbwRk87TgtG+CxgJ3E
qpmE8TCS8tG7D8fBzX5DV74qfTA7iCkt42I05Nz2iXkpCS824jYcR19BViRHiUNk01XwwTESoBv0
7lHxoOMscDrZbLh4SmtIVRGZhR9jk7lOaZWq2qPvfp/y4y6b6Cx6smS5iF0wF+tIvlXfLnnlqmME
LgWayZVmRKPsZmDtjFaOdmuvhiPuaAoNEDg391wJ66zkHNio7EtPN4yQUuvmnXIybsZP5hDExSF1
sozyn/6S+aDQ045fLmcXZ+ew0mG2jkrOsa4IrSG7c5aVW3TOr6C/Xy11MmLzLNwPeIJ50iOFKH3S
CVbjHK1v4ythn5CUyEWCDpk15Yk8ZtjtgJlnOT36uVtAkJmMMcqaGaWk/pq72Q1uzVf6k5eWThV4
1vt2LOjmErWCTu7UFwFmEO2TLQQgx7aqocV4PP58tSJ7a/MXzRlcI0vPvmSMA53QCBjUVrIRiNiD
nkl5vdf/8i/JV8+e5ORiOa5mi7Jx1/qsSvfBiiy2y40EiEtjeaX3wJmDd/TVElHHe4CX1ex9lebM
lKF40PkSCFe2PbLfib4fe7GMUcu7b2IgRHvqC+jFnMvDGBBKsyx/JOYdi7RQ31q8loggG6dBYnFX
3obGxkFQT5xfC7tDYICPiqZX+PVPisTdH93FJ5F87wtH8rH7NvMPriZ7su8jJMLwuFuZJ4Lnufao
50rbIc1oD0FTjdltdAvwmc87DuYWFLCSUBx9nJB0Gqt+jXULGJSgXfm/0BTDMzwxZb/dPEZM4IT1
Pktxyz7YSHHYdiIUzoSgzd+ia6lUC59y9rInDVjqb6gfhkDfkD9mD9QIOkwYa8cmTKh5PQVxrSr4
Fu8JOPGd1vjlJHMoMkK4ImWkwSv61BslW6ojw6VIiSZdOICEAaDM9jCr52Wq2L9qE/3RA6eLQvEF
f6fiSZ9Kg36GYlxb4JA6UbOLMYS5FHS0iwem7GPTVn6EBGsxhf0Ig2QVPbptLvNJUF40mTk3pzne
Bk6Voi1GCtnUpPE1YWX/kdvSNNjD7evPr4IXL315Gp4vvm5mG2b2OyB5vncMSMMWUldY5ypKRjG9
gG/GxwRn06R/1Z+LevokgTcCWP2NCZG2FMsWCnok4THN9uCVMcWWDgsltp6eAkNRpxrSU0acyxos
bL99ADITzu5YRTyOslqNqNImBRKe5xeSoP/j9d0UQUDy5KeG44Cc3ii5Nn3xj5vJdktf2dXNV5qp
DO2rq8nmIo/nDRLx8n9aLjUWd3t847nVz6NcZ7TUpFRvDFvRdQO5QwCkxcJWzKf7xl4Cg0/0CUze
9dcylPznf3DeNSuQZHWXbWpK27hlwd2B2GVknlttfxUYbrbMABm15B9sp1GR0B7IWtryqnJM/3wO
9yX5xBTJ4X+3uodTHSL03cpIfZUQ2K50dl8R21+9yitCFRDmUmUh2J1p+3K9uwKcplcDkf7nDN8+
rERbi2cRi2ju5Hd53U0sAiXuMGvCuUKQaJ9+zZ+BPTLjfKIrpRdB0JAgJ5kdQJAF/JwF44ZqVPM0
jTit0EgjJXw60bunnoFXsNvfBl5cLpqQiM+P+Voxbpz1eebzQodh78SFX3ypK9rYDHffsdJa8qKY
IUUNO9fg+3CTtyaVkIFvd1JqB/qKPdD+RNpO94elyHSoEoNddUug3kQptoFRyApYL1ZWw0DEeEfP
hfrU0iSWl1KZQeYLm9diAIPyxwFYs1E65KymBp8JQsvSKs6jBju8rg46J7leOmbBtDrKFFhEM+AZ
Uhw5Vjo4hnajEE1uRnLTPW38ht9qrQmxjzvyvuMUALLi0WXcdj+PNodetHOIC18Luvpr7MVtesUk
1+OT9agdBgN0fY+c6m0bKUjWRTPjjq+GR1Oha6+XuFkDlfVwgNdoVPiBjwRBuaciTuQz+zfKiS0S
36J/uJ4b1HPqxuEp8t8xdr1CCzYysahd33xKQ1/+Qvjz0SroDxBAQXDOT1K5QT8mBqeiNYlRE51S
exQallY47FblYi+Os/VjWyN6Vi32xy9agBJVReJTe5asyj0yW6w3WVIRR6bGuNrQLYXM7X/3zBg3
L3n4xEHS4qxO32eiugPnoInJa1xdc31i/NdYTNRd/rDjcuTLaJxwJX8i52iN1WCiByENzQnEPCOt
3KVZQ5JVRUvmE1G5CArcPUgwGyQSSaO4ohy+ZDS7nw7z6gaH1RxtPfl2iNNGmpv2vrLL/vjTYRRM
eTp+NFElTAg6vn8uoA+84X1yuiv3Y/93DoqqnUEg+fO77K4xtWXNjSi3B+cLsvYbL7R55yK2IbDn
0KfcQDLiL1uIhv7n9yqLFn3bxM5An9VXcuf6ksSIv3hzn5niKPQpTkWNuObe1DKHNOjPPLzI2ExL
t3NOSoGmZQUSciJ8Z/0NHh3l9S3w3o1TVVStaQ0PU1mzUZ+Ho8hrWpZq+A/J9tssEFNDs+655q3k
y//jX3J8Ya+O9nFKWIzWJd798BQCw7VC2QQDxZsQZWoZZV+Fz9NbBRTqFfOgbBCYolpWO6Z9DYE/
kiryjRZOMZJ+O0OIRkvSjSZb0PUgTbPZ9He8jUM4Ai+PC9vAVB1xbqpaZCRO2+IQIF0jfgK+qXvO
3auy7b9Mkds55S+C778dIAxlsAfacxDISh2ejTBHWVrt120UjYXdFQGJvMJ+Zy0zNCH3obKtufvC
6o50IVbhUoyV7IEAV9+crAhZcLUvo96Gy5OyvfyGMGUdayla8j4Nkv2XaBnR8x6zGkj8xJ4gYBqQ
B/cJV/0Ax0t35c12qv7x+9Hds0VgrSOsYy7Yql8RrvT+4CYoXe2awyqZyfkVQK2/EufAC4Ean/OK
jPr9fT0yeZqKEwr9vC35CcKzpGBdmhNbVB9Uxob5ZUt6hSGW1EFCPfphSItI/22vLhPvdX6mS8fj
tuBvKMGVKYHqe75Y5azjgbfRxyKdJVLyoJVuU5wJPL/w8bd+kgZmf+bAkpZ4hCcLqsKwp/234BT4
i0HfD5pPGf6luYzLETPGvCYKf9wknHHpX8Fay2oAjFzXwKmO+dr6t2tBLVE7V4DrJEODA7TWQY5S
yP+55a756fCG2VM4Cj0E3jrHROIKmeghtalSUsJTR7b8qtdK5EFJ84wNGkXEzzM10Eu8hBSP9kYh
rASZ4gxKoxoce02g/dVfwpsoazHE2eHr3AtR9MRQ8lrpidmVOKRlfSadguQKGQ1fsmNcq/Rj5knv
4unlx/sH9WX8FInkRu6CCg9dZN76ABL3jn4AruSrhpD6pClFOHe66Y2ziP6ZNzLNzJZy1S+UGF6x
lykp+7UexrCxdpJwmKQ9TLwB9XIy4wnhl0WEKgY2X1I/CIVlBYR07NJ+7kC4mZDADSd8bVEZTvpN
mW+gElWXExQIQ9PR5AwxIcV+QYRi/mR3yJE5E6XcRNYffctairTZ0hw2mNEfNg2t51+7uY+IEbmh
T49EELy8lPtK58hH8klv5zD/ItO6H+qRDyztBBOGxd2D216Lojl/bw12KwnkD+YW9MNekkjpWQjL
cmDmdrVf/26OswoBLXI19LIqxQM1t7YR6BEqn7Q1mt68N961IrnYVG60DdzxpYi7fIaeQQQW7GYH
QFX5lCf8fAUqbweiDwn5u6DGIJMw0ay0W30ZkRUhjS5cwpEkyUzCcfsrwM+Y077ST31WJw5r8U6n
zo8ouRO3M61gcUe6NGQJflpPgjP9d5mIHzmEsghLlQTOLzeyGwUsHD5GZX0+r25DrBtS6qsi+E8p
S3eVicMT/mHUhSx+B/6m/WJo8IPc5uajq65K2XdcGS3sq0g2swrSk6IdJ4+aODxXq7znW1uCV4Px
sVT98B8YTW4bPlgQh8U5GjJt8PhHsjTenPxVDa1FYQAT1OVBoJ6rsPavk/YLEzcKPG7AdNN/iiPo
pi3PmpxUllxWoYZg7xnpgO2cg8YrH8qXruKchh2nSfMAExUwNu1nC6JjZ2CJ/B0OEqhk1rHvNZE2
JJd70Wz9M2sFm64BHu1RZ1nIHHT916OfqlZOBYb2RWCvxAMpVaWjtxnetxy223LOkaKxwZzMV6mz
AGmGF0TWEsQP92Mf+0Kw1NQ7+UE23dgECRlkJ6rgiSATTnsLAF96OLQA2QhoRfDPYuEB7MwJtMoZ
h+BAkcAY95m7nAGwv631BxvzdWozvVuaXkesXpv2iBDcbGwQCHQLH43eSYMMQKUozjllg4DzOoIi
xaFEhMtKrHe6ys1QTB7Nwz/oRU8wvqq/MkR7NjxuwTdEV2Q/DByCCzc45vxqemoE84eN0RLG/1li
+oMgfQk6zluZNx6bT9zB+JH/XGJ3aWWZsHLFVKPRQNDkyUSpCT9XtWb0Pnbvq0+PsUmQlx3V2GO0
YQDtFR+7XtgC0W2zc/NS4hTYmsmOBaH34HufDQDHoj61oNrqUEFqX+m/9Hv26BvZial2XxecVDNa
3ZLOtO+AwY3FeDvgcQvFKV7bNvXz6u136I4ZfryOvQCWHjS9W5npDMrSaexnCN8IDSh+EszEfDQc
G1gSA9fftFBTnamqyYd2IiaCGdOcl4IAUhn8kAC8gYfnZW2wRiyo4trGjyWE3+Es+Qfp3JvhzrFC
VYGfBN+LWnunxbRgHW3eNGYIYJNyu8CL8NYcQMLUT9IRUptX9T5iDA589cTRoWlcduIp3LH3u5vS
1Iys87R7mABf3PxC85cGAu9OSrP5pXq29/qQuxjnckml3RlkDwFuPiHG9XkJSuHpPujK3xgveRCL
O3kw6Z0vpY8l3dTAKjgvbLIP2+hVOmeMRDCZ9fTaOe55J4DbeycSTFRvoJ4Vv9rBJS7JlxtPyTLa
TGDjJUR8yeTI9thvVMnMe43X/d4oq64oKziw42sECi7NXPj9L0nTseTt1oUhAIlY8z7lRjr0fspi
/EszMJy8S3dW3Sob4N+T9OuxlnwSCqYJPmHQlIsf9s2G1pLl6xYJvANQu/XzL5PGe+KE6V6Iu5wA
oCxHgxVjncHK0Vyp1QR8+DAL0Cyt9SsdSCeBdk+Kq0Raa1NDH+lyABsc3x3F6gjMVUGELXeyXk8y
9n8PdUNUco33SGCkbv1Vkh3XnX1II+7DmaD+F08r8B5Gs41pXna8LelbMMxiJhnKhHLXQOHopT0S
W1VVEwz364d5EePQf2G64iV559tHU6zBgNrRWrfOjIjZYqQQt18r/c6S8a0HLYeDE9Y3OQRpC9uu
zGlsVo4AjEMw5+Be0gXVOXjdT1qOQNbCwfS7Y+7gJgSE1m6pZ1bEvvsRLIwM7c0O+NA9RQqUR+Rj
rnQcqdObWwxz7BWbGm+y0VE7zPg249EZ3RLsaOPo2Q0ON8dYzzZFgVUwDnWFXKzz49K6OyjUEq6q
CjyQxRnO3sh1m/OAPEoh6nhn27QHQAXpVjpZeZQUL9cs6bzbZma8LDvaBXcotp7c1tFb2IsM8Zem
9PqbtBKj0UWKwZ8QJgMzqIR+AuMLMy73WDlvdKzkT6aSTVySVRKGslN96MgkeDKL0dDFnRNY5g5b
ERv8CrSzoGd51R4T5PHXvc0Ms+P57QLkagM5IQ+EAlwGHmmd8NH7m+Dzj5xKr++Vbz6tZRXnu8II
vpodNOkwkWgrAcmpwPpQotkPW1z9d9lXMaJxhsfVTHJ0FBk08KJuvWr+UrWUkQE0zwG17b25Wlgb
dw08sIg+4ZiSaQ1QV3oYpZlNz2OT4516xkPOZq9fpI1pwFEG5o0K3tWP77WlKgibBlZq9t6sTWAG
05KFB/FQTyqBodDGF/gcO71Llr2ONDfvBcGI/cg10k5pu6ZbQqvH2tayyQJ+A9mpGFqIuKYTDW9+
4jBdPRz2D4fvZR6A4ztWK1gnEr49YsubBYnwRT/tdkIFzyvKAvvdwiiQHd9ggHlfwdLpkoOfFLkK
UzzsyFP3loWD2wQP9LenGt6un4e7jVxxzIuDmrZEAkjChCCEJgrF3uP2U8YfEg0rdiSPNONZWm2+
8gsiv5DU2mhW+KlLOySKPFLN9Z9/sm1jiJeOjevQsj0egNnw2tXlcMJUUG24wU1rMiUq3dbaabfO
4d7Bm4rsilW+4j3FI1SvuRGaNr4EqXqa54xttiCOreEJnN9dzNE9mO3403TfE2hO/KdxDOgjhjXu
59a9MsVuK817xnLMEFBXeqPisiw43ZHWjU0CErgcn3HYQB7Fh1kGyKpQ61a7pn9N5oAlHViwX7ZH
HSM3WfTxg4agCDb4j0bR0Z1rF7sexSqOvR+gZMjNyuhKzUQAcfrxbBSAkPBkEAhk2pTTt8rOaWGm
kJAFOmyF+PI+MPMqJvRMRCgQrUpFtfCCYAUU6KYLSp7mxGhFV8YfWU06GeTzuVF07xQHUFOhuC2r
lyQG7Vac0hnAnMBqnlMdH3qPw/09M04UCEKcG+vcHCjkLMBo8lS+CWqP4auih0K2G3LzLnnon1SK
fm22Pro7v/Ao0h0TwW195imXhh2xM9So6qOrrSn50qRMV9vD7fbbOuKsMDV2IcQkj1t1WFNqXzre
wxxcWVfv1g52AUbl9ftf2+CWh3DgxH4whi0s2gRypgFP4YsX/PxgTd3MIf3FxBOkROpcQjUOGKBd
Edpd2wrKivhCWo9dIgPnqzBP0m6KC7NqjsKYH4XtiR7T2loGAot03aWBWY9K42klrxC/5ESbGJxT
uiFmbfbYp/VTPPufvLy20izEavtIFb4TV7nBq67ZwaPBAVgQjTaXdGddTGQ/IhEWBuXv2o9IFYNR
ER1tNiJxBtvIeRZx/XUfWEQDmO1oZeOyzoHXoqEJ3+dwN/bAGm4MFAteTEHB4sKnje3lj6wWiaWT
wJRUfG1xRGiQh6t7965N3o6SyhIymW0/ce+aAbMBadPRBMeci5NdTprH7bbS97XeI2eAZqcDDiov
VCILZBTux4FUpVAXFe5/HSQEvE2pJkAkuLQJ3oBGPz2SC+1STZ3/aeinX9kPCGa3qSgV/MioeATZ
7jw4bIFOV1M9bvV7ZZAx8iZ3ekM5On/gL+YB26Kvzr/mft0LAFPapgz+3tPOR9lAN4zRBklgX3cM
yGke3F2UJllrBk/H7Ise9e5Girhqv1fWXFh6HkPp6YuiNTrJsuhC+8kBCRvxSuCGtYk4aSU1K4a+
naqR+RHUoV3eDR387t4hoWD6mnKonfUxTf/8dnP2V6KZZXRohatlmZgH6KhiJr5gICeOhMlyzCUy
JkKpbtZFTHDAS7WTxZLwaoTj+fXjWs7TfEy/aNNN+G66g+BxoyDSyp+EA8WpvbryDwgOvjvndb/8
BRwY+mGDdSbQS+w0ywIzAjgkmZE7KzTi/HDc0jpVWdR4ObndnXBv6FFmVI0XsZHMufaprdE12bc0
4ogCGSXYNS373EqmtzZ207QuQaRUzw21jFJTUQiZALgtUkXMWLJDIVMOraeHKAxLJItzUL35xzqD
6cCM3mebd7/TEf7k+TdcUSAmtQClyclLS03srtLJs7Z2VImkmxnrbn+A2ioOn594yS0kZZegesBC
e74/VKbpRoXBMlcaeffigDMT0OJa7vQ0pywuz095xtVi4VnRH9pwo0kn8rmpXpbmh+rer+ULUr2S
fie4X3SGUV8vcT7r0dzTjZ7lXL8lILFDQa0I/l4r7l071u0713gvP90Ixb4W9re+wNqRuxVG2lzU
cjIbKdEKG2bI3b9nSYC5MArOUQckiKjO3aPH6widu1DEn1aO5jnq4OY1+79vtwA0/VBd6wmxsiNi
oDkyS1ujYi2a0CqiETMe9QqFkZWiN30oqwAKBeHcozAieo9X8qK8vQyLIDwFps3HynpTIbrZLAJz
uddsK0VS8qVPCaIKJtSgfHB29a8PE+6djM3lrJd6OTkSQFu8JBIrGoravhWZDr3UeoyagacCU2ur
aMVTJktGhC8JNfQnVGhv/I8KOnG84vslrslcId4OiqBVPwi7G8gVNd8aepYtKqT/SZridjP2kdLi
9zelU9AoQlouXNlyQDzCkL1jbjBZSPgrb5dfijscJFNKGDcrTNZWANplkky/bNaQANkr/0hM2faA
IlW9hhiJ27Gvh4AhWebCoKU1/kEE4san4k8yZrefpqzaZL8aIjOWekK9dbILifSgetN5o23i+aSa
fI8gix/ARvDpmT+VlVfOHwvywFlQtGapPM+2mLAQWouXfN6IycN84t3PhMsPrjnYvQ5Ro1PYD1jg
qiKYNwOwUPSYkJj9c1pt6DGDA4JEccwVtCxEKeF+4lPgZ6+nwTozntRUlXAmiOKmF6RUHgs+slfD
OsHkf9eiQ80fUJyFMd5sbWKh4J2XhkMcrGrF8A86IgSOH9JSvX7k7Wjz24FVGZQ+RhUYFaOC938R
snwFlD34HoQA6behQ9Iep8/NIiVUpB4UCk1116P/s6E0biOd+Vj8AyNNLUlbcfI1tZw+iPBkRL2M
ZOAc9Hu58oYdXlDnMwoyqaIBD76wZPfsL4nUfu0IL33dZdlZPAZv/SqPJ7sgkdeq+Lm2QNuUKxG4
1lsA02u3iDr2Y4Js5LQA7o3EQMOpoZn+81h1h1OAssgzw2zrsfttRY/5gF2tvt2bTSKULE9RrEDz
syxEFxnIBtaMa3viGMWw2fQ+IxWlEEAkzcm2FLyBP0b7k6cdKpDBA9MnKxbEwFBLXT5p6K8XUSKv
4JB95VuPQhzRKNk8ergRFOCw+ZW1OEAfNIgoZ4KreKTYcxgIunNnHgOQBTofpNj0H6w2Ir6rTcRE
mLz4V+8ySMbOjbi16FRkTbpBeUtg5zJbF7VJlVmhObDQOR8vBJ6cZKTHteS13aiTMiNHpZ+LG4Jk
bN55ueA/Nno8tA9BkG8AMZT8QlOrCVF6B2/mvMihOz3kuZBuJscDYt9DuJqHgRW2S5We5abK744s
t/eyKHYUYxlX9sy6VSiQXK7I2ZfXJdsC8FKD86VizRqB72S5WY+dvBGByD6RHbmy+BE9e6+PPaxy
l5F+CamL3l0XtSzvepUgtcVDsqdQLEMWYJT+ANIG2Ki92/lv3q87mm7ffr9odFIBMZzbL9uR9Ybd
X8YSKZIAhJASvuzEq7vtvB7r9nueLEO/t5O3aLA/7Zx3ix4JmDNWgGPmkllFp+Ip7nlXPikZpVXA
JQ2ZYQvzdRi2wZMldjOK3ufwAYR7JVj2Q10UHlIWDTCKf3JGfcjY0GEPvEQlBYrEUE7je1PRz87F
nRVFEijavwZzwcmAPdS6iAFJSmZGVdy6cbejb6CWbYTFbs5v34ZNZweNmPBjI9zgoS7bOQd26gtc
k+madM8SYnP45IwRx5wvJZwfvswXPwBxBlFVHpjP4/PnRxkzImVZqXmLF90B1I/sfZrVIqlvNBvA
tQDIt5YczsbhD1XoKsJIcq4vt72VTZYg+jnBs7qwYUyHwqUF0AvEKFBz1btkDELI4ryGGm1C3vMC
fBL/Ql5IeKFBab6Xu43tFboPU28PRzy9aw9VafQ6IA+3FuxCRBOZeiCdA1OnfHmZisebJNFkAXER
ik+scaeozuMCn20Ejind5t9splXsGSN5/QwGltZbl3x72YVy8UhBziCH1GsP/tQN5u27cJR1q8e7
DzsJGRnW93hFi/8AQ5nux+TrZ8aWDefhxCM5pfukCq5mBA5zrrwOvxVAiRXEPyk3XwXqoBAXU41I
DosXK6lNB3onWP+BWJ+szQH6f1jYUl8sE7XU0ky3eVBLstc57lUQ3XjpCe9WmELXpVPOKTA3Ly00
Pc33GJd+7erRAVlJZRQW+ovFIx2zzR+VLplAQU3xAHCwo5rS1mqhJJlxGOtX1y7gj4QXGbnqaYtt
iuDfaTj8ULAWdDfessDS4x+yZTSgsUlSomKj8YqpfoI5O+80yZ/rpAy4rzNmV7TKsKPR1QG3Og5+
4lzPyrtXwktzN3Bue90KHdHW9DAu/3IPf22VOKOSe2YX5Do1gL5sS6kYkmYlLLOcdIPw0z5umaYg
a6n/UJxz+6I0rnEj+pKxXpQCi5Gb1/oNmUfz4VcYYoFiWtGqAP0Zf8QW6TbFuB2doD3HC+9YiHQz
XYhcYEB45W7vuEPIjXSguRwOhRNF8n7KUh1pKTi7myxopKdrQPYvb6jBRXILXamjgZB6czV9rov2
QXP+uNiyNRJlY75SMA/SanegAt3D+TpNfHAeQzUqAnVaZAiodZou+QWfaJ+t0OZmR+mWhH+t5np9
GFhZixsoeq4lyRVCr9yp18XinOB1FZgeNTKncLWAWzL7YmFNceDmK+d5caBd2GnpkqPeXwXZmn5U
m/u7/7WzkeoaqhnNCiBNwOcQC10GXx3EJzAL4MEgHm2potYpiGVtT4Y0dA55dKSD76rmydUUfRKC
X6LPFyhKbynRYEoblhHl/ILr3lMsKxoV2qaGmXMzCVXDwvMGmlXQ1DGgioCuh+xBcNJXAaYeHs5y
BmBua0juVVS9cp/8UHKyC67vKbuPkfHS0OkzbFvUMe6MLPeXqTDf2TFDulzSR6JacHeHnbEpI0ew
dBm+FFLvLnegIcl15beq+PhD4HOoBNmJ4CvfZKV7K8RIG/wuQZq0q++rqUrdcuNBQk6T+zA5iek1
WeQ7oOF5iC37babS9lgjkbbvik6kM49vqa8BgfvmkKCV3Tpo5hr1ot38msi+u4WiKdDGqILvcE2X
DqkxNM2Igs3tr35G7TmecEXACCyL/vHvNsuisqMkDhzizLy90pyl3l+RRD4sDKamrQs/rtbP/VGc
+bfw4TZtoD89pGZEZgiyLGC+/Y7QcAJETUUBP+/Rpo33cubdDXOoyn1nSpTEMWVR5L4pshMN9hdv
2NaQls7PS13185ZHajUB9NaHOqFlSw5EEQtuJo+7J81s8dcC+jX/cjT3+Hde6y4D2xP56UCCBDW7
I8vw9WPao216UJ3hOxCBswZkNRDlOvCMsg/Px2fumgpI60sAgAxKC6F9jXWSQNpSkJFqtquDLpwT
2+gzGjftWn/PaFAbJ/6UNhkbzdj4ADEdr+WU/Sp8SG4pwwr4PobYDsAReIpp2OCz2Up8TDGbINp3
o15nn0TOzortmdxkuo4ASOE//7TOQem9koJ/WEoFgv3Lht9HWdv7xaBF04sdvp5OF73xJaNVhlpe
8RW+CwDD+DG1VxWfREE7/baxqRO5JIdc4f6ffDqUWHyBzyS8KR4NPVZlULCsu3O7ri6XJwQKw/R5
FOeSQjs9s7B0PIeslVoNaSzTQieRo1o3iwiqD9ZG2Oyfa2nyeP+XdLtfZsIvY248EZOu3kR3d3C/
53Lkdr/jD/st6T+hzG1auJtTaKEJiLagBXyK0VcWEy4CD+eKXmti0KaI39WDJnAJ91O6IrGhfEko
Af2dFknZFWrQQFD9ujXQeFLzajzTMtAxafeKpMUVtoH8IemqgppHsbQV3cThw6iGHmP0NeYpZIu3
XkrRrpY85UtXqmS3SHfpHyLgdpsk5AnWxtdco5LHQW70qR9UskOiJPqd6O6pawnQUKJPzcYHGqBE
ibDFxCpS4pK57RgkqZcaHaAJX72MPu1qTscJinAx8K/SLiv1s/QXkKqkW2ew8vRjAAP1gIzfixov
3wwgjxlQo5FSr4xFPSxP0iuE/BkYLerTxsfIgiA/8E/2NXa6slYb572ydLLHQNEMN/ZjfKFaHjDT
1YTkYU1OXX/QqIvc8PKfhurJWdSJHj7O22zz6tTCBTGYejLny0SnZ0/3jcSY/OMEGhh8+UJWYptU
CqlDpjr2L2I2C+/KeN+ZlQo9jGdDqnzticE5hKb+doGpUqB/T/qGbpB/DIubkxRmxf3xnmEhVSuA
X3fVcG+8jKj4wfElZ3eeKNIjxAxNNGmyRetVCNIoOVb5sV2SYEmly38jVeKC9YPp7Znngulj4WY3
2jCPFSxUFagtKpzeuxGzKIDaYm/TtGtOvCidJtulrNU6lC5rHT6lozOwRp6QHcIZw8PeeUeU4CVB
ChbIvjTLh20bAsOw1T0ZxBQcX/bW/q0u4zZBiDTu5whsf4C6mZqaBgi2PAaZHfS+cBhgv6srnosa
4PPZZLLpBoOV8UOcU5xN+K0KUwtHEko4KpCO5Td62QSc0Pv8anBrVtEu98X5SCDeAltbrmeu+06J
SJQVitwKPajUQv4g3W+xY3JxNxQB4iQ2UIFmWZVw/HS3yIQrr6XLKwW5PR+ZrX4ayT+1ZDxckftW
+iOJb9l+An0/gC1rnYgcNsiVgHIFrR/W5amFd11JGAVM7PYf2U1jM6wtn5TqQnKv5mVcIi6bEEvY
VZufLbgLe5fFwFpmtkiAP9YE3dju+b6vnoaMsW5MMGiVKBUjozOGzdGilovTxp5pIWUc+mO2Fvxb
aqZwTaN3L0tN5e0tZENcaV0hIJkjLjdGWzIT1V44Sw16Xqjci5Kfz4UAyvvQm/NawVkZyKIpttQr
I2M5NI7Sy3YV4VzWweInZRT83YwReRLbu3tLcxYuykcpmwNuPiyjjM1eaY5RB45++5r/5GeIaaIV
2fi5c7OzWumd7adXyu8IeEnhzyZcetPFNkitrR3DJFZFoTh+OjuzCDOKVZ1BPNrICTdwYMI+zmMo
5g0sgN8MxxJ9hvcViZJtTcSbeKpnoHTNPcTJpI1PwWrd3PFrAFR4ub5FIlNIc4Q8SoczNeXKdLOJ
Iw39Q4k2wEOEnjZG6tgZckc0fd2moCamDBD6CFwWeu5OTHiUQF/3qSJ4Gm+lsLpxZ6PGLaEPI1FY
CcQ6j2h64lC7imuAley57QybM0eBscIOsFzaP7s1WFw3krBGCERk8/xAB9tZ0FI+IyjTpcwTx2Eo
nMF55HcvcYo6KLftOh3CGHWSfdzLPzrnWuQqdG9S8LzaW61c4l0AU7yqOOE/PAO0IiBtBVvKHJce
O0NjKEyLtYfhhRhaGMi9ApLTAIyZdX9ok/IQhAwUXQcDHFiUuugyViL6riKCXx2StM1/WpLwZSz2
4rywYTbmtIRdjB9MG4WueJ2HFOow3qkgMRhaXIEVUeeCS1Y03d/ybzh5gu1MgRHKv+2CU8o4WVgR
/zWbaqi6qrUJpF/YJnbgzFnTJEzsdvmRtjYGuzvfnEvpjjj/CiqhyxC+cZ/2gW0kEKQy/ypmbgYy
WyGfb4YCUNQu1G1t11mu/Dy69bwwAen+KjIaXv6cmLzhSmCSrIgI0v5FAUbgXGy5ww/Hs+9WdRZH
UBjRYbC63kZfqmjHHWq4EwP0kqOdWhyi67T9ViIQ8eDFQrOug8c7pK47km/9ZLIiKmZVItG33U1m
fEQKcFASFlJdzrcF7aQDD8n3PvZ7tPiNmAtdql1Etvd26rzZY7JgZtccmG3Axm8mjQSCu9UvKbjg
+vjFl3M8BhIW73ELw/s5dWr/CgYQdPdMdzJ4JUa6+bzXSFUcxr4Y9sTOsyC4h9tB5r19oFLq+L+a
J/OU2ySNZlCnZ1hK8WByVmbAtyQkhGU/Un//vAWHWYFyh6+90QKmng5z1kNYyKnnSS3UZsJpcoHG
6/Uo2T6MoeMALPYDwjakFRg6QsEYNc2eUQSY6Zy6GcLTubKhYlQFAdiGe6YQHGetXNODZdqDIAh9
5Y3mRUV0YCCIWdyfbu2Zj246eWojlc2G8uygQnY6la9gUJTe8x5isTMIrEGEgPtDVTHjus/rkG1A
aIrh+vLeueAdBs1X6SXV8ZNx8nrMmUu9HJYv7VVH5b+/37vCfwJ6xKxwr2GeEuCIoA6nRJd1FTHd
b8SQQMy5VBLevgaqGDMtwRQ899HrYvGeSureqTT9ZnaUMXzTZHGZwmFEQVgj9cDNwgA8sJvGQR9/
okQWYZrSCDHOwmUrbODZtCiOjeC3TvhqA8e53nguceThaD+Qq5ADdj7R5Wz07dSL0TU0PKlpI8ei
W9RrPR41QuJL45+PcHZ0FdDQ/HvsF107heUH8MUBvXlu2B0U3/FIuGcVHW3nnz+q92LcjUXvbjFO
IwvpRuWxb8EPaPu+Ob4hoUp8YWxMwFYIm6GL11Ao2BIMsHJs+XpMzC8bRnhabFlKpqygti2ux3J/
0vgBPc2FcRx0ZsyOlyVbjf3aYtxTNGZUyQKaGeuLspnQNwvPBkaokAO0voRh4wnAF1KKNLVIJOPx
AecJCEkCyj6WrtZffMhuarzmQcWTEf/UgciqHuyJNB/VWtyoMb6tf9ltaU3MVWvomdVUWatrW0jZ
2C+pv/CAHz9xmBeBXJlSHJgEoqhIqclYBAO4m7tJtkWjPidjdTY/S8JkSW1p/yd6jnNQuz1Cm8lK
29Lx6WE3BE7GtGzEhJPT0YGmulLmDcQQGPfv3ZZYYjRzS6Y1sk+mvcs/YRZ2ZfZAp+z5ghgeKYIg
uj/x2iC+/QUNz1nvf50QUgNpC/1GBFDi1G5HHW4WHFHzjJYIQ9ysfK69iqtAy6O5YfYugh7AuaHa
pocAqRyj6kTEmaljeZ8to50K2F9fIAqO5ePjcytE+mjpgua/++8Cqd86ZAr63R7vVhR6uxUVfCh2
GbfbtcfFV0nUqsbRzyIhAL0JA4uVxzCG5luDut8Z8eTKjWmppEJ3H8AIZy6DJsrMwuJ0MoQKXZSw
D0xI5MSNiYVAjTVJOXOvRGE2PqvtFfI0bvGZAzsNIrcwhrtnaNvZrrWRwDjTR6v5c3dI3b0/xzvj
AGz/Qesb5ZpSCzsrr2qjnDBbr3Y4lT8J83hR8fCuCS7+uZYTpTii372cbDJiw7x9yBUSPhmXq4yE
ayyTCZ6Us4dULDOFwvnWdndBTUlQcUom3rXNunx4CJhF3feFfo+M78DLvTU3QuyYWiAav+A4ZJho
OzCtcIqCkvPA/5J7PNLSfX+74ybClj7HGWBxnB6qJxIIzKTLUflCz9PSelLrt6o0zlYoVrmwKI4Y
/ZlBd+jgVaCyttTTF8PxJUbNn/MIT0eQQslIzOcbY5DhfZgRzMvqCAl92zQ4LVNGVK54Z4bn22pP
soA74UKbFvF6mSsyGFr6aNXmk7xnlAs471cYoyubgPhNlcrEylXDXhs/7CdlxeT0sFjdG0VCAHg1
bFyHWav6pQiT4slW2INkGz1Xxta/rgqoRUBrYbRG5TZMc0g74gVKuWKkkODe+ypYlKuhCMlsDmJ5
YF6kDhU4RNm8HeIMKkDAlLpMZGdNpkQpE4DEBOxStWJSYgkza00oCVaLSLqY1uK1PAIRq5ZFfeC2
bpJrbCJ+JNgAlZHfZNuhikiaiEpFSdAmFZPIPekGQfEVrwBqlkm1TcT0Q3eKplbSqP8O5EWXlpCT
o0EPSs/IJz5q4anqeqlqLL25AT8kViW8sTzuZParoOASmUA2cmMcmrVT4hjzbVhgRCMD0Xxm/tzY
r7aXTT1+ah0o2jNJzBQgO5T8j/K6dEXgYMHbAKBkjDWQAhLqNYsU1vQHG7l1UibUIT/GpsE7KDWU
wijANPfFII3T8/Pv2YII09hQY39sNDeyB62rXY9fM4BcozpvOXPViR17q0zMNTToM2coa0/fKtmc
pg1JHk+oOKIYKpSQfE+vI5DnWz1oIqkGgfh39muktqzO9cK6l6Cn8WAlfhiKdQ+MgYPhYLnFJhYX
WA1OnuSpfNtqHGccmaYU7pO42hrW+Fx12DPsfTT0Wjq4+BesuVrOsTkVUvcQGweZ4kLISXTUTLxI
fKl+t66iQvwYnPNi0RoEHtwnDUGmwDBFyX7m4xGUYix40hLg8kJ9ALQmJVeJDkiyZIvERQrxooyC
0jJeYevQmoM5EsYFd1iNDHT7nevJ9a0waA0+Hx2RMuCNJic1ZxCZ+sF5gR9k4juXlN2X/2PxSmL7
VnowVGojJMyCKs4UUbip+DoiOZJV70eMjdAO9/93xKfPlDAGIkNOtWWUhOJWV7PQa6a1ltQwjZ9Y
pwNLskTkGXe53/Ve4NAIQTNkn5GvgWcL6zAuLUsT7noExW5Bgppj/mWPaY3Kz4hknLY4Q0KGaKqG
y9exore9WtyMYsjBwoBPwXA/TuF8hBrCv8Q5Pl7EJIrbEwww29FIi0QhWwT1tW9rOZZeSHdJiNiK
nv87OgeEVoF0IcKG2f8MvDrGJRtD3fSVgrtKGBNbfmJNPWrmMFzLnIU1AKSQ6dRmRm7Egs2b6wYG
cBEvT0IVWNjFAs1dwYqijIaxe7hH7OPTjvdBJeynU1XBuPkh7YJFmLsvv7QNCPJb12o2TGh16arF
9VYkgTrMBDaV8ktRnCozeK6FMSeXAhDPbq2p+w7gdAZviXjuNEGYSUCmFWELU5xRm0YxbLjUaH4U
Hediaw/3VQucP/jqr8ZMcIt8QhCd5JX0YwIbl6+g6AFjvuSropBnGbgrySwn5+A/V6lZ6FyjwhBq
aKaXZvrL7NXQugt1uJEFPyr5EuI6xP5gs0daTtwYlow986qUAxCmkWj4RLL/c+g8CQh1nMZwO8KA
76zNwb5YGZODQ/D4EhQF7YxLS9MfkDQBHyShtxLnR4rZEcCRfsiIVzdqugDnfWQbJPNdK0NdjAjT
lQmppY0iuW1Kj/V3EKYdugSnJ5nsab/ZRlvXhusbykiI+73QVqLce4aMeJ2Kr5beA1jI8ozXoTLi
t4aoX3dc4OX9iDtn0wdAYBk6osuT2Goc/WWwVuiYxNZpes9n0ar2BdMRg/mUdRq+c7LQNHVzW7xw
spn2Q4kB9CAKoMh2evhnV/GMLV07Qplw8fgAuNUGi02KQyikkZ+A4STcJWYJXUjs4Tc1p+Ng/LNy
hFvjDE6K8xx5PvYYwI+hrTYrw78duwyD+i54L+ZKaq39OammHt5+jNj7KhWSicsMKjYGalQiNPDM
UyziMqlIEAeb6j4jqGxM+dlOXJtrjYskWVqMGntivyb0Q1bURPpInnq4Xc+j8sqYCo+khAwVuecb
3Afz/Ck+/RcXNyCtBZED6vbfJ7oCPUoQFiGj4so6nNBnHycOVdxqOtZhBwy2fOh6O0DJBlFAHYl8
PIjcF1FUB4iLqMLeKCANRT7Wby4KVuRe9j/OjEL0gaG9iiGFHhcBnf95lwoqjifng8Bp38RLph1A
4QlWjG4jj8XLc3OgI3lSmNo3XihDGCZDWAd5arqQuwP5zRFyycuWwmmKxJ8YhNNHKvroI7HTB7BI
hEGyOjPYqx1jrNWzDR85vfqP4vBy89UQbk8fOxPdW3YHLZLJI4zhxJUV+5Rmbbhfe3S1DGYVTwIa
+XN5u3lF5hHWKBxvTdylCQzqGjLvjS7xgVNGM164JMsvj/K2BXOxZ4rY5G/jHO9JhNJBevpbeiQF
lou7Nq9ibPRGZWhaBpv6ABaRLWO0P/CP+I7VivmNtivH7+Ni1Vms16Kh02R5+PkzFBnYkr5soXs6
I9TgqfK2rl1G+lZYmfhK/PdbM7wkU5hFNejiJiZGW11ts1AMiIPArYcD58vCBGGebY/pZtJtdl/R
dm6XT5jyUtnUyUNzbBT0/lL6zT4XA6x/5VNn83clhivTsEPIPaZ2dJ0tM8AoCl80lBZlLAC488ZM
28zqgkweGpPhF2EuIkiFopM/MfiVB3MjJVlgQcguVlOEC7KKRauLX2TawZIinjq8/cTmYgVIkRcI
vItgllFBERQ5FzTqYPFSCFxLdruHIBuAxL4C4zPp9WSAAI03reRulT3c+bnWgMD+/79OZKpBBgzG
CpWrK49vce+AwSNKw9YA1ZgbgbuDOQxDjUTI5PVwrboUJm09l6VbRyXQDyRO7e5qB3ZTX7u+kqWp
CojNTrdeY7MDv1u/DWciBeI88tCfGBi2ZZ1zSbPQR+a5YkBWndIY0D7L3zenSYw6mLHcWfFr3rpH
jycHIezYXtAo6nBhNDuGY6WGk2IHj6/1cs7pK8THw2JbibiosK4zHR+a26fqlykIO8qSeaS0LJxb
meC9gsVkCMPUd5GqR3yC3pLuLeynYvatZ+Kw4q9jhNbXTq1zjymmWc0tu2MNQBz2oFrl3LTvdCwW
+xra9nOx9w2TZPDo6FuBYhYqqgMAo9x/7lSC+E+ENlJFVWkyZCYZnEinYHqzooF9WGyXW7qPLYyV
WBv9PYju8pHhbYFk0/98YK62IjgV5J+UtbhbLe+qolQcDuC+krhU3lWMO1to1Du+Xob70zMk58XY
2oC8OWVHqax23D8IY2FeCrokJ6g6qxPBBoyxD8MfIs//HHHPCBk40mvUmKv9twlXaPciSeZYrYwg
tyUiVxH93UwOXgxrof93WJpXntypS7Sb8sM7HJGOAK+UHAnymr0AN6xReIjLUDJfLpA1lr4+rg+f
JoEB8Zkx/xNhpsk8CW8Nlhvy8fVApUpajAUPVflcf6USQUOZ6WtgIytzgFLgV31H55tdeWDGe/6S
IxaP2C5dhaKAqoqchwfLLEXEEWAe0j6/H6J6W+EobagqQF3d1lMRYmKYcS+NKwHp0+CaLIX2YLzi
st8t/eCNDEAlRB1SochM24CJM09AmpG+d9OI70WC7IMzmdCXu0V7lq1VF7cSfovwx3G41dBemGbQ
sKGasgFuOIqF1Bdmp0tDVShKSj/J2iYHT6ayP0SBCkzj4nCXg+5MV+1dSssWKEscejQ5WuYPsHXf
aMiwBeemdJWnKt5HefyKfs376Y94/iBDZYCFdV6vyfJJ9oOKGNYa2LsjAG1UWljr2gUdoubSJJzi
3IC6jzjzaRNMqQ+WIWlK7LVxmyVj6aabjl+4GJna88LRmzRMvLShkOvd2uI78V3Qztga1gnEqQak
0FHA0R/EI5fq7ofJX4U8RSappsJZGhJSylnud2eiHVt7MpVQAmWzqfgM47qUSlG8Q6K/SuhWH29T
caqOnK0YiL+02vy0nh4a68/n0rkMKUKIAfYi1KS/Z/tckMEq+Bc6HNOH2YJy2jdDSgdimuqyVspF
KiD7yNQyJvDQS0TEHuf5XtKeQFUeCloYKyUNbAf8Glw0L5p0gLBbOeqatcIokV3qRSVRu0O9z4qs
wTiAkjVZEER4N6e09WZCc9sCrWRbFpEaYBYCxhNVK384Z4aoDq0Ykb6744JgygmIcYEzjFeFuBvJ
wLZHhdSMqpnJZi7cZDJ49lxarQpzLh8L1BtkKJwxdgR3vUvd7L/sICz7k+FNQu6eD1ftfVA+hPLr
KPCtK6w7v7nQTADVPXoNGrDLSEwHVw/51z0i+qq2pC0m4Aar5kEOVyQHtA6KQCtg/4P5w85qlb/8
1RUS+Si40D/qRlVRLrmTsVbTRJRY8VWU2z2/lvbe6FJB/K1Jow+7AEzmYSuVfmaudL/o84DqRUac
l4d6aXRU4bSYCyrFAuB4brLKYYMhHAjl04Yup7pafShW50lAHe8poGq1G/IDTcJf/rGZ6Gnw5ZfQ
88e3X2pUJJD6p85uKMOfC4soxzVJPUJKmh1YiOcF6hWLpEZ/BckbbqxOWCkTDKu40GAEi4Z/Bj7S
Gq4jOJA8Vjfd3hTKL68JM+o/ym88EbocLaiVyLF0+9B+8LEg9Fxc+PstHs8ZHK0ljb7b/FUOcebM
1GheMQqrX9WwVVUfWCaDOZR+SOE1YhOq2u4VhzHkVrQ3XjdM+BuqdXNS4dLLlUi82jLfTUiGN0gf
/GFNuNBhVbmcj7IUW1zmzl6Ldy4xuoBgp1dN11PwIqT6LJtrxIgoc5TdKWGgiq/H59BNcRfFywEZ
UJqnhS3cp+jK47kF65BU+6VRxHbpJN9MvQXPt19T6ArmXGytOqEkgwgwZ62Q+zvAltIBf+GmXdhM
Lx70kuUowrQ0hRik37Qvq8XzLQnDnYOjhAPbIlZUmfjnxA0Qco1H8Z2ubSpIC7jbmKdkQO1qbd2p
L9iAm6UYbkBP9rHtxKccWvp5erO4o01IxaPRwIzf7NWs19M2rRqMgy9RUyoE+TuotHl2+jTlCM+N
H0LL+F/LxncnUwMaLJImV2+AEYXTsLsl0ue1nsQNYiQ/oej1yVZlup1FrO5xDRMGzZMGYuSZAeNM
a4k2cnYw7rOz6/rrQOyAymQu60GoLgDVQ7qU6EnNhpi4u/9IKvImYfxUealj+iDZM3hzp/u7fc/4
vgDTjk9cOJzrsWWRsk/kZVT0Om7KBXC0XBBUWhdfD5178uHjY+GaG7ztQ64hMS0UTQNosC1ljSp3
w7b89V3Uwpt6feXpJGGUXpc9ABetwEwaPEUoISAlsVDG9rmKAX1wx8x5Puec6YFHAZGMk5akWuO0
G4WglIGY1cWCRy4LW+5V70MnZfZzlAj1NOw0iYbtHcg795sxz0PxLyQIiaSkCUGp7yGU6O5aexIi
9/ODAVKh4hLHHw0XQEXWB35txix/zO2PNHKmp+e6G57psuSL9+pbMHcg7E7fvu/nuhwo8gfCzfOg
iUpD9Iq0p735l/Y96tQ+aU7vqwpPEhYZBadU87gZdJB/24z04ZZoI/Wyxbsp/MUXut8biReDmt+w
adG4NosvRmoTx+3bZq/cfOMCnZvhYYsA11jBcGBrSckb3VB0cz7AYxNzp3pTcV7tT8MWRSVwyjh9
/Gh136o1OK51VNBcte+FwF2VxHZULSmdKvv8sM1h+ZAVo1sSX1avjEf2Qk3NjHo2uhlddGIs12X+
xpUjx5pW7Us13s3cIlLVNnkYY3LmtpObikQASCNe9mytwxy7NDe4kibrUizwbhHKF5RbbTv6vAL2
G+HoS0/ZA8o3XgnCHUGZDHUkK2qvcxTI6GKlWfvAn5i2XGxrkavGEkTe2/ufRBquBYOnvBKBC8EO
MNizQPsEHThfXFbcNRM5zdDtj2uxXqSpJqHd3KJtNS8eVEhjpezDOIQRuuFoNDt1NtARB3anxmxT
lWK2sx2wN51gWp1BHM59ph5ZvozF2APIwtQ1Nas6e3nZgwDaac6CXRrzrRvaNuPWF8eDLiqKCR9D
j4j120nw/Q036TSb6Z+Wwigpg03vw+Iuh3Jl+N4vb4P62oqn2YiIB6u3P5WOBefQKY/AI31FHZhb
YnYpdDSi2ML6VmeaxjZ/kfVKhHPyiVk+8eTlA5BnxXOLFJT1NdJhoZrCajZoG7+cCdYQKejjBCKp
5k02Z0qZEAfIE1w7qJThd1wYXVQukqRfK+J9unSjLRHmnLrB5IqQQmMVyYbLi8KDcGVxmeq8wjGs
p3cst3ehMdxPhbI4QYbM+gmbodvr4+/gStdBy0rYJcuNYvgG3zpW32Z2cAkByV0M5au+8rtIar2e
QmN1psU+VMbCbxCAd5OJK6xITcW/krSYERUX8wLiUbWh1GnlVdamX0C493ZHFdllF6RnjNcL8KVn
RjRM7mBBh7lPm92gCrtT5/NVS6HGvd3hgYHkEfZ1hHADbbFCl8fwxhjdibDlwZPZAzebzmW+mMBu
QGZuD/V/8T5TnXC0mSv5x5AgQTCYgEMwfGTZ4sVPROdGk7f8y7YhES9Oemv88tGvgBrHhIDKPCIp
xBZ+FbpfrW3tbpp7LOqg9Abc7FDbZpz+JgaLvzG3Ugyj03l8vLBuKJEF0y9SZAK5aUbFYW3oV48r
fB82ltLJgkaFpRqEhhfvgA8eumji8iq8ziO6RUEsc+asbjV11ur41vtm+3793kuxWWJx4yusaaM3
krxgrVZ6ls63i1zq1VRxl3YgWjCNXDjKOi8ACnW/5uub5iAsvShzkWEUhMvEOYtu82qYYAQF7r2R
ufWY6mb89iYYNZbZ+XDEeJPSYnYmw2bZquOG+KdBF0OnqFHe+ITY9gvGkm8Om4TDzuQylle+IZrH
mB1dMf2TR1kAnFRiQ/nhNOd5LWmYurWDD2cO5jDHgM1FHI578CobacihZR8NlTrevAw9ZEGQvy1R
zfMBXu1baBDeR7pTN2kT33sLeBAInxhhSbe+rQXZT49Ec6TvfpCmMoZv7pRpivV6cluJ7+y4PF0F
ysp47+HGa5Hze6/ON7rINuQhamnt9Viz2nS9FkQC99ETRdTAoOn7H/jTImmVoKjdO6FoG6Sd+vNq
Lz7Djn8DnO3J4MKYI//gS3p+1BCSnOJx9n8z6dDlJLxVctM3V+eYZ5F/NqfFSxr4KfAUbTt7GB5s
/LsTulwa3/WEV3yRiuu2ilnOfxVMV8Zf6M7Zo1n0ZGpkDMKdkRrvNjgTIllW8zLX0yvDabUkCn2z
YJ7EylbG/ScwdgsXewlAixF5EFVI+XRbpp8VVlSjdtjlEzdzWarcGI7xVLeX38/nvQrfwgFcdZba
JtbZAmB+x9s+LrhtItb7KVHQLePYhWvusFqpJ2ncrGpFnoxgAJolfS6ncvLwSe63RWoGu5Xa7Qfz
9fDXxEbcUgmr7EI7Do3S5tDd74Ma9AZYDkZ2JT8x8CpKaFezIhkb70Nr4r05faV7JTlrsDnLIniS
GX8RrPTaIFgTJ6+WNqe7s/vx8uuEmvxwjp7yhz9J/HJYbIkBsql0+dG8woA6k0Ybbec428Zd9ozI
k1e4tUihxwyY0vdxth82WD6xA6cI9o+UtlIFHRh4wwcM77UltStxGxV3Qn2lT7GTmA50ZGb4/331
tciDuw+8p7dWuPIhGDeV3jjkQayqVb7c+EfSBVBa5Y23HUbpd/K3FBGK9DV/tE3ZT1kzZHg8Ns3C
3luEgF/HcpylZzrCd0Gh6kJHwWQ3+rvLWUS+wdC66jeSNfaMRIoDhTA0bgt1MHU0/AC9GmStxSqw
Ya9zAfilF8eTeU2NrnqZm8JoHn0QHzRgYYaY0Hz5/d7TGmsGDxCMtGS1LDiBED2FqXcMeYiisadw
exBhvKCSt8oSo7s2l0U0vmIO3MRaZBf03d0jIaEqJJ6I0f/dwltxHVgwzvdjJdSRY6Snt/OnIn1f
/9vwXe815A4IOvk+5j1QUjR5QPY903xK5wUx2L5qOdrACf3E/2iiV930VFKEU7ajZ42yTXti8tOV
6JGRjICu5hOJgqIcItdAdX6yWAm+1ngEBWhmukhUCuioFMmFGCGf01Ws28CjlDJsBAGP6I7LK64j
bxG1oUqDle2QrTR8yzFPIUiG3iON7xEGYfa4r6S9Zcdd/eYJa317DA1QgaVG19mM7diT79U0/SqD
GlzZp+Su5Ok6gDMqh/4dGjELfEpJZchKMsY/gNHWZHZUFt66XFBMSEpuWk5tC7DIlSkykb8N0+9q
q+BVgsdsfA7Srp6khM9ZoLCaFNkvyvHu3zW06Aqi9AOJlNLiEl9WvYJCtja7fMz2DboRTMI3A/T8
MKe+I/ecnsFyhu8cO3/xGLfsY0nqFxG6gJK0YyuPu4hmFYxz+9ubETAGZy94+7Ye2VRA5RRya1t8
wl1D5XydNjV7cz8beZ6XGV4/CZzoVmPRhFfodBK0XArtANs597yHkQVBOK7o+StW0sV0uBn+DQjz
oJpNBamqjii7XXds6KnAo3deI/RhnRkRJNCYYW5MXI6NHf5Q11BqEceUCN2D7fZM7+qAnWef30zh
+XyY3mVGvt9GVIur6UgolEwF5AEIb8ao5m3gIqq0wr9AB0sv8A4I71yIIsM1YukBtCjBV+ScgbC8
IalSNPTLiDr57BFm64Bl5YjEdNtokBzjw2bzjeQ033142p1zYTjOlKszLMJnM1N/YK7T25N/QSFC
Mf/FmeesekDwpdDo3c+2KedqCvfIai+lLRLRGLHOCP7etb4DvNWY2UU4GT1+iKlXyk2yik7F0zcg
rQifT1WaK7PJQ5WB8UL/Xapipndi4yWIUWjXmZ2CHtgWwoI8jvLLQ9lPOtNjMBPStFl4cvLyB4Dr
ncGkt/GPdJDj+Hvo7Xi4ToPJ+lrK7FhG5Aq5urBprHknDliw8UfKF84uofxvmJck8bZKtkLAGosU
aNCBiS5EgxK+nJQ9ExIZvOtBhvxfhumnJxMBdfeT17NNisbIBvkBQcScIpcU5QQbxNtXWtVVy7xo
irjPHYwoZofyG3Rp0+kTL95yaalWc584uR0erXRBh8/fOpoEt2VwhgHYTd8mduPBo7Jeiv/PEjIJ
GQw8USLJfBJVZCb+3hQZ/u9HZB27dzq4o8+y0/vCtXlGj21U5JW8CguaRctbiKwmQUkoxBn+4SPA
2V6YoakNQBs1DyFMvhbN8l79oOAMka8Ib3Xcz/W7s8nGgzx/+OkgJfKU1OTezSBRRwsc6YaROhHG
xI5J3A0YrZGcTEP2Loa5gqHayh0SdNOSc8veU/1Z9L82RAZIlVRiRUDMADuP1JxB/H5w5vG79wjI
V9hvpn2hx1IyxkEREdH1a0OlN+duLIkbLe9Jrf683YVYXbcxFKKhPlRSf9xTCtxbjsmV9H7Aj3a0
59LZ/SmtGzVKbxnofWq1RZGECFTSXB8CZL58JbjlROgJeMItyC/zVizttqu51Bj4IyZG4a6p9qB+
Ny2Vrd67/LAfuUJrqdOcLorHVTE5gscNmC39pNlBfIyukzbkoUM/1R2tCzLcX6uQNRH0K5PRxkai
NywMc8TxqY8S7ZZFc81guD6uq7mMzf80k09hw30eaQ+Ci/hMz+bbrPNAR23QapepMJQvX4b71Soq
t0afxtS+tO/ck8jn0HZ4H8HgG78MFbv9kSaq/fdpU5AlHFbskPvXjRGmr+Ns31mDXX/P4by2tVBN
Ve+0ioOwRDgOTnts4OJv2MiO4i0QI6oThSbQB0uI1jl3Q+VMDt5KyqdH9bN6mufEmNFnaZvU7p8I
JbEEIIRj9FVoLfInKT6kZVqWBgKg3ij2pFKvMzOLV8SeEZLO9XN7o0O8+r9MWNhv32QnBm8E3x4f
10sJfRjO5JZj/W5JfiNHcw8OvzybNRjBwukBXQ9yC5pUQtJ/RmFBz9NsdJ/iV2qsePAcg7uAg+CN
JYZnTGUjjucjxmOFlOrOQjemVGqQ1/Z/cPbzY+LWUxWbXr78TlkIKwg4ImkP7ywgDbT8NQ5yw6Gj
78eCHffM7v/WzCzM9gQt3UFyouMMroTc6RHpboQwK6szmfCO3RUMyBBUEAUAnsaEN5pW6nooAP1g
OQg0IncTagjK1lZoK/Eaibp6Dd0jTKc1+QhF723pQRj75QkTVOrSMmvO30otLFq2PqV5tZ7PRAxL
oljYT/NjQqaylRkEwtGtzhIG/CkNAFxvd5l4cXFpF/QEVJOUEbLY9rkuy2lscPTVOY7PFBoZy/VT
viaHR+Kji0P1cHW5tsW1iSK0aMrHeDOEw82jh1oorbCs50pGdDoVIUqXrpBmw3SIv6wTfwmheM/5
ySlzwnh67eI4fuL7l4fKmojZJnh2Og+H/uANDwcYWSI7zJ0urFmLZeRSBfcANTDh2co/dC0xAoRU
BzCuBTjYN5Y/7AQjHk3tJCim+O6DRpzYpH9LcvUTFJISgaOIUCyHnxaZ/AxicV3w1gNiUEwv1Pbr
nkULLjwLomj1G7psMs/5Nfjm5G3zGmU8BE9ZxR6WPzHN9z/vZDZJ1rN9IJq7IqwUy4k/HDpV//O9
+814fo3YwGhGHYpkCh3sZmXuT2VWMvIJ1UHQ00uwreblyjibjKZc4uBaKLn0GiOIs1V+MgsUKQ/+
TyA01qwUukYw8MhT5gNaJZXajpkoq3FpaJPQSSN0kOPhot6kYu+jR0d7ekbSee0sgU5jSExMZBUN
A/dOWv1pkUu+508DmZYXrsME0NUePGpvvjc6bQ5CmeMvVmjT3VJkB5yVFizcgXcUiYtxhjlfLefx
QKEV2oNYt4c98JalFqiUd4SIM2IUbA1NZta6TEhbgY7KZ9WN5Ng7L6gjfql76XLUYJWOcz0rqRYF
JodW8s5ILvZC6+ysvK6V/+q9T+3SafSNwF8XgR0ZLlBXjqgnNbOA9uEt/1R7BaTRtPK6x/JHuYsX
RTrEVvKrZvgAeIq9X9fqyLOVmVe9/Mdbu4aGNHVK4LxQiv7Kp21pdbad4qVD28pQvdoCPz1Ezcim
D+/kprkpN6arWXpTbMl01S8kAF0yQ0paNTvWKjBL6yJ53jPhON/N9fqOT6eWsj515m2T9fLSbqPs
iT/vvy7ccwMF6MN/CY0h17M5X2nZP9r7hMZtRdKMDFS4Ss52SFg+RcnejUd+RjNq0XMglzhd3com
VK1bHrQN0Y04aFHPV4uNgMWzFpA3A96SgJXNHOvxydD2lw/jwqt+AyHCNKRHj9Fsba2wvH6jfXHg
OHLhTVPf77EvGOxvY2xjHFho/No8/tJAGEM/uMxzI9Tssy6ubv81zPANnTdcWYnSBWCePcmV8ICA
HUhLN5ygIMZ8ZyS/SQ1fNyYNIyq1Gi3H+rapBis1i23+oy7g8MavkCdCXLAp6YdYix5wHAzBioR+
Gh3V3KFC+XYnZVunYwVX7WxzpsYbQr0FoopXupFUDBYmoYEjAGG79e5mY1HDJyfA2MjduX8Jfx9f
mPnrrPhgvsz1ZnGCOkBN3fXVK2iTzCnR0TEUUYBQijwjqGcAtwToJaHK/VxNF8FsSeATuIk4udAf
nbi6sjE5asaxH5UHSW54yve2l45uq6O1yh8Wao7+hxjdPj4/ZxtP7RhWgXb+kpVUBHwKkV1j0mAd
HYoT70cLS3dAu5P6vfr1eIyWJNGnzh5+WMUxQsVJzY528WXvz/m/e905T3/Fw9thEgs8DCblYRo/
5otwzBSAgJpfsVUBBjUa3QH9F8VQp1C+MCosPZvU8hvzxF6E/vsf+XN3mXu/L02Tz9wdZjAxoWCH
nK57Ow4M1NFGafvy4ygSzRaB77uDkD8x/kBotC5QZeUf+gWh6C0ArMHLRzZUN2RLYY1/Mgs4EIOk
FBKRgeMG4yDMGLblEHLIkRQUIbjJ6GXX1sYzbtFszlpBXSOE31XCFmht9yCTLebk4Ts7DCO+mB8R
9vFkOWaxmjMpIgGet8M6Jhh2mCuYvoFk6lt+ZSZQImsE/j3fURWWPcBYySc5Boud10E6YikfWOU9
8mE1J97B7+MGp745NoqPDLV6dovwoyjKN+sfPcTBUIHJz2xAtLwuXW2YYsoL72qWxuPnxTGaV6pK
HRij7shTQcSX11IE9ndRbG6ed8k7CUDgfIuVlpmvOqQXFTLOYWWYhWh9aXU7svnBBfHNw7enftYj
SUEIYrePgaw6npyDqbbFoJvjnvbnLYf1NnZN9OrUq7Ubux+sco4GX2qXXlFgj4/sp++g10ZA95ng
7LUvTCHcZ65Km3q6BP/5Na71tqMyvm22cFgZKqjR7+Jy7OM3Ai/UBZMVV/qEQe9RMJAxbVYtNXOE
O4XCpVVGEYI8XDAUus4EF90+ulRuil4/g24GDMUi1JNRK5bcOFYDV8wQFAq/7GvEPWZyyxtsUV0g
xS7zgYgzwSQSQwSzkF9GTOBxt5SO0kvJ8ve4mDfQYtoDpAoR/E6RqgHp8itU4RpIVH5sfrlq32Iv
vfApGcNtucOB4b7Y8FFf4qW60rj84r46qsNoCBWfOfH/a8D9z6shbX1vA5SPgDN+RWy+Za8bNNkL
oRuytiLrInfIeqrqDfwvcrjLd3uiITE5LkXmZJYb9dgXZeuA4dBUBaGVCBPytO+zxb1D7iKwvrBi
QjKGafMUqxv1c+46EWD234QICuMwBUTjoesZS4dQ8jxKaVD259dJfxZgso9SV3dy1CvciuOiDdB+
JNqaxbTULLbUpz+2gwVlgnqazLqr4yl2FK+NhAqpsWiDGJFXzV1tY+YdEGif7uQe7k0Ltsg/3fou
bwwaQWWLQw4NRSGPDe4xl6o4gVKVTDfHS63lpqIYgUEXShD+GgG/+n7NuWe5UQfJz0rv5KcqUGs3
ZKNP9fFMGvp4rlVte2ThqHK3uisstjP6n5/qMgzPhDV6Cd7f4wLteWK1Ng7Bmd9CXqiq5dm/l9/I
Y07wYYEnts0yko2Z0X3+YERBcqWnM034YGePN7wa4WM7FjnPSfJ3nUE6n76RHuFmB6wFRaCQDGX/
BBGKXToXsmY3qQOPmhbUuDsdP08hiwQIRPwiq+2lbxaLeCJchlu7tYhbjgxF10R+gJK2Gzoey3yD
gI3hV4PaM9SLhzOdoq/N89DXvNSytx0bV68qpEOf6qSZcYYH4sVmaRydBj2LP8Cuk/7gbWymDCQq
Grq/7mzKB+8XKgiVeJKwzOqHqf5vw5+fdRO++mWVZT9tEunH04hS7bl1BvXRHrsdD1uHYG8Dy45k
oVx5uWhiVtSd43UL73GboaJt2+Jec1BoadIato+aIYblLnIcgEcwUFczoUEXY2H75djvv+WDb/4o
EHKNHUyV57RP8ETQANh+JjmWqZdSlmVCiBWZUN+OpdRCGl4bbi7MMWdzBKXurWjd10nz3PMWyoxk
MMv5utzBDQsESaY1BdCSD54psV7njbB4VetlwkMQVveog+x72N3cJXUNjDB/aW7ffGm+iyCmpVzo
2b9X3SwjhuJA3UYTw+kImDAJynLP0GIjLZYLXJhbZ4yN4bJrfGA/QQuS7Wn6Fx4YTcnUIPCGt5oD
wAMZZNsQa+z1XbsSvk7q3G20zig1z/2hxuCjuO1FDn5ip54Bd3xzZBywL8hlhie8iwOh5vLrQXGj
G5hU+e0xSPlAWD7/g7/DQdnPr3V1zcUY9VbgzQ2nhME95nHEtExDFutSbfzjDTDmL+aYSXWSCL2k
c+vrv8JJFDk900tQuuAQcMaZj7E0OR8iPU7BoWJ0+GpH+WlHCKM59wYpAwVwAK8ifUZus7oVlb83
wAaUrDNF7VkLtH4GFvSaO2VknNtN04LBU8ZyCzytLByHcImdVbx5GrM1tRpZi73JzlKFr54rDEMN
mxCWCb3l56zG70buMsEOIyeWMVf2hICOG+BJ5E3vdu1zhTi5eU+VA+qPBEMlKn+c/MYY9tNHkGLp
KthFZwyVmqWj/k+pU6wDPCJYUaAZCP4eRCmL2wkM/g8w0Sthf6NX4EW1RE2HB2MV0IB4YRklTXqN
EYoQEePQXEreRobM+vwFVEOVZ7Actpn4qTRWgjdaBokO9LcZA9hdxvVnJGv2ifN+VOJ2OqD2fb85
8Av41RAhq3lsg+SxVUGcntWUhVYRlAlJaVRhGdGP5cKFssRCFwkWe/JrkJPHf+sKM0ws0KUUcKYV
WTLYXc+b1LHJpRoBAAUDCrpE1FthyM+/SYrmPH1Q5UJpEHkauuveiljAx7CrKCEyPJTS6zfTH176
vo8JUK7UDFANSeWGg0YBmD2qvzOMJ745fCLOKF2x/fN6HcdcB2UjkYyp8M3lDVs10B6ZaFlXtRg4
ttqrGAw6Nchvb34AugqAciMdeHXGIfgqQmXvHqnIc4jEqWk8gLtYatDInxjES3AAbgOVhcomiITR
X4TqXMYVauqBeIGFsLNeZ5VLVEpzgoFcxXTAL9rnzktGexU2B00jMOEXa+rMactvNkhk26OO7TjL
3bWg/WfKrpeBU0dPBHguyp65u7ynEFnv6OqfoLl9ZdAGR3M9cB3S6+f3gy1TgVrL9oRw30Z4Oimp
/cljumk9PI/V5KHSBsc9CN6S2BXcKCO6VWTS8PN3PkQkWaTmmEF9iDukhmXIPxRw3227vWmwNem3
okEJkvpegBHqeznxph1xG/lbvzHtfAi+dlsjblEXY/O33Rn8vtR3tagcUGbDx6+w641wqTlFfsuj
ixkVt+7mdDrd9dcFZU3ItpqKcfxmMMHywtrBZOwJj5+KRjrDqsdfUu8eatoTtNj6ZkeL99Y9MP5i
BEEckR3WZBSJfNIh7XkkzHS+BZerjaN4lFVsi/z6uXZ+HcgW38VgIjJBHK853l5HqKEFf6TVU4ny
ebrqawF5wruNKoWzxu+Deu4UmvJf1q+fuQbZwLy1JKvz7Muqjues3NSJSltLioFXRUETcuXCjhd9
Pse2mAS8n6dkWe5u/EjAj/0Z7cgj74tKIsh8WylfBe2kF0i8NNVmHDrUICWxVkcZx0hgcLlJoezJ
fRLq0TZsTqyuJavSrgZCTOvgTNMKf1ax+1x+LZhYMfsodC8IiGWcBrRSLuHuskO66wgKlBce0ABt
gk9IBToVU4bSKxnuMXqVXgvybV8KeLIlmEbN90uHTeaw6oYKG0wRbGQigGltzwfDttuVAfV8QNul
faWYWIh+OZxq4kNza18+BpYWMmf2n22ENMo9vzRnl6JHyQUVwnLe98wJj2zVG+IWnjgYB8QhYe44
y9YOGKqQ8vwZcGiwpnYfwmJ5sylQkTm4stYyivBrsHJ9yvckdHKtmRpNyTzeQO0/TSKA+MtqTYuZ
BEhb+sR6GtZfSS4UQJNIG2If52oYW7hyXRIXTnSSqibuXLtDfdpcqvxC/qBy44Id+k3vPN6VYEE5
KkXLizGG9bf/VCgia4EpwnTAU9WlhGHpyzRzg5u2AChaibgfk/HAV/Bba8yaJrUbYA4ZbrDLpo5T
Bnqxi6nzav6ywtkue0OMRZii/n3zBxeHAK8apGIoUyHhfC1IIey2OMRMRLObzWgEDCmGCMeRfc2v
QgNjii03PYyqkTXTt8X9CLFilyXPm64HUUw8CQL4BXjGZtpOBFnN5OcWBT1t+943Yd5ugjCJulaS
IBD0bkap6OWlswRlq4CheAg/GCJNH7rnCvVkommJnNUVtfS9rYsq4GZiAWo0h7NJvmQmWmqsZiTS
miygxoWqti54YZAekYKuz+kuNOtEne3BWdOD7sYy81JnRTzJCIvMBYY1jmHKW/vmAI91zWaq9Vl4
WTPUkopj/GlJwnhXogaHsiTFZ/ZBUE9EnMr2LIYGUaN5adBhixB3mhnxBukDGCNDB/Z/Kvd0//xn
bpP1RSLlGCL8gs2InynnGtBy4uG/DgRXA+lXqcJwJV5g/D9VUDtNJU7cID6k/iUxvXsqRmpyS55L
fshkeQ2/FVrnpSw6ZUn+bkNMs2lpJw++VqTtixneSa4xnq/VumyHLHYcMjeEZlJlgErMSPlaZEXA
gapPrYJaaCB8An33uBHZFHqpndRwS5YpifBiEFUnfehTt+tpcPDoBeQ8qFTNlfxO8BU47v45Ra72
rpLrBGala0yISdaMO5Aq9epq82P4aNbomgwTyT3pXI74XcrswHFu1792N6O3D9NDzLW++Ilk2mlQ
gptdIFGyfzHRv2RJRKpvOMlwUo55Bv0DWT47rV9iaDdrnBdAtNocMBekOGC6KypkLdOxvtaU8QR9
aLdBfJyAuDbFy3UvOvxNm8jeu681BVYL2+TeiWlCfIPXL94pZqnWsTA9DOTenJWEwy3mqscwrzm9
Z9mibxi8tkOl7C3mQZicBjGmyeznysFGbTWK9wIXTGY4EJeoCLKC5sj5o+Yb43G4hNM0mdrXNEO9
BP49VGdg5UahoKOQRR9F/TEijXK1Tyi3uzrc+D7nprGSQ19cHcGtAph/Kffp7yOqCA0/il8y66Ml
VxITjdvruxdJKJagOVR8HHeMIjRwfsZeIDoTU2ebbUWfIXeGoc6hUIo8+sEa/aXd26mqCjcLRElP
0V1vqPupJh3JpidGukxVW7ZwywpF5yVlAe/D7gfXDr7eXMMHQgIg+EixEYXdxfZTnsTVtZjoVs+o
epcLBajvXuLrbqT9wCiju5kpV+w99/y7Z9AlU/v5qMQY3eJ2zuGGW/P8ESfPKlkudISNXy9X2yC6
V+tdb010wkgxNKoHbYYO8a6V/pufLnin21io2BfQNdL9OJHzuZUmbcz7hO5BHIhtldBvcSqkig9Z
/l4O6tr6rWwWDCsANRgK0algLwq6i/Gy+wj+03T87/lVzXKZRS6p36nWywz+xxj58eVfuFHOl0Nz
7T/W42XW6XpHm5NTEjET2qEcMS1/YHnniP/HfOBWynAMPjl7yobmEvdyGXpdRqjE+36QeXAEU2Ml
wkYqWYLwYH9iyAmfAMOb9NziZ0LT7XeOG46kMs36XttOLx4mexC0b5TV/39Z3mtDB35eF7J6KE5d
zpBTL4KfSHSAoDq7Hi+pZu+cVOfRDYF1nLiASXI5JF4wlL7zlPZ0fVuzn0ECqX5BaQ+w8n6OprfA
ftkvCvRxW8h7P0GYhbp4QrLULXFlAuMt86mM0jbyggO0TJb6Mqlijem/fgYChJ0DNwQd1Nr501on
ZbVnC5M3Pb5Grbdr6+to7T/gI3XNzZnzQLgK7Mw+I0L9X2pSQbNJlns5rqcOEn6i0Fyj+Uq6wJ+f
gDZIgKICh1gH8luJhGLPoBtqZbwpPCQJT5w747oXzIo8+iMjLGkK4wL+32VMGMRqbpA1E69FH3Qg
l4N3l5hDBEQfYw1u1bjQVhq+FylVXTtNX9ZcHQpoFpHLYyOiNaUWI3lkqcWu85I5YyC0L/urjpVl
IN4PDc6SI6oV2IUwC14j9BgRtOp2xEzBV3K6KsE2AlmbbFG0B8bT7tnkGbRO0hqwNPK2o+CPcUEL
kpB3XhJ3soCJmUMtVef0uvcVguJIvnY2OfAy8ON+LFZqX3yOa/k1KBZkhSDrzJUVQWaGp8Dg7Djf
LzLZ4287Uo6BuKD+FytyEPLe/855d5J7mC06W1gna3HJJ8cmDOb6tISdHvDTP1uuK3GcMakKX9ye
lFJhqXLK5p6+crw3REdhTSFLlw3bpP+vZd8Qadrz8q+UovQWmf4sqZ85VpPi/5papyG0Nrn/CZ8H
KFMJjzRU/Fxt4Y2S7wYIx6cbFrtY71EIM+THrDFps8HT4eZfUXADv6c6WJGQw3az7Z5UGXnrQo/v
mrnutR6a+xrN96RkGaIy7MsWhS64J5rQG87t8LmtrV75e4fa9ZEdPLugsCflowSXMkxPPuAZj0k6
Qf+U/MUenjLzRIFex2lH64zrtwK2zo/W/ST08n/mwjgDCWQH+aD5tqm7k/VeOKMr003Cfuf5McE/
pW/NtRErpRhhTi8ifj7cPz5KdeYcE7KUEe3Dj0bauLYYQuaEz7m1tqmrgnM7+NdmgKzdCNN+UCG1
YcvD5tyoVVDrGG+ahjfFl0nJyZgIeM37Xu9R1Ata3b5nt3OuRaz9LlA5Ln4gcY+wpi2ABGjEnE2T
+Wkxhxf+rbPJSMIXp8ztmRTHzrph6h5W8HMsKYEEglHDJUML8SBHo2c1Go5TZzgryXqTVu0AdhQX
XYsTc9HFslluLFv4BkC1YoWhCVELBqLQ9qw0lJXAGC2+jvvI2HJeTk6xZmcRXEKoesYrccUoanGQ
o4v6EiJXDZRZX0yewFVSKX1eP+bZqf0tNitGU321sdlBJVQKXqU0138oxWfOFCrtRgyeqdArcNJj
063zpgF1e/MUy5cgjmkZvDlHSw3EU/hCL5oEyGDBCOrOqeSBCtmATEj7pGg8t5UlGaX21DXtGimN
FA4o0o6OgSgOz7x3VANFULmdz1b4+LQLrX9VITeqYK03e7OPQlJb5v8LsI+bHaQ99EwwSmJIW8fa
oVk+F52/6EPavZ5yXdGDTQuOfAKWpUkR3RfMrap/k19yR33kXa8UBYHJV3sHXgP3jAyhmH224+NQ
ZI8OH6eaIbfPBs2ognUO6GO3w3WBwsH1MFFT0VJmd6yZxJuYRK/P2aTA84w+788mfqmZ9pBf4qTW
Q+kxAJ9yfIgXUNTpr9xZxYIhQB80zK0Hjr8RngBoQui7EcMcuG2h+OkOAJcpI+hI9F9KL+kcm0c5
q5XBF5OBLWvK2WSODlw0PAEQhAjIls7oOH0wyB/d3fkJkTubr3BwQC3mGefcJF0g3UOcEWPuh11G
SFYPuNYzxz2EuttnTRkA21pY2nVKc1IJWb4wccJ9gkX4TDx1zLUKEwQe1QDr1oVetTBlFkixSOEB
fpzxP/qU4d379OUs0ffxQFKoaaaXItRpzCdtxusZwq7jMFC291DhHMR8aEj2avIsShnMRGPyU2UC
g2avxt3D7zA9qycXcfN2ltKMSU61GOyP+hD+inY71BEnvm4fS01DG0yJ3Ee8EnxaanTQN0zHZk5S
xxyIzMzbYxDsa6TyqpzJ554FgezzPTO0y0StFrGz8pdYNlL9jfnY62mmgkGtqDGnb5u6iLWRk2Ld
Xc34CNAbsegfMd3U3gMWfEMknjrXctqj0YTYTjFKa1lpgh5XUg1mWnJNNd63BUkpAmVWKScRPpLB
D20CurmPgGotQQNRVtXNOUo1vnBSGozKjZek5pQG4EW+yoWv0xE1VyTyZsetu1iL9mNrB9wnq18R
CisVCLe0Je7HAxJJAm0lUFzXqcJpVrXpURmdvbLu/eBxh25qAFDrcxmPwPWaKm/tosWeIr2he0dO
RacjBoMqB2i816fHpCCm7ld8GPnfYftlLjrm7kQyNaLSQNz7xMp5OV2uUWjB3a5M2MreINvMTXih
JEuYZ1NRbiiCD1VfDjYJ83YjyJb1wrhrKOhzNESWqJBpFNNaKYGKS87SN92QRiaIxZ8+qJ6G6/70
EXUYoPi4f8Yzw2ewlNv8MjFgx4qdRsQdOc+SWn5dHKpYIIh150pCPOvtWYGnL1xhwi/bVA6ENP6S
jl0TfYTS47fjLcdlElBZfsIY6XK2HJRdke9McKaM7XiMbNZp2rf/r7yqDCST467syU4lQ4FGo5D6
cXDRilRpEcllTx8zYTlU83DY9IRH4EcPCtZs629bNwTawnTdqdgk6eRmtTmiz9ZUsmmWV41ajIsy
DpjpVFqEp9nPfUyQJcFvq6aSa7yDK8o8B2ViZhqas9UeN91x2UhbipZY4oUVNiaQEg4Euv6Fp0X1
YaZ/BHRSp2rSjVwAobANGz/lGVkBh5fWMwlAmxXX7fjSksq9uYS5EBifQYfXjENzGnlOmRklPG35
p3cNVHmuvYUkcCRZndhYqE7mrBC0EGgJJlXEAl+kgnGyjQN/x1uzyTdzGrr9YMJTgeApJh/3gIWO
H7qx2BL16ExKo82JLr4za9Ope2ZgAOIRDNAbxd1n2NvfTepZbWCE8WLwyqPSxgSq/qX6DmNroHIm
+taWbgza5o0bY2ROXhi8EomAEJ2RKiqWQL594GeqfDPbAwzC280lwJ4Jk5o/01CmUoutPkyCSNu+
KC6EC2RlQQ7ZdWufrOtgAASYjbGUBViDZdPSL4AJ4jdL6KJLO15HGAzJ6OIPQbfWHGcioAKkg5x+
qcu6tj+z6jG09oQyThlcm0i6Bcfv4n98ZTcYQwusLDEnFyBNa057J+h1VQzonvmF7LP6NTkaHqlg
vJsg4Mcr3sq/fo2jcCDInD8wPAe1v+bT6b6+iOXbebAI1oMWzXg5ebrnuxiIelk/WfsOIiicRXj2
10CAY04bq1au+jGULgQJ7ohrqsZhIS6zEWju3/ryaz+2hBJ9JMq7BxQToPG62ciCS0LLLd8B0Evr
FF/T6awLZRdl3W7Mp2fMXajPNOvdGfROFHNGOK8Bho0q4jzORw+ZhP6XbbElLXXRO5XxgiDJf4Ql
SLbbl09LEZO9REsIes/f0Yhrs+IpQ8Ys9cA/wTajTzz8JdJDtGCtgxJwKXPwO/WsclollZcP1+L9
PNzNFosyyIlC+/YKAo1HDdeEwIps1QSh+1fJBgA6vO+lTK232+7d3Qey8ATDjeDnKIQxBmqjul13
D2l0WdeGyTJPHCGbcic7y1sYyCjSVsh//ORoUKYmWSK/CbL1TX320NMqXNyEbKDyE8lSDutZ5dKt
WKk4WaGVxAmJ4J24jKV7xWdTdqv2NO+AaS3ec3w3yHxYOkTqlQaZ/BQmxzk+aiu90Ymx/OZcuVp3
zzpAy7LayP7gsP5OGuy6cM/YwnJQrHNCcLIXSTd3PqSdcUolHtR0va4dsI9DKypyi6ApXNOkDCE1
8yR/F+uNd55O/yDfbtTTDDNmeK3lOVcjwR5M/M0Z7oxfjE6I/OMnMdcKeAMfTJWUlikQF3HizoEG
/9xZrm7HTjoHwSqnw5jib0QTR4aG9WO6ChyoyemD6rZrnA0I4sq+hvWVD/PDHau44vOXO8/0Dyv/
4nl1a6d+V+Ws8w4Um9SU1ktpHZ7pTYlLi5GCVriCy/E6NzdVIHO8ToBAD5UrpWOhxWp8X1QTFWpR
n1ytbZ/nzKZImPj+Xj13F1Qf7M77gBCQ+aa5jM9ZXUfgVcm1yWZggBBQz6J++79iBzijFqUKw2DH
dXWoEqgdX47Pg9/VzJlGhl2wyvf/Sn8NaPMIQ6J5s6UiAWiafmMDhP2J4EYQ5SL2KRNRxpsw0U3M
a+JgbzC7HFfORyFBfeKs4hCKE1oHvrDmn81fMNX/mt1vx5DnHJOmc0hdL1Paai5v6UFDvW4uklLu
EjUzeMfYk+t8VLkiY9zXHHwOaYfFFKxWeMe4kpF5NIv0i4QPmoRCqRFq1ZE9qvlt567xPvM9tNG6
nn6TB+F9q1cCZmRkER/xmcriYe8/OYwvEHVnJRCQ6QqFgx5aUOtERMs1TBqgLyH2kigXn6lfOoye
FSi+ugpISGwBh+MQUZ1lPv+ZWNrTRK8ygA0VBSW3jAhQYDL/XBMopGXFxMqsnXEcFUMXBzxRj1U3
vVmUm6QBdJZ0wQhXgQl1TZsNhklmdP93Z+4VjIepNtxHYPnPmndp6YdI27yfpSSiLY+BHAxdH9iP
WNrBXCYLXjiQ+qH6ZQyuy1N8wl0QWtuT2e0l/HXFwpG4x2T57cwnLMTNfHjBNkKmY/nDXEs1WkrA
46G1jed4BasikkAyQVeJitbvy2lSwXV4Due0B7PPveUueX1iDtHeIk56GPG0+BYLVuSvlrgY+lum
camkqGcsuDohof96/Oc1AFqfoqElQJGoypFD2RBBlJLaPrv9FDZwzW/ZiLIQN6qBfAqcaUTFWRWm
1btajOoLruC0S2IWyWVZzTZs4eL5YPcM23crLerUJW0l6t+ZToji2RsInSyV+FayGXRUDPRfw1wS
2+JhUa5Q6xpjnhgnQ7hM+InWqzwigIR2DEkdctJ3+c/LZhA2KeNxUQQMITsYz6sRuZq4IPmiapEk
Rd1W2wnRqy7NpaqGgWAQSso9ssX+FpvauvEpeHg476shUvWYzOSfvaYcVVz/VSTcQwLJeVO4MVhp
C+olE1Vj9doukG+UHOApGXoUV/73xVJQcJ4dNOyGprcwX1jCuWc9SPzHdJD2YoIWWCgm9u8i6hXO
brH7W9/wRJPlL0/bcPHW4mh+ckgrdDLHtI01O9uuwG3OnlKV8AO9tidggESwkFW2R0RmyEgDuBBj
zHNWgAfMgvhmnZfd0Ui3QCXqvH2rV1RYSGi4QkSR+Unh3k4mnf5Gefuoi1TfGIrThu+miAXG2oqI
R9NuTLnBk882o3ZUDHf76g5pkNkLZJkhXqNvNQznxCEYrrGVVgN15LuYamrgWe1Gj4pXnnryiYgf
wIbFzgSm9Hvv/NRfn/mtC//Va9Xmu/XFGV3uzT4gofX4ZWJoria4woeM0iiKy9ou2WPwNBUNKNS8
BGKV2cGIigntC1TEYJh7WnVrFNjV4XGJsztyy2VdskeHgG5nN2T4TpR1ESmDSTmPdhoRJYkfAqRb
KnM4Y9tDvcuzrcOQQoi8iUr4vJfrhRaX3/B6nWmbNOFQi7IEBss6nRkJfF6EtIG+j9JfSJmCO/Td
vOS6v4+PQzp7vLH3PUln59b/8lB7ccoxBz54uTS0Fkfa/fkmzWGSJaX8y4keGh+4XMnnkGrLn++M
T5srxRwQMeg/6+BVfmn4F25kRzsJWqQud2/9Z/kFeFLVxNa4q1cLPERD6l0G/lDyGVdkTUdQr8be
lPq1/TDw9h4WgHHXgQUG+ENfLdh9Ic9bxGlnkOjWFBjXKwhfoP9gQ64e9QWs+ft0AzSuNAg+AL3X
eHwSqvjSfZXXA/uHdTzzXylvpr+Ot7mVwZBorSrl3/7vF5mhYaccA9+LstolvUeSIUMF7wO6WVbs
tiZOLvIH/5LJaa+Sl8XXbuEdIRLX7co9lXLSWLXpUAUVFZwnXVlG+oM0H1Kk/xglaQvZnVxNgflu
+YCSnnPY5MH/nBzgZcouAFNh1ras3Ci094wwotxwRzMs3XbxiS+dMrbhJ+ssZV/9GTbWZzL5LliO
7k+6oaa6UHeW0IssVKIT3sB6dOQNP5kycIdrRcxl3hSV5gd5wqh3Bt8PXMnM65HmSSxYBWwZ/VV7
oovotllVmcPAahPazd1vrqnJZfjtbn+ualUHwLMI3p/GiDgt3tSqs8YXv6UB/SIPQ0+bJAiuViPR
rbKHM+sqMCi54vJxJUJgQBW2UrNuFu53Z6+fuajjfDxDtUzMkY1HMlafThP+ikR2dvE5m+ypA7zP
c0mTmQR4wPqA9crPxj4uHZe8ilnGefMURQSyV3ZTwrk8xSvVdnD+/n6sS0h+703+6hqJf2C2hobj
cgkoOg9R2jCeE3gGvum6CmHC0Ro1j6OEqXxS5KuXN2Q6Ts9BaQ67yx1RsP3XQmborVGpAvwW3ed8
Ha0GdQfMbS/9byYbW2zJdCnIGj0vBiXN7WKPDi3NtGBabAuL4Ri0YkNp9ouJPwkfdBpI3RuM8RUD
msYbSfunnkxAHOVB82tEFQUyNQhOQ90ezYJVKDvUKBZqV30ORNmFhL+2m6khRyHXpgdTFg0CjUm7
A06rU9eHQZIKANR9REO1xk4Fq41Q5gmWBZUyNB7qUek4A/OWZsno1Ba9l5Mj0zJ1LV+6MtLaXlDH
r98FcFxF/Ev9m6upC4DDrnAv8GYDT1VQnHGUBlIpWoRkGdBwiv0ujDxttY+VWxTYhVRfWPzfCGhU
HQJI2tWmGcQs7ioFPbjL3201bIa/nILcvkyC1EQ41BpZYg+TkZue5ohB5Rvtw3LoWucO6SbtXyO6
xM8rYxA/kaObmJqWnPaMDGzWaJ7Vu3JH5l73pJMgt14vjeIYpsAHl8vTF7zpXELjKWMHTlop6JWX
/6Xj+D8AgIfG8RKRkNz50FCo9yP63EkqLqv3DPRN1MWUyp1VjzcRJ9rPAMNb3Hr1yvtZUUKSkKOD
UGNNjuRq27nA0kktliNm3EpBnftoUeZ2BeNfn8wJ1rhwcfgzoLkkZwJwhkJdOkygbBbRj1cOGyjR
eYeW5HbLoat5gN1TlShYcVaKsorAy6poxijbnIaGwYD1tc9HallNAkJHwNTFElk1QsC/+u6E+5tE
TQuLpx0CX9+vfiRLIBrMETy29wTC1FMTpbFQMPVvcRN7SnX4eoIIoCJ7E5TpP27Trc/YlqrZpAlM
i0dyTC5ahuFQGiLyaF4pCmRLA40HXAvFWdvTTSDGK+Rrg5hKJFjD30yL4W939W8KT3URtoQqB9vd
vjbFxEHU6JQfUGNtb4LdV3lyTu16+5aqieHs1ttXxRJvwcQQ91pJkAhb3ZgtEm9COQ5v1WigjwXF
VkIiCygQUV8EgTped/kP6bqeUXAaLfoENb6HfP0CikLn7eIwVVJ6qNVyucI+HJK5T+Qs8TASzAo/
lwidfuRekTj7FpRGFPZMkFPxg0dN/waglSY+iiUEZzpOuJOfcrLWE7rT3K1anHacoBwpq1Sh7BCk
CcH9rzMoifVYG2zocdO8839ncMlWyPnYB2CL13XrynJIHe7rCeOPMJxp7fPT7wr8DjPkfvFFC4zY
mZ8WQflwtuV+qXQ78mpR+souZimomcCXNbXiPZeilaofotrTnFDys7mA/DpjoMwnjhJ6LW47rOC/
wavs6ei4p7zLRf8+46FRXhp4SI4QBdZcESrEfztXbdhqwBmbHiEA5WKifMzTqaxQ6U6E8CDED7bW
UIkXRQhjgnkqdXthTVaq0mafLeEgi2NKLbkQYu5NUntI7B/pKJnRWRljhQvEopz+6l2JGp2qBfnQ
SvhhZNKKlAsqx1+P9xRstV5yE0SwORCvbyLRbymloa9TeDi3mMwiwrJYK3J8eWv7rT4NVoOZjk+n
XpXOrq7+23sAyr14g6dsRAmBFBhlUr1GIiGvfvc5OEx110EqjWRGhzpOD3lQVHgEmThK1mWbBuo2
X9tfa2qKOPjo/L1sJNmkwRBksAAqXLNImoawbH2KescXyXK82VP8njVTbTxzPE9siRAS3gU0pJaW
n53rV6NNq9zBb3E/tCUvruZMvoOMvZ3wJ8Old5gO59X6L2+qYGDcd9geGKsdcYylZI+6/CdScQ1x
h+9iRZBgCLzv2+XTHFEs85E1RGZDoJ9QYaCKh5IIBY8z39q/srGO7FVo9XJqTudDoPtbGPpkGwx7
5uDp0WfqmQbRJDfkPA5PyBSFN3b5i55wBriCY5bMsmqTByvunnDdlKdPyuwsdwgUh1waDX3WKFdW
RxHhWDIzSXZO4I3lSURwTwFbx6c6pX4t2Tz7+8rZbtbRlS1vlYiVF41UHbnj7z35ih9G6jvWaZTL
X77Jrk5pRAPrcz8D3Xw0HNSuqGD3KwDp3HQ/urF6J8UQvLsgdw/+fnGrH1EI/y4kzI71N3BNnpoG
Y/zyss9yjdBjRZfBw2Oqwsz+41BKzh3tBuMKIbJofr2dr7cunnNHHUhcaOWianJ/L3Y4pMRhoFQR
UQrvwPw73bBmGtCy+2kEnwnvlwQVRk0InhWHOgdoPv7gqiM06iuuE+LbwiZvWHh3Tt6RgyVNKIBq
72KOveRk7UxPDBpvmaI3N5Pw05P5pjyYLvuWPdfMVtfJE8HBi833LuoNdwT46NG9PhLpD1yLlg0j
qktUUG9rTHEzEMvzKbNvXJ7zXQWqSObQlhUt+dTybhDK/847cLYwwqZ9Jkn2flVGdwjom/7w6tuV
UNLUbGbh9LRmDWiTQiH1CDj7DPjIwr53e/EGXpT6YPV8KTScJUZRNYvqAhgQC4ssXKD2TnhUENUy
WbEJWvO6jDnHP0lfKGJR5cqwnIikQ7KAsEC9v4XmMTx8VGj0kk7Z4p/98ktCKXl3VzQOmyCR2qfK
krMCbD7edyQM54/6Ua/+fOcXCuLSPeD4ascCi3LKCCHZTg/7wIl+Nv/z4F2qzmmdTu3Wf4+hCBp3
rud+ECvnY1WQDfxyQ/OUXY3YHTX5IdU8Z75fpi79624bwbYBoaBCwQMIUDeyM5v/wiSQ2L9Tnr0V
PSIsMuP8r/hLUVp4sqXoWhll7fJhXC7FRvkkt1fhX+jjHybYjQ9uDlcrAdWIRxlG2/BdAx0pdyNB
4toBDXH/Wh7VloU/CqE780MpZi25kzsxVzO4/SJnyPqjaNbI4fUxfnBS6jY8LFBFQkiea8PAYdfL
WjDVBEJWiIOPqnACKEWqydBfTEBFBBCdjutPmpSxMeagSTgE7fNfKaH/VduHbzaljLLiNNuty0Qq
YqVUyAjT7bwcoCxFQdyYEo6SSkWm1W3gKCdeFyQyLdK7cjWFpYK6vDx/qu9eamenTQTi98FTRYG4
GqVWuhSPBL5kijt8i/aZRojcRapc+hmJgGMqCrhgbCxHf9HnqWsA8Prtd/VGnWBCBF4HOm55n0iP
txwSH2A10lnGFmmj2WgUTbt6wg3OdNW18U+EmejvfnQZUqcqMH++om57/vH5DlGazd+EXO/u1bMH
t7Usuc3DrN+mM2I94joi3YGCtmE6DLvzdMDDBxLZhqEDlNDr+EbKJp2dMJK88hhVvPfFZCvDU7l8
y55fs+IDswP7y/Xjt8+qXF3T/cApGVwooYuRON41Gs+urQm55ufmjNTGVaROdy+w/MlgaaFmkp3u
yPQB6XaAHGJzOfVisQkKolNi+g1vonteczo9rpTkgOvoNxzTMZyMxQKQ1O3XZ7V6sr0P0Z3RDW3j
/JDdmvpQpc4MF6cSQFtZVlb1SohxH1COoaRWtfI8ApeubfpxJ+SAn2gmqdAnLFgSKVBTwL/WR3WF
mTRAc/y4o9wTs618PQS9+cPVkKCoaq+EzkNdr56rkoC4F2MnBrvnhjSZPuYDQP2o7WzaiXh7QTtT
nI5CUUeV/ahvIhx00bGuohJZJQwLlNnMp08GZ/ePq8rxYSQE0mPzeASY7xUwT2Vy+g48SDJMpiWu
PWor6kF/J1LY5yJSXp0usWUlSAOwyzlBmUWeke/AdTuStr28EMNxv8zkoaSuranqE1N4ux8r1ytY
xqvshee+9JAcgU3tJfukL7inYkXHYxRhOECHrWPD+VQ8+8dkTxIiw2LVzH4r0mqwqo5axJ42E0Nb
2fTpK70fYUpH8q45dyNhcSanLZVTxsiQI4SqEClRlLJ1eGyZLe6WBveMKEtaV96WyL3ktJRB8E0O
zIKvFb40ncZaB5zlo4FFNeUUdGKyJtJ0B3NOwGkGDuznPEP1Rgld0gd0vYQIIMmcz2eLNVpHf3CR
Zp4bigVdvrJS4YLLedQk99p8jtcgbLtv13olziXC/1Ewk0f84KXhVAilA7UWDPadvTF8+hoNFkO8
hu0LUjKKm/R0g1VZhWIRmSvrUXN4jhli6Js0UvMx0uQs+Z+m0XG+Np4UnmfdDzyeIlBHlwCTKhjM
dCbW03Ao23eU3b71KmxxooRmiYrOFaVlXVGtq7G63clW0vB5l3xol5N9MqQ2HrcwUuFFVvDPUM/U
NK3Z5KPvRBDaK+WEtm5Xw4WsUF/L4eArkJVOEa1tnE4rmywhSH7UMfc0R+oJY0AHAKN9NFI/mUry
eNWWNGzR3XseuKT0b7TkHzKKq/vOaqfaQqlTF/X1SMC1n17tdYU7J8X7Iu27u8mmvl4EizMfUNfz
T4BNbt6osOk+JN3RFItUASxPjOAAwzFlsnW8HGiwmaHqv/AWUr9yAr7fYyKbS87+kpt0r8kTXZcJ
6OY7s7P0/VRKwC7zZYzOuThJNosv5VRFmZ5lqMVSnyt55qk5BrzQi0pH14591efoSTenEZHPDCUW
PNH/JDgQb0J+tTSRN8FPxzjun4Fw9xvhwqpbkn6xqQjgyTAtwy4UU8dRseh26QbzkcJQAg49Fl0m
Xx8JUOXi766hACEMmr/volM2zTY/6pf/dToShwpUUHAH2tE3JXY8eX1UmsMKAFDJiCx2CEqi47Ov
JEj0Fmu6HeOMq2sZpemIvM9ymAJnsiXchGfeDzPMXcYyiAzeLMTB7HlcbLwH+Fb//w+1d/Hha9HR
PbFHqAy2g2PzqRqOUz8fjz8I5bsF9wONBxuZyvVNT9+HdI5kmR1PA2UZ+Vfc/9YPUtVZdM+5sATy
FeVu3C2FPhJoBxL2csShyA4ayLFKPufRIS5FzTZEFGW+x5JvmER82jMHCKOi0xev470NvRfXkUcP
OP+6k5Jetck0b5t6/1LNufUsSbaXH859MXNb1UvJmGD1vdLv6/b8BkQlmvVkqbQ0+iEC43reePqL
sfX4+DGH4pm5dYNdKHARqTJnH//vXlOIEVVWolS5uhH/VKQlf35vrnZrZDAbV9Zi2GlMKW9/dtYE
RUgn5v7aT0/4/djtLENRcZCyz0za/vIvXdOEjBNpEq12fRBIPwGeyhO+jKBeUdJKswuzGYeQf1zZ
DgcBJVTcAEGhOLPetd+HlOY5eYdyKMvRxshQ4XGcblGctd4F5FJZLqgLR4fd1cAK+lYKz8BIkOba
9Iasb84sEtIG5E/Klo/P8Bgzo8ePegHhKKmJP+xwflOxCb0oXYlronwz23kUbUM+yY7prIxpALeW
+MQesBgMndrdJW7XuRIDEvGFTAw5TxcUb26e41pwELSn+DujlnRl1IKB2uBJjx5dm8uPmZiZm6hg
GosbpZElVQEMbMjSY2ZywyGIcDS5HnQyPipQjGF8cU2zuuK3hIeCZo7Gm1lLrV2bY69/iFG7qcc4
+aGKlOkybYq/6+ZIVqzMDfY2guYDNFUz7OZQie5apfDQ7IQXFMYb91zaifhG10uNku8SDOoYmFgV
qbZka7kvlg/0KVoIgUf0lUd9ymBNOWnD7XRUI1IdaaOREeFlcad0AHAyce1hB2iV7qKIasji8ySc
BlOUQeuOJ64whwmD3xP+h2RtXvXDi/7psCj3cajs+3CfmFKRyJHvhz4jVme/gefs2NHmbdr05YRm
UbOtbzsyp4QTA68GPcfg5H9SsqNHEZDYpEMQy0U+Nx8muonXiI0YUNmdUmXCMfu5AlUJkn0NxW75
ctMA729uxPwf/VB3FtsZE1wmRr9B5V2tFpQPo5wZMiWVedXB3C77nmZjSb2FlDqf459HDhJEYOm6
+9akD+OaUAtiDsGaHmvxTXxrLvLdohrjqs/Mc36AQV4nRqJ9UxP9gx7z/GYPPu1CUOiJIuNm3prx
7NfS7Uc2q7zcHm/jVvxT1D+TLbu7UqVI2lG7FgYuIwHL0nJO+XfOJ65LjVPZBOj86X1GO/uQKqq9
QjscpCO5DOdarnayFTRfWraNz3S52lrsxGDrzK/O2G2JpVr+DLC+Sl9qSHgr21u0PygDGZtovPGP
EzDLsY/MJCe5rQPKSUewJvvV6bTkiL33If79fOPzduvpWMxLN+Afo+h7f2MQKCMyhjbAppnSJ5Nz
fvNfwdiMzYJgp0HYh+NQw8k0cI+zaj5dxINkn+vFRzIor730oEUEYYsN4OJiS/DrKWCqWCCzC5Hv
VFTpHJdMlTqtA/iCwKKjBJpxMUoabrkQqP856bDGeNEMFVqHfPcx2Mzr/TZxSwK0geIqxRrLAa09
BOfCj6FkjMbTg5I3UZS1NgQ+f0dJo7aT47DkoylHYXp0bIttaqcCsIMaD8x/Fp5OT+vvDga+xCqJ
0seHu+eJSlVztUEJSFu+8LLIQq7Y85D6DdWUlYXgWzrbYW8w9b7xc8UkBY5e9NVsu1i0+z5vc1dT
R5xipqYxhzz6OCcbAn/F9BSW1W8Qd57jLJn8f9Pg34g1rnSIEni71RevAHpVLFTEC6PzcGcyTeSK
s1muUJ0+lp+f+K0je8bQ2FJWydFs0mXZvffelJdPeXjdlmpAu+lK7RWaQyy7blXZFOAJVOwklrow
G0xL938rXQBVQWTcmRoW+xYKvxfuNAM9dE0JkHKNVA4Wm6DgfwN3VUzmQD2I8ZYgUtdcZnc7l+ul
Agw5xb7O+OnN+JA22jd94FEMoBweey4ZhWh6q3+2f3d+hQOBzxMz9ddv7GXrmDy83Pc8UjlB8dh2
CGRz9BuCTq0nFmxThlxcJIGC/XVT5XsRvHX1GXjDiAXl+kXVXFjSPaPqsMND/9w4NqV6BSzCHRGS
rt7uoajDdzTydnLowWkNVNOb8xpp17FoSWacSozOLyMs7izcgzJWX4o30/g/kCXeGrtQpaTE+XV3
FBQgfGIMBm4tk8X6owCCpbvBFkOBYI+Icn+gf+cN6ayyTF5uJAt+nI1I/itGl0qC28gkTqSI49IH
qmRKVTXj/XGYaDh6Dqi48wLDTX+qrqXkviaSDUbHlOSop65VdYWr5rhgTF5GqvmkGBkdD7HvW/N7
XxwxIh97gjj3WK62DDy5AExdFCz4uevXhHByGKGULQNEKqNgzMWqelt+/FDSgyIHyGoWnCy9Sd4j
+6eqM+Du0ZPNCvQK3DrXt6N3DIaVaE/09eXo3ug75lS2W5bH7oCUH5PQX+zU9gctNdLAht7YLFi4
iJIOFF/fuiJ+PMfYGacpBqncbcxfEGZIlIRIc6y5ZIvnx8XgUMm9kxFUP+LnFl/iliPrZ/iR47d2
H6n6JZRrAIev83M8KTWvhzjzQKaXOm3w/NwAl6qaLpL7JoKu1ml8S8giJv8ONWXufZKG2hcZvEVA
II8Zvun/CFunLrh67DN0ZNauT8iXhJfjNSix0UizZLqQlhZO6LsH/8IdSfDp+6D2/lcsD1muf3Qk
deHlrEnOttoYgSpoSl3C7wlICOBa2y3Ygd7CgZhxCcYsqjOqFsQnvgGntTSEdBnIPZ4xP53aD6zp
MnJSII0h2uNcqVnIQW8Yx9P4kDq334mQTsel1w5DG9cr/xqGq92+niGpSV0BIrDCBGTzQDfTWrLa
1Ih+CT+4wMSG8vm7Xqv1E56pdEcF4oVimENAM97+2hF5VQtVpSD+FBWsebSxxijfduA/Egu6e894
lsnUMAHwAmyAmIsvhkqiBoVoISEejOQ8ik2KBExPHx77nm7F0nbqpepXTjAWfUy6fv6BPxp1vB3s
lrxFe2LlK9433iqxcd/W0a2LIghrqPkL1ksNSSCa97TFFLDA7VdeLzhJPPrAJiUwHjHfx9D8F4yS
taS0WWTW7I5rqFf3HeK5viWNuF3Akt5irCvlyCq7AAfDzq/SQ/SEG3OgzcWQEfAIMuFY1dsvSWIv
aoXpC+2FKCQDqLSv81uY9uKhsv7rFOquCbFQz3WTyGnrBicvZVSfLTVTxmB1gFcVfV5loAPmNg4X
dVq73YAI2QI81A1+4uN9FGN8fj6SwhuUYA+ZNyfntO2+n8JPdgPSlRKZpyiXcbnc+aEs7/612Qac
ovIItUkMAUH3pTcM79ZrxFSgedpsTVOyRHgAXMLJlAG7iH5OipPongChK9+s/+eJNRakiF4v235s
bo+d48b2ftM1LBOMm1rLQN3sNqXWnLAt82Ig+g8OQEeSQypneZXOvDtCzeIUl58Y7VSeshwl95eY
EDgj+dpovlyB/98Dw9SCXkmgu8vmNDroS+srPRHRJAHxKdQYtWnLcM556aCQDCnoiifc1h457EHr
XVv6WMqCDg8bpkJzFwXB2dwPhQ2A+Z+MFmPOEXBo598xu6M4oh0ww1UVpGuKGLtriFnzAf7StICv
l0pKjh630H3pAfJjDK+tTVqplGdadWwU+Lntmlcn1FkXwLT0gkSedxsJxKZqDTMJLBM3VTfrmgtc
2Dir3/UObaG8Iy7f/+Ofz9LOWfEdFXK6GVydCn6fP0C95Xm2irdTzu2AHZ509MXnhipS6w39wFFb
fHmZU/yj8yCrvhmW4Y/+7gsXvJbYFqxw75YFTJwzg4eI6vnckbezoPo2y6Kg7uE6j3MslsGknnF4
6oKgQP5iL3OKQFV+tmfBu7c1keT/bXltlhCP0XCsKl6e3H13BTLicfMxJ+oQo44bdqa9Y+ElRrk4
VxIn1SlxP8JaIOZc/x14Y4z4bAzWR1DZv8/4hUEBp064z9QLBiiycOx5538x1JOecYARP2R+gWqu
NUvCCOvL88v6vdfdnVJRy+wQPUUrSw3c/drmmZUm/CPvjoeU+GNUj4g6sHzlxaUKPrFiUMkc5IFN
D/oaLJGon+uvxaFJfd4cdpiAk3PJ7pFr2KtmQ5foEjtPMLj3Jrf8shCnmjeS5qo0PePICnHbnchO
4WIxQ+piGGU0hYiqlvPn37DXi8lUauIqo4Jk2eFhrbyKZ/VMzAlBitUvkjucuGt4UiHzcO6crL48
DOwu5KpV7nKxOHxw5z8L2ypwklj057+wWNn1+UDqXMbkqWqYwlIkIOSpbBqx1mPzcJG+Lucvzldp
mjv6aWkDTZKKrl8Fnvr6UUeYhB+IOZiFk+BIRUdeNt6Sd1yc8Z5pWfKTVWDorTWzjc6S5QjN3KTW
q2qB6jJp8xpMlvlVus5GpgDAYhHEU09VBorEHz/pk2Of343Bq7roQIXjSKNlNsSa1pNJnnDlf+Qt
I6s1qI6UEboqGY8qprU85qmLBN99xhfSs3j3P0FgDKs9VAhPV2X1Eayv1xHyxirsZqXdrytghrKS
lhKRqpubyZasN9iiJzY70dFF6D2XIpwhoZDt7V6prTd5s4LD2xiAiMyLZwH/EGHif7DfUGjZ8yEl
BG0voPReNyRy/AjZLkhbpafO6nRKTR8XubSEpv9conuP+6d3uADWbxVXumDkLZP9UE05NjpEexdf
ixR0Cmgb2iAePWXnHCJWb11d5L8NiEGTTxjik4Pfm/91RfMZtJZKGtotVPIZTixT0kouGdrJT2C3
PoEMzq9ycKCeKk+ukRnkaEqMuCV3IudpbdzBuDmxG/y6OofpaQ27+8jPgjTtEx13kPzZhdCFmsm2
Nb5QvnAfwtcdZFSmGI9Vf2GepOn6rAJ/rkbAXIfOvMVINuwQSl38tSucfBhXkC/btvwSG4i82xFm
hD00SgAsQV4IQlOT+TwdvDX0/+oibqfwSwSSwyRNIc4Mfsy6v+7XQPyLDfj77ODRF1n+fvLBFtsl
w/4oXdkT4TZl+kTvDotiQntR4QaNNCre4usG9+AkSkprEQTYJOuJPBqTBXL0RnMT/E7fewVA6N4b
6oF1C374YfbzfWpgD2SQv8txDTnTHKhKAsTL4ELNgAPMd40KganbBee2ETbt55vFpAafmgaw6GCd
DAHMCj53lefZmhtNsB2tpiIhMVLDwXOwjxnoEe1MIoyMgcK6OzA2UzjhHt9EyIRbmk/ZALczAwQz
ZmdIX24S/x0qrGYD/nk2UhMwwo1VIoSeapBIsTZ0iEwkx/9ELFMyjrMUbRAC03xuCzL7mjOI005x
ygNdLnaw6OQsZGw8dRLDFkJJHOyWpykhQePfQOeVEnztSjIJtiteR6MfKDq8wOJkeK2vHBkTk+3G
RjkQ6eSIJwm6SFVcL0JUPPQIFFoDcbq6fBJc5FnZ5TgPZfUBNEg+xVugj5XTIqLyEWtKGb5DurLL
zTTh2r3pXXgrwTP6CjNhMUDS+gl9QbR0rd3ixDQ+NO0SyZa4nRNouOMbNk5sZ+l6pOGP4lriQ4Df
BKZuBkZQuyS91VvbgAylkHAKJ724C3BoRtB5Cmod0f4fv1sfZ2aH4izjyivoFaapfEz3rSHV9G2c
Q5JYkjYagmLQzEkFX4uU7CnSqrLIeVnl+IPbf9w8phktFQH5jpbEGQa9Uc0rpB7+VgGoAtR9zQKU
rGEH/S2dhf2HSrTa+urGjOdbHpd709aZbB+4jJ1nwgAV7Kuc3clzlT/36jmFPv246eLPY2llESh8
spRfeuSQ71PfMhHe00ztqq7ceu1Yg4Bwy/yBAitqMuhUElE6+2BoK8N3pWmuS9fvYb6BetZAi3DC
tPbkuI0xvo/DzVwTLrbOfFZT9ffkTPISd81gQeNQLJwysXXTHruZ8EgQNnEm/2XCCOwN903Ctw/Z
B+aBUf9tIT7jw+sXxfBZ+ed6pyPTM72rWtFz2zxjfEqLS8E9JR37m1GBLxWHGXCrBAKRz91YVNRl
BvPC8r6t/b7RSe+dkIdJa8IoUukWmi9tx8Hmt+7Mni7/jGCRDhNZ+QpOgjnXF0cq7XETheDJNQU6
ui2E/2l528K5fxWWCRtkN9XQDjSYlICU1SIXVuqSgye4xyGx3l5SxhUrb3GAen8MG5s8VfeKVUL1
uw/i0wMmDF7vaLajkUQrYmufppZisL3/Z6jIXCtx376PpJ9F5HZnhhUSLfLLGwzXgnSNQRmTu9TB
o2ut2QMxKEv5Z4PDvkT+RqNoumnZFS04HmsYt4LuaPSsJfxjI+wHyZcju4APHOVa4EFJ2v4i9wij
EIQE3iXG/N0em9Kf/ux8FyYz2Zna2kwSF1/fBGAsCItSwmYwTZmJmG9TZZD68FLtkUFV618K2rK8
lyw5j9+TAV0qq7Jf8Rtt6p5XBhASrolBvCDhkQBZWXmTkaTbBZHdtyt00fCukgcy020QwVF6hP5Q
kSzDQPX6XFaTfG5c9V+NST7uhNI/MMtN77NHXZUDlqUdbwjzzQzj3Fb/kmA/xIQ0jcRypLTxvg/4
UZG9Q8kV7dLkpkZBPHt/TxsWYAO68FBuCKFwIYRTDe3Bd6xRt5K+q0rAfz4/TBN1fXOUC736ApSU
qQNugytrYms5vNuKGE4cCJDSdPkOH08du7HCZ5cqBBv/yIyLZG0z3xFhskRniQuZtwVthjdEUnC7
Cvz4mGXacrXCl+WFRKCrK7Ng5dKPaSltSAmFtAMpA9WYDvK58tQYltmBoLYsyuEpijsWU2e13L2e
T1dkQOZwNxcsqJ5WBlfR4tFdPm6LZrcpigGIM0xVD4ZrVEmwm9KyIixayQMwjMerOLus29EWbxuI
5KFIkweCwj1riHbohnSegDabU2A3DXNWoyc39IaWTcuUSRncwe8Ct/XRVJJ4z6B4BgFdd0Uw7ZUY
silV7nc9ZEEsxrf3fdT50+fLcadULAj8lSUwLKytCl7J9WI2DGG+Ap/2gd96Gu4k4McjWS6+DMJ4
TDQum/z88sTB+LYTATh5t+QoU0FqKCB7iHvOtniWSwxdiuNFBYvcpgtNK0OC4F5lLFAaoToVzTDC
4VSrSmIIInp/AaTwen7a4DIUx/A+HHixXFVUkyqzcXAG7FKs4IygYm8/24FvNdG51KXHOy+kwBQI
IinU78l8yTAv0XQypATgD5oJRpbSYYvE6XrWrx9ojp5CRlc3eQ171USSeYAH44UvAdoaoOD+sEbF
geSX0rwhVhXVcJ/EtV/xqENKxemUQ9t1dX/yzAXEIfFPK7oxjV7qNg8mphEgkO8pYM1++IXh2zy/
xTDlBBLO7BgMUllP/CQVGMug0nZZArZnpb3NhFSPonJ8OqbWpMJc/Pm0rMddZIvVni6n2DZ7K8/B
waANRnY1xs8Gncf/MQ9ffQt78/tROtBo09uWooRD6j0pQvE2YOoSIU6xUea4R32Y0ef60UOgsNhB
G9TfGCpZyszogg4w00HjZzEa+7Lf6WekUmMnO5XEkbZH8alixv/APbMC/HjdihHxXfrbGpB6WZI8
RiDM5J2sP8x22KafxovQqmguk6m+ZW81dpg4WkTOP7f9/J3zt398ohKSPe0q8jYZ39aXY0wZvYCp
5BFYNq6e9JA5S4iCnpt/deGboH6h4Kov3enPFBUbj16TgFycuznx6CfoXnV78co/A6zk2J9OcfV5
8QvEISL6Arz/dmqGxy71xCBik4Lp0Z6AwPvIiVQ1qYKhqscnYoThCqWx4CWngNUWuvf8oHBOIadV
LjxqccfnKJAahOlCoUdPV4xtGferTciO2OrkHeW/8+LgBV4Bvyy1f82EypsfiZ53vh0/hxYV7TcQ
wc/ZynpoTRR9S1d4/FQ/WGMByoEQA5J4iYSLKv4OifiY7poGAWFy2SVqgkXQKSi/iix51rpIycJb
9qhE6M+0rNjn5fKi58LqP4Jsfm+dAQSCUqvUix4Rot7OIyY6vy+FkcDGC4S5Dx2ru1goQ5fM5yqk
zC/wxXpZHQPNVearspyCA/68KRPVEx8cpA1QykgN1qj1oKyPkQT248fqrZE74Womw9xtGTkRzVNi
+0+cv9vJEZnIFqM9W++MUCOms+mzsTBEd7jAwcq3ssGE+oBtiBdgfs8GcqwluSusuSTYtBtB3GKU
pmZx8Bg6bqoew70aIIGRuFTW4hBjsMZlZcdC1x30PbNlqvuHecmxGb2LjUXNOdDUJU3QaOkvZGug
rRidkrRRGGoOJxcqeTqAosxgwSD0VtVWc8zMCd3DWgwD6+cmVo6NgaT59Vfte4hJVf+860cFygLd
GYm9RD27DMJLCdBojG5IvM/zHKwlh4N2da9IKwfamsto04wEx6i0Br0hE9y4SN/1oSNGF+PqhSug
F5vKozAylY2Src0dcrvZUdGgqNggJQghILkygHmCQk3wxxBkVeQL5WRGEHOwlLEElf7ZmymIBX9/
sC7ClRtmBx2QZJrWWzdykg1INuMMDemCM9glagDvBbtUiIFhhnvj0Fn6yiXNWnJCDvrn9mUbXRdQ
P3wnHtN57WLoOY+1FJw3kbhIFUr2NQ3gLWQNoB9xNufD54FahR9b+glm6Yw3ntV9TFgGqrCoaz40
4vm8yo3DfbRpS1WWDNvbgkvlavbVN3fDVlIY1Ba1yVkUAxLNK82Zb9AcVPN+Su5I3nEL5eMljIJo
eeXuYrQi8rtTezbPPd+3uoUywgpu3/6fY786AKHURhc64E9KBWsBVZrIym4ZqQqgSw+1h9csGhh3
JvRkvfBe7NyQBQ8LfWXEPzqCOSazHO05RyfzIa2yiK/ovGLtqeuJquBae2WKVesabTqcqGsyIzHB
MgbUYWvzThYqXxIGOM0GPlILvN9YZqE0EI0u0h2vXCXGyMWtpJD/1dEWlXjtZ4ztzjwzkU3wqf7w
/xh6tNIcNGUOvkkvQGE9Igul6LhMY51HfSGDAs7iSPCcRMWhOo5FH3SSP9cdrLBQk3Bxy2TNUluj
mXT/NfxBTeMx6lUNdL+Z/gMYi5qnMFOuDeQd2MjmNoH+z+LxWpK2lpdVSLIfoUZ4IVxOU6fCjETp
G7pfuqhzq5I1kqrNMSRbGj4WIE9GJcAhjLGRh0y5QmWSNksiSVz5Nx/TlLWekrzS6TrZZN0HF+gU
mclbYlcXmLQ+6e2+csSGblwzK4OiOy7pTWIZa1IV9HP+sZ3H78eWOwFgVXTQ9snL/n6O8PK4QM5C
RAudPLS8BoJl4UcJMT9T+xf4aBUW6J6kugMWrAl2e2ACqL3aRqxj3mkWHIM8dp8pCQltJEwnpw6g
9MZRRewWcThsAYjnhdqk/Ay8FcXlR9pig969TH5z9v+I3NwW4LzDnGeYHA3cj1s2li/GW+3tiFLO
GjPacLjjmpYnraBALXLOlFdK032gf7zFyfcU89/NofZ1C9O6udXncUpS4+WO9c+UC6/O8CFpe90u
Ndrx9GZIxpYZ7at76MPjoIjeM0Dat87qfgPA7ZTjEQ4W2t2XYt2ZY5WFPh1eSSwAvw1Ner0/TxKx
d8bt+hZb5M8rLp6Sa+5xDk+u1wPWEMkAhTQCUTteKyDptaGQWtN0+Bi15fhuWvqQT8M01kHqjzxt
OAc+bRnygFWDEGwMger+IzZ+hS66cocqc7ToBODWDbeFN86t0AwCN93YWxq4BdFK3dznIRJUGWyq
CupYJ86BDvmLSGYXbcjFNbowwUBYxAhGnGnHaSXXiBT6YGl1PYC/WzEQp9LoM5ElVg6fTHwPaQ+Y
vrMtSyu5a0abKftp/wJ0dfgZS7vGrYntQcqd6+2bZXazvzLWHgFdqRFGacv1lbte7o/M4jemQFr/
nNRgK/z2Eb+eQaSgD1PRU61NuJJFFLYloHk42IdxVdNuhFjZ99q9qSdIHPgZEvXN+wpmYYXs3vr5
L4QNgokfAh6iMW2BjnmYiRTil5zr6S1DpGh7z4gZYZUJ9vRdAP5TV/nZWgaCxZ3Xi5U0xL7rWP4Y
MOqhFHGuDAXKVZKHPYg0qKC+Q0oRsuaXSy5VR4PJ53OcuZ4zBJiBWMaGOccFH40iemxJ7MbdQ2Rn
bx6+xg1R7GlW7/GUR4+6w55qVUF8EfsosNmicH6w8Rdvl7VkSZD2RoFKpf44FNvpF7OqJW75hrm1
eUZVdEirtAsl/D52IJgE3cHWPC9lSl/5Euw8tlCZkSVesjpwnwNAU+z8QAdwMNOAmiDUdoughs7U
2ZXIJTuFBry2c102MEu0IZQs+SD5wlndt0Mrm+zhR473OmELssP/xocDIg7FBTktsPuQAsXxKh2k
SW9NGWBSy6o75kjZoqA368yTvDBSthpEzGFtuOX+1ieB+lOFJZR2T5WS5rFVHtAUGWDfEa7uwb7L
FMtC/a2KGUevkxC4gC57lXKnAuW/IAnbKL18qKwI27YUVl4hgITa5ZLKmoCLhy2/sEA5G1bqkEHy
zS91E5qHTl/KNaSQPpzVGFh39RRdA+AD8OIutmxdLjc6nUx6zsxeRolt0KWSPY+2ep6hZaD5juOP
lAm7Sp1CoLtezTQNSWLoYwCcGum1Wg99PfNpYsb501eGCx43lwjcZ3OMRMkgkeNbnHEkhWdMM00t
XClTh1Z8WmEDYi0Uz06inRzCyfD++02XJS1f6CfrWzgyJKpFwLpbtCw4fY64w6uTcsxjI68pneQ+
JjoTSm/UZnV/AMTZR4pjYXdaHt1Vq8X6gXbpRxQYgjTBThKb+IYlnL+3+k1lFqGqBb0ipfhtoD4f
6g42/OMPRJf7lUhzE9in92o+esxMabM6SHk+h1tR2RPlLv/R8YWKm0WRjBCYoARM7qHX9yi1e61x
ZeQogj9Ka6DWzZOwj9X1pFNOFOtIEUNV8fgU7Il1XY4S8hIH7qHCmxpYaU0Qm0mgLSsY0sXJEahJ
Z3LvVH3vw1WEggICi/ptnJ+DBBwJpBH1EDy8Xv0MYvjhQLDiAFcZdHjh9+ebkPvCtoNt3Zz28y6M
yq0sYsP407mEHCQ1f/f0ERMxQI1XRFY4lYMuL24UdxSlZz+tlRZ5QGGcd6FUCER9KCjkZ59XgHai
pCmbFmQsnyHTBKYq97gfO1M0J/8GXRXDhGa2fe6Qxc9kCrkS3bqTPJR9ab2abFNEiyx7daqWic7C
2lniI58BxQqpEv+j8T6WPZm3rB9owHJHOE3cZ8eCtwQMhWhhrX28956nPBzmgYi2Pr8Q2G4v9LFZ
ofii2HZg35WT1wBBsp/IYeJ3nGIU0D1GBNRPiH0FpMEdvJlgkcuogpM5VcpScsZar8e8b6NwBx6N
YslVA1ITIiMsEC5Ohh2CQJsGaPMJ/MOIufhPR1eZSY64qyLb3ykZ6ccEMpE/+SgM1szzg9XO3F8n
At6mEVRxNYmM/hByERYW24EccKCdhrpxVHREEl4dRWnKTkKa2Obhf321img9Z8o6zl5pxK2JmmN2
lK2sOKtbEgNxDM4a7DCjtXj2XTXY+8WBg8Q+vxnogjV26DJ1O7PLPNNJ+/DHAi7WCA3B/h6FHVeZ
u1GO9vPSY26qaCGZGsJY3VWxnliFIU2rM3WKcBSO4DVLD5yJZbeLBJedfJfSyp29deS+/rPvydWB
E+g8QiID/HUz1k9Z86USsEERSnRMqe+hOoBcFqdtgaLDxQrXtucUrYfLkUhNzwWHaYnWY3q4HRT8
OctcysgMEVUKXYgJWfjzy0t1PDn4XROqkpiuayMf/R4I2kVopx8P9JV67RlotVcO7TBIM9YdzRLK
8BVZ50G5sLnpi4brCOsp8TCoIS+DYHxz4Htb8AuF+G/ZxGg75F8VVWmhiHlz+stK2Ce1jVtz3SrH
5pH3UQSpNzUiJ+DyNGGBQi13Slp6mLVmg4Dq0h14MHOWtL9QfYNh4BtxLahkIYlSAK8R+U/JHAtr
GlwLyrMgSNwXp9YF17U5Y9p0BKtL0ODYf+Ja5XrpntZeLbcBwT2kSt+wQ6T34lj4KxhH7c8Tz3Z0
RdNexq9k2Q+k5jwO6ht80/o5KfC3otsN9tSM3owYgysl39tbhDn1WFlEPaA3PsJd3AtBtM+eXkhT
Qj41f2eKQKnsXRo0JOURcufFrsnrUm9KYcXpaIYKY+1NJQhHWjJw/WoiA172tJAXOvLhHNIFF3CO
vcpAoB60PxKKMkEVvwFIFhYPBhQ+kQ8RxEFW/DujGhg/bNCpvdZyppejmNkygxrIWeJuOFLDCe5d
lVPfI4WSAFVtAue0EiewRqwZdtdIUAFwgPFwqA5zlom1H9eiUc4sy+UeiGWRFCrAQqDWqPsom+bo
DBaq0bLhiqLhjfl6KQjv9p934EJ6pdki87xGMkiTyH01CMAUHuySa6Gl6XE1k4xKImwRPCpwFDE8
0Eae16Vueels7XxabXzTonIT1Qg7iGmguDvCLmua5STivaFMV9F27Weye6uJa0Gklwkf13mHg8ww
ZmipfHXIZU3zesZJb8EYNpzDLFiy8UGGR4Pz7j8hskQU0KkG2a0n58BwlhNz5m7gh5QUymbiaZdd
EWHS8EtOARLaxhgqLuBNw64ZBzyNgperQuJfnJBhlunip5ciXu194HzKk2654LAg5bki76Zze/o8
5iRIRDkSaDlN+CZ9oEp0c3ORmBwIuY/sprmZglnqzXauix0PIkeQRvwSb3C4NA4EQP+unuNfmf8S
LCPTTLDxDLtehVnXoJzdw4DQ0TX8KadTjptPSNJUNmjWLA6oiUySAk2zbE3QQ/AAqfaZB5TBBHfO
GGdZAZ9/Qcjr0D3nM+kuvybRkqZyoagUR3PSgp1t6S7uLtmKh3zWup0wlzQJnGN2Zgqy64N+szcA
IB4YP7JOXK1kbPsCZw8CoBlZsN/Q3GzYEPzztTDDOeb21psHRc5Ulm8bqyXE93sFbFHIZsg9UesM
Qrhg+qwzAqVQwXRY3OJxtBCdC5HgPeCRF1nP1NnGIFBJCJnn0CNTCNSdnq+zCYFp3ABqtMU3HNL+
li9EnMFwvUjGKPphK461CkgBtK8wb/8t2PrqhN+C5dejiriooPj7V9qfp0ohV0Zcv9PdOqqs2RuD
OXK+dw0BPVzY1YMYSGpr7FcfYRLK839m5bPQQF2a4kYUD31faZvGpmoHYKu02ixr9DfqTgViKMTZ
4ASZTRqC8YTwjTdTvDw6D/fZTFT535WnBTAYo6ivymdIYJLxTNU8FD1ra1+9Sg7fdKE90+mUc6xw
cUparyerdzTA7wfgv4y/Xtgpu0fgFBUTaSSadZFQkAw9k1AX0ri6DSPL/hzMxoIhUzPalvgoMCXa
n6e2Q6x68SAUxoy5fzQ7yZwB+t9PKfEhGKApdmo04HO+p1/inZYNWkaQvdEbjSdHznJDb18bewM0
TaimXe/R4GVKWyI2o/w78g/mxeB+PZffZUB1gouu4ap+KWjgmfFoTvb1hsflgrlpUEdGw0RxJmPD
1jG1yuF/zFTtyT6in93ZiwGZ9fO2/mOlJkfeIPCOnMhIxvkfnvuI64vwOt8SbT4alKr55FUAPJGU
bFb3v0opJpuSTl7BWsi6Me2kZpiV0igmTIFtTetnM+9ywCJKc/aNvzmQHczhI2rL2H3rrjZPjlMG
3nWMAgU2qV27K6A1KuW/R6c9O1fMHifz7Bbd+f7PzTF6SqSyBCpZL7ZKmOOC2X+c5MwyHTo2dzOe
HQOLY8iF0AbdBXPMPsrQZu2HQXazQ6YVm5uCxPz4VyzMG6B2MPsdBnIXOrG18yG/y/QhApaQTosz
P5m6fA/eRbAHhyPimksIfAdOBxwnCcwTKgUxSK6uxh8n1h2AQa76xk9eUX97zebsO0/qJ81yZgFr
ml+wW83gkt+s8ENf9g/jTzZzn860eHipm3lKb38xmcRblV96q9pg1urmIIBZYGGC7RLdkkfMItzE
Zwh4Tk+jyy3rBu+PkQKT30Kvhwtmggr6/D76Tp69kkxSuwMhpZWI1I5gRunu9GMFH6x2GYs0eOYs
PA3YGFpMCS3QgAMDNDmH7k2y2cnDUZsed3SZszR/lmspY7g1tmta5VQEEeje8G+1T5oXGtsFmz8A
+2JmMmwnSG58V007XRRUTDKY0aAs99HnjXApYkeHDy4l10uP3PZ8ftxO/XH82qNj0lVrTDUYj+4x
5e0VwJmqsVH63sUu43zlbyxKc5YLeZNIaXMwkfKSviwSaU5KyolXwcmQTxG9z7aI10AK7orkulwA
e8YmyjwZWGLwz4q/heoHol2dvaoDNDivQUck+jYf5/Vr4sQwKWm+chXHRML6JHMg15regxJOi5/6
p5pvOJmdYD70NhosCuoEwfb8sLk4/29z8NMN+zK7mWAqiUdji5GHCpB+x0Us24fIxJRgDA1yzGSb
f4+ypNFE03zctLmNA/0IILafTqI8N3Q23l2xtmPsqpmwyKIRhnqjx4ZNT6II1OJyjbTKJuoFSmYt
K2ixlNzBsDVtCupg4vkwwLzEAmocKLiRICUwmmOSu4+sTUAqdCCIDZ+gRTl+5JmmJyB1XCBOQZOV
UFoOcA0F7+HcP9x4aSJw9Suvuw7YLt3jKOCr0QDEvwPmnXwfv5PQyctdCKvdvEdN5BokSzoU8uy0
ipfv/L7ovvD2cPxRTKg2MuCjfJBkLnHaC0uF3tLek4cjI6/8NilEBEuJFVKFREU4IrPt6I1lu5la
Y3xBpwGfB7PvapPZuDtErf+eNkCOXOcMp3f2eosXU5mPpztjpuTXnC8NVFEC0Y+KjA683FAsEMc7
uy9Ve4TaOnfcjbsAxNQJ76+m+BceBzMrhuX6gc0Rjij2mZIF7RkmHzPbay+V7wI99BOcfwiFYEuV
4BH6rp846Di2nZqfxt9+AG87yTllw39RAdJWk9SOk1VE6rfIz6Dtol7g1PUuf2y/XiheaPAnZft/
/FNao4qIn/Vsf6W31qEpro7VK1UyVwPjtTj4MJTPPHzme8ogZXa4daHfU3k1VZT/a9iAS6qTHaxT
ca4nSa2XQbPQIeYnWFu3wksIVnjDN3JEBluSREJpMC6xmMVeLUbJB+8z+9FdgTLgUbxjYt4KHEIh
qOVs3ooOc7hcYsRe5v3Tq5WzLe+ISc5Sm+QRod6t2gWnDCeViQxB1gbvMgs5Ed+vx5/uJ8GP8qUK
9QBp25Hgq5GvLzYtTwo/oEDILAncYMrWsR6IEqSt+NvGnP0eWR8WR8Iyx6chl9W0A1Wp97EKkBhc
cRN0BNRc1yNUCD+QgzjpUXM58yKFQcSb9vaPKS3RhNT1Wz/zvIisY68jTq5oGiSvxydwuYTda1JO
4LRxwvZFQ5UQiWY0F79ZUlm1V+fwR4Tv0aQrvxoYKF0Nyaab0e9tGdSVrdF5wtXiDytj16qJtKNM
kvMN6CTbLY/QvTOczc/cgaBGXSD2xhA3xFxfR7BFPhA7h0zOfiXisSy4euNdvHRCTLka8kROH/Bh
zVHk7ErVloth4bfiQ8xW5cqNNYozIsr9w9bDXp1hSe1lVFBD3tjv3mo8l8rI9dqst5feYe1+IdWV
2LQxD/TgqwunSnmCKun2RONbt4g95sSV6yh+TIACDy+FPfHGArb0xnYy8Q2Kbv6P0Bf5bZR6Wy/n
z/whiHXZKNzeUVrW2Zs1p6Ymmiy63i23Xu4G4PIpoIt8xSztDHK/vbOYLAXUtdBkv2elBTy5d7Te
hMNV6PIxVwkxgR2VsKx6/90V7Urxs5/SVIHtZLmunfL7YydPT8R2zLi2CEMsAu9Yx0H6j8FlW2mM
e6fW4fUr4RbcpGOTd6L/rqoi0PmK8ye+kw4l4H73VhXRahfV8rdPbo3MNgzdBOQJhTiJS56QnOjk
YpqJaex6ozSrkfTtFKk1lbVu0gQqWrO4Z+2Cm6Rb8Q1Y9yMBCKNclmfPQlVVW1YzrHXg9XI4T2z/
icmWIFMFuJuZqNNBqYN6YD60UKG4tVjRyHqfsNEKXL+8oWwwyT/v09WKwYJXP1hM05Vdx8AfXtoD
/dqIB8fMlP3vYnCQF3O3P6xuwzFdgq03tgihogzDMBOh0q3kBBKiC+VfQenKMT0TI/N1iBH7H7Ug
q3GvRPOeILezaciBBYMs6hJcrqGLbQ2EBJf3GJY3XOGYhOfvJdMm1/OCGvAmgrtKfS+VJ3heI7Qo
e8sfpnY+Ut57ujtnZE4hrOKf9a73JxjVEYbPhfoZrIem7xf0GBa/JCmwQjyIWE6wOAts0C+0Riq/
cUPrd10DVmfmG0mGHr0u8dW7bFYn/27TZbi+N5uildwOTyhiZQ0gN378bWpxPTwuUcBaGrxTSiO3
iH2fxj4Pq2ZALZaPqJIVD+ER6kjNf6FCF1nTqoK2YPbWI7JeMEN0XzqwU0745fPtjv4S0/75U1I/
ySAAmOBbyhIPUEP4RhxQ6hHNzW4r0SomT7Ihkpp/M9JDgh6EzeNVM7d3PXfkFVVnZrqqTbi6mg2V
NT6Koalqr7FJZX/pff6Ia9HC8zpX25/A6apvb9YSFxvvOEpjyXW4RO4IYCZRB8UPpdYrlicTQwBE
c0lZV20S1xcRhPqo+pVGoTS1lq1OW9z0F1gAOGU5w+K9RopCLRNaxzKoeLUX7yRzYABLCMky2lHt
PjOy0Rghxj+1diqPLtfozBQ9UZzGi+nm206ATWMQu4KRRs/LXrBdO+FQ7nbBDNShrBOWEegHyvGk
mOdojCB319lAV1O8GWN4CypL44nw5Vy+mJvt9QhZ4ow8QYfz+0CEnxyAfvL5V9WVCOBqgs5emYg+
nRhsok46rYAITPeAhTnQ1so/UNBEwyAooB9fO4NG0jbP+F7c6cdvmE7WkwCArv+ZAzzBWLZDbRSM
u3xkp2FE3WKwSTaPupnuNqLdfT99/n+SeRxRi1VlkhgyZJDms1HybrIuo+8VmtXyYDANtQWakuht
yzsVf2YbwSrQd0bsmZcqfsZ+9W+yS3zQrpO0vG61oE/ovhZPWkTRy2VSv8Fnz4xANSiFvfJDyGUT
sBlWFuhCFjkWUtiN1+yrN+etMvt+Zl3Yy+Bdd8zEKmvAw87UnH0OKQ4YkqLYBRSeosJM21M3M+Xn
I9Db6YCIgxf4XouCj5q8Jq27J0QL/eyuTJhKqMhhTKIGQaY/g2+mI3yDgWW3Aui1nUz3CcMELsBa
vtEfb1lUFU0enWaRvs+KvteM0bX2B/IdMvh3Liw8DuYvlMDGp9SIVJ4SWKH09VRK/ft87zDaAkeZ
HSRHeM+4wiGKDTT+tq4yGGq9XQcOlc9+TQro+0zlTSluxIJYjzaskaxrEWUvoS/QLCH/ZRBNrqHE
FaYufenbQM5H1DylEBkuqVcg2F9e/2nzoM0dUTNrVW1ZwDHNqGwePMD0iLu/NY438xc3AWDsple1
a/0m5R2wYL1YGkXevYDkHL5oT1eP6MJBqLB+GllXqIyypDJKoJrL+kO3JuHZAbiI5fGIB3cQjjMU
wejMvvUpwZE4t8r7lrVW6H4q7CZ3kml9Z7SwqogGvEZ5XlktdQK4I9fJgi2tyjM7dLDjXwSYGh4/
K1SDIZCxzV6/l89sFjakDHadkwHT9/GyoW74c+67LgizCG0ty/OXHpMMTn/NmAShikol85pikqq+
8M+e3oxYvqFyIiAGPSbUaHfFB4JdJRw8NgIwq/RcdisWVvCg5KaTBZQZnrxESsyujFTz5U9a5FOM
pQgVf8YvsR3RaRLaJL+wVEFI7866J9ZhpZ6v17XPOPYObuTgNWKdXOtv5R3knzmTWO8GqYyXbmit
rfC3VqxH0ojQOqnAsSv+kUihXzIO7AqoKgsUwbn/hGLbEkFWLQ0zUji6BWQps/vO6ntAl8maEyH5
5vyVPNhCVKSxSLw4Rs7djL5kPZZ3K46YthAqQ5vifdn3TsaQGC/AWjk8jTFEWEM9B58t4G6JLR6+
dCn91ieuy0Yam33kuA+RAYUr4E7IOpIonzcX2KN4405Q9ZXVQ8zmT0liMoDVSKlXkuWoo9IscAlM
qDR2X6unwdQbZXR1nDQSsIgOUGAbEcsA5QZbObMofnbwEHbhcja/lhEfhZs3DM1ZTq1egDLH+WbH
Rp6PdorIM3KLTAR03kg8ZmrkaIYZhAqNAsBufvdLHhqCMlvvgwlGyDbaceth2JdO8vGsRuxxZ2SW
If1wPwDVXr6fxG2R8q4+znpBYdK83WVVQH1wV3Fbbs0x5+au2gBa4360dgnQ/Km53eSWJRLm3kVt
f4oXVITxXbPTshUjr55NhTaAZCPc7eaoOD/tnQUwSYZbOFff+cMoCLHLq+QVsp5Zw8IcXphhnlEn
6OJhoJpgVVlAdU096ytStpDPG+ir9vYIBIp4MHf49ERe1r3XeEyvaXWrelQgifOrkQ9XTKhIKvxQ
rXMZeeSQFYBO1KiDWN0e0OT7Z4AIc02Gsdkr0N+ciL/HteMV+V1KnZzU8VHRWA2CTyafVr3zrsDX
ytjWSErINUwcyqVdA55ic1cC51/yo+PpOydPsxsBg09wv0e0FJlBF09I6/L5PJD6X3zbCZ6Ea5nj
HyoaKpsUn+5JbrjB237iMHynykiJEq5xVxdt4MPyHJayVf5gzFCxVxPKGlFHQB2gv8UWEcUd8eDy
8QRYZtEwDjOIQWx7HSphPCuEgh+IOfVw+jUF0BjVNOzdEoFKUcSZLJ6zAnE+EtedqjXO9+lFfwdj
dfXqz9+90H6qmBWRmegZwyxVWtnjAHJI9Mw8nO/lX+KkX7ImnMIiQiYCDu7lu9pa9c0/0cd63FFc
zyEaNrZbTFGJnOv8K54pDunSSX3xtBjtgkd/L1U3mW4geaVBrGC9thcP501PBvYJIbyv9B58dxiX
uD8MEF35N1f9a63xNS4pLKhFZi3b1W4yJB+vWvZ+stbaivX/mVQMl2kwyvM98UbPge5jpb/cvOPW
QMKMi+N09qFrDolYI9FYJ9m35jCPjyCepE6eckTwFi9T9VebRr5nE4ZgEfVbnt8FOyiAVfw4rUwm
4HLuF6840weVZYqjs8rSuWTorNXDZ3bGvLuM9bAt9U+igi7R+sMEiQucUlmllG+SpagZYNrPydNV
di1YE51/zbIt/TLI7KXiqbnQQS92Q8u7QiMgOmoOB51M529L6xOHtEbkNEBgUJqFcJjt7q/NzcJU
aQFWemQ2g5XtxsXBMyLZAy51CI9TEJ+yWAIKjTm9Te+bQQnLSsYkjUlVLJEp6r8P64iVPxXvieNg
5T5weuRvLaNtpHyR8mXWgvwBCZ1IEctFrwFBXxZu8Mqaq5KbxePZOTCPNKZ5vsRtaZKrM0hXVLdP
EOAGDDQ8Y6UGS8syBv4QHUqZbCOyiygtdYpd/Azk+pnt2BxJfzJVxuFBdPyx1tj0tVWu0MSKRVTP
kArR0qYNWhgryLcSDAqoJNeTuXQqlbqKkpCXbUj+30Luhk3g5RRlQ9wsNwy+mp58bYMXhnsKPHei
p5ybBfqG/GlOSxF0lLw+o+bAmf8D1qH130x7JtzWn3actuYL/YP5+y8P7NocJ9BgrxhTzMtTwPsl
5K69QdyqBAj51Inl04GUaFjHd04tsPCztllG6vaMTlTXBCMpxDhzW+12k3W+Y+cxVajVGfpuSVFE
oPdye93nt2YbYx+vMW7VhaBb184XZOnF9GwNhEIGrNlUn4s+yzS3sXfdqqqyJULTbLodpv8sdull
dI4LF4xd/X1ypCpYON0fnNuQnhhUmhVCWZc8GswG1y/UUGoikIKGtigG/Srt58yGn3M23MamQajv
lhhrV0nPWm07qYE2A5D2qBWnryyPUv5gWVWcCaEC7mX6FfOdvA8gQSK9pzF30X/coQIjKx5L4g1m
i73c05K1t+jn70lHPwarhgOWudxx3+88DfebkTUAXO8V6p888Ow54HRNYNMXE0SxngyDdJ1cqux4
b6tBy6YRkVe6blOxg62/Wi0DxsqBlFcoNXrjCyup5PaRqLZNNII7zaUB9qAQu4m1TO9AC3VlvSWE
12CzWK73s6m78YOvWuCU3zmktoX1t+V7Mm3GhGaOtbhvZZEX4ODGUH5aGVruCRVwbS3kY+tP94x4
BA0K/KSWbEhjL0u0BbnNocwyKD/aBB4G1+SpEfI1dTHExaJtBuvsuzd17sMe1CVkqv3gsaoJl9pJ
cXoOTk3iz3izdqWrydE2L6XZvzm1+kwjC6iFEYg1nQaJL+GsFkCAM70DBQxfetAy/6SjVkV58Diu
dumlcFXjPeQ6bbP7Gj3wtEO1ZQMMZLkrd16U5M4V6Q2iZd8iCvHBmheZ/pMatUuV/vv3haV8QKlO
xRM+5b//srmwN82TuTdrZT5JDnYCd1u1BCo68iUD7OynIap2r0E76iv5ss/ii8/9v5HT+NbG4SP/
/owj+o5Jcle1HY/WLMl3nPlHb3nHSx0TIlbbP/5hW/4yNh+OUxx16AE6nVrnixkefE+8c1aHTV4D
6JvM7Dpah0DHqZ55u3FdA4CQmy+9i7mNCHBjr8XoR8bO4tZRrZfSERfkPYaeQ95yxxbUl/F8G1yU
yvvVJy+wcWE+Ytafh9fTsubyheEXiRbHOBDdPAZvcF6+3RcN+RuRTvFZH8kRGX7vXYgUw5dgrLGA
rcX1fsTEDLsx8q0da0+uodgGObLOgq1FLOETPG/baRVf/XUofurhQ4l6/Ge2Q0JeZbttRscrEsQa
gEmYI+atyw1TznknKqUAhnW7Rjuk6PiAlhZa+Vs85KcfRKDU66c9hnzyUggaM6WgjEsAaKJzoM1l
S3BVPota6ZKtwkU7sDxOIVgM2sGJXfTqCllHv6PGYPL2KpiO4P/gi6KIVmy3VbjNKxnsBRcoD7ub
ELd9jnBNc2MqxceZiJCa+OB3orImiPWgaotlOZcIAfLjVBSu+WKHjnBNf5nTI8lrIpyFhTcwZ9JS
Nl5qul1jAVgm2vJJfNwY9WO3U3p3M3oL8B2S90phuhPhAOxS9nXi3Qo2grEX/rI6dQdVghFQuVQE
FuhVYzHuMrkRYcejYhLDMyaJFZlkqPlAthgCEpIkZ1ZgURGPBdE6x0fo6tqPZAFmZ7/HVE3vNvxC
2M4+lKCsG+CztErWM48jj5kuUhYCVebN7hAIh8T+x6pvDHkr11VbnFee8wZfRQnjDU9KSgUP9NWw
C3VRu7aRmYkWrP5wjkCY/ZMJfUAs608taBJwhGL4fRH4FjO+gyLxTktjsgiY31iQUCqr+pVHK/PS
njXHsnfwGRJ0EqmIzxFQsSbvYei3pFx7dJAdlopPa2mVu4MeeOXPdXvX8sziXqTwHz8dolfJlaij
o2WK0LPwt+gbVeZ6IkJoTY25VsoOtRYrQlq8AtJgcFVSncaeYG3wGnPUEYOd04ZbqNs9vk4NG7Tx
5oLMyLo6v6yNQNszCzCBX7Kh5Emd/PHXsZ33H6sHH1aD/JvQ7fBGpT/DtIOhHieNP2A1RUZXnLP3
cP//LeY8G1Tr8BGYa3ArhDKJuQtc2rOuIQhYK892Ek1vnzwClRIfkoHzhqchog9qfdRhVUbvAd3T
VcG0sQBZzm4NMFexAmOVO8XD3aocNKcPfdLflVy6G3eHu3V1c3V6PvM9LYulfm6OVUeERzqG5rvn
uaNf+u9Nj2fEJPRB/37A0wWBufWoYU1Fm8aEBm2xyxX7KHvVAYuiXeKPXSUzI/K2a/IL+NGnpfvh
Eh3O/2HZa9+cGbo9WjDGMcoNwv79m5U4t5MfNID9p6Z4XP7bbMxGFYDu9Pgq8ero2M32qKR48+Ji
AebpPoP75l+fsYtFyrvxtWMFzTr0KF7yjuBbhvjSibRpPlRyQxYViDoCe4Wm0ooM6Of9yJF3Pf5P
RDWK8YZwpfjgWX5v52W9Ryt1I+IP0yt6Tm2qqXEj+uEEwdFIHsAlFNQ2Eb6VDX4PibFBJj889rCt
VrfcYZ+LoYaKOErmVgpNvV2IJdhzE0WxOdRAHX3AoHUxsPO87HAcwvdJ/608pMJid9VFpPoVWXyA
DtKZFCwQGEas1M0ucl6PvV70TGgh7ENWL+h9b8dvHl0L9+514iiHQnmH+DJheBbKnSggjc35Ucdd
EpZ0eCuWy1NtGfYemPw9jtlkZGZwuiWNL5vRxFExqsbAYKNVtCFU3ghu8a4leAILtMBzz+9yWGno
DuiVmI8yf0BOh0+h9cJxkBZjW5gWH1hI/6Nz6j3rY1eS2q28OaQAdZ6Dbg6Ztf7jG3MyS2qpGryx
QlZ9LZItRehrrRpsP6jNqg0jFBEI1eF0YHhMR5HWBPLsKVQfAParYFnJMpvROghfAGnKycPreDmQ
ESCHVglP+4gctGZdjFgqmwMw/R/uc5ewileE/WVAcmGfLH58hZMfvh782JSrzrdjal/eQ9bDX++T
bvZErXBx94ua5EIdLgtq2dFPKWhW1xspoT8TyTvgTvhEpeKIDePnhLElr5U+OBN695aj1jckdLzV
ePe6o0p0sLMIh2cHpgDC1iESXzw+IH3yWxilOSTKC8o/JzsdSdB6Ev1mZ1BN40f/8ajpBA7X/XXl
y5Lzxdrfobwq08daSGJ8SH5CvGWWSq3lYmSbzIS2e2DMnUHN1Imfvt5cJfOEud1ClaFlegFF4yC1
UR5aBD0c5f61KulQDMwQTmfe7rz2MU0SvBk7t0kDCRy8b4DW9S2EVJP0w26fAEpPrUbGphvHvDJ7
i44QR3XeoWY27SuAfvQU+haEhxBxWkLlmGFEr7X5ETdx7s7te3igc5OP+JHMkNs5vo70XmHyn2OJ
zVdPtjAiElhJkLTXlGA97a3iJ/XW8jPVb3s9yvhhVMAxnSOCym6Oom99cYFfa1MnduLgvQSXGxhx
ZruQaItvVw5003XzgUHZ9JYEMr9w4wkLqsin026GMl+QCvFZQL5YOOWB5BicK2UyRVQgIFBiQiKF
r9uZI9GjgyoC5RtMtyC5hofbLkF2EA0/nlPOZIWQHZuLKGfhAn8XwUdZLPp/YOJ/36clK3FiAHfM
J6inIFknETLBEKj/VxpumZfChQNOjvrY/unCMB0NbKWnXxheAl3RYxkUDOXWVTi5FmkuJ3By+R2w
9t5K7h6Jhd+6vKdV+hMSnIMogbY/a9IAZPSfzOcSIbjWnHhG5sRjtElNKzDdU0vY9QFaHl1ujcEr
Fhfvd5Z0aSEDL7SQoJmA45+frgvx9AP5WNUfs1XstpXjWOtqexdxNFie0ZD0Y21OC3HdnP0/qPHC
2fjfD2TZTLnBnxrfJ2s+eyEK6cCaRDIHBgwb0+PN4462s+ylSZQdXY97unNNLNbnJKk8dlaJ0ru+
Va0COwZKE6/Z1tfVsbOdjKcIQwNiQYg8LVeSWLnNwWfj+GsvWGRk0RA10ScCweqFDUiLzqQSf8Rr
iOebNFoQn9q8vrl27ZD8sHLyeOdqZ7mDIEaSpFW+WLepNFxq70W2crtue1yrMaRenG01DAx9docR
SxGwWp8jg3T6pUzDHJK07JqcnuKaqCM0B5wjNStq0ZN6EHIPVOul43KRXx96VbT4R20Q4NqQTzFF
PDjsRqMwspSZvWfUKqQGf3gK69sizTpRQAyfOenzG5jXwn1v7QpO4t5ZwFyXPOxumJ9M6nIWYmfS
oNe2D2z7f/n6rVxOsmcB631j+X2f9NgHCWn4yfc6Kjn8Uly/fh/OQMmmX10zSHf5KJ/7RIiUfT3f
srQ8ouzaKY8lZX9FOU9UlG+NvwNOk0HWDbXXQ757Q4uuoBLTtpGo6tu7VEjTBMO1r419G445qWVE
kFAvuF6Rmmv45xha1MjShoNX9fAl7HAIYb3vfUOLgLGR4FrKIEDAd2w3R8s6KlURxOXZKKVotlJ7
9+fyzN6RTIfGL1TdGSas76QSpCHYLm9Na+Bj88nCUsOASRyw4yH9ghgwP3CBklMqkKsl4qZqj++M
PvAh4twe2d3Wp8zqgtwE2Oj4mAVxu9wCFXM7W4wDT8t7JIFBhLQ4OASquRO+ebQBYUlj/PuhjlLL
XkDsv9jCHRV5a6Qj59L/ClVfH0Xanj3Os8Yl9XmbuiAtL9jj7bEFzzNUuEsMKLcu1kZFNKGGQvoC
xhbBdm5jzdBIHB6zNKbucKFlyAIjuUzKVKwzkXCG33zfcPxtENdKOwJnnYndCLL3tIR7itLLR7WN
jEhwQasjzKp7svETciKuPzGeW7yH6hvV2lGgNy5crfIcPhaGSmrgd+BJs2OlY7V9op7W8zARbz/A
UKK3u9jgGGDTXTopYy0tzXJpInvtjGhqfP+E72W7N3BxrXqwSN0crwKtSe1M6GMWP1r6e+C8lLGb
yE+hVgm61Hzuoq8c8MXQuIsLxuiFzzSOmGCdrbAAU18f0SMw4MC7oFUnyBbsxU/68qSUWz4KKQCr
X+Jj1HQxgezuWxZ2pD488iPE5cgYddNf+QzUmtPMe36EeGMSsUjQLKZxEZZT6MukfKkBz/doCgr2
Jb2leUnY8EIBDbDqtoMuQIFfvWIdDX1yAfqCJRc/K00qZSNNIMZ3CACkUQU66Q8xRVLT/zIBBdwy
aLYg7tQRJKmDwtZCQcKZhXu9nlB0WOPWp3DDJ/X7/E9IZCp0o72DhSmVEewubGYNSshK66gK4JyA
fm5U9xJbdFoI8hDdev+d2QtTF8ErdaMxI00HmTpxCfLXQ6Wy+QLc1fjN4mCtY9OL1a6xigDz0tP9
McntkULEAewgSCCVLtxshlKhy1D26c/2/W2kscUoWbsH5V/z4UhGlOKUfko6+u0noWp7Jho3DITG
kZcVS9HFV9IZ5SIEKbEiQlOi+BDeVrdxb5SU5C5B7Etp5WIBgL6VGvnSeGybhiz6HBsV+vmU0m7C
V+yl5sseI/piKYUz2r1lat1Kob+3uvZvkFXOx2mjdq6sDGMHAbRo7/8EhZAA3+HHm97P7vlbzmd8
zqdUA6284ZTwENM+QbstBFGQVNDohJG4SDygceEj5672N8gMmui2p6rwFrLOAL6HEEmqItR0g+Wo
J/R0t6DO77DZ4gaWoSjUKI9Ee6iY8+WMPevCG7MUUso5WrcrXAdyFEon8iEAXlB7ddqydr7ZempT
1vtEPd61WtvR8npUve5VsZeRyaZZ+/tDpZp1QrSw4BHCH8VR7/gySJor5HjF2y2Y8RdF6qezZmvd
RrpaXhIvbMB92Rhtzn73i56Xe5YEdD8nX4JbrfcB20gHKxxYULal7ghZyJemfETQYgNzrwvOWzpp
d3sjtH6BKbmu5ViqFOURyQOu7Q5Dk6kCKFod2A93wuEijzBEPbUbnX6XYZgWYgh39+7kqXMwz9qB
ZPo7ZEusIUFWnhqYzSnUBKdmCt7pdE2taefVAxNpLAE5PeKEgzN4Sv3DzQnKLxlp/9MnnL4xykh8
v4uA8KRykqorxdpb72enwxNRQ+cSo2EQGCdPAeoBpmhQn7XEXHA3rqCcR5uHZQXgwKMv7NbmXBAK
U/C2VWf4q3CpN6RRVuUpoy5Yd9o3IfQQYd0W1ZKZn58PNPGp2HiRqFUucxUvgzG20vQKkr28Zifs
KHLBIjohNSZ95XviO388pkCcdyfCBJhtADq1WlkvSEvQGmfcSDjF+6unOxG9Do6W4hG6qAhbMl+M
ylqjHUkdGkoRbRf+vOjjmyXYncukzIHGBC/+bCIMSHBeF6/ocybOIlYHRKt5d8J+z4slFdqQEFb4
Gwj+XPzTzbZeU09A/isckdTC1kcYZw2vvQDG5EGWWkaLekrHoxyYZN14XE5htvymNLn5mgunG3j2
0jKCJsnBBTC3lel0sJMnWIWqaVb5pzxXpooJ13Dm4a533g3NY4cAdPAP2guYZGssLuL7WhDBRnAZ
XdpeE6a0oI+R5q9qZM7HFQyT/W3SMRNch+GCIlxL/t2HvPS04i7miWYpb6DZ9s8BmwXEM3LuuzbN
UeX6aEyVryMr6oerZ0el3jn+Ssgx2Qy/Tz85Lf6d2xJ+CnJtwMhjHYVLl4loyduVy//49ZlJwgb4
llrzyA5awQqEDa94Km7+3sNNi9Cj1+ZBuQBGIyd7Jg9PC0osdj6ahmgwKD3g/hcJiBBy7OSIFq7M
pbfueEL5xegm2HtsaMZ3UqncdovxKvbUbzxsSOuc3gPq12Ue9a8yuDSWistx8FktSFWSbg9Xn2/h
gxJYiX8YQ7aAux3TalZj/pVaG11aWDVPkAb8vKjGOfTyajtskiXV4+y+7QaC9e41Sb0iK0jnQ7up
QkRmaoOhSjCBB9nbz+uN5Nrg7wONKUdKu4qSWiANYp1gxdXqMf2SWs+D23tfnBcdftRDSDPS8MzU
tVwnb4pTuUllJBsCr+NuYgVaiir23go47ASozJHzWx1UL3tKyBV75WEIl4gHQpkQb8Ipe8+lNbKw
HTEVetUkgoq6YcrggWmQsWQnfuBbOZ01gfEI0L1L0WQNBUow/g3+roVpL3yb+fzw4jn1qQKvDeIH
c5xIwleL7QjL9Ka/f0KDKbMuz8aZOHV5j4wC/U5p+4LSK1NbfgtJZ93tE2Uatq0oA2V82tm/Mop6
+tfRol+KqnOEVOo713eUS4rD7zKuaeJ+RkrPVnv09bCHE0jISLnKcsLKZ6x79ycMT6vijxIhKmWj
6IXRXBvaRk5Ii/Gy/Cmd7+PqgoPzLodoLCO3P7PggX6STVVtHEz+IwDZsxciKqYRknBJfgnje+ni
JwKes4Uj6wN6t1lOiAVlrH641UOSqXSkRofAl7Bjx7OZUkOChxj1xjnrWW2092MYhcmf5Cplz8LB
djyy4uXRpkr1JPCpOliqjxiRQIu5kzK0vbuJVxKhh6RqdJ0JkHMKIvYjdrFZ5HhoSo0jg0O4kvFk
Pk8tMlmFBEf1JuCgmR+sNz9Ep8gT/oDrJQO4ZOkLID+xbdBI71iznFG7iV8ODOaGuJRIE+afk0qa
K18v+mSf80UsCmyIl6iwlpYCQRdwa0C6UQ1hNQxlA6icPYJ3y1CQ7gOuLw9lXHTO37LnYGNC9dQK
HyWx202UOGkTxFhq/fI653jN72kpo8yWLxcDbYKiqkoRzOoYcYHwlAB8JnQHlJQI0pY7C05IMsK1
k/KXcBTgkXYZVFrV6Y/d1+TRm5ztjBaSoQLgen3zKBciKzGPcjeke6wqHQWUSQpMWX1rVSVws002
mtOPYGhLyinQ+jIFICMsZDT7dH8KJ+QfntHtKJpLdU/3Q6aho0hOXbOGRmJWVtz0bFyCPT9xEPH1
hScenR/+MVeNg0tRlrJHLrWj8N+GCIEohgFZpidtDbdc0x0MOGduyxmPKxrlwTv43IbuGTKVuRJZ
9KybhQJT8kz0o6jXwgno0Ue8bDB9qubO/jxkSrwWbeQrFRRGhTHw6TmEJF3iRf3ctkUO1SDIARFg
yOPUdEkcicPkK5SJ2hVZ2J3LEeLl+FIxsI/Tu1dTvF+dQ/Ib3GdrrOWihMO5Lv1o/Owmlx2eiHNV
YnUycoF8T9PrCTHAyzver8sS0SdR3JdhMc6hD6KHqAj9Pd8RsJ0Kh9BKQc3RCH0HrZa72xtuw48Z
X2NrMKiK1cUkxHsU3PrewMEEy0Wf54J3m7eCCMlzoz/I0ecn8tKaGEwvP5DYW6qwM9TnZOe5DTuU
WWLDjc0DWolOb7+2FxMGOFCNb8ndoEKe9zLfibroUh8CAkLqHR5dgj3r2ltazBJ6zv7/Y0NLSFj3
PEiZIqjN+QFSA9eoLGHHIkjoglFlOkBn4eu1av1yt4k99w3Ln82CpCEZTf6i3nLie4EkDT+2lq7O
rcLonugUiKOaeKLZvP/Q50j7AetDwyxOZdnntQCbRnuBT44v8NHtVIzV7lHDRlF2/pH2R8uUESN2
2IunxvtDmk4pTQsBm0QocL5AuybIAdF3/v1+q/lHNyVpOG059Cw/kV9yxpxVSuac6L7ESLeAvjde
2qlp5puUJ3bV3aIsLONi2WWI4D4uq7Kgovii82QQKQUG8VGf4JiHJZPWO62MJb/uLMACAt02E076
bs2lpaQj5sh5g09eOlGhurNxGHSfqdIUQZmOdhYAG/RLy5ZFoF9GFEqiQsnTm1GNXBwfpKDhSSJn
W2Gi95wpmYbU5iyzc8itPQUTVuomxTdDqWctWTAQzy+H0VfZnX2Y1mt/0NjK4GiFabPzDNg/1L1e
5/lY4NeNlYhpJ7fOXI+581MpSHIqmu9y6Rr+F443HZIniHamS9kTRD3X71GcwH+gghV8QUwwsq/h
wekjFqptkIDO/nzuTgig6iVMXqIU4rw8zS4EVOHml9k+ryIByX58XomAVEffZn7cuRtR21I54Ef+
RMFCp1077IlpvXE2D4awG9oePxKRgv9tsKJtYR1o6uQEMnsORD4l6S+1c7zXrASgfrQEm2Iaszeq
M+EOO6hwFSPS+oqpe1NgJ88dPa18U+gzr+qh9+dT90gkRxbbBALfnvEagWwHJS7dQ3u67oQ90byb
q29sD6oUmLaH1Kvvlf39LY31mAR/ppb05AxS9JGgsu3q6lj7/tk86hGp7weyjY3vl/WuXR+8AEOy
keqG4wkzAF6JrmztnDEIc9pCDNbQh/I8MapzyGynSxy5g4qSjnT61BeVirORa79wPoftdPXIlreD
4ncgv7v7OxiqiUFTgq8uWcZV9hCJVuYt3wYFohZona4f1gZiR22HgL4SDPE88tjWp54kyew8etD3
FZnSCLkV5/QuHHkkZ74nFcydhOuQiDrzNMfNfPWCaKwW53nWS3x+ptBvZ7VKXvlpqN8uCK6LKVVb
qvb0S0owqVYN/uhx88AY7aent5B/kpHy09fHCC8Ah6EYaRIAiry/HAooJ968YYFLEv5efuVNx4IC
prmGuHd4MSYC3vWkCmW4goExSJNCa0VTXC4KM3aZ1RLrppzs3sA9JV/Q2PT67R69ddIu+f4oBbTB
WTLk0C4/GVv71MCOOWo5DvMtN5v5pr5DG3aoUH1sLvBhacdBL3OvPZrlsvAoXnzvlBfgvyy7IbeU
zsMzkS5tVz7tosdXKt6DiJPhOrd/ejUhYrGmDcGzecDjbw9TuugGkexo/29ZbA52Hgz5jr/C+38P
YFDbuWyiVW5O9TuO2HOlKGsrd8UByj9JCLIgA0cI8NFqMlJyn2sgBvaXVALkbL6bk/zepm5YbXhI
QdggAtSphBatHckyaNbwfLItSV3Diap9rLoys6dOBwYjLijGzPBu1uyH2AywfNiiVCmnEqntMCF+
wPxZ2DmOvGXVvPvCu5RkfUPtsnrDhKOW8syZtbN48nCAeUi9JDXenrSsNVTMrLgdgfhXuTmRB1PH
h38t0fDvA2s54NY7aQbZVHt8NdebJvgp0LgmFSe3YRcI0q23HbGZ9zNqd+T3Q4GFw7ZLS5pB1nZs
ezuO2NvY0ExWULJe6PZBGSbSJoKgTXPEIbh717SnYtwEje/h6GLElxhAMB2CD69bku80lmVhxdEl
fPBISV1HWAumDjMaCxSNsAQ9sFj3A+HhN7GnKRj7Qm3RBG/1WjIjMbSXOwyOcUmqc3OKDZO+6k/c
xRNRLN6XXOJVTvA8Xa9olJ/e+9ieQqTsyGmIb3YczCqGMO4FJS18RYAXUfqoII08gbNMcJx7slKR
ndpq3jYCRx3JKDiwQhcbjtaEW4mP9OnOjnij5cfuUXJJlsAb+6Q5Z03ul0qNyd50Kxc4hYyQGhp6
XxcFIuDJnWb5eWtENowv/7/9A7n03Ro/DSeEv40z/1A+WpGOoC/7YVtMz0DX2GPLNXf1TQzSpD7M
zN8LoVZdf2pK13B9l5ZWhUzEbzu2o+23SpYq7XUOO4WrIVCJ5JYFKQsmaChQyYySVkVnMzQrviTG
7Kg3BJXdLtD65BamRtYqul5GJyD3ejRhWmvGaW0LhwwKeBXB2LcNePGjneLwrE6STVecPDwMQJ0L
yMAf0KYL2K6KvuSLEJkHsn3W7lek+k2wDEEFYEzYYwS0HxAkfEsr23vaOaSYbeUUUk98oSMRanDB
z7FADfXneBz//eItTth/m45mPr3oRzXWT8aYVX+izZ8Rtbd6ddhp4txTW1KR3+1z+VP1Kax+tSdh
co+7I/jglhXT6s/we89psL8wsk/3gnoOjjNWmX7M73v5K5hbnj4uZVGHrAeUypYuU5T5k3pMzMuK
SgSrTu79IK0zOHMFsnfPWRe6smGacYYi1EGrxCBTUWRcbYng6udJ84yztyoRy2bCa0F8fEu8JlSH
Tt+5cximLgd8ekQjqighHiPUf15Flkld0g/nSRx8S46WvCCKhe8wzJjuB+hqYgz8ZyH9hjSe8cP1
XOCXx2GB2iS5v53D/pSwb2ERF54FItNhwRRyW0NlIZ7Y48JEb9ypgffsG/lv7mH/jrAbdU5lOZEN
mdbWThaoAdXNo7nvrAtsZbBIYmMmcjBtb2Co9frdO8kj6SrO8I6osUhcO8FU0NOE6nEuOvmNMt4a
gbeJ9UztcvR0XJWliBsGcWJTVOTlsviriJV8ABw1+b3er7ssTErm5+sa1//tonf7qLdlrEkDRQ5W
tLobBuXio1Q0m6Ki9uyywl+0rkyL1UVIauXA9Ameu2s2FXvlZY9JkC6p5fBTaJWreQaBAAZNBNUc
cU2yzDI5fjDGIbn9By4cELlqYb7XhsDHZzsZpsG47+NZe7ZWXpy3iAXuAYLu7nXW1jv58aRwHb79
/kdO4nysQwReCPQGLSZ3PeIA2a4AK2clcc7kJi3dAjOoJ9JDBRtBUI+0BIdoPWZM3MQ8wZu4Nn3m
NL/B1LyIogh2TSXJJmwYcI6WjaCo2ByA4iIJ4jvmRdOMNneNdoDgR8uwCMak+qfyEF1S2dTY38Em
4b3FtlmUBy0M5Dg/ypCFeUcseFWEHtxa6Gw75HEEwaEZhy6UrXFQWOd529TYzG3gyAasWK9e/eox
8k1KP3GoFFo3FYKHmDJjEurIBfL7s5iknlgJ/QvP60F9mksOrJik2TZqZFropr5u+uos/2Xy5L3x
Du2UgbeHXai2N5n3+GzTc8FsMYn3G7UMwWeUYukI3ryDmVfsdSRo42W/0/L/VAl6QBsjmOgE1cnh
4M74CSpTTBeQjJMpf94yY7j0tTgoBvjyO1Se3RJedpOyQmhSKIishfQoSDORUy4J9h/y7mpqk1q5
v3LdAUExscPZmolbN/F+QVy+Yegj+viPN3s6eoYeor7Zsk2hy/kV32ctMQA/qHJdqXUeffDQ1mAc
xAwGo79bRxO0xN8QmI+reGmXh1DYAYaFE09eDNk1JLTD+nnP0eAkULMg/ttd51J3s00Kh0yy+lUO
gwSMEgIutbMnUKk3rr/AKDvE5/r2JPXJun2qq3pwN7IkmlLJPEPFLtRF/r0NHQu5iD1z9tGqr85I
FqILh4io+xgiHLJYvJnF3GwPkftAyepSS+sb/CBoTz5llJaxlvkLW8gRsCr/lc57qSQlg20Ew2Kk
AX5fBzjhTOMYH0OeH++taNWS9daGRjpdLBdf6JygxKoftiVpYni3Ewx8r4QI8CoZy3TlHGgGX3qu
xBpIlE85GuRC1dpCx2C3JtCubJ0ly47TZBQe7SN+weyIqnu0e7FDp2qP1msokTo8pN88IdDE1cT/
DmHcelItjsOl+J2NPOmG3IZ0zCNRRkrMnZghjxtmVSREoCNWa+7gbzZX3qqDOg83wHNayscWnlse
RduI9WQoG8wEc1B6n8UUh8dWTZ/8QlEYSUHE8rvJVSsuLAnzwojakMtj7sJ99FOZ5IiEn4f7J6mz
HVZA0gAgzNxUfzLnCmS8Uoudmi5hCThHwOod60cTIJ3WFKNLDFnJPxUPO0K0A9j82GcpAeVQgPVd
mvvtMxCElcEN7sY0T7vBRp3udFoLjKZt59wUTtPAGifHvP9HLqvuR1JxZ1CzUht2fYdm8KdTz99T
a15G0sOTIlLt/SmC9qLOHKCM5x8rsN6+TlgO/dLOsqnKe0utVYv/UtYQeZG+q36jPHZ3mWVTtzT2
3IYigE3zYaJi3R70L1PvD8RV6kfm4gA3biXVDFLMkO+dktZxwdug9HIMwuTDwhDrHYG84lz0cEw7
ayodqpH+6X/sFhrhmrvxFb1dY9Q2XgQW0kKXQJWWCjDejLlf4sAF0k3wOHzaRZ3n5KddZhP7Mbt4
K64SvoLqrkvOhr46Nsl1FpAW+adAag7FMIwRn1/Kuu52kvKixTrJOr9MEvKVNMMPbzePhk/7x39P
EdTwUTDxLjmSwkfFxy4gEHm/YKyXmiyPtk0THrZ9++4OIkrGglnLLuMchNbEp9Ier1AbTGMbT2Qu
miY8Kq9XrLTL6dL7o4jbDGIq5mOfklXHGL2XB9cZBfZzHIR/9nm1LlrVj9OLpxbOakkk2LLeW7E6
9W9Xl/u2Pxv4LjY+9zlMMI8E+MPdRzaOFYmMRL/0HkqBvcC5zFXBO20SWeH74XDL6LHFoU5J1WJ8
B3v2tWwBy5U7ljo6S3spylxDZECxz1IEwthLtHHtQ87tFctRTTLEegO/slb8y5CjRc/4Gbh6phZl
XYVtD0j0LBPxdZFnuC/c/zNm7fWf63N9Urn6dh9tMKNUiBgR9dzPN48xyqLRt5ZAGG9t4W6Nr3Ko
N1dXrN1L0RGp13qvmiSwpoKsgwfKcfDv1cJyLM1WJldTYFi2rZ5dnzvoZUgwjzRtn/G6ZqLSIIvH
TCVpY3/mZPE5Pn9xSDXMHYinHpiXHnGB2fLfoHjrEfayKjk3OGzVHpSbc0gi3Bkley+jZT5aK0Oo
4K+ojQ0JiZkBpl+7bCrPrDxfIll8tzO7pNut0v3bPfja+i4evimhLhQymaJxgZEtEzeVW8p/Ij4Q
xh3PSla0yZmUozBz8vXlbm8+0SFVa2fbmpRwJYpXXaECVuPqp4dhOAyM0hci8IPCF93AN4IJh1lm
W8GjD6/VaDsZafFNxWb8rHNNupI0IEvPkHl7OK+xXhYpm0yFw15pPFfJDWjqwsF1ih0AmUw5o1hn
xYj0dUJ18E9U1T/4t09F2+0Ue2ZGCAqDCxdwCbTomYdyCSkfa4sWyblW37RAOqrIIL4o3GPK4QVJ
EXlcrBoc64fQNiOCV1nlkbLtnn2GVFGWsSBzG7o9pSjjZyypIzzlcWfZ7q8u6QIOa4ZoW87Np6q0
enAgVnEcmu9tD07O6V7P7yyYU5UIfBIYzM3BeVOR465kLlhBnOT/5FqljzPu2CSiqGB0Bo3f9Yr0
1vccjspRD2F3ErPMK1erVdoo/c5NGlkhywY8gDXTkvgT+AVFiioRtfsfrIIe2FEqRVWHpuDN2xzT
OqydEf0ujYgq5hfPVSjI3yMtsax9Vlt+s4zwglP3i3HccRh8jEBqPtHvXTuUwnxrJ5TwCToFsw9X
m2NdlOG0fPc92DK7+KQ4DmBX3MgO3j0tns8c64nZtAWekD+Yxou4PO8Oep1z4q3zc4uzLuTheIKz
smEAt+knKhWfuPCHv2+rBfvwPWcQfndK5eECwkKlC6z6ORO0RvAu9Lsxyi6jzTRoKC+TPCFjRen5
v6Q7NI6Fulc7pVjpCYitvi+lNP64+FEFN2cLkGtqQZzKuo1r9o7FxfhGCSwn+/L10GJr3z2E62Ym
ywIBuuSRyIzBelO+2c64+uTNMal4Gm9vLjac0xZrKi36uUcBEX3ynz3dSWFqu8CupjKQcGas3eW0
7zyKccINRD/cZDqFwqm2s9FU2MJvxW9IAkMAJekqSdZom7Q5M+ptT7ky58MySA6w1HBLHgnyIREX
3yUtC42ozuA1osN6qUNU6TVTHppAXdf3BJwx3fOxieYlbb67rcB5Gagy1x7sMzAREboF0rjKRtvb
LjyQeISrn/fwpKEWztX+N9hTai9f+HqJvYZax9xlb8//LusO12haHuALPi49fLTyRUE5Q0nILXcb
M/70V7up3rHBTEBLVqNo9b1h0FrSzNTEIvVmQWAAYtbTGc0GCRLtzWHO776EmzrME1Xeuq35jnH2
vMD1zTSAaKLx60RSbKeGNc2RuHwC0Jhxj868n5LadERz5mHm5bzh1hidYyLmXAdJMWtQJuOOXOOv
525w4p18aWKTTwfPwOjS4CKBiKhqmh+d/RzhjvA+yntotCu8Pal7ij0tgZQxC3bGxy9/geGygBHr
z3EdXxJkVVZIFD6xDW2xNF7LJqnDmJzHiY+Lq/cJXOrBcg7lh04WQbjEpVm2MKHVrfOVx8WBF82x
RNK1ZpOyQW/m8/cxsFHstBrhdTjEM5lOdpSXKms6hu9sSFYEvuDWofaEZdHlMvqtcXQxiTbEc0Em
hJhH3J43Aw4EC97ZzctsFfB/yGSD6aCQD1fn5JaejF+r+sWxBKLUJ0ZiGBmdbo2e9gEH6ihXgxdT
Z5Yw16p+9QwC+mMTstHTrPIjJSRdnZ8i6MrWFsFNZlNV9EIS8SJnNigkOqkM3+UEoOBYTIdgvwvw
Gq5tYYz4IE6xstbQfCENpsgA6YRrXcRTcUnVwk9DjFNMGEZposA8yaA8L9nmtLhqB7lqUzAn/ujf
JeE3DODRDf+HJOmDiHVLy1m/AE+E8d3tRUvkrnM1bd5g3mr0jvdFjLJ6k9K5dginTdsjeIfu22bk
1StKKWzPzqN5UAskV7tZNIyhz3TwcGzEX0BCd8r6CBtTR2FWPffxMn0LGziYCpLCRtdXw4qFd9VT
qgNWTNmdaP76Mo+Wz1HvZJBcj39riGYWSQqTNQRQG7Ke7BKqJ0PHYTzBGt6ElTQ/NIKVY3YMkjbL
zErbuBKd20YPAGJd+qfUGE2LfCgZS0GPdsH7EJDChZoZioAEhhUHIvoAFT0AvviY81zaSdYIRSnM
bx+YopxDsRpsEJNfp5ppActWZolSL6twrltjowYlJVYjCHrbgtBtdIXJ45SeA0PN9Z4Gu8IL99gr
pcf43n8VfIKVRTXGzayiOnlzCTTLhdwGaSIM3jN7SCSNF+E+SVjS3+3aJyZXxVOUGRnRJJVkXLUK
YAzm5cNN5x86VGX6GJ4Izm0bp6qMnzzv/XPndQVVjtM3Vk0M1i6k9j8j5t/6QeP7RcMHqoPRcMSG
8hK0uyhyi9ynHONtXcr71rbD1y8AptTiVvYwDgtRCv1ebu48f2tfRBQiP2pL94wpWNcyyQqq6z8K
yX5Bcc514gtUv4qLpcXCHkGweW6/WyOO4CwvmPMXhTwy20o/JF9HDdk8SHKLVJW/Boz9dfUDDOdj
AA6iq9gJk+qMzlw4hMVgaaCFDPRhK4eL4XRdJE8r6kYQ+4VbF4pRC+k4oiv6taeTc7tJfSPvkuVc
wSo3NHU976+l1RUegJEtXar8BDFfaJkmmC/zmUy0fobK0Wrp4Xvo76luNkob3D7KEByZYKKusD79
N3Gn0ShDT6JHTl2qiyfTE52lP1edz8bbNDK+eBMym/f1W1cECIQNt5+hgzzRy3t8V6JOSFDbHsIQ
YVKS8mDmnitEQFe+m8j0pjZBOij3/8yDNntkrTNprHh60aGXs3Lzpnhjn5crbIX7JQmlCOtLqqEQ
AvPWjVAHAsNSMwtm8Ak53wY8eTjaT3aB068xcQsZrF9FRGBdL0u3Fw6UyIVejbgm5grsHKSyvLv5
uQHyd7tryR9ERmx0gvKQJHEMC31wMc/ugC+tEzkjWnRyksXPbt4s8afCEB0Tu9WlUcD+tHrh3p7V
83HckPJUetCnXJeiv3ifK0OzW32+mj9xGNT18A2rR873SDD2FPHtfmFwI7pj53gRl1+WB6JTreEQ
0jpgY7JlrHtaUiPib/62K880MWm58jXeqljIzradS1uqOnX9Hze5xGCz4mCdTzA3LaxjlQTHP2tw
HeAKgOO0wL1+85kh/nGUyASrZXZoVzUsu4fcY2BaOvDb8It7DtFTkZC3B9lV1avn4kktG0X1tmMa
yL7kgPOz98NW3cbY2MDZex2DU6Zf9DJ/8DtL0aUJdfb2Hy8+yBGch9HNlBfVHranISgW7PWrCt8Y
Ns/O1SXVnLWKyOpIZHC1P2qZzZ/imC8+XtNOMa6GpCELELf/ABSMB2GXJvXyQQcChvMexZhNx1t4
tcx6+ZQLs7bEbGdyaPLqhlp3XOEss8GEYMAXud8+t88mpkRUrm/lJDk7Z+w3IEfLdYYXW8gifdLf
o0Q6vIEOMDekoMwv4Zs1jrkl9CihOuSS9wCedJUodB7pKfiJ2DjMeq10Vrb59v8zMOlH1muNI860
Lf0JUkuPGLeBhdfSoYA3X6QgJ7YWOfXKDJy7b87EMImrEN/Aw79EWlyUoGXRPRW1jcoPoUpO/Mek
SYZKpGot1v7iMyN8X0ffKYTqv2A2wdgOB9jcHhPtfHEF1fw/aq9+W3JKoARsZH7NSNiH4TY1UNZD
BUGWzjP07naQ6DEq2MYEvI8MZBUtyTCutoF2hUnXe0KMlBUPEaZ7aQ91XS8VXmFLCc0mvXSPDqIt
TdhD2YwfSnXcdpWD2biF58X3MOSjZ0ksR4I3r/DEpDn96VGf2Dzn+kG6T4nVaX+RX2cSRsxgWnUG
RFtlvzz637VZHGOYqB7Vavis9uhlczLrMCm08H8ihP+zHoWGw3Rs7O+AeUWXQAEUVl3XWOarGQbU
lpl4FQnSDwOMi30r/WWy6fRLdNBmaixcysfE7ZJR9kDhAxZP9j/Mmbtj2Rk5uyLrzbM6dqDsbsJJ
cZnQvP+d+pzjbtaz+lm55/xcxkIKoPQEQZDePWmpZJ8npGAaLrVylWkLxh1mZ/4i1gxCo44FKuig
I0uD1ezuLIjRs4bGVuIb4GTWwNZlc0RxJRNr40FQX0kKXAMshAT687lEI4pvLp8DnoIbHnNr++mj
LdBkBfDmqyDoRiADNjh3FNSpZ2qWI6svB26OsLaM2m32lKfjLnDIhl9IaprujFihl8qMoLIqg1ea
ZLWXisWpfguLzs48/CuQ1P06Ppg/AABrM53jcSYrOi+R3ydWQQd/tZ0QFY9+baSt3Kaa4fh4CDOY
kCm0ntFUJNCYmYTK05LvNH4UyT8FNxF9Y3ldZZLmjVwpplIwtaS58lNpnFmSjX7K8B5NY6kKtvVP
JaySygSo8ZV4/knBVq60e+TxyTzXunE+29fujmZbNXjkoDMzFPKbvcHcnLBDh17p5nqjudSD8cKi
8Vwfhi9lonOuHgRVMzDaLEWrz7K2rRvCM2L9NMiDJvq4+jXm4Yzgh2pHaH7L45o+4Auak7ng5t1P
ha6rV4fXlrci80HcL9RElcJyfmtWTpN+wd043+07ZxW+hhhuC5F8vb+Rr3vlaC/Y67VUkIKAP1oA
MCuyni34GNPcshPEooiy+CqEwXmGoefbWgMNs/5TTx3GE01In3qY0ozBKQ0iauAFBJg130MheYrr
Kxzzt3agUAIk7zXVbmlWJ9oxtHGiMBzXixQrJ9rn4KFwGPOVoTx+JmelItkScH+oYie5WTQPkPvS
PDFxo4vnqI0YZCki6u9vPmSxnEH2aUuVtdg0AERWxlxSkqeYhOiCpqF6+jjy7/2OOlLIWA94eCWw
95zPOjf2WjSC/u/N/vZQMC1DwoIalsooDyKuDDhwHU90+AVzV9xlqlB3oCDVZMQICstZa2HaqSbx
Ljy10ru7PshFRztxvm460LDAcw+buPFz8PADo0Q/5ceYMO51BWOn0zDptypPkbwHhD4Dldpw01NG
5EOucY9c0O3IcHGZ2wi+Em3x22GmwOqyAnoyKSu/+XlOWQEeecgfjgZO0Yd/IDMjRWPmgIUsrtD1
bRn6JDAfgFRGuqy0YZDlfkgYtiywBhHq5maDcwCbjK0AgHNZbVZhKnfhC83toGh1CCdwoMpSpznO
PUx6VCeeBdWPVm0V666CGxpXkMInL4xFANjNBu21JYIzm6UliKRZH7IdUhE09Eo0wQVqphNLvgrh
jRY+h767HqIIU5akFUAqYuQNqzsUXQDj0ztdKF4hPbkPeQGHhYaZMaDaSDQiEJogrO4oPE6yLQWY
hrlpL4QoQtegv7OGui32PBslDBiy0wChbtrsduTwSncx2y9OhYSzqI2eRmUGHaFJSu8BiT8VHLHX
7FSStdWbmhs9x4HP9XPIHar9+tqqQUEMWSj6qLS3DeKbNPstNcxXz3h521E8ROXax565m3u0+baw
U9imLAundMeE9jBIyZJBioP+N3AvF/tscU1g0VSW4GHMo2H0swbk2vdLPd/VoI4GVnRyq9SFuaVo
JhfBzIYgCDKFsgIsunHhZADRdaEJobd4+4fsPkZ3ZOiuKVgUXVCNIAxR/edHbsoa4x6olShF9xdH
86DCOy4xAu+mq9UQZRIn0kjqcDp8htL9uD++jJp78VnPAbbZh1D4QeK5KwSeVaMJOOR2FNv4up9e
8WGTGJtANj+tFS92xJ7Meww3piiqHPHB9QckqGF8d6uku2PtJG5aMMSgryUeq02RO2ESIkXazv6G
XfYwk8Q2lb80vmFMpUOlBg1eKbruDjv8E4FSJBJa6eSH2iQ8gZ85zHGGE823HdSbkdsuVqtAAMCN
Th5Y4Ix37x9oaXOwj8jfGkeWJq69zfQsE0A45JisBF8ea2u+RmNQ01d4AM0LG6VNrXI4Bun9CNb8
kzJupiRUB6v13Gq1dx1mx/6AOfAyWUg/mXvLMqaDGkhb3G86P1WT7tBiNEVSD4HcO2rFOAoiA1z0
BIVFKXRDn/nrZ+QwacC6kzG3bz58tLhwEKeEoGeQ/I/M3upqgr31tEH/orOLohRYshuy9SQfpY2y
hq4oi9XlUJKIeelhnO/pAHI2SrJrvDEH2gzkAKABwcVLyZUfhLS/u0GArIwCF+J4Yw26pTmDRrJf
torA7+iVnLRO94T2nSOBWY2CBeDMaGODNpGnxR293NjFplO6RB6rCZfG5j56tEDxUDmk3wDxVN/+
M2tlTLj8GMKUjgWDOciKA5wlEPpu0uJGSjlRXwzXJkFLU3yFOomHBNoo1L2Kn+725hHVjVjDfbII
wYYfFFgy5S1ifSRc1a0O9KkotBK57hdJkJUlTCB8+XtmAwSBhQycPCUDVmkaF+nW16MaAYyZLQFX
XACFAyZdVHwXNtatR1uBU2t80WAQGhm8vlX8ZWNBzBe3NIvUSUBmzjzs45h7YD3TyPtVVPe0ex/4
+akVDu3gX7mcArk3dbjaUeF4S3MdiTd8giPUXlkY+Dj7aQC9SNkQRsRBZ3Y44K+yzgKDWc73Ele+
TR6PQ7YztuhpRTWOUKMBH6SOd+cjsGYMqqw3G0r5oo1B59yQUGTQDZMDFH9kJCrBSuk1xplqSfBu
oKf8ANOtQhCSlPVfx53Lhsd9mecvOfdLXyY1RJsO23TP3VT/6GgeA2rad6+bS4Vlo2nHUE3ppsnK
VxOmEA9GQIA+40k/C11cuqfhvwsUi2PLTauM2ozvd3PZ/gnZ79U0ZTRyUBtM3iIsSN6sBeHm3KVH
ldXEQIDCRA+LstoWRc3/DcFCN4VpyCM7ImxpGoiFZleX7BQ/YSqb4/Dn52lwU5jwNK1Ni5oJ8wKS
CdTsspJFS5/0Manf4wjwX8Wpw4/vw1njJ08ZOQBUbCEJbZPkAMd/uIJ8iFxAJeZWnCyDeEU6JDnf
HVvBliahbm67Qsmze/P0HSYzRWtA25ISgieltNoKdYB587k1/ZmsfVEUKVd+O5dIvNPLDhIFuVYZ
0wY6mFlWoK0ctftiBYGVgJeRVqG8NxxL61mHEIE38vuEK781YXb8fYmhgtsRPLW+LLP12vaF60YY
eFK6ht/zu9WIXxNKhErnCNhxs6qYwQM0oFLkVnfwpJY6O++9ZCDF5VFLTDt54JukeasjuXZD5+Zo
f4A7qYij2W80+Lj/O71X2WERQ9D2pYiAFPI9kBMwR6qQyzFjikzxWi9wW9h8ipJGymNJVoDwUJDv
cuwNX8gPt65c3Jpk4FPPBqQ+wDotE2lgI479jtNXBK9AaH9VGzxWeAwfOpQ9f3fxLLtZ77UBgCll
HtHSwSk/KN+JFqNDePzpJmlFe/UTV5CI9IAZOzM8tn/9ufjcvjxyX46EQSk0TIZbHMFwZMoTax6G
/iHfaH/d14YA2xHzotgHiLPx7j1AX8DIXj4uheRCSt9S9F/WruONVfxmbzGUSeTs3r3Vc8jkW3FS
QyIk4Y2MSa6F5S1PUTdF3UAPBxJQArDDsl7Ki0sYOVVGnGyg85oKYl5PT5cIvCk84n8gbHBzrl3I
cpEUMJPapdxw08JMzYYRydMMkLkq4+zlb+t0qLdFYlLFBV8Yf/9Qc6Etb22OQNFCCQgCXehqvsdK
JKSUr0FonPaGxBYDgur4LHUNr470uFnimoE5ZnO4yJLE1HjOgLDy9zWzR7qpxKBl6UWsrSXYQkne
nKV1MlGg2LgfhbjOcKImVpCd/3Md1DWqPPNdGSwLH8+cNgPjvhRa8vYV2HmLO5QcVjVXVJPILTiR
AVAvAJQ4t8DS/DikSEUosNYIr8a9UFdf79Mc0bwv3dVv4XIDh5dMQBoZq7Cxv4Tp3wclnGcSpO0f
vjBpkvN9XdU7GtRLZu0nHJxbMDuK9kg1bCtQDJ8qyowAFALbnqfbMl39BTWYLCu3WeE6BWN3jg9k
ONPnbQlAYBksZgzk93agyLvLe0/sPX+ig+2nrV8cwwAajzWA3SQUQe3krp9ZXPpcO9+h0AfrBXBe
cFTydN/3bH2S2GUn6N2VC0VM2aTpIpQFa9ao2xvN9tJldq5C/i1J3VVUXzQ61jZwh9ZmKEKoxKIg
MTsLUNMAh9sz6tEHUvCgzHq2NzRJmsze2ziw8KPVORUC2fUFZrPu0mtWC7yKbZWYLk9RgAxYWaC/
eC7OJrEH1LsvUdx7qrhq/dpErXzKG0YNiyAGVBcRwLENfz0+0PRbzvZprYlflp4oPhVbfen086Xl
ANIxcF55KO79JDV9P8ssHIypLJmW5E2j18yY/KRZgoGEdZaGvxekkiCVkVLJB8nodcWRxkj+3Yfs
PPbCpYsM6aBGZl62ZKDZPk6eNvW57tfG6xSBz6F7T9vnZFV2/F3w4UlS4b7K+G8A8kdBXtCcNiJZ
ClT9dnk7oX+8/Brkt517x9vvUriDCWCYTeIImLB0UMHi7lwWTpCb4q6UFPA+4scPEAJNwy06lpq7
h1qOO9rRoTPjnhe2XOMrIDtjM7abeHFUU39PjPqfqukNmHMbTd+Xj9sYvEhaDOg4tYp+DQv5NmcK
eVrq15L7H6tZ6SHz5aj1GpPxbI+P3JAf9VCaNW+eWhBPhb7k7T4bETtQsfKAZdKlvR88JFSyr5rf
UfXpTu55Ln5HwynoqniQ/UrGKXlYnnC8ipD3HTT+eohl6aI9eIs80tdJP5CDlyUBE+0sg+aYUC5h
v6DqNY5nEmEFsndOlmpBoV+8GrIT0TDPfCsmnVz0AeS/XzQBAOZa4TIatdAfy8FpR+wY19YL+dgY
B+IdoO7q8Uf8A6hA1lY5fhan8IkBZK9vJ3k3AlKxuSedKJkr0G64WL0WmRVrpmi4SyXqtgIcRTnm
zVsh5HOQdyONUrlPyH3/L+6Zr04bULP+5PdsZnoXvoIwCYyFVwgQKwYlPOmVTHbiBVvvsWqIiR5h
8jSyRxwqDY8xvBFw+EWhNEzqIkpwxajQB7gGBzHtdcP25cSw9+LjEs14Ck93TUbpOBrwOm4fLRQC
GlHsm3szGEWiBIYn5dowqx/GNcmQXN6P0X7hpxYJXaA1Q97XHgqxgmoCH5UWnL7s7X2DYIe5zeF2
F5TNk3XdlAK9kipd9J7+ynT5PDekpZvUS2rJOEDznjthEowHJqsIi7ffXjxjZ1WcJvomR3PsP1A6
GVnDWLM5/hgv1hMPg0Op02B+b9wjedTiPJX1Hn3FRoLt4TEWLi/56zGPCzikbrhjfGVoN506no2k
QyIEsgafssZTdcfvW3sb9BiaNOhz29Gzwwd2tyyvKINmgvYUwtgacsEUf/i97d1Kgruxx18gm544
onRdsF1WfBSpMiyWybqswR7wQ+rZCLNrD6G2Gqj8FYvXOxwgxRJUxt96j9yTtDgndWTNEmCw9blz
K3CptuyYODj2jPCUMiUBvQMnhLBHqpgGapMLXVXNIrcBSJGDZWANFWeH+sVe9f60m8BSrN464ihk
ZDuV+OSEL3dhLBNcbIoBVAcr8V12yIUc7A3kMZactip79E0VbMMbZ6hQktaMk7P+F8RfvObperAX
nBj0AueSuRR+tc06DQ7E5GbEb3ChaN/Pk9ciCEzzNju7eSp5kb8uuJbjFv0S8KiSfYiLEwm3iszg
UZxA6ie60g8ZIdeqyS7o0CCI/Upico9APatdVWPy658kbonO9lyqjo75z51MNYtfsoVK4w/O41fN
3pnHKIk/nr/H66U52zO2FeEhoh6JzeFIlaK4dCIOt/pP8Jc8f02W37EZv5hlsd2L/jcazWMQ5Y57
lQVr1+2KZCDymV1kL4D8Jr35bmKJIKg9W/xNUdLJE2Brqg/un4Wpmush+Wr4MWMirGWUntDRR1q5
YB2DZiKA6GiPf/Amk+kkoCXr9BYnYMU/XfY7EKf+p99vcVPWqxM1rzEe22XLhsR4YepO82ag8kun
aMv10YZWHdJIwROYNx+FkbhC2D9eM4NcjvIP41FspfHcALtRU7hLp9xQOp5eVTToMq5dbqRn4uBK
vcX41ju0x4JtUqDMdfPnrXlLPlT6Sd5btjZveIWpUrJeu21syM5hAndSuIKkao/qtVSszHYwmU/+
NXYf2KxV23FeiETO0qqH0c2tFfxTcfPn98cQTHjhj+1eYBvbm06nN0PM/1vX8z/GPF/DyYgVTXtP
tZka8mk2k4PfMd5Vpq19pS9PLpqB7PwYWzNIIHckE74W8DwWj+9keRLLavREfPFq7CUqq1FS7gkA
Onkx1AiZrOTJQSkGUSFfbfWKDhirrqOP08gMjaDenk0yEYBQvmjQ3ys/gePe3ekXbBJsYcpf4x0F
SdUzn6owsFsZEiF+yhP5vw2Dq2PLKi8YWse3dUrr2yq05PcMoQpbkxQiwaaVjFL6j09JdYedl43a
GQC9w1qtIVQ41HgxUt6Y6Er+q6ZmZmn5OEjp7Sv66JlgA4BxgkEMO0eTel0yts58SEcD9zXQ26a4
TCHMPLJYJZ/MIRuH9JxLf9VCqjegMflzwXgAMp9vNtxWKOoeHYgxgG7HJccFcAMt4bqQiqr8GY7A
bLT+Bajk5jv7/5sK9xNZ9h8WFvinwRJwBggANiPD2paoitvH53zUkyS61YOD7PGSnDqxYuApchuk
wuvKAFqf5JUyhqKwWGHHU179vp5dzigA50dS6M7FZ6zbmsb8oAEr4yYrJvgEBKEdDd1ISxotWaib
QI6aQ9zQ3HIkdXxX1Rbbgo15PEfmdFFONMQYrxLq2KwvpWf6tW6zDVPNnSTGZDrlFGHOJsxGE6Ug
B+BmNTk1K/KO5dKfw8DuXmcfW2dkITllOjVBSBjtEONd5BOMgO6IVcDpPR3lE+9pV3groDSgPq2r
Y/vJx8XDhq/PimYx5cr4IO7wNjBrQzMg1nevnNwIzrRk76PEju8yN5dXAQWC3OZJxvKt8SvzziJT
iOMgduGBruKgYRGu93o34AA6yxCmWAFGJZXSaN+Yqc1F1jc8RcdghELY4gDB2o9+AeND/lRZng39
FAYriziFmpAk7IzBTbKEtGOu4u/DT/re3ywO34UXTfnESXgyGYa73vLvrIWmppkqgrz7M/HBtylr
8AtFs8Jfti85RcfNeqG5wg1uJQ6VXu4kqJ0+e70LhAgNwgLXDVPEXgQVv6QFXseKbviqm9tlk9g/
2OWXG1uni/whlPtIP2RZxBCcoXcHx0xKWA5ftj1xc8b8u/VbS+RtA4P9EcQBcJZYvooebi0VkHqk
1GVHa4ZAK8qfWdEb2llks81OmVicNHCfENbnn3hbKj6yM8emsOEvFbrhPMntiW6jUY8QWWCeqEOw
0K6joi3SgI/4EfvJlY2CVe6f17T78ZQGZcLxA7zkZ457h+Pdsj1r/U3jMd9sPmE4Wo0+m0jNbMBu
YVy7wJcUdUAgualCm3Ian3+yv+ls909OXTV8y+dQ62Zja9Cr1jCghZsFyDLBT9UG44npquJVEd1C
+F4GGvIiH4UbX/TMQXXYLF6ksKHEpS9iWiahuI1rfmtXFh6sQtATixQwofdRfDlinmZoBqNrmeu/
oPqUxOwpa6BtS69ZGrDdHiVQjZm4dbP/LbSpGiQHFVyWgChsNQW8rdjOB2MQDemmsCLsUZ5drYLi
0hzUvtYyBq3hoRUm0D0QDeePGwDhLl0vcW9mnmemHYek9w7owEtH8cofQuFLHhTbKJJI1HT76Fbz
/wwQ0lnCd0pudQ95meO5ppDXmHli7mJ9FWPIsoCGjCM9DwrN1qfmPmAqbef4brYCLA7PTdETPw3q
zJJTmfcTwCdwA4M7qBQOGJ4sPvFmucmV3GvlOyYTO3irL9rhEjBlhZ8cMmMOByvQW/Wl/Yx2O9cp
+HAuwsLyHly9K6HPEeOK2XSCGdXNGbbkZRg+ltDOm/gO8mg8Anqql4nFU4GRjwzjuZNPkrJgVfw1
SbKP+euzVKP9zhOWeY8b9ssolRs5CGHJA4J6GE9N0a1htDt7rfqKom1VGOcJPsNPtE4xXuo3+8UC
fLiOyIGgSO8sFjvKLtCrHla5fMLrumn4nc1Z+6hoVUzFY2QDGQTtA7gKSLqrOHs/OdKAgnFaTCrv
SLLt6W6afpLEJyObKCec4qSjQB5/hj0/Wk62ISgTZIEnRRtrNvf50R2xepV0/l9DiGPtimnvXu0c
Ls3euxmcsblkbj9IWS7vVTh2EBvJmCziY5dlSEkpLM/RXmJQIIIhqglmtockytU2oKvN0W7hOzLW
DX3tX6+qvjogEi3aJPH+gG8GgotULOzrpUWkZUYxZDFzVBEM09Oag/UIrMu3gBtNd36UFQCiXP3B
awJr4IP0VqzvP3IYEK0FG01ff6jjkjGgGXtNS5zt1a20sZXOOWUv/KTSjK7dZEGC2LPh4JYyUyee
j+TdgjXQRNvBWjnZorHpgJP3aU6fntAXEKyNOuV6KhO1TiOhniLym1F2yWsoItoe7at6UQ+epwT2
z9lAJsxKuBjvxo2cPIuaCExscARfaSjGkTyspSRhOWiNAEc7/n1qNgU3oOY3oqwJK4BiI/OimOgl
Wx1dNUZIVDN6KfPXVnf6h1VIUQyaq1lmMe8qRguWMJur30nJqm6s4VksOk8JNYo0jqqk+SGFZ/pB
Db0rZ00tWJBATn6ynKkYNDEIHC4uTbmC3Wn5H5sqzWbwq3OXZkbIlA0xd6echRkvIZh+U+QPNWR5
MCjwrJYamYFJEliuCtOJllacRDhzbAhmHHhcVrkDxxV+rsb7XV32n3xIYIQ5KO5jsTeRgYRd+3uU
o6oIxaydYAdQAg3Rs2jvAklqYOb7SdIcQJ/xRyxMi9su5oTIrI6yDzkAgVOMtZQfZttUFpp3n3YS
wJidD9IqMFtG6MUUYwQC4LTTniCDZDuDuGK7xlBry2NtSD/PgnWJrLNmpTANbPc0yeeNmK4yoewi
jOpTCZPiIgrJiO2BFiZSQ1+fvOhjgMK0oUOHti/2xDzmNhDg8V3YvYtxuRYJAKKRTF2Hx8hB4gC+
5UCWLBkZUEu20huBgp/Jvem2GUijkzF9QwnNYC+HFoAa83lZhHfBF7Bm+TmCL2fxHEmLwKy2z6B2
OIWlGLx1wE9uZz9m3NrW5VkZu7D86/SmbKKIN+V5aYz0pfvLVhI0UyH5M+3oVOvHSmaK3EZEhCp5
tWCEDiH70GFAouYcOzimWXa8nb691IcInNoZmZv8RSGCzhlMcm7fD21ynqk8hDwflDvIowsCF1I6
JFR8Y5YqqLpjQBktogYg4YG4VQ/sCxe7dQni+lQMp9t6hwN+9XZS3jW4KB/iliMXX726cPLjfm9+
9YJnXBybkUdiF/olhcWv2UUK86wRFGTl9hGpBqa3hwNlNWPjrKYmaDY73Tbwm6iZXXZmxIwY8o7L
F6hKKGzkjvxBGPbx+JXAQt1lODXh0Z7xRmwjROqVF9x+m6xhMX6/ch+IfVVe7TBx9zTc/Sqc2lEx
C/tc0ATBMAqVBtLlYLqnzSQ6XYl2gYEJ0cPdLrL9kbVi4ILa8uAVy6wssPfkf1xRix2xUw5s+WHG
p8q50rBIAiR3GUVOQmXuL90r/8tk8CEmmKkdINtqogsUrBKiLnJIsiIRdQYc9RusNZ2fDI3lI3vb
nZDbqIKhWKZB3COBlERrfEfIYkty+1WO4mfxW77C/CWP6Zz5r7f/G33PPlFs8TM+Z/+BWScjbEXM
qgCVhBXoiWxG2Q3WStc24h5qtueoY6up1Bg3yRz4+Ga9QJRXN69+lJG7o9Gj3R5GJARqvXrotcsr
zP4tMZl8JNAkosuE2tSzKW5/WoyZDu3KWt3RqiRYAZde9AsYyONLKpvDnQYNsoGaf4BrHGgD75h1
OnzQlvrgu2T0oKuE5W8DfQ9z5IeaJXyaUvtsVXzRrIsNeFYnVXNhakGJsU/VcFS8gsAyJPYS/8o6
Es0XPCHge0Gf8Q+LiA1EOSA5czXW/bumYZsiI9OD9y89Kxp5Lj2NmQ/o7Kmb3ekNOicAogcx2/nO
FoqxWnoph+/rNQCDkpsRf82bv6fuXOkAutzAb2ZPiVs3PZzMhi0BTdWTULslmzDJw90u7Tw48Alm
cCgnjofPfCSXKb77DYkmJ1OPlBKOJR7q7gl+f8LUAR60UyoOmIiPzX/AlRSDC8FsejTYV/ZZJdzW
MKVaeri8PDG8vK7LAhyux0CWIESD/A8yzFaTX/Fa1H4FfEWCtM1t2sulrUuOY3JWNTXkn6jR0NU2
4K7xRMv5WtphGacV1i+dEhYQdNKpwJLY4zKb+N/P7I6bVqq+cPRFKxOFKobxDU3KUZOo6oFfQiqv
zT6813IqDuRVu1XdiUAZV/uNaEFZz1Z7Ec8nogHp2pMAnNeBdDnzm+vINI1zMcfTvvH4Pa41gk86
OdPWaJv18tP1bBA3ERYyH74AZ2wnAacbllVsdXFDA+PqP8PPoKqa9YBIGAMHhuSDDlPmVaTbyek5
Dp33WxVNkswx9P1kStL/Bg80sGPuJdUdAG8bLWKX/xHdB6RHvYGlx8rarQxpydiAwB9Zqd2U2Ffk
RAgEdO3z+CsXFpvnamj0WJU142C0FOkl/01o5zrP2upcWBDuSYKUPpJfuUWvkb3Gh4x46q8ksziP
EfVE9im+YwN9xE72JLbdEXCsP94y19R1m1X+jwQHvvJBZD1aWa8cX5xEpXc7xDVvvfCsdDe+pUB7
/MySqaAhvQRWgqSCRMhCwAunKINwSwDyiTtZRDS9lI7PvGJw2Jyhh7UqSVMzjVGOyooAlj795YdN
iK/0Af5b3AVPsH4SItXjxGTsoosKbdjsjj190bPDlwkdNB00Y8Ms+Ia8Ty2Dou6Ca5NxIgXmQF30
gN0pouoPCqYh1bvliA3GYGssPEBJXRP8pPFK4AqSq1og6PCFnVj2MuS6qoSj5WSrcHIdgYqdIrnq
DdqTxq7SutgmwFSxXAp+FjyJlN0jMgXxPc100vS9HvmC1OFCTyfwH2/9R7I5OrJEuIWlK+uVt/p+
EGO5l/g0Pk3N52m+OEyX2Ex7ZbApilakwR//Jl7S95GVyYRHZKKFeGeVYZ9bqCcKNBhvYT4hunkC
AIdVp/4/hjcEUVzQVDM2r/Ymmk7AUFp/tONIydfkAGWgiINuGVFuuGPikL/+v1GLaQsDx6QsRcXG
g4B/fivr5H8UCG6tmVjIXLk+HePq/ZCGj9AwD2ZNZox1YWGVS6GJkdRNe51zGZjpun49PoDcxkpG
iXPY9EAE2v3vw7vP5bEvauBvzfU97WIuncjYt0ZhH9CnlUran2/Tfx0yXlnfK/0phsCab0M7mH9y
SPGFCuWpzNCTgAm6DH4Qzq8evvIRK74j2JT+zeQErdUPfpqdDEVh1TqlOy+DsbeEhPHDgTdHwUYA
4AJyvhOpIzcOHa7vecL68nRxo+NNMLwicrebzgvDTLsqO0t1/NWQoR9VV2hL8TlrQu4OssH9mhNs
5Dh4rsnvbIxYcjV1Zfw0cGiZpp1jSlh3OTlIul8fdyZCYP7JPiGuohj7jUD6n6lhfWiPM6o6YAi2
61am03WPrWga9tksg/wgFaDRQ0hjhD69CafkDcrmJ9+Ci9EFpwVGJh0wvIJ21pS4oZL72IpakteX
xgPHgmvhN9GfCTK5EtviaVQ78QQ+6vQWLMZETCImR1AZYFgiRJrYBgxlIftMypDKWpZEUsaKyQi5
FSTFHy0/s1z5NSNvRVdA/8MzScDrwSYgek6c7G2j00dc9vTt3IjkFUFxw/TyB+qXgQVUE2jycjF1
cH6VPAh/bzQJYOyyAYclCKMZrBut6IFgGLOSsU72gz6FMKc8a4ZOhiHYeuHAntBkzMZ48E796eWb
CEMD8AxX2rjeYLaG1Iu5En4ifhhG0554oGkEkXPZlApyTvXGYhhEKpJ1sz+e7o5hLJwSfNMIhLih
6tD0J5tgFKVjKiVgBZbokRVdEPZT6vyGMK+Ql9jL3ZDRUMQ17dfmE1UiCCP4gluZDHxDNKyYFqNt
vZdPda8kjsdWDO4F9xpciJZI+0cXbirEJMHtQSbjNuvb/9strA9F3a2ogunLmWrZxvqJH71Yw1PE
wrcuRpGsCP9GpK0tMYomFA9/XELqxluxj4ltMaN8jRJAk03fxRqwAreWEX/OvUgnLd0qDvrnY7XQ
NaxZZOwbHd3c2Zbn65fQfFQnk3Y0lZgFpYpycsSze+vmJnSuGs9fseLcmitlNO/ph/6EZTCnBV6Y
L9F83doaApvoeFxPzGsSJxh+TbGuQjp+H/b2ZqeTs/E7jyLGqWHmi/f9IjvFHZk4imu/IFFyY3AA
jAJsa+2p5a1Rq8DVQh3AtFDbwXDbwwUyIfEP7+jfxh522HxcIlbZSPv2rw/gVJxKMbB9aTrfTHuV
TmoQ/lT0GW7voRWPotQEEeUGIqBxWw+95VGDTBfdPcYDSpo8lJzDxouwQHTPNBZAeqARF3gjO20J
+Y+uhMmq8Lg1N6DskGrWzlQXpj1RbDm77wT8PRxmw4F9CKkuEjPWPhPR/r9816Z1+JDLi2v6YdYF
VX3EVbuRpx0v0jzI8oOnfw2Wi5/LYF/C3VWJYls8kI+ofnFloPUwGwj05eWtGMFzaeqEN25a1GyV
lut9LhBib/ftR2hH26FhGcn6pcMhUoJOnFXM93GC3jpi9Hk3HWpCKAInz74LwVJAft9Qfhrdcs3Q
XeWkjORYH+dMsXW6JYFbQBt9OS1c/31b9gQVPKBLIVxBpFfUHIhhfRbWiS5eCfGc4uDZPAq2NvWB
FVnNqJfGTGqnd3EPn176YzXfARrLeZwWDO6mgaJtdKoPfh2vEy2y/d9R4CWk8Jc9iKwn9kKoMnDG
Z6M+t+L/+dKLiO8kZULJIB1nT49DMisz+7HcWi+DOivK7zHgx7BqMCXcRhVi3v0VsJ6YmAzclmGp
aiFecCazQpSE0gAv7ngd9sYO1/+3V1wRiiDUxdONoY2mIhc16H/mJ1beNpXTF/iP0AA36rr2vZTS
v2gDKzmvfjD3dhySLPd/etFylnuzbLcfZ049E3ylsC/QJ2RtVPnuIeg3WIDC/of57x3G5N8Yo6hg
zMifz+n8iNdTN+RuJMp4MhupTpR8c6JxTfVCPomXgWWIt3cjhvffsx8fMZsH5jDENUnqLvnrYe9w
Y4i3YNUPU9I8aD4mnv6MLsUC1lTJ7jNNl9nDFhJOvxHZYRDXOzx3kEsdXOEFjTHkpn6iDdXdYtpm
nXrLYwJUwSRAGkFxcPKClXC5Sq7WW10O8LrUu3uVKDtfW6mVNQ+fndMyRoKI+ePQKfhQjS7L/kuG
s7GoYVDEeNYwx2XLxtbk3D4OMGpwi0uRjZxyABNRk7MDZMjrSQue9JggCJx5fwKr3S84T6RDazHW
C2BflvGIYvSiCTs00VkNtCH9B+T108d6eNUcENGcJBQmDcbMBv6hsKM24eVJPxYR8I13vN0lpZJC
VtwIZTkbSvOjFnbru+9+tDRC/5Zv5RONXBuFGQmMx5z/n9CTUpZa7gmqNyqWesrLkSJD0zpEIAQF
NvoHXfm/C1gQ4hyPeOyEUZ3IZx3A61UV/wtpG2ay+BaNQe8igJgC161zfd6Z3zTJJNT2kMue6iiH
4U+K/cPffJqA6R3n5Ae6aC7tp+aBFoDzwIVZI3YmulfN+KVGpmimLbirVeVj4pv4DGC0MgnzJCJd
KeqoM8BGWIk6SUJAUqYLOlVIL0n4S74yPLH2HSOav8FrWox3frWNULE5ZPuAgUagYcMuHVmpF7cN
YU/l9cBKYzEGLFP+hFSdRz+9BHqFzno9PRAsNsMT9m2XHHTY93bDoUlRLOjNsK3gayYf0sUAKxN+
SUHDElPkjGVdeEsYa7Hhy2A7aMx4eX2CnQDqZtB9uNFRCOkF7PVefRBpeTz5AECIYsAlYwk0WeGi
PWzoxcevhNWVns3Fy98nf4vx5Ke35KJnt7/sOVhXzW9MfOkhGUh5K1kAwQ5kCgFhzEb/1iVOmfF+
Dpt2+9mteuQFNGCzDWRXyY/KAGcmblXLk8Wgq3QVG79zbf7Ve1hR0fgEdpaZKYrDoGUKIZFGZdZV
q+OFVWah1TYhxg9bIDakkH6L5tgFZiBHbXlur5kKFkMokYhblACb2r/M7qkjnqnCm9dUoemep2kW
jwSH7V3Eem/if3Nib/mMyXDGFT/rVwGmxlPHY5stJoesx9+Z+uvNbJSqiv/nnG8rWTYNNppnKmuA
jYhecd/VtoGi6jHM90Eo/WskfaGRNpZDpJYDe8ZvDGoB2rCja17e7RT4GB3SBeoOoP0Ky9LbvpBI
asalhWUxToOpM+L2ea7ywkldTN7UrIh0eUNH0pP0+NXlXxDybyqj6wt16WjvASLhMqiL7lLd3HMz
Xt2y1lsK9ciD7AHKDKdAy5gt+T1GQAqVH9UA9zMlsR5cxVV2rslWGUNOB9Ekm0Vj28uYHfcGDl1i
Tr0G65difS4vVjuwmk+iCS/KDQ7phB9WHALhQs/vFMktcX2UXqYOa5A0XhjNJY8pKoPy4HaniZH7
Ki0fQxz9qmWnORLH1Ytv0549VoIKKCUWYtjBpZggVF1otOlAXBYjqi/XypQ6V4OoEVfpCMVxnjPW
dKoogHHR5kjVPfzXW/hgyGnOqSbkBsBAEJl5G8/K1JrRl3HWbUY81Rboc9ihTCauDX5DhNYlQi00
oN/Clu8xXdr7TD5M9PsNdM+xqOnkzUXa7qVJRQOrCQO1UAK8vOVE0luQ1qjYMp2LTqsSU/MixwVy
APjmpb/wRbG8nqkyhBXHrq/11FEv5opo7Db07B7d20DPAyVKcIugv94kiXDEOvyLwPYo+vigtgvU
2umVwaXSWjw34VQVwRvzDAMrYhpX8BRsg8XRIs50u15DF5ELZWr9Alq1wVvwECFH0QNUf+mNARqQ
gDZ8diAbkg6fZ0Us04fc5/gAasx9kLI78pNoZCeP37WQPFUhv/3G7VQNxuohuiEVzpPMygL8ybNf
7MvzU0nOCk4FNFR5U6Yq+AqWxcNwijIZNxFLpYU2/Frneajv1NdYEuH/+m/yVHNVaF7slI7uIIZS
J/HDzaN4Y7U9Cev6Wk0yB7xtmbCoYxw/2XiNCuk+e9Y6+g7XA7+vAs8vkEHPYhe57AiTfwW0bzuI
jmU0LIoJ4VfvSpfFa2RZ4zN/LK17q5jji5J1hzd8rurur414UKvO1DJ+hYAlYO1xrGIiCqQsInI5
9gRShWUh1GdLvgb51KU5ihcUAYpPMfGkYQfIgOVzxis/uQTKaECs7q7FUaDqCx0YtHWmbThGl3Wf
fzxHD4pUXiai4yqsm56MSEwaPBuBoE0HHwB7Z+um50haPZqYocxN+Hi2obXOf35z9/LxVU1cKGfP
p9rOkKsf2uQD0A15gcVtCidpzGAm9uxI/znUwyPdsfQTs92iMLTcPccgCVEiV9+VnHYmqxa2Scbb
QCLZkUpyq/rHxc9a9Gr1Y3lEOQU5K3N5u0+AbcokoD5lQ6LZ2qYHI40hN6mVyIZ+UKLH0rXbXxFf
InxEp/YmeY7HJPVLq6lTk9+R0GlDlqkfXPgHGST1TDF/dzqAAoLpMKGJp6vqXEggoIoTlQwYKsRq
tIQGjwxBMQFLrUT6vDG3hbXmbjjpTeAGy2sFsrrpS8Ehv3oBQ8WjBwPvwUNmimAySz7gfCvzh7Pk
6t3oQ5/A24j4Qz1u2O3iw00dArCxogmv5bDVIdWBqd1HAcp5fkLiNt8Qh58Tuhcw8iUjm8mume0g
L/cCLFYXen0TGRqsN1QV5r2ejbq2REk/NJgODyesVpQCYGgFbKzTFqmW9AAZamo3+ui2R/wfSvS4
vGjh07qlYST7Pv3/3W18vAxQkdoJZnPWPa/qEwSYZe9sgxpBmmOT9SO+oL8atTSHok5HY/sa9edA
cscsGms4Bc+a9SFn2o3gl5oVHl0eHYAZKIHkS0vciSHGo85oJZGa/Iz86BfJCOzH3Dd/62uDzRVn
c6w6HUTrLVnnqGrNVU1O5ny7qZrjtQl1nW/vaeC8rtYIruadi+7TSN0o+QGPG3lN8Eu71NGGQmZQ
x2kzEdjmE5bC8ebdqxsQdWc1tag0y3wKqEyooIe3EtAjQzV2MFbsam8tzn1/EnKdJ3c1cYCL7f9X
W4Ci8CmGrFGVzxuXJL2y4SxzNCvdQclRAY4rkErWTXkfc4EOYRMmZYGPFAoCmGCfNw8Yq2QYfSWE
iKgnyQLMfgduG2NruNYO8dr8c/ufi8GSVCDXJQpSTlfqoc5QGYnHvtfRXFOmQvtTngL85wudUAf4
PSIbRaj4Rzx43o2Emi57pmYZgPYD2vDtWwRnWrKpLAS/MpxDULP4IMraw6bpocOABzZiyQoXjQGL
XZeD8CSF4fLKzYw+JNNkcegNB4m/INNS+oppzXZRSShJQ8tCgcS+8U3BrGgfICWCDbuqroDq5MVG
I9/IEIxKJXGbtXUbZfx1phG/t4w6dR98yWeTS7ikRr68JUyDX+IoZg6FaLo50ciimK0b7FWXBCzM
AAy4sxpKi7CYVi8QhTuAUiaGQuHO/liRdPCV4Gx88Cl8PdQfMw/eV3HiDy9sQaq5aVeyLfr7i/GT
pbSr97XG2sZWErQ9JCmpui+9+BroirXWZkGy56Wdeq9RPSXbdv7q9/U2tZdy4BLfzRLJHEonOZYN
Pw/i5PEjNHfdoeFoRjnnlv5Dhu302ictxbhZBuP6awf+C34Bs/I5/n16FWU7vuXZhy2FE6dryhG6
d9nHOzkEqohAg7e0WgiV5zLTDlmWWwYFMNxJBn26oH8P7HNUAGboWDmsQXvrgzD1zWg+aeG8Dfee
8tjR/Wl5JO9K3n0HZ5wCiDFtmFSntmLechxl+YiEiOS6aPLNguUSg+cte7+0j2uMj+mJhKAzqSdN
MG5R95MDzOMCVsZt2XAK8uVeItanYDifiG1jIQv3sIGsZeh6A3tt65GsdjRBnu6Qg8LEy2BPWhYY
k/+rlvFNTFXk8nLMV2lmyw3Q/W22b1lddL0jn5IZHZZKclP/IOW3mG2vjBCDK3XuOPkSBUFhZDOs
Id0EVW9a/Jg4rT71sMoLrB7SDTdVrTUJAZUQ9E9wxF4iJrEsLRGN6U4jEg07TvYhur+LsyyHW/HN
1xpask4ifFlRD/N0pD/dxIT7uww54iD53M8IQR5IMCsOmOd4/tQBkmnRZ7V/t+OGEqVhQH4Bo0Y/
PxL7H8MTX5vhfdK+0c8+VtasvqZFQmJ6zdZgxEk1z8EVc5I1sL8fF5msh0N64r7bLr8tTjCNnwR2
WYRmNTOx8HZpb7DbYXegCmgZz2bL+sa2kjmWnzj4J97BitH+K3oNHmLumkT9DdL1ab0URHXy88ji
+Wcid753X32URKKZ2LdTJdVhlovNl1On6uGol3RgvUUx/3bt2yEzSnLu3uS/FlxhAB9IWDZk7tC4
TuwjN6MupxsuaB68TUU90IkFBYEUYx48BP+NVboFiS+d7Z7OvM0E1UdVWXJ73xi7K4hUCGT/paKe
GY+eSwf9mo6UgDrzHhXExF96ALxndg5YfUf1tAY/FDJ1+kPte9MkfhM7/vkcCHLjNFNZtv24ZuUT
/Vn7tCjI/wK2sl0dkNcJyls+FoquyrqNElbpk/n0f1kg+4pudWBEpMukdxDPJxlKmkhFEMq1ArZe
uNI1pkLPGpPVNVU3u/22A73ZU/dQaRFGyJ/Zx3HBHrfFWMSumO6kwqOMl5T/o7FytVZeOnP8envx
2fYP4Y5KE2mbHAGSUhZoZ56kXKbHJIyR151/63RmN4bee6baxR1dF3qSupareLbDEVELAhcLxgHJ
5TplFniLz/s7N6OTNWM+A3InfVtvicNURglHfarZnRZpFWf7TkrOLvh6GA04meoRTAuV9YoJYmJJ
fQb4S5ltS9X5zRa5wqPnHUFN6IsfZ8EezMzlOsNlxlPR6aJH3d0MD1AINWECMAWRtYC+hC/gnwmI
s0lxV7aRrZZsfYCNbIzhoEod/ovK2cbywaIPizJHNLKcW2HK+xipYLgF97z+BQ40fs6ABq66hWek
t5aI0r2//fa9+bFeEK9wks/Ev094WW+lGzxWOQV9YPpuigMg3sOVIbFXlH1+QHZsagqyn+MZu0zA
OksXv7iHMsgCe5rEnFZUwtD/dLsdZ2/n8T0cPwHUbtVgLK2V1UjnjwadVAfzZeYJHCEhoOxsxU/4
bloL7ONPdzhrdSNFlECnHbjYI/WRycN5JfxalCU8f/Fa3SSDO12vvqYEvnAkqHgvCF5G/2A7cMGL
JEEXu/cuiQthNAGi/uywcMHSoHcCra5fMbCd7HRwrc2UFy4imI7kYs9UEy6Yj7K6VQDeyaVgvE2U
KBdPx5+9T1+BNASvpJnIZIEDy40wHrd7bJLcrdyFIbNJooLQGeHair6cECXkG0f6Qw0lj4L4rJRF
f5ul44T0f39qs6zfDSF2vsLY/SbKrHGiHlvdKP7flE/JXfw/xiOiBNgBuNQlyuZF9aGD6z3WcnRF
KBicHyjgXqTLHHrTvYBwA9HG465tYw8kVz8epgaPfFJDfxlsEgEsM34e/7488H/mZqc9+b9Sn7sr
j1P9m6R/O7YOkjArSckah1GcGHcsvrgzcq1rbfjrpr18Y9FRAWSmf+tQoETZtSuw9QG3hXSkwhr2
qaqI2+z3RGjksa9Wk4PV6eJv4oVUUX7r9wy1SZM6O7p8WItNgjlS4n3dVk/ndvIY129pA2vXJJpd
TBvHqylcD1vhH752jNNn+gh3QSq96YLJ+ptoLHQUSaxgvL98Ep15dEoCN833FAf8sJFo3spJnZFl
Y7wyvgWBVjwQa89jGcxgiSeWiV5d6dukYip2eUogTzZ9gnELGyQO5AfRe5Czzai3utFfr33wnwQ0
XLXDCIZnstOq9EJbpa856Iw+IsDh+MZARzFA7Cvkmsemk4wFz5prUCOojPkbwu4Yj9oS9njM013h
yrzfscDGXno2R477EJrikHoEb3FdhhlIAZY5xkqe9ee2rg29gdsum7bmRpZac5ugdiY08Mx4ikhZ
NL2J6MPdouKD4nv2Pjv0CdJenPEJ7YBaq3FL/fwufC0mFOqchouZpDDrf9abbuyVlchMNuwRW6eN
JjBG6ruG1PkPfOzZoPjGCVKch01b5BxRazd093DcmZywdBZOcIIkfwMBOHeGgbGFzhwnkKVPn6vT
cVImiKt+QWGpRw6o8yKTjAO6kNJdUqQb0MajupgPHMg1Q3P+YzPzvpI/5cj/RJ58HVbvcsePjWKW
HPan1VR/n8vWhbVvdoOt4tCzx3AXXi+h0YZT+2ptYyf8FZ2TEgQen25mhgvlLMI6HnCNdB566QQW
ZHxUld+z8/6XOcG7CCA10W96AweNSznrZGNtcs/J3rrt/LAJJpF26FfF8R77dnm3RVLZbigNky46
AaoWs0v+1XFzSyePVe3l7f3z1sPl33mhp826878dFFxJKaW32MGqUkpmDwWeHZ9kjkLXXGEePhct
1jzOkGYFiyo6rvK+49IynwFQOQ24LPMfY2te6ExKaaIlJUEYX3BEWP7ZhIt2G7IiS98oC2/LZEup
Q7B4KfQS2lIskIR40OZa62oZglBnUKy3Oiw5iJ8aKFJ/3F5GgJVnWP5lclMQW1Hzk+BX00lG/j46
JNRzxCZDkM5oBTJbx4jS5KUtvJz/00v43G1kEEtc0/ogOoJnjbqH8FBoVbVJUKAQR1Br50CRbc0R
5s0wsKzNvEpOjVPrOymU5H7nOgcRuEBurtjiJACpnFg+f0USSyEXQO10Mr2Pcq49c1dgNZfDgW3W
6wVtm/t6WMjTZVFW2oSNjkcImIJsX+yD/CdSZf2hufW7ClwGoo+x/G9nzn4Vcv2Z6TXhCfowNG9U
ZMBB2LuWHvt4WRH3R61ngiSGXpJ3EWoFj8l6gCJhBu9jK5rQjSOBlYlcjGDfrfjsyzO24TiF4N5g
8JXP5g1ywZa3llyrruCONHrPu0I0S0/pkRhvVF0ohpTFDtUBwxBiKuiH/zx4xIiLT63HukZZA48B
aJLN66i2t3Hd3H+V8IpDZQVYiorVEzB6MdmnwwM1Oh/xgeVTsxDcD/GbsAhgCtK9bzhSPS55q8vB
bqf4a6MQuJ4YK5FMJjlfIj1nbc7ARvkqb2NL/nFBPboSSX2Vu/UVJ57SU2qakqxJM3qjiLswJQDo
ho94YhXPqbcyfz6d3jpuubVafvGYu1X5/dBjWZep+csUujI2psty71NzXG3jAJsim0qLId4MQ3VD
mhfLKpmfh4YrUsg+AxXNZB8TICttDuyVz3bdhymy5uyrCIRlVyTNPuf+aZ4R/jKbYK9lOgyuiYM1
fzyEZ4Z0S5q4DOGARNJlcQOZQ1SZe6cx3/A7Xme2P6gjOFSeDDdiIpGw5YyII/eXDSNOTmf6d+qx
7nrt3oqeFiq2J5KjVbmi0nYkgKNp0Gdd3E9Xn0S6Bt31QJ4j9Tm6dDKpFEFZetbqZqRw+SfK9Xnu
KgXCQnbqwnLYmALWE6WGXFp1VxSI2nzQBxNnDethoEDism7xQmqqpqXW7ePQfEz5VfKrDLw96s8r
+iHxS3ubNAYPN0iLHIx0OrMzdoiiHwKtL4slZeWByBBIm3v1+6M2g8rodr3GS/V4DRR5orpAPcej
MaSyGeQdTPEbTfqSDYPUDc0rwZHZYx859TbPDLkgyRJhgjAYmtUZkrMs9TvI+3ooumGC4RV7FDCd
gMyCBZapjooz9i0baIf6qUyCgqxaooRcMDf9raOoqhSnwlY50D/dPQKHSlAMwG265kxjYV4I5dO1
nEhV2a613NhdYnzavGuJNsPdx5xeDucfkHaG/MSfikhEJQVXEMa9rHoA6BqYAcN4IAu9ipjnCl2e
aMTQo6x7TDg2pxd5UKYVtYB0f1LIWO5cUP/7OgYwzp22LG834FQVXcvVAEBUJUbbnykGd8BC1v4y
qBHIQ+sc5obKga+sJZ7V0dkjXha8RR4eZRZnFT7AH5XRCr0J5Avf7RgR7rq/71KH0SKQyoEJ1gni
E8XURvAWoHqP78xYbyO3Tlv8RyZqmm0ld2D2S7W0okSM4JQAZbdHJW00guQsPw6ji1v7xoRAnA53
hbwXVeELUt06XzfvHdK+2D82uB6SPZm8suzshftX0r7x6zx8SiXWjKYZhC7Jvvx0vibg/Qs4+IoE
1Xwp7N3vFBUt/96qkfL4RkB1Hw7Lg/w2PvKkive0fFltFu4kYbvzkT65Wtj+bLPTuqTmJQhJHbGb
qFvtR09/5nQ/vx8VEkGuwCOp9CckF+Q66qY1lz08TPMt+X7+tUbhVrw0LaeyPfTEyWOawFnCFUH5
FJLkSq+LVZK10y5nb93AScCrV5o3Z1uDqCY7Vs/euwWCnFaW6fdC8CDAyrKwp0UmJB6oFnykqwg6
oJR7QhPjF+7YEOTEgipT8DPi71x+gQ9GGj43TqLZl3jBf4k0fHGh9r6lsE0VPdq6Wz1P+15EunXV
QGmq72UqjGmH2tvQdOajA79v2JTwx9Y6VDsBjndx6M+C6IbWTi/W4H5mXfWSMUO7S2r4u00s9nO6
WWpdadDXWUyCPc/1dFtINzHWm2b7Ctqm92ub/1JFcxwMrvaicYXHxSiqrkMMarPjBIFXfRXkRRhy
06749ynbpM82S+dqkHBD2XXLTg285VXUPxJLDYZb0arFltKS2HKcZKDmiDMvghKiuMvPhoSDZcaq
ILQpZ1Q3gp/Ixh+pCyraKtAOXwz6tnH3DoqoQUkjt+WDZTaOmQR4S51a6K2SE6byvbcdFa0qX3AA
QgQ761ym6uNZa2FyBA98Gdq7OyvpsbAH8YgJ2RFAbM7D/5bBOs0lEb63AeK57wYUDZe6dDJrh5XH
Fe39qsXt3G0DJiKL2QP9IiR1iFJHR7mJHylXngIyVCRIiMIomEgwh/2ZDE6MGJ9BcAu2l9GGMAia
hEUG0dsJnqONcHieLB0dSc775dpJzC5Bl6ddHgpel/dYvyGT+bB41jgr6lBZCEH40K2gGsptymgl
JxKYGlw2FFrWKRyqzQpR7Utt6NjW+e66gmm9l7KI1+TKygr4Yoq6FQj+FMXBjCXSDWr2Xh4QWPcO
IJb3idcj+LCTrNc02S9J8JKDK40W3hnu/aFJwRR9Ald2j9LSvlDJu9nEnzIqeO26QHUuKn1EDjrV
+krqjSfjsDZv8Ko+0l0mE19UOnuwL/Vv7mYm2tKjr1rZy+j+HqI397NfiL6L26ZdluIcUJmLhcXa
r49KijcdH7d7eFZVAWvCrwtPxoKD86ydp4Goayiefy01WBVOoanT3xn+EcPpmrsY71+P8bjvLM04
UADEsTybwvX9b5E2yMTKhkZW1clEtL9yJkGbZybMyHY5WALfp2gLOqTxyxAzxZkgEzSQO7TAUvgN
SjEcHwFioVPZaXSFKmoUmW2MNwTX2RzwQIISrafpLBLlYdlcHQ9Y4zdYy4QMQVEprqBhAm2KGMVy
G9NY2eEczsLfFun12CTUXQ1hnVSJDYnYNwr/C5UP6ShBPc643COYWhkYbbSIswtF4o3Q6utXDo9t
oJjt66h+ehO3nX2/TwFU2MtZP+zTWSgE93spnWxydh6vOfC34Q5GBgxqW3CMU0WFIb7+waoPn1YV
hUq7KmVvc6LxG27zWJ3JaSaHTXGQaZ7lT5kA1gYlFSFEd7Hj3/J/JPODgsLFNinIYsy96DM73GHI
Odt1xlZVoWcaAL+jBoVaiGmGHs4NanUzrD/WkUlAcsDlmwe+WsJGHXmdtVRYh8T4GVYr1Qf/xHN7
oydDr41N6qG/h/K4/bMiLf/3Z4y8to5Pu6O1hvxCJRQtsK16GSsxdR8oT15zzmRxZ0VELjrQqnKO
C6YZF8HzFVNrOus1g4squfTy8Anh14EO2kZGu3JZtC1UOXNzIY36iuSvTMiNZI5r2m9Ob+9YHPoi
p0q+jS5cKnJoW7t8SNYBki/NsUVca9DYVYiP+FfeEWS7BpXgyq3V6QxaoecwfnWH1fuwlqz7idDC
ZndcZ2C4Y0t6X8bDaS+n2+eaHLzsJlzKNQ7WU/atBTg8gz1vNSvq+6fLFv0SpTcUxcNhEtLLqwXh
mb6fqgzvfyKCu7FIuVmFbBChNrZmzi+Ch7f/LHMp/yikva6J6pnye6T2f7UfNNRU1HRd8hIEDwq3
+rwMV6Vb7D69gpB4EjqsyBmPyjn0nicR1yMFMgwrJhGxsE54ovoYRX9FonxpWSHomkbaIK5gy7Ds
t9EDeKj5ZA+QUUAylCU25qBOKAELns9qsp6CKuf53d5QBk17WecSvgySG9R7fQ3cQRhUlHB0oMQl
1RfhbBdvPZkJF0mAbXG6g04U6MEQ7tve/ciGs8mRXyZWKQrQNKP/1aF7dBIqKka6MLGEMNKc/oyp
Iskvhpgrwa8uo/VbpKvhhII9KC8E5NdO7OEW8toRG+jN967LTv8u2Zfd+3nlFTqg/TJnRqnCsK0u
smMT4BFLBFxzc/vAUXm1rX5hvBvIWSQYH2fSogDVA1U2FkP8nArkGE0P470R+jRq2/k2tX7tXMkQ
lQV4FXMu6zD5yK+Au1t+ZFqtxiIEieTlETt0qQG6maSfiYqnr1dVjI8nM7p0Thh2/YB95MPGFgnN
qtU4eQdBJbRV8E4Cr/6awRcaugya0m5llM+YBlavnoDujFRbQW3Jc2IzeVUlU+j/557wDBoXi2DK
ZL5df65AqXpK5GosK43+DEzsAzX5rEgAifIEwVXHhYtAegibPtPUO74LST2PhAtOC2JnLp/MSM3u
tMe0pbJ2E18a7mSWNPd6d71jPkAdAcm7N9ioPmySbSxqJbeC8Eblu0CZa93d3PlFSS6VC/Rq2m4k
4msy4dPMReyhoPSp2v+/u+7aORSCd1vKKRaB0GEuQnfbNitctNJu5VqBomeK0Xcvyrdlc9qCd97q
4EhiK2vk2lwOASsmt2BbJiiE6TeBwUqWimBwaQtc/MCMtQ/SvzZp1JgaQERj7Nq2Y4Ebhp4kAe0f
6nbC4HjAo1CMonTXaxN0KiJ0UaUsJdKyadQC2gd2916EkZi1g20LJQBmVOBGLaVp9zesKx95Vf5K
qrqYRRh0Kh5NQ+oRB2txx4NZlQ3Or5Yj5fzhTWp/e7UKIRtIMqdt/bkLRWCfrlMaLsmkX4Igg5yH
PDKPOx9yz0n0vPovmEuvQs0uD8gFTdG89+Fn6hYKxE+n9VzGSjFs+juwx4iG0qu6u74lHuKTs3nb
zOGXQXMPW9F2vTVKhQhs10IzGzXlZOiC62rbGqVRy2AXsDb44/lFljZRynug1SVk4pohEd/ppgv7
Zt5o6arN2JqkHTJGg3+MvWF2HDCrdIABTg9g8uEoGDYhkTR/lVK0EcEp2Negapb5cG90vHW9izUo
zgEJ2lQrkB1sQ4uMKiCYpQVimY+6hawOOejWvdVvAIO4ThIa2RmebnZTuPjuBCoW7whAHeDM8T0A
AIlyeiFoe9KYjKqOK2ZzZOZqzPTKB8VChWpDGRx8aknBbE85Cm2m2vPvC45vbzKdGkU6Eevcnnmn
htF5keOl3cZrM2moDao0MLoJW4H78RJW5XG9d6Jqw7a4UjpdYCalHNCKydI6+Ld3CJGB8T5ujbvu
SFxryqS/ETQHi6AqWCfiQLwCOIGOPeFco8CiB25oNU03egulSxwE1a7hcUoAmR8jTCo2SzY6ffP1
8It91mTgXSqBIOdZCnb8uXAQ7OL6C5qmtlX9WYKhFR1Wfek4unINUKW5R5v2VybsYb6c+Nn/PXAo
Zye6/dTgcEIpI+ZVb4I3VaBfsfWZlX5STftLHH8pXDlYoHN7BgPF07l8J89sAuYbKLsGwMzGWWPd
NuB2k8F/WruCc3n4NbYQRCutgIPiUZRv8KHZvin7WKA9rN4eShNGsye63Bljeupuf05+z3IrkFnk
m5lmY/39wT+Fgt45X7DWEgbHwHbrUkrUOb9eGwt6YtFJ3gIBm4TIdYDDiGjDRbW9DfMtsH7CseGz
pOlh+fMI/7mB8JAbJ4gW5p44VLZS/xr27MWmUNBaZYEgvGkknV4wM9xcXsDuC89pReyee/lAkboH
+deIT7GE2XSahE/drwuYOOg7bLYHjt58qMYt9xOQDwkHIiTO5BcQyWb6225sDx8j7GE5bMfchsNV
rckG7/pltJhxvRWwH3mgupoe7GQmHGtaP6ErV4Rxc+/J+8TSPTkWKaTHU0c+gqGlMXUc1NhEGYBg
INTGEp4EtqMJHErYbCXiNMMW/wODmw2DNIEM8pLSMyxEc0nLbT3zaJ07MCwgZf4pxVFA3wGVO9L6
UeEB1IeJcXVv0IPJOhfkS0hSpmE1IdOdzN7p7qs12pu4KJvas4L3dfi5x9rUsaRIuc05BUGEHK7E
GwceMo0gRNRUjjc68iEqVFbypzXe02KKpUMhr8DblDqrVVzXHZECUoXkHa98t0CfBfUwK3tZ6udA
8XRcMqz7/aIXE46eHVp9dECQI4DU0RxypOuaifiIOBpI2O2Ux3w9Uf4XMmhSf88dHpE3788HXjVE
1x6+R0TYXPgrgpUXFTR3e+jBmRBphR4Us51UwEyXhwbXSRYYGi3cBhuXiakr9mzRGP40w6bwGFve
fzEFKTV0A6E0nO2mPyFLy4dmYQtlsPZvQI6FO7T8pxAwruQoqBQeNk13D7UFMPYU1233Jwu92ETR
/sZqJYw8m6VSBqIdg8g/4w8Iv5+Hjv82fymYwLOuX87Ey3+7hXhxpFIAIqfeUdL3ZnTD8YkY5A3c
Nf3KZhZ8CMVr/P3zsmg/nIBrgCxyK4Su0qgquxqFnu9Ou2RHVrh9CN012UJoP0+qhhUBBVX+O6Aa
jgOPwmqHQD931YAW9jUn3BfqUm0hKbt90iRXZMNUIlO6Zb7hHqHPaysqbZ5SPpDlp2PPP7rSd+cu
TzFvKmnk7MREvYRitSXX5OyGDU5OBCxd94VUqJCUzsZgr79BLKesf9zPCdtnMZBUD6NiR/LMDIlp
mLR28fRhFc3g3wGACLjIlMDEbz6r2s+G2wxgvB6CRkPajM+WEtdH0t/Z75NqOzGKXavKpPJeA6aQ
kppeldToiLZ9xb+A40s1CPD3B/6YkB/yAwhrQsnSljcTWgR7WkiIHiVp6c6RMxcJC1VoPUg8xw7g
AV+WN1wO7FBOJaqdq+lDFzlcxSfUK9tKM5qdRfcINAuwbQCL5XJeLcd/f++eIEtNx7A9OGxh0KuL
8nbzhkc3j0KZN0GkSBy73DOihN2K4nRIrKXjl62K77zVBkdhWgXNOH7QgHuugaIzEcrOrHy5RFAR
vVb7qLipQZHA/6ITDbaEPLbxK5tgMpHJrlE15pcQsqIXCmXNyOEcWxjSdXOO2r1B3bDcCvK5iyzh
+NGOglvTIz15UOLKtIUxTK4fTSLV9A2Yd8mJBmhyQv1jStnmwXfqvhqavgitq/vIqGLTUlqSm9SW
mpYwzw8+4MDPSaAPXWINK1bYux9K/vrrzNJiTa4BzH6DzghxeD0AZtDV7Ol0s7Y/hnfIBwjTwpFZ
Hko/5PEIWYht8FHfRl9sgscLNajDZ9c59q4fgc3OIzeBVpdWxuk+D5Sjy9tzHilzTVPE8Sd1Qc6j
5AdxlXI67RQWB7pQPBL7/B2ZEIgC9jkkKeSG+8iUZk+TgKEUbtKemY3pD/ncMyEFkbFA6dulx3JC
XPuiGwPFrWJNcbzVmN4KbmOIS6tL0sWziNYaUkEUFpy0BqUT2+MrfjeRQyGd+57UKSnq6ZAKSYQV
jR2PfRX4uxEShfRNdXr2qbf72JQzjkHCW+tT0SKdw1pCuglnmSWSmpwGr0Lb5ShhB0s6IV4x8RN/
fSsaehgkBPPr/AxbpyWArmJeSS58PG7sFl7XEMsPSdzaVhNiVlcavKFalSQmLnb9dV3B4+9efhRJ
zVgzxd5vPkIi6H2r3XzxIDeyeU6tlG3j1tiHP9a0e3TNAaOKyNr2jmasl72jB/gWqFrKXog1UDCz
1VNDh6fSlfzwITHlYiXuBzuee/ro9Vxr+KMjO2gr0In85Nf83uvNbfNKxtMk26Jac1u/hUaf4Qbh
PNOXF8MUPAUeEY2i9luq6f+93lVVeSZHLoeXDl6yZgupALNHu0rvwTWLbOpn7pp3KNheSZCD0EHJ
SiBzG1IlJTdDYhjDpVlxmXNqlbKz2im/vrQ5VMYTmt6K3Vuq6FUpJHJKQ1znviIvSdnCRkgnWUxA
2hNro1fsPZ7+4Ao6WaI2jKDLWr8I36l156LHPKbEzfRoQ+4GD+YXdHG8yUhDGhvYfrowbD5T46Lq
rjxv2bVzAfo9Cs3BMlhkKUzZ4Cvlw/fboPIobTGCQ52j6a5dFz+kWb+mWhgOXsMgjjof7Di8iN2U
5LkU9Tsnnm9kOAhKHu89hMqly+Qjsu+xejoozuaO4yQhLdSlkPOKotu9dPeP4yW/8HuWQhbrcOxd
+yj5iDL7f8AsvRrxnrGnZEXC+rXmn7M01jR7ojo7igIctOyeU3Y7dh8CuPmHEb58YGIyai4xkUov
9pVzyvR+BBH9uGH5slNIpx/HywKaqG2MgNmwVE+2HViZMRhr0nPhf0gONPBzvihpPpXBlbX1JXFu
IN2aUTMghF0cyI1Lm8gZhZ7+dXAA8L7omM+6D+WUrmCdufIp1zrrY43giJoo9/oFymge4pIWTbIb
mlR2R2ECDsZ1vwXZYdZyoj7MhnNHInXeGRLUTjnp3xhNc/99is9suM4hs/OvKMWJw8QsZ8BQfhSj
u8OSdP5L1p7oYq9/V1TpueIe144X+SyfOKb2P7zIF6M+lfDbkM2GbnQLwmqUJaNvHSS3jk5XFbUw
OlETfAoTzqgTwDDWfZ/X2hCaDJIwGRVsb/dYe19GveRNCG4eoa2xXlUDfnBt8M2rEDuYpDpTPx+d
pDc2XxFyf5g+aajYWnTETMSeUROIffpZXx1MXaF2upcdBf/e1B1Qff1n2HRmAlA4lfqVnpZZGNTj
UwYMTEkBuOUKI6vjcvlu94hgKRNvnMzzNyqZWcEhc5JMiTWBbsjFmV3TuwmEilgtRHt3XayJU045
Yvay57n7EDs6l6KcGBidc4o2GRdr1D1icQu/9FDMh0wsWsRK8tsdG9Ul5tR8ylce4PCgkB7jNrZr
zO00zxID/P5YB+KPuHMYC6S5T1QOomT0OONiqpEl9svv8BQ+fxWJzFR7nySvUK841lwXE2O+HOk5
yeTK58l0IQkJoIXwD0tYps4IOZisvNGo89IospnFk2ApAbG98+F+zFW48bqh1Un5qFHWlHzkAxw7
f4gHK3mC5OqUspi+Wdkw3lj2Des8iVgS/IQwURvjRQnyBKb34qLJfBUibaMFvpFVCr80pSSm6vI6
MUe/13mltxkvxD2UWrywh0/YNmoZffMHZb84toI8G34XCYufGTAwKiBboqz9LEulQOQfCMBgDw1s
4Vz3qw3ieTaQNJKpG8lIZ8jM8cRgpTAnlIms7hfTvf6B60yAQbH2epqVcJ+dIC3vvjy+YWe0/XoC
kuPiqhGiJR6eAt7ouWPwY+qEeYwB6P4/zga1tHOgv+/NyyhshelXh2zE0ZJcnz1hdHGY1o7pXEUf
2T0ufM3whyLghDBx2jprLiEak+Xut3W9PtW90LX449cs+H+T8BF7nSmqjhHytIybNkRXfI2TiMBC
JUCJ+WJdMPZ5Fsvtd2VMQWY9JbshIzrT85ixMvv/MvP5mftVJreZsux5kDOaxo07itDa9CVFJmcf
GYcIn+1OtWjEK+nzFOfwl0eglrd7os5Fj7RM96SC5n+odPPaX6BwPwEwGaoKQp7uxKAHGFOsYbD/
OIFwXL/mu51b/sT3SyrYFUztvEjx1mVGOOrc3jjp4xKVkWjvKuqb1BC5Mx50qaiWwRNJr3xv2TA9
qiUZ5pm1nNbslYX//wBx6bI0ZNbuKoSfz7NBGmnW3/rQ1fvR3/DVHbnetxcdv6btKMhA8Hewxog4
YDx2QHu0hH4jG7Syc1uWLK0C9btiow3WrbMf5/fW7bYGE6D+uiwTs5TjILlZk8kgst/JjkCJWnmL
RUGw4OQywMGcmhT4EGfrQN0vDkiqPA2CO5GnpV414kfLjpw3OL6js7fQKpE9StTKsMwRcmv6FmvU
sU+8QtpFp6VMicxghRhlJAt7guWSO3swHrrbuCgOwwkNF2/uHQLMbzrlC3VmS0Y2MwmD2+ZwGkkJ
zTv5/FV2pnaKKTm5tGBN+IOckGnjCMwV3zzuguTO5fRhqBioe5UqcsDCmlqixjyN6avMqdqSPe64
mioKV3Dktr9F9wS20u2sV8qr7alrsJI/sTRVEfH6fJpqLMZsij1U+TkcwD1Z8L0XPAI+PK5y24S5
LEddvg9PiPjPJS0McbnOfM/GU+z0TiX/M+OLIT9xa9YTdnG2Kbcrrt1A/uvDj+4RKsi/UrWr3fLH
Y0xVKxay/LLHAX+LOgH4ZxhfMAUXJRM1klImfyD1iDXI8sPOeYXcEgKpvm/3MEL0iP11300QF4Q/
TXpRTZd8g5OiDhVCtL7r3goaF62WoJR5U1B2d5VxYXr1IJ+YO5abcmhnbOcD8S1VTMsy9JhW09+c
4O02Jgqa6CbOz5vDhZ4YrKkP+lYIvOxCIenxIp7vnKuJ42YTosF7x8nBBfnN95bxd6RL99KHQsGY
2AM6VoTZ9+bx7YEYEF5AJfj21SVYTeUq/EcBGFsM5rpbrr1RsyJtXc84ifCbHRs4I6SvkomtEoAU
JInU1iDypg6DYR2ajYWyUOrIXH19Tia1C48yO5/pO4rQqcBQ5fSyqW48Ka4kuGeWm4Y2EgzR3Hr4
uCGPj03BpHlxRXplavnzo5yI+O9RVGriDsGn+LiiI3KKEL2qqDrMeir4M1hRWOC50Fcv/wkkLftL
ancfiukVd0Jnq38DlTLm/aHy6Ft/iNw0xxqvihxKkpezRXaDQLrgi5lg+1/e3vubA5wJPC7TyCuP
YmnNloiOj33kWeYqGZNfuO78KEQ0ZEUyb6pXf8ML+raNHKV3Uj1CN4Xz6vaVUWfETZD9vxkg/4o4
eqtaERpUMJjIJcDezHH4fD4C5LBW/y8xZZS8ULeG1S3mMqsYjRO6msHInLUGXM+pVVS7pIOeT2Fr
dLMSSJ6GfQ4t6PkaSBxgoLji0FYDCqN+7vMqaJESGA6se+1uTP3kcBbnvMQC0Rap4GZbMQQl0FoB
6ty6vzZsR4Sgfpw2RfkfAGQKIOVmy97tH5fgA2poZZqQ2BddYf4c1cGuYbAMSC3Ulyoxh2O+Gmbl
owZWHdvdxCGKEQ9PZ9Wp2ZACoAKtxbywxG/WiZiTNHyMtl+WnNNYqKyLrVFXpzy6zhLkHjs7sBcn
VipAbkbuAXxkCRGWno1BrPFYBK+uOB9TCRkdgh5gujU1ZKa/gA7fjCTAf/57C856/Mc1ttXSdya8
fGaSPG8+RcUETJPbmXGv3gl1WlAKdMgfF0MLrF39qXVQUX2KWy9OiPt17NTzTqvcl2JYSAJ9NEjA
PMeZkiJ8sLA2hnUtyBPxNTyCIC1BzLMC5aMQIOhw8wdzWP3EV8KdrbkGGxqLyfykLOeEgt15FdXL
Qgs912rMlN9PElcCohtV1jK2rhld76f1dE1npsuZab3A7X+VZAiLz7B3wpvG0Ba3M6u8rAtLCTV4
cSjSZbz7TlNeq2DdequcJfbX0SYUKF6keBLunCbO5qC0Wl0NY42OVGfuXE2bMxWJQam8k+hKnJEc
F2dzNAWqBu5AXo3kxs0ghudNb6c/8NFhe6MRdFYTabTdOI78z5S2yWB9YOPstq//qY4evtvp3MWN
mYqndX3/Xc3cfEszMLu2XESdv6E9CYswrPn7wGued6/3dyZVQ6lMCNENH2EhDHDtY4AvVQrN2xMr
y5i9gr2JsvtB6B6/frOQBys5pUd0RUzuLoM0SR8xl8I/lQ1Yck+8bCIrOXM01ey+rN7M/+gbUrjU
jQN/UzpHu1pI66Id6ItMjnLfbksRUnvWaMdOau9xE/HTGV8drazVX6S9K9nIED0bVOp2TfHpQEKo
Q7FSwULn7qJV3dMtxK07sS0tcqiRPXxvQesxChgWZiuOkDaJmvWAU3aCgoi4USA06pZeQe1IcuCs
5VWfE32kH/3if7YFZl6i5htZPUftEUi8d0PzWNSZxbxEVc4DK+HXgLYik7qE7pHoCtqddiJO95BB
Ldzj47EmGObh1JfQJcOhm3Xr6Axea4zUhkb1GLWlnDVOjFfnRHBcs0uBOACEhDlSFGKXBDnq4Qgb
pQE5PQOzC0Q2R1PbGKRoWw1mrGTZbOe/NmWQFs4YsyU25jETC9SeDIlwWMY8GjzASJbrew4RPBQY
k/VvaqgG2eL9vmcSTVHYhGYWNmPKz39S1EBtNfrSwwYIfSRrbJzF7KmtFEqyaBlbgeknWFgPv01+
Pwnt1VItIHkUuNm9CRlj3hkDU30u85sJz8xQBHGcdi3r3KXrtveX/temvijDxu6rRMu85f41jGgn
EIp8mB781L665eAQB2bczxitv3k7Fal/NL+InojpYjDy2tWLsEdrHDcb3QlUl6LX0T8quujAxa8X
NIEq5UoKprCcjaYetH+uNiglWmmgfNbKkv3Z4m7xwuGIbbd57GHiyrmy03qBAtSaT7Be7SlLRrHt
pJ3bSKhnwjZz0T6KDGjrVk1b47d/KjFafbiYipTHL8ipWdHyqUpN1H9qWe09Z8eZvG6JpsHJB2XM
5x4kYq/8zu334bJD/+/wjZpPO8B8+YDKotEelIv0kpM3MzU1hGJQnvxoBfzMH4jDf2O4meM7HPr+
XSxPt7BeNnZR5kcGuu1scQRAOC9HoLWjNnS+14Capv0Hmx3M6MMqgIEWJGe8D2N8LQ9+9IB5GIFa
VyyDc8zbOGtZTd9BZYV+lYshv7x5B9g56IxP9KgUUK1Zqx5yV2TORB+mZ7VD1TRQyAlA04VWJjTn
EvEj9/aqC8A1cOsaQSvP/rnNZgV6mDzxHOZhFX0upMUH99cTZ/NtrNOmNkodH39CePueuWY8abpD
DvmGdqrjD/vnQ+3GI+qq+UAw+rwNwYnL9LMUnLqXTva4OjK5QWaisuSY/sGbgCXU8UOuM/Cc4KZy
qit00LXNkv+5rBK0ymTioEbHVjORFL7vMRaP7l3UE0S0CKT6zblbS9J7R0nRYFCp9c7muLP8pyV1
qlL9wgi+hhzmg+7LmaKFzNHwLEYwdG4xyZOYtSNmW/dBpkMClMkk17lq0SG87FEEjha6o2bo4JbG
6hGz6pdSj+tw2fa5C36e2HrVFO6DE/iUphGszz/qmoGKmxtERoOzBqXQWtUByLGAOdS8dbhrlJlp
8VbVypbBYeNZ5A/qJGuBZeykq8sxkt1IZqBt/T9mg9mHOTsokkvz3MTQk1QV0WBPRuCOVikVcpZZ
VN2UUx5eULFpsJevjlznBVVNYgdUUJ9JlLfXBkYmbfHaeF8u3873NDvb6J/2eoTV8o76U2cnwBUH
dLWQr8hHkmXMc2i77UNVFEQ94Uy4ssgBlOwfnkJ1LPAt27ZOVttGKw2husH+CoeJm9mKp+O+POed
NgoWCMRKdGaw6V8RbmPI2lMv4fA7JOBwMOQuvHlzdEOc0kz2mx+clW6NChSWC+bTyB0L9zdQbjGD
qbPemCYljjBsnr0fvIYM+JrNCQ8bc/qjH1V1+Y2xjdH0cvcSGcr6+EHmLNkGFMlgPhYei0e19bpP
vn+Hsiu4f/Iu1P3JVQJxZCg3nadIKSswjkq3kXwW3WYTO/MqgSRKT112KPKpXctx4Dcn6hBiTqeZ
C5TmY2vYz7QQfVDV7SLA9oDQlYoKOmv8wVYao2ozGXxrdxwiGliTgC/1Lr1Rd931i+Hg1jlJ12sw
LuopT99InwlNcPCrY7iPp28SVL6VDPZe1VKsSSmh9SufEtJSfYgpY5ZAihBOLq26wkhSaA3vW240
7NEfyvEDBbtrIpPDAXNmtkLFY/Jae/T0ZpN1h7rwjFxt1FG93lcOdd0AOW15E1jCaT4okmQe7fgZ
1Jpko/pXWfZ2BtTjMGMJTiJvdIPLyRMu6uwYQXQ0svpAXKkI3+YojdgqHm5D6Ms+jyklDNznElwZ
aPdBrnmOE3YT+Ery7g6D3PCqJxCoQmW0NpVRPqNjZtqT4joZewOwI0EXMNJvoP/8NgxD/8RK309K
qDPsIEv8zQhqG3uGLo+qUtDWBRtcEWAdEtrsTyOxdKiNDVEeBp/hValun/QJtTxmNMAdxF/+MlJy
oGZqwknFDVVzHxK9o6R8AyS9udXwEDxn9Zx1Zmu/zU6WO9zaqC+a90vdnjfb06LzsPjalnHlB02S
KVA56/qQP/dm/xAIycBKcLOzhS8O1HwhZm1jqycXiL0OFxdEiTaEjnHiTsplUIJ1MksJ2FidM9+g
V9jLySUCdOFjFtt7MfA/DzYri1JlaTacqOazmKl7PC4QBnSvzNxFEuiHA6Om4XV4DQkYgOl3ea+0
3QTOZsa7CmIQjqzglJAhsR3ceZQjsgQEe0D8MhhIc03toPR8pkX77GksJsCFxs7lM99EGitrcTdn
IPxD/KCivx9svexmSpr2wlPzgJg2pPwQsmvlD8PoaZkOQmIDO2aZjKbmQww3YhQihDVl0twp2Pjp
31PG+YQ3+Dj5hQa1ziCV9b1/lep3R86tsP/pTbEPUjpVYZDuBgDbN3Ykn/zAZSB5B7K+cZpO9LqN
uFSfUyhQzcrcS7g8GXTM0bW2wNtRNFChwu3w7alBQNiXufFLRtQySd1l1sF/fzyl62BqWO2bVVCB
zu9b1OzhEw0DQHxrCLSPrMMcQFHvduXmYpQK5UUaqm0ULWTSB2uj4SwntAP0EU8kK/DkTA8mxB9E
c9xRxOj2P8zL4QFsMMsJvrfsPzcHyJbWO+nZncmftoJW6CvvwOUBuF9HGE+1AbrPfLUJ50xUkAXf
V3cFFDCsJENIlVYQ1tfWdam2oQp15OwAztTx8aMUlGARnAfLPVGkj5XmKqS3j4YAP/odfjqjqIqg
qMddDuyHLZ7P2pYtf1D9YEd3tlp9NaRCCq8DH+6Yg+ki8vVN+4Zvfldn5cnS6XU50QgG3HFyYT3J
fg1oXBeZiTT6D32KIxHOaT3FfQh9wFMfvss/0g65ZhuhYbBTk9H9ORZbKIZ0TDhYNzOdtgU5j6VF
fDdlYw+kVHEzupmHwaqut8+sgEIOP0UmVjeNvad8S3mZPn6q3dkgZ5Ct13WlZ0x7zV7g2NOhIFkm
8ymJLlpVAle64DHrnV2Y3rtpJhpN3VSoG7FEngYsX00tGx4LtZpXBgaXGn2o6stAREO/cyMFPibY
s2oeqzrmaDqWBzOOv1NpGZu4bjBmF5Zwxp3Xl0H5yw+9OhWf/i3ioF8VvLpgUtSeLD0pQxi26pLp
IwJEnUWYXObnniXSWN9AuZjQzIURuUMmhlMhb+lT4y8BgvNIqKLAQ9pMgSbqZnuSRqNz6GFa3YZ/
yOeRDmHyPA3uzQ7Bt7m0vA7JdpX6NuTn6gqpyF7QPUe9MkCDm0/kCT66Tslf0vNOnSduliFuE1jp
wO6Q7VoJDxsPxEkXncSBX6fBOnfuTgslTAawwu0SyheV8kl/L80bHGFOF26lVlML6kSQ5ufApzis
i5knxCHZGJ2NmdRhguoy5df/ti0DxM6a33rm4oiql7+qBGGQULSYEy9Q4KUqWyqQ2rkd/0M/MGB1
akYZmQbKoMF9yT2zBbDm1VbG2hlKub+vQlYSN81qIoSEeNhGj5TRbq17zaERA5z229PvIhOskVIz
qlUeXFBm2WZx0jj1smlwbyK8yFX3LuKYctidKxgozx3pkE1o034OcEECX4s8WGx4kpz+PDK/oJ4d
+rP/Sj0Q+5cbRlcs1NAgHzNrgZESXhkmmzvIt1v5VaMhWKDHjrZDiVT68DPXtsI5yge0q65VcGu4
Jzml/g+UhLx07O44zGp2I8cWRS99iOY0xd7AtI6JGfiZP+H5zBlnFEfFML9IjE/o6bk3L00CI6s9
hB9stsn0VjJ59X34pvdPGK2EUwmlcnOHeKvAgcpZ4TXwdYL0ed3j+RyCdmPgAoFeGInZMF502420
7/y4Mno+2MKbd3VCjt9Ux3uNpnsHXYwnJ2TupGit7qKvTUMT/0XZfnDsoqpMaC8/ET3z/cVSI0fS
haO6GRRDsHWX/thgqLk4REXQmbK+lAAdq2iAi9YGEqQ08BqgdmGrgvuIe+KSr2Er6Wb4pFn9VCrf
67XbTIjj1eBoOhRTdyRvJJatv+XfNAWUzDwrAHYB3QZrJNRsXMUwASt7/EIbPN3tXrk0TZBGtq30
twOTNeD8ibWPqYCLsgPDrb54r9BM0FYj4kCBFvSXhwaiCToaMxcgxbrPVZwA0woWzgDIobRnicWP
/rNwemfJ732WXbvlaSfWzibwg9vQBQdyxk5C+wqyydiihDb/tLeXr3ckspthweQreHIob9Tjxwes
ZV/Ru2dQbpTXF6Vir5AGrlGUbR3EMxPS//pSAnfOOTmyzjcWBZdfwNJiJwBxZLDrdxgoOAROtivi
wpvUwGO2iU2qC+Hgkuy9h4tzaOuEYsbxO0flw2t0nea64ds7T517qy4CIhNS52wDnYSSHyqX9Qp4
0hZGt4jDM0vFAgbvDPz9VicQU7mE+yV855IfcFTXSaMG4aflQo1iOT7UIwvHNXoDfppV4YKK1wec
mreB8XsASWgo5DJU078ay47vCpoWUUnWp2VUyS9KRPWxoJOmnKofQRAl2z7J5w6x+426+rWsuuQb
05BPEgVUaHI0MU508cNe5LBovZSVyPTYs0o3vxT5kLedJ2b8f7vg8+thJJvuyCfYH8qzDxC5W5X4
eUJ+Y2ajmIi4Gz3+fwBJ63rFCE/kM1KX1jLFlj0IbK/VIIsOXPaPhBTnJXb4PoeuAcaT6TdnysnE
purqZsaTUjVDrRitTUyZDUagH8yRg5Kk6fSjBblrlIa80bM1Y6AuCgdzbxbTIGxkmAllEQ+LsJ7l
nGXq/SeEBAbq/zzvxCYv4Umzwz/frDHIw2XZ78dH0+aTbRsBxZa4ml9PNbUUecEdby510Hb9pZEo
/zn/1j+hYK7ryBu2qKFJLyybd0ffrzdWDtOnop3KrQrgriV0S0/bS39EoUNJtjwPLftYmYmLlkPq
/UyE/7ksfm9EjXfjEcYH8b4QrHcg7yPzRL12ph73tiPWEIDXRSroYgyeX+GgiBxLZjQHNccvgooP
30RgGxlzbMFnvvVvzg8G3DKLo3YV+lgstDU1gErtnPW63CR+AHLJhOjSXzxTxRE5MeLN9G6kNZx2
3cGifc1e5iZy0Dl6BWZdGOp3GzTL43Y+j/3qpnQTXz5QFetEvb/qhfGUbbqQTZAV2Ij6sz20gM0v
korZoAHWX0RFdx2jhGQTF4H8tvAAwK4qgA8aDxRh9fHS+fqJm47S24WDwykak5G/UtjK/uPbxnAO
ANfkx7CfR2Nl5SYpJLqP78LlKHwYbatRr6YzQH0Jgi0NH/V8lQfn20psI2/denWo5cLqSpqvXiGh
jsIDE90YSRF5O5j/VZdNFWwFZCTMaSNzq8lIg6m69N/xElbDoJuE8asomAuT01RJWVr8iTbIWHFu
Ax6ph+/3GM1t13/ovOMvb9pqyLwB0INRgCrcTVg4tkciaCZO52OBW+xi3ROQyY4TbXlOs+xzqbNp
XmdT8ctSU8CFoyBTQEcuyFPNhxRVqp0isfgMVZQY8PcxgJ1Gx5tmUA/6fA0OSuiFKL+3qYCL4+EM
yfaG7PPL4Sv9tKGyy8Gp6rDpM/uiBpa5mPahI7SVhTzboLxLSVvCOZSxRYL7ueg8wDaQj40uGc6X
JhAhHwf7ZjB+LFEDPqg7unLaDmybwgrO95EXIO9f8sTz2sEUhFKUVUjLCTGqd3XuKloYaRkkd6d8
F3sAamlmhJWOtHr59G8qJUuUiDYouoU6ToSubNzweVPj2WlLA/rweWnFwPLrK3aKQVWADNawZAzU
exTF57D+1mOYno+8cGbSlK6ncHol3CXErsVfKC5hRkC0Y8ijUYoaoP9CFrVSqOpJDYLkoPipK2EX
rDJSG4IP2fvGIULRlGBTKz7e0z+xYJaxBVCPIr6zu4dit94eke5kZ1rV8Iqg5T1A0SeWKYdIl4zw
aqMAj/2BufSNxhtWh9/UthbxZNGMRvm7QH+Tu0CQwh4elfpQEe3TbYmXU9xahlSUURohWgK5vWc0
f09O0oddDs3AdPvk1H/c9DwczjfCZTfWzurvEy0V6hocgEbIxdvMRC9u/dXUaJ6bqOYniuLDiDuG
P607mRZ8FurMYQwvHi1e/YxZXYusQyptEDlNa2+TSQhSV7t2hhk7yO9PaXZ3kEvKBPXaYazHIlh9
CRv6jO201+jI8t15/osi6v9yRDXlqI6Jq0u+fYUhUn3M4tRmsIAsEGHK06FmlUGnRH3bvWho5zM0
62KkDloKJ7F5Oi0lF4l0AST0EZ1/vECUyugh8RoW9BQjeVFrHVPSQ862C54sW+fHpNJ2HTEEH+RI
XBlTLIAw0jviETPCT3WACk0DUQ5NJZ5G9LcGGZuAaKZWtW395Tiq7waOIG9EOxtGdw7KS0s5UGt8
aOpzO6MxD9Isf18ZTs1iVEX0NS3kLVRm2Xuhk6+shdOc+H06x10sMwWXPAPI3PEVZGwL6gTg/jS5
MLKTqmDnunABKRN5X9tjdjhCmlVtcRy55yzTlXIiFkgl8ERgJVDBm0o0aZ6UQwPWA5/HDCmq2BLU
qr5z73kw59Kt0AGYu0NnDUSZti8nEDsbWa7TDvTA15BU2VVTTxqezoUD3Qw7DNbPGOMrcGEv9wmz
WuflUWrUHkcne4nhPje9NHzvZvPRFywVIrtv5jPGp6jRNsI7Vt8lLVHK6vlZhgViXeQQFWwDXHpj
v8qiUqzgDoQdLFV4SVYMXU4vbIOR8OpujLoijrbgAESSky7UAtVFzZnn8f4+E1gIUz5ZCw52yfzI
J4ToukaU4rqAIyXKGPBmcq9ex/fJLm+IN02egMsmONd6JoYdmeHU8ioVT50JOBz4+WLZvmmxL7Cp
vJR4MJWOBBZGpfEMa9wqXLanLY5dTKGBZj+UIkmnqUoQzyZCWihod+oklnVl1WINcqI5XUqacDgq
jr/a2Mq/GQX5k61kGsrgdJ2d8LMK4EKQQUNtYXLMCMuMTkv4utZv26yldhpe9xkqoTJZ1q7yEGuk
efKFYX9pCCdEJ81QobP1r2IcF4FCbB/qrtsW/fZhlkzvcc21cr/OewQJ8h5Tmaa1G5koguMLELbv
EKI0/fWVddkZCsdiizTtkJPJawr9iLkSRgtJn7sPxVrsbT13wq5nfkeBWTqht7sWJQo6WR5vZFGt
YfHGGRZmfdrnnbrav3OqBFjFGJ6eTOHbXDjpf2J9j0xkznO0gN+Sl43xTWL+af2wpGgZRUIp+ad9
rBKK97Jdr4W3r1hnUnhUmzngMLnr2P/XzcXgZkoOOFZWBIVdrSzXFfYTp6Xm1Md5xyMTJBHFOM88
hseL0We/qFmwVIs6uGMwM4b0S4oGxnqnUcWohQbL1SWftsaH5rYLgLsaz5EvpAYE1hhuzFL7EmaS
OQ00YXMNJCOcg2l0zDVfoAz4QBF6JOCEuscVrIRhnToCs5AuHk4ow9ACZCW5kgOG1+WEqX1zOrzr
8Ww65N+t3oTQ2F0gCSZqgDtiVbi3zD1Qucb+ZDjfMNWXUUmTvrrYGZdzxViLx/+0hSglWyOp8bHV
qOUH8pThySBxQIFlqHRLzByXg5JuhKtWJCXZuz8+Zi/KPSLPoiD9EAsJWtyKItaTNe2avRJ4wP56
qLpFvS0ggZ+zS0JjC89s1Ndqan7Rdb5MI/yLW3J/Ias7PGhq84647xOLk9/HhW5siGFPo3tjTlzi
F5WHPUaSCRYIHNt/NP7Db+Y55eXvAo+4hEp9gtv2FCavORjiYgq99dmCK3eBhSOelBEBwPz/NBQ9
Vyxyi+rTemlzChv34zYllYuClgB+OixGeur9/P1Ms+mFrJEqXEDC24e6QedtokUzxHQzNVXIO4BU
92lrMwcC/wH03QIFocs8BSX2rGPpK4OXPgm1YPNGDQG5vuzapwsZ33VHQ960x3NFEMzWBCXa/rs4
jtDqRiZEHAqkx2yQBbrgyZhuf8WAG8epHrGnpUINsbIcHPb7cYw/c4vlD8RyDKP3LVqS7D/vIrIn
XVCW9W29OVhI6Rdceq+FDx5rwJaA+44xWO2EfJhYPEBAZ+yZ0Q/dAZKL4JR4cnUtkKBVH1s/tVkB
T6DOGnuP2C/XDFljh0bGFrY3EjpNjicOTZDLIwbfsNXqk5VSDJ9KDz0EH/LGGHoFKcFowwN0MHRA
r9BoIunMQ4rcdd5Yn9GbK1wh9d1di358pFCDdAzsGIopGznPXOked1itVu2CBjTW4j/IDxQCu3bx
KU6ymi4zR2ZEBGec1VaT1ITdsT0wWwSqV5GM+ziobWRYBWY5EO2hlt6DpIMTgHi+xwpnYU6HFZpG
VOtKIx2/vKbpGCzTpfE2uT/4Bd9upk/hMZGJLCywI7gtIYk1kFXTAP/HwTxPB2xf/KBHPs6SUwu4
xQjgwIog/CA6OLWJsgnyBzvMMq7xfnDRxe/XTsuJAxcoHzKMFl7gGlqGVlWliTO5pfN45MRDeNgl
nUheXcN4coSV6P1k0gMhzrRrRHJu5XOAXNmGwhwa41Dtvhc8XR5SqhGqCiiPrjFW/hxiYmNJc24i
Myz0ciuEBJNEEap6jaKudh2+0hyLYxmKcvh00rglDzzpqoPnqoP7SYU957H8QwXZAtH2ah+dYQAi
Ufj/Tk1vpHqJhSlM90vbhMF4RjKBtV7asfGn6UtU6cS2mvMmR8PjFmHiawTm+HGa5aY6HPClnkcM
wq1RRgdt6cNcz2KqcdsN+iCExuZMSPIRg5Bum8JJYdFdEbU3uBl0GqJRvhffn6uK8h5dMvgyyVej
5EJA7NOrXVIvs6inw3GBSdKkeJ6Nq9LoHPmQUIaNUSWiS0+LjWo3JRAVu0HDxLIY/t5kBJUs6XSW
VjdDNHLDFUohfTwOzU/ddPDszrD8ZXze2/VPpwVx4lDcL/aevXjs7LeRkBb4j6FIch+OwoyA8LqZ
XWpWdWKbI6Fi2ExOI0PvO8rrDyxFgwHkN3TVyo3JDUfQUInWz4lQ9qpdn2f+2I+f9dzmacrd9R0b
y9/9XWgoEv7TOPXkzroD9wE1jLXAm9YaGvBC7Ev2VhCDrzx7sNvao39aIZLcDSZZ2hCqS9YkQPSH
WcyKYt61nqSjgQ9WZ+f5zVOeCLCnQolDzcvta14/FrAbxgAq9IRsT+uobdyX2/VLTrzvYXbgaNG1
dS5KKVGLfPBW4ZWaJwY6/7W9hgW6hDKHOnGzn2fK+EGDIhF5aQdHOSiE8gv3rCaktC6XMhXDUSiv
fHvLp+KnwPhDp1vtf5YjMYRdaIFAlstFFg5PajgY6JeABqIFc7TG9YbskdbkpESE0ybI8bw+oMAd
UNNz6fptLeqAv8cNFcKLh9Yjat3cVESJsKeTBDD6FqJAYXt24EV1NvOWpPeEovSQrZGkHQ1bWUX7
ixKUoQU0pBCEKk5DppUFT7LUK4B6cIZgm4/kAczL7DyDkZ0D54R6Y2/Nb0QehM2dS/ZFSUWbZd4e
3cp18AV+trBzv3RCYmwUJmTiCsGjYQYcLLsgtDcDAuejTi16EHGjy82/AUga/z85F/xOQDcjuVTF
7JcpVvxEH+XKbFmxJfp8byMUv49w3az35enxsQcDbo7FNVN8jzlpMCxcCHo62+TTqytSP208LMqK
A9cWvKp2J7EGO3CH/eyiV8zrsERBTopPAl5bcLiBNArhsWCOXswuKvdXpK6b0NZ8BxlwgOrQT7e1
O+xVzizxFn9t/meNtU7shTjg5tIr1syhJRQviLYA687gh5kqyAgQgkIrkxDKtc7SFtuelyeyN8Hi
AoTJ+qHh4MvyjTUzsXc7wDiIxcguJZs1h3J051X29rVoaP5m6AHIlseb9jvsdTSyRldUfl30824v
zie6CJjB+Ocya2SWBwo+1Tda8DALh2JPPwxZq4EjVyY3vlXJl/4pxt/8cATEaIaICWENksbnrdq0
eU+sAfQ7EYhMHspf7IH6yEyNXasWcZmiizvwhzgy+0TzN0Qu8Nh6MLoJgD2fxzxxNfP+5BOP4j0d
p+QyaM4j03RPfcigk0i9jTvzUatvvz3tcN2ZblGpPl/Od45811RKPK5wfZhIScIv50547WBjU+bD
8t+KXp2LO93x5oRrcZ2Xqs8iToFo8iuEA3Bl6Pota3tejL0owYbzUrutIWLWQZDUj6ZpPAgxfABA
ANuhPNQXWY/2z+rYfDPXlAcBRpfQ/lD9nCetE3mf3D1+BOonZueM5HO+cBgQKyfrBDDUvMrKgh5h
YZNftFZdUbefZiqcKvL0orRgC5cnlsi5LuBhCnrZp+wzW4+yiivJz+BQ1htKNaB5rG12Crl5dbJU
FHjYDwhGYvbWdADAlFiQH7tW3YMoXZwEi9LiXwcVBgS87ObTiyY1T8hj50PX1aJY3HxPRVzM1Wfl
H2Hk2/6u/cng0Kz/rGpLR3oBsUpREV6OVj/yiHSi2l2xsIbfzB+zdYVxonCR2sGTn3Q5kFiuPBrL
4p2wE71ZqjYIZI62VYzB0WKiKKIOBcWr9bCeuwG1TPQGhglpC7+CpCfnh+R3OCv773eKLYoiok/0
TUi55JDKSlzH8GtWJ4ADh4CRS9kaNjqEvsIpcBYS36x+U0+t2Mk3/icCe4H0ItWIFhq2gO2Xt6RH
zQWDk52GgoQFUpb5EmMsc9FXhpeTXuyuXBC1/KCtUzbKz4e1yEvInaop3HUZOuALzJMbKviHa25J
ZT/iNj3VkwKMc5rd28qy2NMsx+ZgFp8YYA40fKCjwwz4hRyGpllPa25YwiPzFsdYXukych2W3ubt
jPW4L1rG5bwnyH/ilLcqu9p1A0rMYYw7I0SBHtnm+50JqhfgsIIV+gGKoXZ6uro67+g3/C2b18S1
KAxJOS5pbfIQbkATlPaivG1lML5lERxD2yOJa51+i/e2WGqPB15IO7yKWbmCNuqkaWSg6so9wYAs
CKhknoUqzoGSwD0nneMAC2U2ChBUIgCywDUn94PiEvTGx2k6JkXgn33GCT8SqA8LKy8qd7sxXpJV
fi6KrVEmfT+cjT3RNRudPoEbcCBDVNQ2fcpFPpCwWa2ovcJXemCNHipwieKqSAnm9NbFg1zDgcxK
L/tM/p/2fbj26BCq4HH8EOHRTfnue4JBmP2p9qsXlkewkn4Z++wgbAoZ1jD9Jx6lgetzS7c1EDuh
HcmhQIKlJJ4S0Laf8eHXr3xr7RYtpyxry8/aSq+SihoURcFW3e3RzUt5W76qQ8rfCyINTxuWMcOq
IMzzxVE/ShC3nHC6iL/i9wp4uY3Uo8zjSjTrJYm37+TYFh/30QB3xQgP09i3foZJ03OLMgT1wB0k
tb1hUJJhCiks7sM+oSxFDIna2hG0lyhIRjFz7oat0VYOohUXPQE6llDWJae78drDfWbeZWZB/y5G
yGByobp6Yz0ZpnKA+F/QnRQAP4ikRJX/hHNPr/Y1jA7ED2Q0Ctfi4RkdxlhINdwmVgJri4IfJDWq
0cDxkBFHbmwKb5ipQgyr18X5RjUE44wIebjm4UEISs9Et4fPiVJ1/avac8brXt5Z/OzJaiJtL/a2
9zspRtS0X03ubZmsW7sbiOQv5iz2Bs9oQ3XLm8GB1AY5VjbXNtrhToqZru2AkGMfrsIHXuDzzXNy
NTIM/ZlU5c1SJbtwkTgLvp9lYzhfXWlU3i16qsvR7nJa/A0MzyhzJK7XwLpMM6L3Y28GI9PE12m2
lfmrCADdoxpmbYSg7pdOUkjcKofVrSDBL/mpNjVBlr7SfIdp7nJFC/1xhOGb/v0K09OdGT0Qc8Pv
o91f6kp1QuLBpbvGWxhh4PEpot2gfDPx+tjqDpugG4T3pY9NMst6sBQm1Q3I2kOlvNgO+jwPHu04
ukv+W26HYRmOIRnwcmuG8MZFHnEczkedWFu1biMVl2Eq2HwVckM8zxXEllUItaohSR+ENpChXINC
xc3Htqgt9BMajRiWpNofhQ1cHAJgyk5clnpwgsvZBbao+2z18uekh89qGRfj5R9RRZHDTXzKoATz
3rnsv2UUvBB4hVXK+XCG3R8lDKWC6dAFbS9Fs08P/rVpu2aWNwJfkWkXNhnoBAKXQUJC/wnQCG58
x5znx97IbBbwwY7EtsX2gwC5i7h7Wr8lx/FzNrUjn1jc+c4vrPTY69qwhWeHJfuOzkNmLKrBF+3r
YR94egEVJgCVu38ufLyCJcl2pyUyEM0wP9iYiaf9yCIfXt7mRf9dNnOWYwxat49qIMqCbh4lPJiC
O1L/BMAoKIDnf6H+vtjdqNaLbqRfLeSRysaHJxLtcqKe8M0RQVWkrNPASLB+7WuWv12i5vCOfxni
ItU2K29HRrO21/d/120HW6kpPaFS5qSeB+KRJXPMGsAglyVOJRTX9vU1PYUz3MZ91ZYNKtuA8k0n
og/NwXO9EdsHzAd6uTwlMAqSscfGhYNWPGCdr6wj8W8z6E0RAHmRRPzUfj2sFPMhluNDcXxLW3uW
38fu4R1FknSw6SV9M3zMIVmaJCcLcp62TnboKR+DfFx0W5Y9/T37nD3Ck+3w2KFVn8FVo6S9fYst
3gFWtLGcCAdm/vAXY9WFzEvQ5XziBef434t2Tydq1/D1YOeyzyhKFivAgrCBnadv38TneQCyGZTP
QaeWbDZdUZjFFwkhAXOBOj7DljgirSL91D5WgoCtiG0ISZW7LfDFDffthoEKPEl9YQuJZslUb/yc
i1uAa4jjtI3yyFTsH3BdU1/3FwgVUsBUpS+k8oSpy7AbOGZshaK7jy17OrUwuyOHPPWNuN7/36c3
5p4V1jRP0mvaOPVDD8mx5dwAjb48Xw7HrwOsPxc4DtsTqV782GyK68R9xJ3LAD0N9DL4DTrrC4OV
DwUiikRv0yWrrwCk7N0SsdVMYamiBeO3hOKMn2msgCE1/mrIYz3ELguSG2C0TZNOgnwuHhUUYhA/
rwWiXqGxIK/w3bXRTBmaWAJ1TAkrkoaKlte4SeAD5EcJ12nVsCQCcpA+zKPrbxxkN7myrkqO7Gnt
6vnu9I4DhJxPrO0I6bMto/Iq9bXRdyOXOtNJMZUoj2v8A2eMDfYQgdSYneFpOx8tsDg8H06Oy6JZ
o7pdc8+/3AO8NxOhSP9UY24a5cS0dfmc3HTRY73bii7KYvyTMcJltfoXeDYaQgXjG95Cs7ihYySX
8k4NeZ4eSigIGGimsVtHmoaley8De6KA6+EMobxJzj9uwn1Zlp/2TAHCCsNrIUnb2LFaaKHNW+qu
dXk5LDCKebWhLwh2kEx29uhqobR6B9mg8M4I2RHjPlcVu0ij+IHCQspuau1yfbQEHqR5cbu96plA
+GV6HlrhoqOB8vPoQzkEi3qfikFyJmG8CyTXwV0q6W9d2PQ4/u9bInyCTdMxK/+FhsUAOVuaoIey
ppwZhxDjqjpO6cOKxOmOdbm7nDVci0KU+WqoV2GlV4VvUDWXPZkMHabkHnKzKdTqpXyV7Sr1mLLX
8v8j86CzByoQewLJjbAkWKflwFdI6PUVIYi4PCBCnMtR9xRI4UdF/nygVyCXyVioVzBa8xXN431+
qsFCPwoDBqvN12AakVj3ItUo2rxf/iUiI1+5vAvpUJgOZ6+AuESuPnDrJmsapls+9fOKL1CMrgpe
VHdQGW1KdcHEZfsBpLnIs2aVqpDYd164W7w8XpncB9OdDnlWQ6Yw6uDmc9HhmO/LS/+WQHv6y9yr
54WsivGdyDBjW3HHSM1135aCZDNYf/CEwqA5YhU9ZjmxXtIx66m3zBO17gNXA/ZKnG5zPE3dORFP
QpMMp/Rpewppt1oD958WSvFSxv6Sv1DkuVLs1/YUjno3Ib0QOTqpToBUiX9PqjPtxwDFNMcfO1Z9
Av2b7O2WN1F908axSKZ5bhJLZcRn/L2sXMVjUtqXBebhQe3YUbXqD8syANya4ae+3VMAQN4Ue7tM
ylF4t/HJb0mIMvKR+gZWT08gra0PzpsIvAn1Y55T9QhkULY0pK51hkNaHSSVAc0yorueMxqMPHcO
yhZyRF1bPz73Sjzt/X8U201Mx3xlXMOy7tEH0AolzFFzzheA8YOo/RP43I8C8MR4q0XIUtVzwdcK
iWYWesZo0ZeBCw3CHWqVt21hs9QfPsSLU8kpsTyBeBEJWHN75Fq/dh19L8SGXI6xlD1Iwoj1BtyC
yX4rergI+VJRzy8fZXeWNzBFTs58qsdSzoqtIc30gb4cn4oQKXRqMIPayWpP+n6x1fT4e1XVS5Kb
6OpA7TMniBinpVPK0mAA6ZumcQxkFAcMT3oMCszJGTWrG5nVSXMJPoPuRusWYUEQzt9XXT0F9Kiw
hqORB4wNcM1vaWo7DY16IUJq6sg8S1CANCqSZB2pHfmpV2dWyglN9xe/8AtpRiL5M9uxxj46TaWW
NuJIF0FGoBVjNEej+vrE1BL6CpCoKZmPjEBCUTHBUjSn6X1YNYUd0mW8BxxoDK136xMydAQYo8Pi
Vsyt0Sg6WxFyktwkmOuAVMoUpMOS77k2PIcXNst4yfly4YvsDGQyhR7J9valDE+aa5kdP+i2cqLC
zaGhk9RO3XhEQg7bznF+N9eVs5eNwM/tB7/+ChBBga0MjaDNqeOkvDruabYXg8EuG4DnLpU/ty3r
2CtWE5g5LFI9KwZD9/ZR73FPStjvn8hcT7jiG5BT3ZgnbkTtcF6o12XIzvqBDdfNF+hOi8YaF6ff
sJDVd+Ajri6UaBXa+tnCyIRItByiymWX/0jdRnXhSNz07+336uzBGA7zE/kDfGpRXTIWJQZa07+T
xPmxBFZFgGlVggxgcvGO6xwEsfLGSF90drUZ+fGDYYUN73xCilDCWkvs0Cy/gH7KOAoxF/7afB0Z
Pdvt9e9MxB9cIrv5dkN7+MMEIR8zwRS/NNfCFDoLt6L0cc9JiRn/MCB4iqfX16Gd714D+pBOyEnY
rx9aBUh5m7QjgB1SHErt+VWURQlBnf4rW5PzJa8aCG7H/47XePFj/Hhflhe2xw4Hx7UncbxWLZJq
NuPgE36MggqAFP4DPw6NTlVZZ4VC65wO8xxrkANmnSNpYtnywhxszn/fVEDF2J2dIj8uv6kE9goe
P7pPK+ewoEH4Jh3FZQxPsa/FuqaallBIxxsiMr5aRm3b414bQTEQZpWyvMsuFmKlkTqSMbyovNEH
pYNFX2LkDUqcaM5FI4hnP0HS3m6yB4Lo6yAFYwhvan66/qrrkSV/Je0WXtYyJewY/TChq5V2V4Ae
4Il2ts8pK6B8KDMXANJRAvR2KshzplJfMbtgCot6FMvdY6yqLmbz02lYTfqPV84LtcgcWGZWJqqs
x9tpgU9QZ1fBX4sYRlaLHYAemqEON9D3NUQTzISLHzmFfIvP5tryjVP0BfET9hff8R5Q88g7vYGF
vtKM0Vgw5vvT9Ps3qB8OML5ZkI/40htE/B5ulkVcCuteeLOQTI7+EfmBcs+35dkKOl5KrjNDRa6X
hrtU+P9jsca9oPwSdSfHbPWE9SMjyN2oDPHsLLRIIu/C/WHkSDX1Z83A4Bhi/uWWOqzCUkhghzGX
UY396RrLhVCVjFPiIg670C5XEvqW5KF7d3eLO7P78JqGMfjn2O1hURr49mZutyOMc6QwjGxgHp6B
CDpiTcWSv4nyGZmONDnu/sviMjn36mju7jL/eOub2yK5VxznhXhSElhm0IN+KeIG3FzOZawB7Ccc
tDnMZzMmCQHF7IG5eHzHXvvQ5G5rnmsQbvJKn64H6vauT3KaeGTM0+jWNHVQkYPyeF77mVAG1ZUg
r1Mga5MKGD87cvOifXauZj5bSwSEd6HcXIsOm/XYwpQi4IHzH5zj8Fy/PD39ntQkyQKWaBydOsO9
DY9e4kGza4vwkys0jWLhP7oj//soYlEaD+DSCm4FAxacSk8b0j1nnicpyjb6Bs/2dsuowgiafbbw
pzW6O0JC52Ih4uAGf9rclHocPjrVGRMHPQqY6B1mC0buGAdTgde/fNj3RqSKN4fJ4rj2mdhOndfM
j1YarJINffWQ8I2hpVPFucO1FAhGQDoO5ZtngGLffYcT40p068OFYGXEd/OFoWlQHmVQzUMoLgW5
7kKafo6pyOdLSPRHIKkuHV4dpr8g8DfAPVx8/EFDNTzJwdH97rG4d/bOe1qAtDIPCtRjtZThSoUB
qAPd36S52p/kcn4Ongw0+PadmVPX8sYPu+4HIo8gf+QmB9+aKeELhBSF7JRXHiIJaNlGooNAV2KO
EFZXMRGV4d9y0+fvI8ZQIarENjLlwYzjK+imTIiT0iHXXUThxBmjf8JRaxC1FwPanpyF3HTTwlTk
uM6tVy95fINmpr4DNg7WWU9P4/3GhniZ+8deXb580YnF9H9v5K7JId9521MxtRhwy4sbHNRblB7B
QoMt/1N6Jxlc04g8AucvO6LShptlnh6ECBE6G9rZPP4TvNVIm8woU01lpStI9hXeZP/9B3aRWOF/
RPf3K+dBBaVX5/5LVIzT1RHuQ35/WpOctIDBkxbgaHcK3Ql9kt79NLvW3ABYTC+YubR4at7uX/zZ
IQUdYdb42+KHXkUySqvCt5ZNwNUyGqH4SKhdngEwEcWeEdEPRuTzt4Op9UyGqWY6WF7LVbckz14R
CqjyXMPJtW3jqQ/SC594idSoX2muBBpMJ8MGWJt6GyAA8ulu7Lu8hbNhpNm5001MBHn333+Ffsnr
IRC6gXM2SQz9yHoN2sa1ET4XJNoYsPq+W/5I7GuPyKeEGCf+TDoC1zkR01vUJj4cF7drqMRb5HXR
C1zn8WQP1ABcdo9flMPZSTpfRLs7LgEfa3xhwXF0Og/fpF4Wqv8JwmLpTlM5JaxoyCe0VFVVGjQR
G2M3TK/n/jlbQW4W50kH6GMWHTjRxEbHtXUVDeEbe57J1839Ab0xfM6N9fPB7/M0+MCnDJGHA6ia
MtRjZ9GtEf9xWP+C3ECNMso91+GZ70e/zLzgjw3hYRl1Px1kIp0V3DhPIGl/oaC8RCOe9XegcybP
Mx3YuO4KfDaRbCWkA3jP+/D9nUcjg+U+5B6R71ptRDy8g+mm379Ykh9uRBcXmpfXDMmX8Em9IEOA
NEYTQ/2x69F8vyiSvsLbnxMq/lg4Q1hPB9NbvhAZUD1+Oymr9f8rRkIpYsGjSDFDEU5VK4t8fBxM
NH5ZMtPIL7Rkh+FG9jTML6YdMvQE8k+zSO1I1qUzSHDjpw0GeQyekcWc8iwiqIHCCayRun3i/4cW
y8ZuzGHdQQVb6kCLPOIS2MUQY9VK27wjN5YCiA9z11Oa0vr8dqop6nMFDVtNkXvCiceQGlO7K8v7
hw0TbIY4DIoJXPsv/09X6JS1NdefDw4CkVv/qgdJIINE3Cpeti1U80lG1E3K7WixGNERpNlWJQZI
JVcM6zWDENdvu7Ny9Pg/bwrUVKHoeWFPZ2JcjFRZ0WYSs1KM+sV6g9uSrjQIV08TOdIbcR7TYxqu
vTFxLhWTnULVogwGXEUl9KHM08tXMwNZSKw9SJ59ohOpVAtDox9bUo4AIQTxNUnwAwIk52TYYZyj
MsFkq5yZHIzVYF3e9157L5nGKH9RFgLHIEOqsetufB4fWF0veLVID4vraWGHmnvzNYB8H5GUDJqV
Hvdjdayv5v1yc0Zx1QtmTLGyCv6d/tR7k79/boDSsbKBUs4rVg6Jgw97UCyBfJObXtw1t5TxAmSW
dPJKhBV/14bIypnRU65YW2biGmpvIkXGg+HSf3bnGrlZCuEe7AGibEMxlwuXHcyuZwDM8NB5ud1d
vSTS3St6+ksrli7KP9oqdK3CdmzhphWraE3l8XbVHJcGjmu6WEBdTdEePktBrOEvHCHmQb86WWw3
A4CTc7wy0hlOAA9R47Pq5sfdYe3JvQp2OU+pXGxKASPtVDxse+B84Nh1dvw1epfJTJXxGrwqe3Ha
8oXZezAAouoPXOe4X1j3wqtDsgZi6c1MW+6ZFv8GpjaimSMUUXYxswW5rqWbvwjHU9rTdPS/kxl0
WRA2wmtHFNwj+1fyoULx5HnQU9HczAIfppkVxd+i51SVKPXtWTHYKYjLNZT9FcbmXJk0qosYrzUV
m/ZAtJjukxruJghB+CSpJcXToz/g+RHCw8CUnk9zNxg0XGRl3A8QzVv0oodWvNiOqdzgctxkCvOg
WG3vfad7NyxBncLwrua5SKgp96ion0pLTbvsCyYqohZnDh9NAJKsiSdCk/rt6tnQ0oQFaakF9kiL
LS3fPLNo3wIiWpoAn+WycXGP47Bxh+U7ptx56Q4I3ajWZBisqGRzN/WSBkOsg05TMGvm30s+ZL0x
mFVb6Mjzh0lYV+THeY3eMxHAvS98CDfWHX4HgbCcwpnncsTGI2en6p+k7Yd29VUZY3da5452xWUK
fIjEwRrcfMba/aBNSMOYEwyXH8RC8KIhkyldhC9+oIrfFIiaAbcmp8J5EGMt6iS0hMBdJAGJz65Y
qvGUn/NuJn4fgezw/p0Oj5meogG5dW7dYqgLfgn0vjzoJetOQs4XNGOGW6GIR+jS1lH0dijOJHGp
Kkf/wL8ydq0/JuWmQOveY4T5EkD1oASQHY36csD1ce4ZyBtZ701v/FB5bcY05h+IBQeb/ilcrAMW
nJc+ra0NNgVz60KQFa0wQbD7DiX3+B2L0SreZtxycA2bxWw7WuRb+9K2/0H4FsDGN14pSPyA/Eon
DbPO1kT5m3ge3OAeN3DB0r4MP7NFgCkCgxgk6OoSttTNGBL0CrNd/9grGgocaNuDaNZCz+NgvSn5
49zfqDgXDMxZeWytH7uZkbNlZ7oVhSwHPD+jtGW3B4rv8i/SAsMeMsnr73uOrc4CDQ9w3a2Z/bj/
e9/1rVo2ACYT+zLVTQQLmjCtJdtecmQGTIYedpovS7Vw4Ifp2ouEU/AN4q8tT0L57NIGXYPvEPOY
1guEIWYw3Mbq6WWSjY5wFfBZUUWqvmMFaJPkSRMwtZYrIjpNKvGkEmLrUF9p8ovKUwW9wKyCyjY0
2e60MwS7vIEvTC0FQzBxFYmydmFWsmbH5z44akG6LXRqgsYSpBGpmmwR5YDjEP8463cAe4IZlWx6
lcpbywovMBqqnwQnDFIr/uEJvTk0Wd95+Iviq4cWst6iO2xUevvAdWXh8BECyTygQfpewrFCXQpI
KWTrZQP3I9uKFcnjeWA5pC9OfsHI4E4kaLiBDD8V/3JUeCVP7Dr4JQQU7n+2srEJhX/qLOZC7K2Q
5xFXi0RiYH1PkHbo1EQKHYR0k5QQB7NowPPPZSCfo0MdrNfpNqUbNg45+DkAgiqtsjesENOAifSP
IRv2xzG1whfu95BIdwsFwvK1qc4CF9vp4rKZjGDOCFdiZuAmhkvxHvjSB76wgUBgOpj1gnnWGLop
9KO5IxR/rSxi9YfljpFiwyonmdJwLNB3GYmp911wYQAi5NQB/0uwuDuw7cFNasvkAAHPhvtWNBlG
LIl8zFJ/Qwh52HKcEOfk+Yxo7iWvqq7OfKSkVk7pAmaJqFv/+Gb4klCW4BevVCNvQ2hXDgHukF+F
1Kb4aPrnvNIkew6QxdA++Wi1GBTOL49aNkab11QYFLfyRYSHrfOsplUU9mAPLBJIQblp2wcYkGDt
bIJiJQ3YgotIxageNQYYCjOuShwGoBAyxipcH++CXSFPQ4u4gAMgSh8d8ZY6SAKYaEguuSpINYvL
C75OkOMjqMhFhB68JYhXJWTkY33w536zGJHsWMKkHTZ5e06TPsyXRlF/t0F0KeR0BJR47RGYeKkx
08kl5zqHSdc8JhjdV97Ejvfcg6pLKEF3iFgVnYxleMpLTkdC3v2M21EkKSlEZUPQ2cqfGF8eDLG0
tOXF/3/0bayMk+jXtFj/z6NUkd5QdyIqEv8dVjEg+BSxFu4UQ+U7gDPNN6+eyM4avVzt8Ach+ZrG
mRmjX+lIw2SSodTg1Aws4B1vuoHz0997o0leFdibec9DxcG4DmSGGpUY/U0/X+/Hj0sy9MZAaofc
YzwdhCzu31FfpGMASlk3Pe5/mJiljfL01QGArETnsGMQGRNQD4OOuboOfDtMMm1e+5dnnpVLXCFs
zdyrDhtpQ8upeYYAFCVegcwuCNv18zYc2sA57MF7FoA1nMh4FlDTru3f5piFW19zPBWUovT5qcJX
eO7KiL2nUZ4BB8vBBZls6dW7/jVxhqjh1kC+2yi5olPPQRBEG7W1Nj9/9hNr62UgHzJ1VeC3CAaC
tYs0doWRFy4PuIwJb0PvO9dX+xnaORbeA+4qUAtfm/beX2BECnHjETUUN4Tv8/UErnbLwl1tHdCY
Xte9hqsFpbw2OFK59JiaXXoRIRnEIWjWy1kcnYwgwIsCcv1igbZePi9hCKDZl09s325a+jpKlFrO
uKUFh0O3Xa1R3qvfzp4tJCEwkXPtU+IsNSB026BVwPVdw8/GCpEUunlHl4yjgwG4XuvcOT91ikMH
1Zz0wEFx5Vjz+o8raQyW7spVrMdNMFqkm+cOUGHdZTzk6H4iX//+HTw9R1iDJZQ+Eurek8hOvxQv
tLBoLWN65SA2jmV+lRZ9+nGVGIgNJ8pnvEM6CV9XlMGrZnw3rP1S4UWOkavcBcGi0p6ClPJuDIbZ
mmk+lL051t8bXeqUwW4J/p/NZv+6UV0qvZvl+rmL8Iz2HxrTE6imhIAqHJrbmNt839YwnFQu2r+v
ettifZrcri/RAFZsPfeII/UowepqgisZ9D54j8V/OFuAyL7aVZjUT7u2/ab4F/01eBr6KHMHW0Lu
ZemmI2yohuUUE+IKHVFyJkIcksky83qWF+RVIP2FaLWxf3O6CWf2MNbRPMDp/S4SKSXzpoxcTcK8
You/lLO2KOHxfh6h67u8u7rF+PchN1ZUl+EgNj+f3Ypb7MuT2VUl/X1kJSShRt14xHh7KWR7DPwl
nnVphG2keIdIULWU1goJNP/BYX2TdYehSBPWLTHUOEPEmIKZ5d+xGsklYhAreY/Bc4IZyTkIdZHa
YlRwOy1oTCcmx2oDNaUir5gmIQ2FojOpMFQpK7AnbzlSJeQ6/zKY5HK1LpzCM056LpA3EbUvzLQ+
y/2b1SMMcsvqhVbtiYXVwIuoqmGJGPwyX9Ni+U1If4nnBWumjrXEWPb724GGjWWKWMqHdUcFFMjC
Kh0pHmT0VdKkzcgp8ONKT4RgT3Ejjy8WsIHzplG9mo+sBOLNzEe76DBxaLNPKfo9rtNUh2DfBw3k
CGhM1rOPBzg38slEfON+ZE+NHJl0idbppieanwtkL/kGbu8HLvEdRrj5z4MLfLYnTQb5XSc53dWz
KhgGBMyCSr4A31HLnLOViJ0zNxFdRJb9rggly1FPcRFer2cJpt9QZ38JosZ94BYC4upl2mj+YNPr
2gFTdpx0Erug0gw+v2xsMjTV34x9T/O5JCzcsL1wUj7ctmDMwRuS87u2fsqbSeoa/yh0Z8AzZyO5
TYZuwuOe6IC+DPWXn3+PEpJYazdiIIB5JcxEOPUC9kgifvr57fsskTt6mGRWaVmyZmbmlykHr3fr
jgTHXS0Z2PprqQ58p/DdApLdYsdhJNAv5RTpE4zXYwnzXh42Cq6Tj8ASeWx8j0CGFucdqdsxJo1l
Rc+Gr6uNBHVNuUFd0vREgPWFhhVxYITxUZtlYQbioVT9FcdXoWEi19oKd7yrHsMK6QXshFyexATV
4kq4S8gxVx0qYXmG1lTpcOw//Z7gwjL8qvH8e7uLIftd2fMbUdyRsnn+0EXC40dLhGBvcrgQU0ym
PX7PkPAWxZudKi70naaDWJTnt+7SrlcVy70/S2Fcve2XWxLzXmFO9KyWIDxgTysFErLWUnwkpEMi
ZzThmyl7gPNQVusBMrgHfrpM01deMV+IzZ0oxzHDSXCC730rZsUD/Q/y2uyUNl5it9Hk93fRPYh0
ANWVfCW73MC4qkL9UDRy7IdPuZLh11QwCEYeTLRH44r8cSayKDLHGcu0DBN7K+BU2mNrMX9DgFUr
Jm8aNJSDFk+xxd6+t0iqrmJfs7gI1kv5/XKmQvfstMLnsYCYXGvl8nkMgZE2YqVmKYWGaoPN5esP
pTf9mqLGGmNRu9kSq4KXm8Z6RpwBY0TZW67GGuRAInt3McXFtNkalXGpR3qRjry4g1C7yW/D4NJI
/7UOoXtu+lUFtlLzn3ZEX+QVtduzy5ZXIz9Ih9oE65yn18xz4ZvHyUpL2mhr1Tl62HfeFLp0AezI
NUa5LlVYOIRL5yl+EJq09IkAWAodV/JScnyXaDgymZYpIJotswbqVqGwY/lGY6u5ZOHgisT7prHG
sBRHSbFkRaaY9xu0JZ21ei+HP3z5cuslDpqM95GNVHuHDMbUjm4uR3ZHEj1fLNzr2DCZM+yAQ9Mo
HaiWayN+iIwuOv5Gbo8tIZDNaeyG7OEKquObtI2P/2KJBowXUcwidbrNUX6n+QIxRbrhT5mdhSGZ
tu8cvLMjzuuEuWpI4ZrODetXsn2rn+w7vDziIfytfE4pEmpnkMis/imKZw3Xs0UHzhSlymN3xAHo
kBv680EA6J2VDoAOte29Dq7KECw9XrWpadT+UvSy0WmN+PMoehUsQZDxngpWHMFRmW7Cb0VOqcAM
AhALkGWEfdTEwrCsTexU1ZzfZaCNoIZmQaOT936Sgtp6Jh6CbNy5lE1OCkgyv/U3XepYSvoVkBcx
9jy3vejTw4VWFsAVrN4RYdTZ+ImTLC7WQ0VmMo7UaIYaaA2ecbvY+QGqYT4jIIw/rSVpzGl0T6pq
7pkR+mLw4eKXt1FFNGfPNGbldNjGJLbDi0PXN2pVqvCq5/3HFSo7ravzk7WAyCOa0Avv4X/B4oRf
sHz7NmFmCzB1WZkDu2R9qLmIQ/0bqksjNWjlVhuSrwGeOIJ74sLWsyoyU7+LkN8ANTw2/05Gx4lP
PHyM7FxEe/2SU8jV9V8P4vjGgkmiSyv7NKnDXjb6SIvJR36iF+IV2ktVev8uvev2c8Rry+ETXx5i
IqjMhdv+T+M1U7WC5ozd+WT10SMOu7SS+xrTcteT7vjON+5BPIqpIsanscG8EzcumHN6DnMOBQHL
fa49FEj1oSLLW1/IybqRfGsHamCtUDKVRtLkOT8/q5sOxdWvt3m/iQWqKeexwfKsfj0WOjQfifBz
IWt1DaBpHVHqyiEXlZjupnxtqHB2BDeMl6npkdTUPQNvJY2EkehbPQLMYT3MhKINKp+UaYtkJh7k
UjBVMRw6Ll55z5RN1V4+dTSc+YPDeajIinbpYg1ML7pPkEQAERJoBBd5VgaaEtKJsmbBXGXddE25
KzGYmpm28GITc1DMd4/ST2p8o8KwbFScGXWNSxu4ZWCCVYPQd3LqnDhFWrSNG+69grFMf52lyY39
eOeSBShFLOlA5+bZtiTxA53eUGVBRpk9yEAHBDgwrb20VXASh5oZjrAD2GN2+o6v4NzgRe1q0H+t
F/Xu+FHDePcWJihfKbRfbZOv8JY8w+PB6t2+iovIeDiIE/9f7wv9XqVij3MNF2SwLbRo3IzP/yXP
0i1+a7TzXPsDtXuY9AWQ+e5VWIuCkTB0BQ+g1TTkuE/6rvtZW6JnsAYKU68Oj+M5I7yV3lFgEft8
z4QiT6bnlPzfjR4RTu2S/aSUaiOogIcHEeLX6/FPbV4hJWZK1qGSCAgDbVyJq0VT0tqp9P5FsDFK
3/pul5vNx51BaaUe5i7y3knG3HdzonXLWEYCB7aYMiSotp3kHM1ePWJ/p4ABezgZ8nOmsfFwX7lM
3FPs6ow6SNCCJ5Qdf5rtdwLdRqpRYB8huQfOdCzKj3MoJaouXJ4MJvl+Lw9xCTU+CcorG8CgGL7w
smyKgq3RkmZZo4UpDtIVv4M93Tir3erBgy8R02i2Ybyj/Eh/Y+Bb1IZV4QM1V7In19BzIGDJNAXH
6L/Tr2pRrnWrWqoHr0ajIFKB8ZySlOd/dwCf5aFzi9FpugE+iaPUFDsjFIrGV2SCzd0DlkBXK7+j
Ux4A/j6evgRKNMKrPFQuIx+AJuEij6vLSO0hqH9mOx8o15PZ56/3fqMeGgp1bL8hnefRW7VsCiOj
dLAmLljZt3kuwSc+NKJHkOL+rnE9yPgy8Oa8hvXBGeBNVV/tz6NfS4/UgpTgAuTzFrYvAXeyOFSv
kD8hdDHFgGj8aAKiSpKZzMH+etHRLiSBke5OthP5IZF/AWnt3j+PbOH33KK40rA32DUHdDBOUw39
IbClfPOCriG84vJna1ol5HyhJO+vFG+kcv32pTMUjCCwECmsHlbhXA51E4/Hjb4ximxTN3QQFezh
IJQVl7mtueA7tyst4KpTkFZjBXEhjBaxez1rvTVw2tL7apkihqw6L/QyX0T+rI3Szm1XjHC6/6vk
sf+RSDgCQgOESD7PmNc3VBafm5imvCNENovGakLrbebRPxREbzhjmZEcgSu2zVx9CBmPp65O+t3S
yoor7rjAjCVLbhzCbfvaKjzC+KDVqUfzV/7Y2LhqHyMFvL0iUaN6MDhNinlCaqaeXU6f+xZxZh2M
yBZCn/R+RN46e9F1P2Em2zKiMcoCo/LuDiTZH4uezOpW8E5DuSwssA1c+UGI6sfrwgLptdY0p51A
6/zJH4AxCm6FIE3e7cmsn7nPsbdJN2a6orCcbbwH0jRGpiQ8ue9Hu8vlV5dwV1R10rnnO23EXelD
cF/X4H8D1D/2z4NyGf3mezguABVR2vIVkR5lD34IN50sTffP4d48zjZlS64SpYZqIKOZRPx8sKmj
svVlUjjlKimTWHiaTjDADrpUpH3Hbd9/YiR5OuJZ338fAnij5BY2wKiXUDtOOCcAX5wIF8JGbcHx
FTxAu9a52Wyh+/T1sI637ZkLY5+8RDiIvT/RW5GEddVshErHR1WFm5YKPUi5CwMSmr5SQhxeCu8E
HCUyHJa6H6rhb352rla/013GJA1E1sGaHTZIlyjYaUc/C3Cr0MIvJ7Rn/oaTobSEHdg9lvCpDAEM
AqS/tnzHI3EI83a54dJWZU2HTyAcnW1v8iZlw8ADWpjHD0PG80l530U/GwrBkWN69o3pSEQkZBlD
Xq7La09HnE2saHFo0jAdYrzXNlT4j/LiKjXYzjr9LwgbZWTRTLtxxir8DJ3hptfuV8nov9gwh9kM
eP2YB0m4Y8+tFLf3hjN5tQVn8fExDLmrNlFP89OxVzjlIlTDWkaey6EIeTIPAkaI633I1ypXq3Fh
KfamlL6LEFaoWBhColVqkF7ZXlhKkTGBvJz3QC1xdeJUQfttIjioVXGkYelfXNnH9xErChW4J8nz
Qu7h00bx7QaIM4R6l0kkscTM81VKgpHRlc4UgPWGa312xuwVoFkR+uCnM8TaiNc7V/Iye5kciqVp
JlT+V/zTmcNmQB6astL89d/uI8EAhnL7eFMFSEWpj+scx22s+4UAbn61ynIUHbZ6kZeYB9V2GmmN
nvvxnTc/JjbIFoEadPbEw5rzd5bzTZNuX13R0Cvj/b/BTFKZAzmAZ+0SZI86yCEFWrdrxzvNwQzH
L+dnec93xbdOrrDsdOa7SnA4/gYUm5iZCz+vtFUsBcN6Pr0TylBvxeTtdK/rkTJB5/cmivvE2T8i
pnsDIxf5SMGoiNVWGzk3tpJ52h4nnPrqHOSdSFFGEtAaDhaBPVXikSNJC1+wnF+woQAHhFh4ZZRG
bOH5m+iPTP0mRINAh1AVk5NrIHvy4A5lmSrrtDKfdhNMzJ2Qyd5yyMZnL3MxJMhOXvF5S4BNKQfh
tUR9KJnxFE1uBiY+rvq+cNKgWn3BGfyEAkBBE7cg+7g3itRXC/K7M6nIU7ZDNGfrv0takvFIvA1x
AuNOJAjYMEb5Gy7HPe7O2Hz5Sco7tTSwArAJ4A/XPfQjlg2j1biGLWZtRDN11tOgH2G8LPxNO+mz
BYfL3RPRres96SljoIK4XBoxhNjx/WsCoceYPhI26qxuSSg7LyraSV44aNN+Qjp/SmHaEO27DBSY
Lu2OkOXBtzosTmTzsq2NASOsJEbA43yKbwNF3Hs6wQGfaLRBc1subXmvgDKpKVBEkvYuZzocIwQr
IIVqOUEpjWzJkWPkVSTDOeooBMDehr5FQkoBrJ29qQzb4LSP5SmLKgHlAuSXDJvJ/wci++88nU34
ZjDN88UQgFh3oClUCqGiQpwg9fbq7mffmsrbsAe+h1S8/D600duf6CrPjE51bFjbgjOMrpIdsgep
1yoQyORyyUjhauZ5Cyb5psQ2uuPWIBIfagFA6WwJ9los9glGtsqyIffBVjcxukneJmpVUsnkE3Am
K4LOZBzQiVHOjSUgbx+iBLyVRXQnvP4ald5i9qBRqCtnERFY6o+gn2dOcISxrp+0oDPYM31adnO4
egKiVTw8eSY0QAM/MESp+p+Sxyj0VCZcY0CwUu2n0QHrZkjXr9V17et4iDAn/JNCQ2n9qOd9c8cK
ovUdPx44dnJugoyl7rS1G9yi8fKuQGvzFAh9rwi5biAG/GFYgVqmTzMGUc8oei+lnnA3LEraeYaL
krYaT8SVP5rk/d0nNqnS1z8uwoH+4bqYgDElbr2l2orBGTxAhSsoM6JgCb6fZt0j4cs1NudamRG7
XThnn0hAaCcQc1dyoNl6JZFaI8ICabCchUdJYC8popSQhJC7L0YClZwdL7hTO+PuSf8RZaAKu00X
OCMVSl2H5sA/ITfG7ILSSaoiqJk4XdUOe9FiIlu4PEdUpi/rQ1qq3+TfwdVS4jRPBhHQi0VQHBuc
/F458n7PhpNUpuy7ecPNgTZOCg4pUS+YJAo9qAsUZkFa8O5L3MGVZ1AC3YNa90olo6yEnio6ziXs
d41Qyyl7hLm4sd2PmXBFRkBbONwSwSadLThg6GeBWXvVpFOmNlkLuZSuLgXGWKQHrczZHpHPTMB9
QG89g6Jz1N1IE29H6onaTlvLvhI60UosueX/Cr0dw65m2XBoX0gzJC3aBE74LqZVpgGhTBrNrGDU
4koNG13qXirHtynRlmS3mgOMayvhfbcOsqKadMMrNQGwCkBvy8ehr3H8JeBuUnc+n/JzDL+9B3bp
cb4gxPvC5nEuDRSRwtRWaf/mxgHAdQIoiowggkmIjClnuQB35niELoO8Q7aBhraJbDv1afQ985xB
XvS+oncgGDUTQb+OQ6KIvDslD7AY5qiof+O68KdNxMp/C9bIQQ1TSQqwKvBV80NIFmxBWRj53AAN
8qsysMpEmIad1uscNJvCqQ4ikGDSzrCDoXtthWBTIjSl4iVdjknzpFTGZqr+yUoy24XBAeBC/w8P
xrTdMTJiiwqGHxYMKmLyRt4eVXi1rIHTV5Ku23egPWKFSZiDKcxZ3K64mqACR8ObWX06S2cCm42z
xotZGR2GdZWIroikDKMt74OkcQafqQTlmvNmOxaVz3Z6cc+dVLtDS0ljK+QdtqClKcH/0Gqel20C
8lb4J7FMRGtpWvDT795/jvwZcBa6kl/HiaWmbMU4tsq6Q7XCkwLrpSd2zKvaGCrFVM+H7IHSrASe
M1/4olc32eRcxphM9nUY5Tzx8Otb4xUEfocwn6UFAxH+OM0M14aKrfieskGV5SWPkaOyIJ6FoY8H
nFTazAX8kUimcZSUAQL4hj9SQLDJxM9F0iA7Ae57eosVmqp5QegmhARRHjqAYuszG4f9UG0U0ST7
RY2IWQOR+5VU8zzAGaNb2WgrkCkVzIUXJtz9wh1ADdVxIdDoJbpWtkNjF100KPDpCrU4ip/5SbbI
odLlB7CiU+PkzLyoAD48SEXHL1BVVYaQ0NjYBQYH3AeZeHaFwbd20TRvHqbb5MYec/ghMoqFNdtN
bgmg5ZhIHHYlkq11PRplcmv8bf/6+GHMNp2QwkAHspyNogWgRtIBs5XT61xvZ7/cOQ61DIlIRna3
MBsWXwLRTpOTiJFhHA9vguriVlPs1OJPG79JZWn7E0FiWoczXQkaKNa7HJ4SYJb26oxZaeoAm/TQ
did0GSdPyLhW0Q/M8/BnxYK1YwecVWJHyr0fDs+EV+jRttYj22BdZmw34RaYGLuF/cmnPwonYk95
5JSu+9KcxLoBc1DmtDQ6iQsjk6FRRdgbNS+UvsqG/Et+LOJ9eDqxQo1GSj/PL217GndzhH/CAPv2
rkp6fqCG77MTddDcl1TnFzjwJnm6Chn0dd3KlpRa1eLyylEP758x/0rI3BsoY6H+4Dwfwv36Tatz
BRHlv+BeeoQkx1ya7fJXlU4Md8vzHjgM0KnMQN3qqtr278rWVwbGOW+eeUEjLf2XB4By/bIAnuTt
f+di3IaVc5VWSuoP6IUfX8xoNJoRvSVbgXHfmHKCj1HdbeuwOEwpOqj2ts3TxeQj5D8JfdxwgNKO
NkHFmrO59aZIu/Y0zD+Gcn4ecI9cQpDwoL0D4A7g/AxSSlIj33dnrhkRexzs+SEXm/F58haj5May
eM8PbpaRJfeFoI7Dh6HFrgiODQXHHZAGmGkzRMusMJ9RZWOlXcWk6jnhcHH5xT6R3GT8WXtZKb9O
VrO7Ob5VPc/uBX4CDxNxsoctCb3QsByIwSSBrTw9X0HDRGspkdXUuXUE9dijbKU6NanDNPFXNFRM
3B+KbYGxPFM0aekF33Hwoe6KNjrSaMmCT5RuQuc4/FzCjDB4+6SvHFnBtIz2Vm5uXOQsaiEKXEan
HsJT7WCSDHTNTr82pqAWBHnKEtqDwGrGEL7TGHkeOt2+I/3WfVDCt2rhX1XP1Wz+gfGDlKa0e1df
503kWdgwRr5LZwEVy6UkUwciWNBayCLIKXGpulhXgzcLTHyMsKFNUfAUSxZMj6Acbt6MAmUx2NxQ
v+GYz3j1UfofEj77iq9cmKdz39AASDn6/x33ycKjWm4zAOSIPg0vKDZRIslAs27vazy8OjejP6YQ
MHqNGlEeqAFMOvQSlxH1GK6qYKrSYG8/fI28MWTSFa03UblZfTCAkDfHyNd3VcKaRh45DN3aeWT+
tIv121YqjjX6NyUAKljlZiYxdYM465jFdJP3+vnJoduGxo7pDigG6cO7imXrC88WF+nrT5bS3bZP
6hBP4X+yXxSF2hDYih6CpnyDC4J4mYTQ3kfhSfWvRRpiIDkL+LRgwz3GB5WdgK95pb3IrhJpJBGu
nu7NdueXDqHY1etKgwov52ak6/AHx6WrBWM0/CNosrQCnKGblAD7GRS0tuB4hl9MuTq3QRN20fxe
9RHtm+EUJ7EdJqbDSSffdnnllRF2Tt4NYBDYMMX2cLE5O/EblhlWljJ53EWKmYa+3pTkO47mJR8r
S6O0Qr6tFjFeVWQRgZ3IRqzcUk7X4tBdJys7z+u41F/Rv4uo4AmsGKeZPVbdWPazaLOxufzMXxxR
Iuif1aezWCnF2bioBMSyGie8UwZMw3KX5HQaI6YqLWbi7+N1y0p1BuMg+rSxuzPe42lMZbfrU0p+
EJe2aY03YOaPijojY0w3ciiYgS9hQ5yetkDCLvEMEmWahpf88pJnr0LIYyq8HPuiRzHA5QHs2aWO
cb37KIMMz1GLvnM5MEHQYTKjQDkVDsRIY7nVF5PgH8ncUtKVUZr8kow7tICmw2S10dHlgt2/0ydB
b5dx+VFcVAUP2CX8zJTSINrv4VUbVKOWN1iV0KiRsFyESWXZaPLSB2OsksOy0KeVU6ezZVG1WGch
Q4fBeik2S5RA+K0f2ADz/7B+S3NdL1a04T6mltM02GVyHPTgDN6tlRO4FNRCNKlpSAnnOq2FlrP2
DtIk3WJGLqfBjZfCtLxRjdTlJxz+m8L7hPUmF44UIR3UeR37INn8qIm5+i7tBHcRRIKCLODgbtlN
GcOUUtyiF8/pHLVLBtZ3BiSGkhzXHhW2fzs4Eo8mebbjR+xXaf1GRgqw4j9WfHeQHIwXJMQagJuL
um2qdQ3eciXx8njJaamzGDPRJ/PnSGvly7mppfgrxAfdbkg8U4P94a4Dobu1X17WdJpTLybc5HbI
SyItTmtD/LEV8ibbEQNqJPMy278MYXxwqnWXseEIfhkM1QM+ueN22MjTFEF4qQICd/yNdW+Jdqy7
35wgNRFFvws1C28NYvGd1r/SQMSbY/VKm2lFjWCqCj3tCWO3BUukg/osqYW1luCeo9GXiVPxssEs
cA5dEH3yC41ZgUxo3YQzPZERmlCEvK1uUb5sq0R2uo+FQ8aO8qkEyTrrhicFmkDdP98wnx096kiB
Gmhk3SLKiTq6T0wc5PirRCsJFEhQwIVo9sR0Hj+0P6XlRwED7586GqtWAbWZ+SWOdKUS5aCLc4oB
QHA6OIJhznA8kywW7c7b/6rMbrDeUU//x3KSbrgGdIADdOk5sfn7qG09nc6nGQFGLCanh2LFzxPh
opKqC15eG/VXnz8AjzGwmpWsCpv+AhQE3U8ST/HQyaYjBZvKLLrkjvq0im9sSVPmGE54U4Zkh8Pf
rbPIXBbm09IhF+jsat0NR/nnNWGw1WPRzdMDh82218bbTZSw6lwTNwGx9oW8txXoNK+9Mx4AKLow
tMzbMDBgvL1qeOHEf+Gp2liEefxmklJLm4vC8FZGpSgKwpoiZL03wsSltOLX5NqXKwjP70mpX2TK
Vmvmb+QEK6DeRN52DC+VxipT0Oluvb9nLvnr+mfGQ6qd9Tg3v+9iDPW77TOcjYOkB9KII5fk8T5h
Gfk9zrES/ZNUbmh8zr3gA88VzFltd+xYStYfr7J9+2MqR85w/J/ZkdyoYATCvLH1T5RWt4nlA1HS
aNmaZX/xX6yrEkUEkoKmWfrUda/DFL2WDcfZSS2rTo71uw0vcL3UB5DuEXKuj9wNcKRHTd+3ivxE
mLBye7qRYeZRQODr63F0+4b+HweuR26OF/uac8H5GYdPE9jKKD8aCKsgwNpnnZmJuaRZ89UvTIAE
iTmJ38SlAxCvC4it3aIlNo3UTnqrdXVKJdRAwg9zKjD+goRY/aRP1F9QvHnDm1LxvBRaOGkv22a1
pkF7SeHBpj0+PXR6SoXTVwDKveKbfsE30j7bLS3V2MKaoIle69xG1YadpCnb44NBvoUxiQ1qwqqN
pAJ2mc+Ys0H1HIB1teTv6nEN/7Kw7P11BG5qlRft3VEuJ138Yw5GGj9HqEzk5e/8OoZf9iCIT1A5
DG0v5vDRPSQ7vJx9u2zVbRSHZuItAfGB0KsDfus4MVR654BMHnPHm0aMQNRIAMBW7RlIBWmRtjHB
5DTSU+8tDJ2Ekl9UhUd4dZP64uAxRBJOxYnuvKX2ovVp9MF9XkU1adPYU01XAUgWR5rq7tPnWLix
dTVSxcEUs1k6NMy+XzGy9GbWuTfT9XjIaRXHMeQ8WXVrpwu2qmIA3XrD75FZw/wEkX8ux8bkRjAS
PHwbHjy7QcaMwsqRh9qBgCFGByLHRqX/Wt5Qw47imcI2lBuqgQNXXaf4QLBtg/VNwRca74Uwzpn+
t2G9DVpxscD89GwOGrsBKmGHlsz5yyVy2PY9zITQsQjNcntnr9EHdwuLsrxd0RfRTwVgOPx1Clx8
JPmHtaiKKQDV94+j1AIeAs6MJp0QKVtynYHK/ymjZjjW8/KqK854lnbdf6l/Pw2lAcPm9oJEYCqD
eJib2Gb3Ys9dNLnEkKQHq1XF/aGfo29KEgbn7dOWHcBN5IUKTVfcNmcAN4vEC/byykkoJ4t05UvG
A/fffJlta6VWhjnwmK5BpQBSCv+lYcLbUcD9GkshGwoAcWKKlk+GbBMitBJAuYWXNuY1JpQDn8YZ
xw6vx+wDkjynz3TyB68OQGdjEIGdYjEgNHWXIid+6yJHg8cvTX4I8/g2ydIHMVfO65UyC9BHSHE7
pqvxQ4Y2zMa8t7jO7Jj32GrU7gOiLXTq6QAk7i/cljt/goU8ztxiM/OGIIjvkLlkV7mqg0VgeUU5
Mc30vxZJzlOw/zOmFCpvtAOkg4YCEPDUC5994RfJyc5D6neyZx4d+Cc+7dqa6HFtZCc3NUMGnCHv
7y5fkvhsvfgKtLZD6kH45WB+HQLZtUys1fuNAjgK3WNhTnROSzz81evFDsyt8x4nW1kZiSAdCwwT
R4rtaTyO/4Uwp+B8e6wMr4UCn3kCy2cy98soxMCDYQUyjrabmFoMRcOn/+NRN+YeOYz+AbImUuvB
FATp6hu+ootQn6xG0YfpIOjOc+aTYSucFH+fZ8ju5kaeG8MQEN6xN4IHOAPoO9J9N6VgO+ePgTZf
sPkwHNwZM+kBFnsDvQn4R0FbrF5QB01a82nkW2/GYAoGGXg+GN4PPSoH/e5KhXFCFJrFDnbNaf+I
BoQfQRUhWXPMA1df7iNL9jqvS1JSW0ipL+ON9M5/g8E27wMqUESCnHdPrgTIvYkqJ6s1PCz1GgRT
klNwwcY1pCTCgiuEk37xTqg77RC+L1Esq5o24AirzfMDM1YU0yxvrN07N9KxpdbBamDekUE/Dvfb
T5BurNhou5pn+GDoVS83mjqB2mgqdkU8Kgyn1TS8zWZ8JOYYFqr6M0mzWOwdnnutxUW4J4le7Vjn
0xdXYyMaDC158TtjA2SdO+d0mC9DFRp5eonpg39Nv3xu7XX+MUlncXO1jLkirlcJ0jJHNLrpiAzv
jCvIVhU4IY3K5hKoZAqOv3ReyyshCmY6hSvW6lUYufk18wFlkhu6ukdXf6arqXgDH67yqQpNXvFH
EvJIjuDvFn04VcSNE5XACuPjyEAgn/p2Ia6jRk6Vm+wpaMHGY9QJkxVCLWKLruKRJCR/JY3Hmihg
FWDsDKX6i1hTVyk+K9ira/+999DT6wIfkC3FkrUW49WOEmoxZI1BzL45AdEs/B0PgkSflE7ukhXv
1cdHfgcUgIoSlz7UD2KE9W2rT9uS8nA8LEjbQ7DdEeVE6OG7yDVBCTR6xSjEO5I90jPsvgV7H/tg
DtzpTvMZqgGr2WCxNgNMyN2mVkWMpgrWzzs5U7TFrdIyKiovOT+8IkcoiG3mivneY3o9h20vLqAH
mU97yprPgO+/nHVwi6RmhSHRjIosJHI/H4es2PO/CZolqho5AuFRe87gCAJfkc0CDN0R8iEPWcW2
dt6/MofV2U8+ZTu/rnMdWH1TNMvdQqgBx0Ho70pyERCIL5vD5ZBwR/IKy91FokwH6+4SrjWtmUfy
dJIgSlqa9fIi/4S/qp7kLGnEMZqs2C9PFcRvxPothbv9fo0JcsG2Bdt4Jwy+ZoMbmD3Y9dTjoUuV
1EgkhD1n1S2HRAKeMbnn/FCreFUMdLaoadxz/emgmD5prmQt+L9u5gBViNRFYFCvTLFPQbUUsdPD
R9Chfph/Wr8fyLMxAKosZTq5e9xKSu/jspM78WUdzMNxHlcxq4u00ZaApaRmR7fw8uG7adpvyp+H
42OLuFTyAe9JIJzfkcdZk6TbvYZoxHW2cAnyy4IJzU/zeCNTVMoHuH01ByexU12ffigNQyj8lRrN
6ywGbJZJgTmfl0wA3eOKBLwWCRc3aCmrlx4h2Ll9nm7NqGddMHTiPvbDKx9ecsonUbtEF6HuS0ax
g0lvJI1LL0Zyr7aMdefeKxq3iXv3s/rubfCrdFzNBpSz2hf6XAO4er29Zwu3VFnWZrJ+3r44M4qe
m16V+SXchyFA8f4N5lBN3kMJtj96Ymot70xjFS9uugLL1vnBEr3Xuu7QXgsBa1kZsZ0NT/48UW1v
tm1pJJNWJw2t3ni0mnnoJ07gMXw+/KHTRu40dwOp4YnpZ/Df2TFxZ82rKDrVUtuHIJvuhMqsM64N
dQHKjX7dZ0RGSjdJ3h94hw9ClEfB4icgxAbZtTvG1TiYEPcfbTIaecSpRT9c38Dwo/3u9xKDzjX3
9yJDfEKtjHihIWzOL0XC0WN1t8SQLV4zIe99XxJpxRGO/oJlV8nZRCZidA21Ke4HdvFI197m8erR
m4Ea10PXCbSja0x+kghkbMSBFLrFTo6xG3kNeePHIjgY2Y3ENpHj3e+mmPMIH1CXXvsr5XCu74Cx
wsbmn7H3XIGypGbICuBmfej5BF+KzG3Bb4INs5GA2DHll4oiwkkrcCndRnG7iVlNA3exAvpweIu0
ggnU4mWOzcYf+vj3PREMCsVbaq7KT00vUNz+8m5KfN9am0J1WgJpfwydjZmmbCwQcl7NAVv6OFlO
RWxYYV6XeC2mw3sF254LYUKEpIOWIJANbW3n/g5rlFVqeOcBgfj7TLUVU+SLVnMSGBeQxMfR01EY
Qsj9mlWBQgF2oaa35x6C6jW0IbsKLh4t6GRfHGa10ZiF8oOuWb8MywXi0abSRBJSF+yB0U80BngY
wslQ0cO4rppW3gNk3yy026glDIrMN6ehCUcYDYgqis8jBDxObhPutUO/LdxxRnMGs0U25pzH0Oik
RmvGjBhISAhjrMTv2BiMyi2tKpqmT0SK68hTVnne8Ro8pfaoQWOiEJ/aiu3gV7i11oj56wPlgGWr
YUZp1svkia0icsmyEb7ykE3KYSrFruoPj9R4RJxevAXFpKodoOYg1o0zMEdOi+j6lfi/MNCQu6XK
9IrvZXknNIno7FGyWHAxFM7U5UqaCWNfKchGHL7iMJYT0/g1wIczN+EjEnsMGRbYmGAHBQEiyv52
0mYpjqxnxvUxbgkkvU11gMrybAJEuV3SHbs/Dv8iS7wsCyWHUomZis02vRFhJSg5vrMyvjg0wm8Z
++ZINlgyN8ly39mC2/E4D80PhjctEYUU4jQFdJ9i1r5bGvI3MBQIJXh1oOq8T4j84qslGKZxqJYm
tII1sQnBRvkfLnhEPgZVHEAJjNbhp7y14Uz/gV+ta1yC7ybPofxTH+SLWMn/Ch4TZI0W14tqG/jt
xUx7uK4RbWe+eW7HroFmQbNksbtQH7o5Z2cTEwNbtv3T4URV3Kf7zLyARjurPFDM51JREFDxwDyd
nkTG4+MHqo8nfXctUgVEtstNLcUqbOAlzhnrFsKDtVxnX42GjguPTjvgZuUNE/6pgicGMWILTTok
iOgBv2r5s3jF8ebGg9M0dSKgHwJsQBpJFgHJL7U/ABUAzUgpMhq2yt97daFi+Dke6zYSV5neD493
WJaF/y7q88w7Y16cD0BMo+t/KAL63PUtI7BZBgPS5/L3iSTADAuGi4QyPtkFDN5ILy8c2PF2mh1h
GY6JehmnZVPQOPGiZyc7d+ONbQtmZ5pUOs2jGNiMBCYjaxVQyhH64Yx+60TrMbNhVaJMsnF8fSmZ
q5RjS0CHrCsMYCcOMPPq9397DkENi0SngeGpEoySQOME/fiN77dKRjMMDWvX5SZZFg+mQaHyq6X+
oi8XOXY+bkqzWsdIu33i9B2q9XCOhqCbyCmuhTYr2T2kUyM3ZHxmoERN9vKXh2FK2VnF8k5faN2T
R9JPlr2uVhghraFCj0FDyMfAGeFrQYzrszM0r8DwWa8pbWbWNI+yXzA/TZZRZ8BOX8A6OSQ43sKr
hwmg+U91nZhZfa+uDBMOs2I+oFu8pJr43fqDQojQNY6mVZ4cw5SMWgKEoHvJTGhgAozml/TJrJnA
EsFVbeK5KicNUyV9NCupOIxUQ8KCOODqzNvBm/8YuObWHnLQ2WV+Ib9AUgQU2vNXl27lGhj4D/hi
n+D2FqrZKhwTYL1PfUbES3HWoTrbTSQdUA/BlnalyKhMO+6CTGVi9ccwY4zPksM0T8t2lLxZroR2
iIEPzwvk0z+iXWd22qePAyjmwgQbqeS9dGnnALRsiXfXo3tOHoh48bZCBY6MzNLWmmhY2MZOrHDr
4c3SM6lRma1W0N8tk+cbccohpefp5ouLBKZwS9hG+X0ae9SRCGjnN8RH3I79SY4NYj3PZ/1wFWkp
81YUHRj2SXKWvGtnCJQYI3b1A2BAX4pM9DC3SNHbAqqxFUezWwmdzYmI7Kk2dvhXg/uHb+zMSaFR
XmB/Y7qAmRgphdthbsWB89YSb7aeYbXKavFgJCYQYVFuOZj9Wh9/GhO1ztdmrBaZtJaiOQ4gEYr3
RE1I21PCeCBzDd7CZlvqViH9qKDVgWvd36h07m1Al20iyTl8OVoryyAbBivuXqmGjgFNvxr+EUGo
PO8uep5Evn/OgsxYBfPV2TfNBhULFzO7yeo2gpJ7Ky8cslsI2N2LN/cxuvjVY0oQDqVd+N0acLFG
TjSnKOvuxyZp0J+lK0HABOIEK42gW1ZPO8XXO/VRATYQtKKhFiiymPUCbg/m8uHommS1EpClk0tu
o4fsLSZM3L3+2iD1P9j86nmt+zJSw3rQqYcuK/y93iZqgfD/wnjGQKzRkERfbZI6foq1iRFuAOmB
Dj++/4A+AjcWZCDEAp10rMzX2rOBqMW6eo/Ck/hHyp3MI60A1xE9N/TZlTjZ2DP1wuNIXOnhU+0+
CtMRKjqdd/OYLoTLX6pH+kSLMLIZ3ZzYm0OZS5ua41YTbQxbsQCIrvt84VKf3pJnNPwZuvD/iAPb
xL4kt7Ms80PLRROUZGWXigf8ygnK60WjvwNQKSGnhzD8GkSSb10kjw3p51uj2wn0WA68yjtlgk/l
AEDajjBc7iEVI/Cd0OciKNbH/WO2V1Sg7jg7PFfp/GDJj+Fc6in2vfvS/p26LKXJRI6AFMfyk1/E
mfP3Uky4S8hcQPUazT7h/yaVSE6ZEd5LmL5Vmln/cA7O3I/2vvWN0KnpWWK3shdpRgwDgXFA2Z4U
JFmP1G/oFd+69q9I0XIv2jtg3g5q1GCFwj13ItKzGKQL6CnVDlZLcoAgRlZcvt3aj2WbdJ9j1tKp
oU+hTvqyGJVvRhsNkiVsyOvbu7NE9E6uVjEJkP+GXjKGB6eVJn/fDN8hjeOwQXSSemW61ZL2HNll
jL7h8f4MEheYiHK5V2ygBuG/HqdIIx4uuuBlZDem1KA4AvPktsoX9QrKcVRFb0pDdHbsCQcLtHNp
GrQVkCF+TRXwI8PSTYXW43+gBxbrYzFye3avusePXSNaeOBIxTo7JCxktwgExAt3jzvJG3oMfPKM
z81oHVOmhYjvuX/J8gi6vzRAg46j44n5vyWHPTf3uKzFzKZUQ3al3iWQk+qLw+C9umg7PBSW3EOq
gRbnJWan0E2yxeZnMOSJtBPa+PWyXycKii1/RuUoi5KoIm72ysuItAB99XSD2BvtWirCC6c1mJTO
ibAeLKmurtgPjn00kj8X39H8zwTnX8jPI4Vp0+ESO5+i8ziB9N9tOUtM31kQAyB9sWx79AwT15ln
LAEoNC51Pl27IaDGwI1wCdcJR/MHUUrYiKFV1dvfJzw5endf9bzp7TpGdPnq4ifuXJf33S9x2UFL
dnQI7DfoLVO5Ws1ERsk+pTDN3fmjPmrb0BxxqwdwsjHU0hSCbItyPlJYBTCBkglIeGgSFRhuboc3
cLlgvz6R/ddyZ+N2l0eCInuQKjrM4/yPawSth7FdsjabjxAAeowLNaQMOHrkD+kjTB8xSI8Q26Uf
XrffRAB16x+xdPzEJIUvLysIWDPRq29S5IDJw4D5NwD7PPvg6axVsxnScNOerraiB23uxRtqxHIP
Kgxlm71C/5atrf7R3Qk/z/+v+3oz5Dit/f98n5/sITojFnrjZ34HPXA2uSeNVFpKNKXsAMZIOEWI
MJkBJwPfJgWbJn0fvu8cYLWEhTQCpqGRjni8jKJtvF2mSpI5cs/W4vMhKGhLV0b8vrLRC4Eo00dD
lGcZ3OApdSKnW7FG4HAGhIGNcJV1FkV+guM2bz1mVJZajEHDrVRW9kP75o6rUZMSHNAYAl3GPjJl
hIurps+AmZx5+aHa2vzM3Xmdb4sKaA8PvNMFOcoDf1nS00K7Jr6+eB6JYlBKFmZFrKlQcBzXoViD
cL4Zewy+4+NVWIvRLjxBPHXTx3sYlTYLX10qbwaxEt5/9JVncuE35kJJyD9Wg3at9rwGIodyUJrR
EBxx55+7a5IwYnZjiKz6R4tOw15DRJY6UrCm9YG35l24omYXmFnmUkICctgslKNMrdwpHoo8hwG7
526pHMwnEWIseupZOefDAs/m7gpg0PWNiBSeGkNbNN7yNyymsC2nnSrqtL46EQmZat0GhrMTA65U
plDEicl9ImAG2g0zNotsG4pIH+uk+MZpcdZ2GPQ4vC1cSIi7WvPlakZ5iOKGyjCkDuk/gGj9xmVH
LtN7MWmwt4kmhWtpXrXhvlYUknrBaE7/xrVGwHj8a77N+nxhfIHas5/ofl3vU0zQcGSMG83f+kLz
CemDz5jXcMloAhcl/Gl0No1sjR/iky2if6DF5Wv4MV6/xVQR28BAr+x8B7QjLH8evksp0aeh+9eq
bSp3PFoPRsTSOIcO9Rk8HpMfT+r0LIYjzsyf7ic3QwHBLQeRas2XvtJtc2DATW46di17KTFoEV01
4BQR5Z/Q25l0kTqDkHEURTO1RJgKoOC9yvYeGSfb+XGLumCoCx4cfJuzSKfkwxRJLCLIJ+UFiMne
n0a0MKX+n8NKU8MOh5EiBTOMgq2sd6WWtYhCUddcxS2YEupjHTmYZrDsfA6qSspLXPW4qxDzPisp
SAA+IrsUz9+wPWSbn8Wd00Lc1qD1Bl5Oxkw78YBf+5ZF7K2ZqYlTm9My7y2c/T5Z6SMhGfQYRHwN
2t8nqItgi+Ob7j5ODs7hXit8H8qf3LDqvI1pNWX/z0GFQJ24eUSCjCtFG0xjsFWZcSEu+6q9gMwv
SbobOVOQl4zfKRmBkwMV/qKPua2tj0IZRZlNOero7w87cJVCAY/yAq1y23UYh1uwSw3gavifNcq1
HK778YHsK7nOPIhT0NnK2nOokI1uWhKHVm9ohVyiMD7QgTiP8Mz+z6A7nFPTPwNuATJJspgyxt4a
wjzj51zyMDTL5xjEanyprbLNkGFxw7/WE6G2yEH4UIWJekkuCP0oMN22kZJ/t7T81DoBwKEEWAfV
PSbakXSnCAkTP0PEwiiiS1liZVGf5Ty9LTb8ZWlCd9lVLcU/eAbHB9Hbu/dsU6Pik/OacSCbYHk7
znvZZMhNKpeGY8W+7URAZ86P7+YEq9iEETJs47fYRsGzRyDe3kNQLmgjY9beLiGOLFy8/iMiiTrq
fG7yoWTikP0W8TDASvGIMzr18qwYK5Fw6GnUXTpluyAzV10X9nFhGBRBNjE22wbA6Jo9aMq0nvHj
uLOmjTl2D38CdTO8ioSKQ9iS6bFU0UtxDeQfSMB00thrtBGHsWBc2Myqi77xP9xVw5oeXGf3Bf0l
YFAlXdSfdJxuLbkN6UE+/UbqYM+QUmfuKAV16HwmNlnw5dAIsRB5iZSnjeZfSDpUZYwTtIa31pUO
qlxdnyPlbzaX1pybbMGOzR9J0E2zMyW7nAQtSdC5L7gYKXuPXHqJa/obvdj88xMUfpXGt2YXuUaa
STTzOyfRBva0+rS5arrW01lNSORgcUmKOQX4SYqZHbmPf9ArtBEe7ruFNNCwrDglDvanFeED9ce5
KEE7yXki+ZAZPEbxLv4Vs31kKB5xmI2e+rbt5HbxLGqghIluFVXtnG/mjuywhI7jh7caanmA2Rxk
WyAifpDxgwXtjqBSSSwvK8R7sfYR182uXPXLDACsmRjB03pORBnL64XpZzWeYo4/RtU2cNXA5xtu
rAJ2gh5kLsQ9fCAXvyn183VFaEeyUnaiNvIhC/DFqlPDCgyDTdg0uuNQz1Ul2QroobC7gGUH9OJw
k84QCIAlIl3YfzS9UJlvh3er8+qqKg6Y6H3wrer9j5EqZJelKuU2Mr+W1AQHrbj5Um8e9yexu8kI
WJnU+VMiShHANT3hyaNHYXTTPlSe9lsWV3I4b6oJDr+/K+AMaIquDmOvpwlU6mcmxFBxeVO9Yfqw
IPzOG38GYvPyZwJUN/J894uvcznGlk3Bh9oEWr9NVkXe9Y/loQ2r5+OtO5ZwNmFQGPSPb1wxyam4
9GE/xJwiBcIyufeHNbEVADzoD82HblQFBUbVYIEZyNrZT8UD+vDtAYEkCv6VXbTPhysNURKy/thl
LFBeVUeIn3TZPX4fZTGo+Lb91P0PVvjvRsU8Cxux+E8qm+m0s5h2CkEJKXptayZ3boYdz3iZGboU
Kdz9Pet4TzW+EZJb6LYJKBFQ2+w/2dUdTh+509PrMXM7c5kULN4pqHa34aM19rBIcDuDHHW0roih
hC/IA2HwrRSfBvQAMJHRf2N9FdLTUVxRputP0F1w3pAc6DIy21pLdWqOa2iq8PkUtXfuuE5ycdPW
V5gfnO0NGujvWOPR4fhPje2fdFcpsZdxyOYcuGOKEV3m8sTzlK2BYiSavWFioqnEyg1VsU0CXxM5
VFct8Fl9tfd23HF4qH6ALbUdA20OiYOQZZowdg7cYdoVVpS3iaqd8cAHKwmbTnKkg4Xz0CJY+HTP
h3+dNWKlth0F+0JUTTOOwaPQxaGaO0X14SV4AThn/JvJqVtqmt5FyTBlb3EIyS7+264hQzPGqXQi
LiTaEnizg64368wDijneuxRta6XuhQSClSE+hWGPEc0sjNDdNmeKWwq7mW5uzQ76uGjhbMzvV3Og
iQUVle3xE7/BI5siBEe5TKfLrAK+9qUluafQjlIxK6/89fGQtDlJ+Sk7ouFrNUHT25VpQQomOWgQ
Y/6LuZajxtAYU5CGWWgmdKtQb9C4qUi4S6EmUY3MRl+OWNx1GGUjXAqecmyLTLrDghL8bt3KHvqW
+9q074xfg6PNMqd9+LbWodk+CkUhIU7sv0jfuAuEJwu0TLdshnX3o31aoD7JgzwB51QH5RNtBBqP
l3GVYNv/92hwBZXVBn2477dMzxYjqA+hliMlz1FQsC2UDP4kT3w1L5TUNKIQfKP69Kz1rrIIrSVN
5BXUEne+MWttX4Sz4OUcxMXsyfRbQ0Z1jKLGLBkkRqRpRgrJWRfZLFR/1pFhcIoWrah+F+1rxqJo
NliNTrZ/nMzOBRmBvAIuwimKjGt5ztY5X18X0RtFzEcpw4Juzd7eEB9wkJ+IBbl6DrDpqKOzqmpo
y0FYqZKfQGkxzaJbUkmTS6n3/Mr+wj3MQeiP4fKMkfobgu+htyIwC+ayfDdf7emNWWb6aBBFi9+B
bboE0hF6LMxlxVj8pZgRCdETgPtkrcIn12zuD+3Z5VRypEfU8NNiMOWeHrWBWqDP1cCfgJRuGVxq
ZxdTeXKVcqiqRwkNw5ZFEHIsBjd/Fsr18bzpBftyIn0AN2sko6C6ovEO+oFDbWvlQPRc3tC9yjqJ
qGpn05mqCpZ2lvhg4jp2xxvBtQy+OKSxr4ad0yjLIguxOYw1jLrjZwv6m6UA9jGeMY90mC9gFVWf
EQJHIHqFzpVf57qngDWDrNnYgqNkfDLBqAN1xUDTFv9Uya+OyZbk7OV/wyKsUTNP9WpNQDt+MT9p
UF0zrfIyrnpY0gkEXP0eNUXuaDaI9SdcWrPKxVciGlVshOc2F93+DjOxIjfMjulYEGHYCrjIKSgo
yoaEq2lD3YVKMEyA2VjJfratpN/etnn8DnW4Ggd3ozTvr8m1YVrC2EQyk9xndP3LUOHHACFrGODS
b7sPuG7iMvaooIiQtUIbc25XxU6VdyFGCldI1/JBGXJAOrTqDb/GFg6FzQeVGkb0TgUN2J/9H+Wq
MFIUr+yV7DWb7CTXEgbk5Ksj/DgQ/mtzulTU4v1iz6KaWYurfnzwy/UkYN29rSi4fo64mCWL7cxG
C01PdOl4dt6JLcyu37TENuA8M0CUryMSt6/tkfLgNZBp/QBjuetkjmPTin/M54pH0QD6yDHDHrh5
VhIhq//+bkwgB9gOuyCGI2qgAhXNpQruu4h7L7VVpL3grLO619igdcpu737IKxRvB2oALf0l3Fyf
Ln0jfrLRUYKJcggBi4MXvewqKjOZZ1Tr7kuxVxEgBBYWCNkCvZrCdIGvs86GPXcHeJc1V5B+rxW/
4JL6t+74EDVDw/1y6AhSMd0mQT0ufbp+zmV8AH2HlQ0u20iFNe94GdAAmOgEcNGyzh+FMArqlpfU
D2fGYX8DD67ldBHb7s4+GeddzG/poBHnqVB1slbC7lS44LYxYe5pG0ozoJn/JmIMwlEO0I26xnDe
yN2BmBP98vr0P4TmKnOBHf7RIgVRpfsGezEVjnDS1EKh1O9sLSg4k5mLSss2+PgM4JX4mxxeVz+X
sa5vvoSmxVewAu6Hq1/m4w5Agn06xDFNrgsNS2u8DdKbIv7q3u/6tXH+uu802v1XH+yFUJlog6PY
Ep3eeWNb3pXmimeeQYHJ5ByBh9SIUFZ/Ha8pqv/4MIriQ129HEtQsKATcn8oL0IDQ3WSrGpzhzkN
CdJhsPEEE5Qwx/oGeGJMSouFLdhQL/PLgCHkP0CkCoX4bHgdxM27ebGMfu1KnKsm2DUaReENdTOD
l6k8UkacnFx0Jyf9TJDlaL52reJDRlQbRX4xS9wXc9w5bWhdJ/SueJjVOrq/cNzNjHqMZkDRGxPC
XabA5c1N5wlAZ3M3iqG6yBJ1/swvxmcaWpCKkFZqlloigHPHFn5NIbCH4h3ZMb9nky3MErWT675X
o1msKcWzEg9eGekc31VxejetkVSFALQja/RT0e2xhnoS3uwHVR5nRGv5U7a6fFWh1KWLdqqliGtd
ZdbG89qcW4C+HWQD8zXAA51H6xeGZbhIz5lgCo8km56V6HQQeXsoa0QV/QpPQCWtP2ZJXWtQr2X2
JciZzg4Lv7py65clWFxp6/dj+fkSJR/gCV1Z2itPUdGbxPCuDIE8MsfQqa8S9UiJS9SsatWuCttv
kbI7qC44+SoPp/uX46At3YTCMYExkQN1b7U6J1bJiOQsoWxdcbW6SQyL/7aZ+podn4NH7Pq8oKXt
rBddD830YxONLPvIzrof5mTuokzARIk2wZZe+s+eBoLWE9vGqBJtF2QF91+tlQd93+BlVYPsGC0C
faCpUoBCdh9PrHA0rZ2EOkzIqWHZt8SPMYiHWYB3aadCmZFOt6r/Z8Mmnv5EaCu7m77D3iKq5WSP
z5Rx28SXsjhUlW0KFXa3O2eKQBqGTruHdCXX2FYe2Nu58CeaHDtdIYSzVKaoDkzhwp0XaQw+rnOI
CXmTfUpUlhnRcLMN9r6J5XPPQGH92m3Z/wQ+XHlBmkLctG0ieOoLmwnsyoFFOJjRDxP8WD68PQWj
WpuM5ZEsSrKpYSI9ILnblDV63GPw+Y7mDSNH7Mu7MV+7q4jxkERgU1UEZYgz7/NqrXlDb40663H2
/EQeiZYYZkwj2Ei5UII/s6Ej4BdhO9CPVh1rBhNuRFLOPhG4o2e39MVbNZj5gIKLhSLIao+3P3LQ
IedIXIAf+3zCV67/lhsle7Pd7l/QtSbdsI7HCU/OfL9N/8zauQh0dw/FLXOlDsBBuP9L/NbxfBcZ
FUX8Z9x9ejZCmI33OYeBTWEoD+s874HEPq3aryJ6jbpymH69StD40BQb+G1yvyas94XKZ99gAwR1
/qeiedLzTfDNVgGDN+NoAo/Vb6E5qjTJZvWTdgM2w2qWz5cWa+VPzBu6tMY6TPYlP6Ut7LJJp9Jc
rQRLiH/5nqFUiEeiWt+27qJ8tI/Tfl0wLlYP/s0U7LikKiBavYuzWviAhJka68FrA7y4NHIWsNa+
OGw88AgXrmuKvfxWHLNl6at+Jn3nYfCB5RyNABy9EzxivzIYuX5v1M5UxobC5bJqYOqtYDyF7T64
a1nOoOPYt/6mYTpdZfBcJLq6+JrI4wOErKjuQORnGKlzo19Me5M2h9j4fwMAYC0IXDLkfqfcHYPJ
4RtyauUu4eB1H+ypuii7mTsrcZuThDdCY+kYJplU9IU3ztTIq/xp/GjWI5SwxQx+reeQtaWsAW9a
2yFDGGuj3M0MqP1DGb37wsAYKDAAnx/OmY9pdIBkIuXsh+fNfesvAdmgp8CwnMnIsWz3wDG30A7m
AJ7nPbU8kHESDPQ2TOt0MBl2meUE1Gam2Qb+vwjsducxFs3OEFKG1DDdX1KlHnGOF0ovHNXD4CVl
r8I9oG3GCCiRN0QHxUHLRyPnlKwqQV+JZXLngv23xGmdiwh5dXo7Rmmam0cOsLRvaKarkZOSctc8
N7OAXdvC5E+fyWsGEBhlWPbYM6s1CSBVWwgXmbmf+7abI+lmOlyRdrCNpPdkmjptuljjMR77uNWa
NIdxgfCZVf65jPuNzmBLoX6Pa0HUYu6HCp8CGaZ2Zwiyu2SVI481Jcd6ZftmE4qOunGk7sObXYib
VwDyU529dn9tn4mKkZuzu81d2LA5r6YA9rdm5O1tShIXOSSmp8PRuzD/TOXi+Qo0qR3WrFmkUF1J
Y3NSoUJG0MSJh8gW8CTLXsGd4zUk8VPbd+uEY9Uk1prt2swTEO3sONbfvGXzZuQvQphazJ7NYRFX
2gAnPzeA2tpEk/PL/FotOwyhim9Pi4/sVSou7H4C0Z6yVuC5jUcU6GIBtx78NHC5WegUk4jZ1Y8S
ZbWEGR2QLuCfxTTSij1BAq5OJ4ehGec/nR+1W87bJQRqv1EjM84J7eLe+7wf9tA8S/bRfs6hahPP
Z1Pd+reTJcKez4FTjAxNDqr9OduK0gB0AphmJ6KUb63sBB7RNkMWsAh4u375UThyM0ms7AB/dgQt
riDuz++HP326nLPY8sWnssppJ8RHYmZj5iXtd2ClK6NTr1qCFEaFhe8/F+012xnr9NlEHusMOtm9
o/OkuTwU/xaWJAhc3SxmdH/phqGEoOyN8D40pIns5chq88wYLO+VtadKBhTT1hxPiuObfSSLzTcX
4rXvjf8Gkm/Csa5qTyqvnxvK/XtGSwwhPmC8m6PLQTcb3TgrTQO00YilTuO6ociOZhCjnFqq26mS
EniTdQJ6ApIeaZe88+LPGlPhHO7NdQZMPoMK3pV+gbd4kDX51lL8hXyVXuGLlWaP2HuJR5YEHgmZ
o+94EmwWTt1A1+gG0uPzAUtbryAKwoOA4NgsfWAhAZLdx5OjXhUm4dyZyCWrao4PG9/WqeZBRcq8
JaKWoRTwrpZPhT/Lr8VtLvD3xunax3g1Z6+PLwh4juMnSWBTWQPIJ1PoDXiNMTnndaVVTXkmkJqr
7tEvzz7CYh2oHE1r9nEmfX5r/NtPOJRyjHt/OaojOZOYLuODIxRTLZdVavX3WJsgESXtoQItSTVy
72PGdAbAGuaTlnbOeTrbyVHk+3HNeVqvhKv81BFxD5rWgwJuhsiAwmIDQOXF9RwTyiPfQ2M2J0UZ
2APDwdPKC/CE6sZ4dU1IPsLXN4N2gyqrAdGOJuYRLSxPCmV9DXH3a20V24xiIdWVW+vcfs10lrMg
gWt09Iaoent4/8MJgS8ms6WvFh4eBPkafI18qJfyoFJlsJ7TMthWsRkkkUEtANm517rWUYMHOYCx
vZtE1Q8llWerOGmAk/367Re0IaAdlsXbRJWwcOn7gxXlP0efC4OvJq442tC6HLsnhclnzBJS4qc9
XyInY8tM5Yenoh0/ivWP6sSd0yVdXG9BAnmqzX97hdXU9icqbEqZTKYUAaZDOkU6XvbppqjkSikN
wONeZpOwfIeo7dT+ZPOg7MubGh52l2NF2uGHqvMZraAzsm/fvDxCSvzeoGtueUGrMrWDdyqQzodg
iBw5YQ8Zsbn5vMtTGeIDWI40UQinRegZx4sLX4EE8dcXX6AXjjpuFNynaGb3XrNxbLzFYlZMPvJu
486SBqQnw2pSF0dbZ6VJUqt48pLyLd5LeyO+gzoiEKV+ySMHKg/CRv6ZeGchAznRVfg9XZYQp6vw
Ca9Fh7wp/YahnPsQu6LofkK3KrZlhG7NE+Fs8Ee8bNSEfyRlnWtfyRmstJk6tXWzHVDjnB9/V/f8
3viwLqgVlkQHPjbk5sAz+T5G52F5/8IeYXiwY7E096YC7A4/RIhNebSzjaa+L9yfzWkpymxQTRFS
BJKcHAoaq5brR2tWrbH+mM3oCZ42FpKTNh6H5vuHDRlELwDb10qSwoU7IbDqQI/VqxDuh2dvfhZn
Lv/CrsCLPrvK4zoVLB2nMX/6O4qx9nkUMqcOBi/mqAevj2fi3T/3738bO3FlRtdAqe+SgCJEH97L
mBEj+yvNBIqBAz0aocNoN43Y2sUDZ1FFcajnyEKfGmvEielfYV3BjUdHEPVSNg2IATBJXItQkPyK
8o6kZ4xxf7oNGkMvknjxzI4BdNvznTOyWUZoUQQK0Ys5MC8JJ9uN2PdxLACnEPy5sDlUwuWYq2Bo
LugbicMUfPlPYE+b3WGIiPP2A00uEDPRNnlnsCjl9xZl/1sbdZozIXcw5tUCMAyq4Zm9TE2pDzgw
Sl4gsG3Ki5aW6i2qGiJzoHfwCHQ8fkXZHL93naHJGZQRM2u7SLpVG9j5rHOUaxu/6fYVwgbFbKYu
3kmPE5BDOMKUbBO76t2+L2c+jIKYaepNERiyIP15qO5aZdGUCCwahI4mhCB1cr1dvvFxtuoehSdy
0VVxnn/FIZN6K1Ap1DMEiP+q/GUPw/g1pHnn9Kr4LxxyVZqgD+LKofzpvt9T5CcFepNKV2TN2xyg
HI/21fJ4JdPKPqO4VrnJrHxUdePngZImHvy+XIUb9kYwZTWaZFMuQzTbZVFI2XiWZ5rn7JRSs15z
9oJnpQ9RZqr2vxG6U+8eFiOxrS3yZPvDbDRTWgf2FtcjMGL3B3lN/Wna97Fgy7y43R+sIehhz9k1
phTOaRMLVgUe9Syd6n7ye2oDg1jt9tavtFEQSI8TXICD9bgwfLk7aD/eprwqHpXMouM1IZVpGsUP
cIe06eKmiC6AeEwq+CQ+vOrlnCXJFvR0Sf3DcSnrddZChKnVR6hGokR4VsPACafa4niafppfrsip
pPSp9CV3wF+xHo2Ktk1LRk0cZ8xEebDPdb6ihQz+SOwX24TXXeTzDOS3HNv6+bJanJdQu/Rl3fKd
k2cIVBJGA1TnJQuBaCAKS2PDbgTHmHxnA3WjKEL8yRZWAZj5D3g7IgnEPQRyefTXRujyl40d7Yx0
5l4ZVph/+BOgXAswGtC7wnx1F1qe55fE45iL1Xbee2LuWpJCHH64sjx6XSX+PrpT9yJKPqy4ULxG
AkRqDdpPmckfWukoW6jAKmPAbEVUFR5e4V0ncZry51cI/EOpLAM+MpTc0eLplwno9cEWIKU499LU
M1K7+xCatkjcfoxXKXOolDY4D64UjZnvkVVbwsg5CtuSD6R8pC5nuEYTq/bPd1DIyuVyRSQ5Wwvp
wTqtraIF1saxcVVnrCXbG3X8lP3YPJEiwI7G4rdZILV2tjJyAbA22aqHttrpjprR15vhpzF4cbcZ
iJKQ444lsGeKjKihXVpKEaOWb4iLe7SGbXPX2s0AwoGgG+0Vya9ixqEvy9+BjFeunEDD5gow2a5E
2r4oWp1MI0imZ+eGt4encMgvADkpz5k2p2ZO7hdwwLdegdwyN/rtBqA7M3b47V0Pt1uzG5J4i5vs
l8UMVpwjTzGG/MkXa5Xn1Nh3LBYV0uDvdW3eSiYoSID+WkxBPFXE9g/bSSWykKWJMWdxL3TnslNR
hos+d4XkZfvHJ+3MO0Hw+qieKE9cQXqLJZ+Dv0anJKzxQab5MtGOhu/Kr6zVh8AShiQTfLhCLs+j
r67FBTgF7IJJwUfj0s5Coe/32qpzOjWVnhJpvGBHQIJr9GTqDgB0Sr+l3An6ksInYfjMrhBmxEB5
2ENzSEU0VlEiIP7oJFo2zBvo4shqWItiNOL22VCFgcXB5tRwS8E06iW5uglp9X5u6gVjgmOf4x+T
9VH/HtFEAXl0T7t0z9PhYGGMU0ytayTX93NWDj1yVio8Q4PeSLp83ngOpi6yd7h9795J7CU6Ln+n
1WEFVEUFNvh2LmVh9QQEVnNIItFPCPi+4CUowoBtlZiOvF05jHr49I1+/Maxgp5SPkNdBfBBhSXh
TB6Gf5Mq3e8NGsTdo9wUeqqR6+aheYIs1RGQaLbqtfvlgCkLSh3HCmz2RhsFYxzI3YoUD64FKp0g
kMGwSbalWmVhQ/JVxa+sUA5CDIv/LMCWax2fHyb5j0n9KXKXJ4yRCc5fnEIcDGbuvkFbXucEOmYE
AQDpgJ2QCrAWE2iHH8dvVcdNtU4bYS0xN12h4lig9vUt/9FjwV/PmNjx0vz2hrtJYd7BJJiCJAM6
B635cE+FsoAxzfEpcpaBl9CSLH6Zcj1b/0Q8kpRGSnq3PrRjyOOPFTR2Q0ocoqlt3wWWKdkk4BiX
XRAUcP7ZPGiElNubm79xdXq2bCxw622MNonEAVtG4s7KwFeX5tqCepA5Xxs5Tt0taxktwXw1Cyd5
3Xs5HeW6w1mY/HOobqsL070oUJuhPxuMkuWndhLXWUXYqEEBy2x745Ll1QP0kyQplNID7JvIKh3A
nsg6/iKbEDjuMUdSvxrUGGTh5z6hSGlzSyLFQdAEj/MnlKcSHHCmqqX1NXwXEX+dkcEPrRZ5D/tQ
E2AhY56qLQXtpH7WjqlIl/guw1rn5fnWA8egjPfOXuLAru1kOU7rHyuKSaz1ddR1D7OfjiQu8qM9
BcrEkyIY9i1EJw5x/eDVJo6ZNkggFWOfrR0iICMjlvR1IZiUmfzQdGHJS2kwt88sudZT0kefCnXD
CAPi9ih8nahqzZDLAJgv+NGiVu7GPqvQHzFnA8sUqtAlgdVwKXp8HmYn5Y0QlO5KvbHPC8Tcu+1/
moWIiHjSxuE/JQVLMas3dvi6av3/1Jr/7JoCss7RCGMQxmyqe6d8BF6I5Cuc1uMxovA5o94Ymijk
lifqKaRFOr7pzeO3QcvtkrH9NKem8nvfWeqVeqvXw26qEW7TTg5lOGdQ7QTrurFE/gZCNO6obsOi
EaRUbSn0392RV8EFSLNv+QmnIWkbzvEWL+2azitATki3gSMsAnfNx08foBw2UXryxGkMk+k7OlM/
KFhD35fBLJp+XbsWyWydVTh25/LbM8jZsF6V+Sf0cfS8NR39EYnk8pKQnODNMqrAXlATwNGMlrhv
srPU9UrmstV/14zI8xIkZociYIoqq7wEulxhcAvrv52sngm3WYQOlL0zs6iFrKVITrgsjxfI8l2T
TjG42UkpgO+c+Dc3WcMimceAB0pr0C1qYc9WeexFgQYeXPmB3+/ktSniLw3EUkYnJswYAMP12ePG
h+3u0EFhAUkCduLgbvZwTtU8ehrYoW6bTxXpqk0tmBLwCuTgWDsD9xpp9tGSFHl43izSFmQNqxpI
9kYh2sXCZgOd1KnDCMsi00TOk3V2EowaExigyPMu3mkoRnIVk953uepQ5v1eV4QEUCkSAdLcW3NL
Sue6vrMC+pQs0Is8eQqorQCvnnE9dk0MWGPvWnp7EaLSTBPLT3x/LnZ9UN8xALjABzbucDXB03B6
tvl+lH4hiOEVjH+Gqp3y3z+9CMsT9Z0/ZejC4mtUVY6Kfie6qnTAC5GLmhZc4eJKXK9aQf8vD5sI
IrhPF92VOgPMO1b+uxS6Bgc+6739FIVhyDu2IzZFR3egUd96IeqeA6u1IjGYS0EUSf0F8QaqvfZC
aOSImvzTaP1GiuHGU+psD68mm0Mn4UIFkP3ENd223380NbJ0zm8FaEXP+fLVzBAKjbPyaOlbWesG
46PiMeS5+b92qjpqW9tcqrgS5w8r2iUozsoOoIZvFw/lgIjNgJI3DGiHbY5h5IxnKACLeimN/6Tc
2ib9/W3xt2W6j9PSrnWs6AZyTZHG5gW3wHjUQ5DU6IQmWZmd1pU82vZedm5V68lf3ybs185gvR/c
kQUQ7b5xh6RWjS0ojnxwv9GX2ycE2B/LjfVt3cTysbgXbMjYIIcHcTf6tWVM2b2Dk7hDBxy/0ZRV
7UtdHYBf6fEpnjy2x44Xg+vNTB8wMYbZrb50iEWNqmqMF5Vap7C53az7d3TMLlXeU2WPa0IYbrgB
mx6N4SbSqFeHTbqh7No5bZj7o1DMIs6i1JmEqcpst3wjQmM+vq2C8tmlI96Tgfk83Ws04LhL2RTB
e21pAKdhM3GXzI+Z6EfVGVEwIdn7Eexur5c3Xo8bAllCelbRSGYo2PZZxqK0krXj4mSThic6NeMj
7ijyGvtVwYsBZZZvGFOX3Nw6kbtEhq9fe+0R98QDFvUc1HNsWhSMIK8DVjOG2VJ9VQ3kT/nXbrvq
QLpkx8j1Vk+qQJEbvNme8OiSh2yvLUMgE5tqC0K2+xNDt+ZrOz20xp6hvoLKqtO1Kgbh5ivp5h8j
KK5dSBd0IBDCXa7toSyS1c6ZDFP99Wfy8kDj9BvVh3WFISoF17T7n54xmC48r4CiGJNTIiWbKdzc
wD70Q+ykWrM8Vl59fYNZHpJ8mh7gtSI6rGOSvysweOPRfD1Wo8sDodUJsC9hsc0LxBouSoFoTlSI
Y0wPBuir4eZ7gySA72tg3TZPfR6ecdeMRa4pFDvbZy3cjT97MC31RaC32MDbAAGwAFMpwWpz1yt1
ySKoGCLBa6ITnRYZLDMhIZpu4e2q6l3qSWkVsoygh7YjqIUpFiSQ/XdB2PwoTiQ1F5tSdl8SA2zp
55TXvAn4QfnyQRP1BMshVzinuJhGARlwoe9zDonJk6sj3/IIdVOKGVyo9/ZtOBEKCkvTYvmflv40
LN3cOga9T3cRZnEkvYKZi02LCOF/waClk/pDNgB84dRRL9irss0Mn6UnPRzM0Rv4zUSvZdDkIdq0
LR9WZqPJQTdkp3yUoi52Njk2dERe/V7XWbayZbqkeDkztziO9EoR/fsNuCjMOWjJjQ3W8Baf51l/
g4OYmN42E15uI/e/ADLrbAhHNw0b7wYEJiDU0ORQng2B++0tNKsvSksasv7mis4eGa8bxJonHAE9
zXljBb9dQuc6KA1brLmNkbAyhrNiJ9ZMQhd/4dyKHnmAsFei5S8W7aQZ8eviVUH+beh9AW1jP6CH
dc2Vete9yq1Tq0OKdOnjMCgc/Ns9mDEYYmlq6/3TmMlHH3S3VqmZ+hg9NtX9dES1zmIMHoY2B86r
UWw7Fwp0ypiloeCVpVMoAd5KB5tHnu6+twZ4OcEcdhr68jZfVYeiTuIpylXHex+ZE/qRaMp5xa2B
+/u39aI2xNcQFSKPe8Urk7Jo0tc3uRWkunMeL7d5l6sgnJwvCIJZBci7n9V4vZdCIQZKDDgaxkrK
lg7+riOQdNs/c5J9dCRF2r3q7AH0cq8x/mw0+oS+W8x+LbKtKbwfuKZmXuBpKBFwRLUuaPRePEEz
I68e1ajKGbiWXiGD/xF6C6IvWR+ZWxdtbzHjJ/2bRsMTiRFCWUHbn3JctQm+C/aNMN+CNoIsNE0H
J61vgI5VmPgVuuzg6F4E+YoTAtE/LSi+j+UBsbji8t5e8RUlXUZzL2PP2ht9adTRzceaJQTYfiel
I7eLFP+6c9JL63gvOKTdXRRwS5m+podpY9jjtd+1Bf2C+vm+fqfJS2R+rEuJmjEnEG+ohgypIDfn
UZVUIvJPdEbJ68P1iC0n1uSWHLfYt66tDCSi2+aaishYJPstCfthU7pqhTd6FgrfKtg853R2iNGh
fw30wRSNghyMzvOYVRN3ekL37CCuh2JvIapiO/1eh4Tx1eNx5Cac6UJsFcFsSfmS97C+Tik9I+n7
j2JWt7yeW3ivJeOPCrzoF8uUrCbhfthP3y/039BTllYkskRiYHhevoEQSAXmv+9goPWhx4JHnsxg
sRiYlvb0PkGHP4RNsVdElrSZqCGgD/uqgr7LrjaCW0rEG3D2A4EuyJCWCteWoH253oSoPhBqxk72
Ej+sn9gcIaobtOeVESniFxi4lYvV+6UbtYk83IG0i9MxLaaO2F+ufwHPM/r0/slclbgAtttmAQVB
LWxSGuddKWY6fOdR1gRKo+X1ATrw8l+1YhKyumUOoBomG5ek5w7ri8UAxrpgV6OFVIOwdwZcOd7B
dCNOBKoTCfWMwCpLXXXqvPrVZN+CnE/gCwHjAygS3W8wMr3jQeOw7Tg5tOml7o/9blSMo6vfN56o
LU6kWnBazKlpV3mypG6zOe+TYZvDAjoLCiq+CPUeHyi6j/lRlH214OeFqVhdvbErG5JfNF8nPtag
tdtZU+1Jqee5BILlup2q6SgzDbT1EWlV+r7yUfKr8DJ+turi1aCux/SpMHrWqKHs8pqUiVWjkdzY
f7UWz9ExW4hDhj0MyvhaWqTUTdnKsit79a3cYAfl/ZMkOaiNLuC931LKfARUqWeGy/ZsoR3gMCZh
CWvD09MRXEWDaO8MFH8kpnf9HEQoV7jEwM6shg829xshG7HRw2nzIxikR4CmOFPiQgO54I5jNOIC
ZV020M1zOM+bpzRtGwqxQq0B3CjcspcrdmtFGdYN9SesLaEYfify2ICgAX3TlK5wDfT/qqYHi0/p
5pxTy2V/t4wjpttUqO9JA/Zd0xqUQeg6RVbt+sTblm3pMSdhcFcnDxq2praq8pd4MiSyH92ImFRC
iTOXcpSp1YxxYJYebIec4+89xA5m1C4f8uxjRILZyEvlMVLrAsmlH/P7QU5LqbqlBRuMSZOiE3vg
50ksEoME4eLvmtuWoZzCYajBM30dAnmyveeXGrK2gZqwdy7lJ3KKn4nPGOlj1WMntnl6r5Cp/mST
kz0VH2VDtnapbfm7TaoYntHqfe8kdfNuoWG2ZWejHPzzfC2D6nUIcd6JruMGDTSgdF66FEnfxCa9
lgWg+tIpOYikwnSxgH+wNnnbqgNIYvfgaPCL4376JW9qDd9G4XGl+PD2ylPXoH6VbbaEhVfhUgyS
Z4POuWuuNY/PwNJuIS6a3P2As16kIWeoW33IMHLUYR7fVCVStzuGfgSbspTw3JUxrSSFSbpkV4ZE
0YSppicoRs0bkhvtqLAp/fBwP7Z4oworhcnaDlHhpyvEpKZuC++wEsiIx115bizeQIUMRm+DiZHY
PViovAg/1nr5ADq6x/TahRBqyK5A3G9N5lkVwkJlR1TwdNmpQupOzSyEnYuQQKNxPQSfYk5KL9nm
xmd6G+DfacMqUB4m21rqMtNSAEnPF97XfSSkVlczBgca4aYCbuZdjlda26duCBwyBz8uYtq6aVll
ltGpwXK7AvrVOzUO40WTIh4Ud6bF7Aln5v198fM/q5Dh69LxheHqR/zUsQipyN9CzDVeEcdPr/QO
oqo0rL9rV1RPEKoUfnuMsZ5VW3fIWAvoWk+CPGJ/Ef8VIqH3Q1U0cIznkO74WJJFwbOFjEu4W6dI
ZhYfYpXGk3OoHU6WimNekKHKBupANXRu4cieELaBrbN/UxH81mxLCLNwwsD1EpijgzOOqGGn+diX
ceTlfcqCuSUma1sHwsQxbg5QdwTFaSdHpNmgAEMgKXg8DGvD24fjpwNv/PwCKnCcu2tunKakFdNP
meHUFZzBtZM8HVaPsfd1VepPbqmOy+SnhR/AdLoGfDm5ISCQb+K/tKtPUfpHF/CLiONiRSN1b/DZ
3B5FcGQVhrU7qZvkuH3aTLMgDh9IpgecapkCFJfVqYKsa46xDRDOswnIun5TFYI/BHL41pTvxpoK
2xbt/p5fKM39DcWaNQ6RW78m10mjRYfxjR2tGunclYLpBxscYxeK5NRcGF8/yjgy1qfnVqyi1Gc4
Ag/O3XmKTHwPzWagnXBS5ur8sgmy02SMyPKhTo8of5Xq0j06HOjFNi6aXpa2v/lIb4lCshdK2rmG
wdWwmgS9S8ePDPniZE82MO9bwqTK8/NZQY7kMU+43UNgikj6guAUIdeAzPUsHXS2YABPtM4hgEeY
izx71OS9/JVwV7nOdWlfVmXFBUd3xoNkRxgwzYifl5XY7LhaEz30URHOCenwEYrrlLFW7syJFN72
8BymSA7+K0jVTZpPsvJSY/Cv5o44envLbXM7MRelbIxmZbNzkUYkppvJb+jC4FfeKxs2FdfpKUR/
ckhl0V3EefrLUM1KEDOHIOZomzMSEuGnlB6Jd8BSHkLG4iIkybtlCeyK7mk/UK3gTeAw+zgjLeqh
1SrF0kCn8Q1MaqDh2wT8zeXUKN5AuHjgb+ugq0fQVTWeGEqq7QJrj0q2NUmaH3U9PKtKPdCwKAV/
N0lqChOD9F2esS9QTip2Vbd0m/XtKQjCGULUSJJOQJ+xDqO6wl3UGuSaL80IMqLxcSOrAEjAYPts
tU6iOUza66tvqLXZmhKtxJM24QWkwUNj5sKKB6RGJQzql7R/ZEfmCGRkcnJBb3seD4pEr1VKCwlv
uPrn4A9iNDgBitAhQ0GIsT2JSgaGjCFFg4/4x63o9I1N+hxXdw5817HULP336lIRMcq3VHjPhhRq
aCwwg8FpKYX7bK8fXDhzcgMhdzxj5ay3UJPE4FZ2YSmHdKPXe005xe7dSFWm8/+viE4t5CrkEspl
l48SxOUOgld51A7qZfYWJnuDm3T/Qy9Y2RNGPaKRoBkRTXYbnOOrG0ag17sx/lyj6GCZsbU7UC5R
npEQ0Ewbpul6YqPONtmC1l+3MtFOKmwAVnqjH/5xXYcDynEsUnoZC6jtCxewaQlatdcG0OvSaILA
SJJ6EUzoQvGmGcV+f3OZoKd2Oy15jicFfgpfYc6n50cQBi0HULaaWSmC8J9TnYYhoZK1PHDPxJYM
idxnqhnLGcyskg7aP327DnaD7199B9QBaQvJvlhUG8MTGRvRtHernklJ48AGgZhMmvSaDk2NGJzR
d+S06HeJ2cPiBjz/hkDpAaNzfSHLPWvxMRVIqRzMibL99IXEkW4Ud6kC6nyVTuoNVwEqg7fmh5Pn
/zCX9djeRojgEr//Bg5PGp7XjFy8uBzmcqyc2JahzhDqizoClgg79K6YIEHhJCs6+DzS7y+cgQ64
f3oQKZ0oR7Btib8ATRfqwLbgfdnkZUy3bMn9OvdTgVPWFlBcnW6U7RPw80KHukJ5bc3LcLWQRw/L
SMvNxer0FTBo4ybmjJ+DHR7kotXcQsxc7Ni1CHpjcXIqUaVQr0FAxcKdV3A8LVTLPoYih7PrR/5F
wGN6FTdnv3IZuqXVwas80pBHQbO/B8uIqvX0KO3dCk+SuVE1gGDunWdXjCu6wU24btjV+tbAdgA+
Z3aX9tQlDhSvTAPshrAQtweN8ltvjWLSoF1nAbRzcd6vmcz1biVv1uWzeAiVv28iMzKnpUrLzuBx
qWvZHTQf5CN5C+xihxuXyCagj0J+Csl2FoGq2gZJwxQMJBlmxdg5FAyT69sjydKRzu7wh4XoMJS8
56cP2KkP2EBdFV2Y29hVraH5sPh950EMkYqMnwUn35UeJRWpYqagKWFV8fuUWiplZQxrzxNO3Yxt
5xBGqcc64Pe/wtr6wbAwLy8hAXChYKAwtqUwRHIGmF2EZkf15+XY8CcDNO3dBGBT94Y9HR1zszE6
R/eNAquwEdGjXKUFc6ybvIC0xpBre0FvsPDFowCsoFU+SrC2vobHHa9XrtOe/3e+tI/NWYn5t/ld
PAFvCKh94+5kN2BYOLH5lD6CbilXycYg8Zo0XnGP99oTC9UAIt42eTJk0PelELJ5ZyNlbDER15eu
pLnPHge1MY6Ig7vDoehV9AJtsgfYF1rrZVhxhSML5jMDV4EeaaArve6Vmzp2wUaBOjKtKPlYhbWo
SbAJHUI6ZxNvyTU3mcruBhqGa+83oiudFmVWDqXjtQMpZ70IEZ6DUbsqiAnngR64xY1K5Teeyoft
krXe/yzwyAD8u5r6Kdi2Ub22q/LASSlCTcKqg5DEVBCYfO43bDByXmLk/4CGdIJS2k/Czk2AgrEQ
LogkwWsE7b0KBqFATtgtxYDl9TkAf9F3Nkxax2ks+kKSkpjp7qtFgpKKBsyATdTBklop2mJpfPJo
9Qf9hH2fsr2mFyuMgyFpuWLwb6Gd8eznYTqDA4iyPpDFMtTNIDFGjIw48L7O9XQJBHOh0t4YCH5i
XQ0rt0Kmz0GpCBMrOLYl+Do0s/1wP/D+gKhLIBkdavvEdxb4M/ixPA3lB0G4cQ7NRYh5si3Em9vy
2Bn3Sq7rlx8lHJanShdEMdM19pvQOqZWZaBSgbtQCaGp/cjjtAM4uWu3D8OczK0z8xPeaq6kd0/W
vzIrk4QECgjrj8biuPIqAZK2uEJaWTLZuDD3bWNagATK4goLrFpuWPYaCPsM1y0Z4LfxHQoea+4F
7nYr2u3O3k6LjCrG/van7BgrOcDwZqAilaSpJm5O50I/3jMyYX/q6eWGKtrNziwHIq+/vy7O6sIh
GI8HovuW7oSFJEgDjdpCg3SRMJdR+7z3ph7GZxktpbDebNBDWG7h6UAy0IBNkr2ACK2c1ybRKjMO
nBHuaDSDMhTzHc9gro9Jju9FGmH6b39lTJ0z1FMCyZjulF3PcTWUaCq27WEeKqrjM13pRzzp9XJc
apP0Qu6L0Fx1sW4NY9WjsXuDC/AvCqhb4m5c2xLi5N46Am+sF8IeGcI6PUomhknw6wLm9uzwJe5+
i9ivzOvzbFZmYtte3BKHXzkZ5F58gxHkYBVNUaPipAHcbomT6O2kbHUe/7SjSdV82raQOIb1C4kp
eFg4D26ejKy1Xw2nCnmVOfnOwZHZMW35zj/YgNClaov1iO5BMB6ht/ixJvvpwCVgq3zNicYHsCc6
2TQ63oBgfjYamQwO3Kg0COPtvUa0suRidolNL1UtKOcBdjnsaE2pq3LP01o/y7sxUPTk09Of51qV
vx7zQt7BTiU6PdFygQuxOqveuuY1YV6I2c/iNMvXAzB00Pk7YxQE6qpQcvcrXxqcW1Ge3UDibtK8
l/+FEKWQ0xfbbDfzZxuQl86IIdsrktfn8F06aDD51D3C5mE2mV7pKljQiqwvQXYjiokRvtyUZe40
hL6nqDOk2OQOjtUnPtFD/B7864Lw2nzQjGjVM4gdmiyHy/hSHmRVQeKJvSlhBr3u8WhHlS1fMAKU
Bi7SI5CZ85seDhaUI5L3nDvhriqSxS0i9YKYAwb5Vz5Vln4tSw3nSEvMwC7FqU4pd+bnEGcEz8cB
JMPrEjx/OyuCLUlpEDni27DGyp4s4rw1etvDedlgPsIhrn8nwMEc9U32V8YIk01IHaLAj+yNrtb6
dhRvt4HG8oxKS+coy8OmLNzWRp9/zvf8ho/VF7mRlLlWIaR3t/4qfzwr7yGCBjcmIWpaQIYUvNit
aqMBHWrGQr+xS9vp1uajobB+RoNAs8E1HdrhYHewuJ1Z2PcbEIyA/KHltdAvkHBkJfdinOiraiGu
2Vg/rcLOt1mDS1ngSsGGi2uXu8lnOOV1byqLtvjti/cYwNOJgwTgbZ7aiGxxZtlG1fXXRPxDyFir
PA4LxNrbAqjPhWFtSHbGCPr2jtgcjMddN0szq30nLJX48nnZmy/lsf3OVCuAApoUnRE7Gfga6bGk
c36atAOwzolJIZleYciyP2csSCG/BcNZIggEmv5GBccWDnTdEDmu5MKwwaQK3rDo8myX4Pk2qzaM
LTge2S3/5nK6/qytmQFN6Jy2p6Byk9P5SqOt0u3RIA75IWN99Jwy+3WX/TMLEtF+QlzWCzW4jTt8
V7W/ONfuA7/m7OSSiJNkncp4Z6xwy1DblJAw3F6kzyOb/IYHKyI8bbXSf43ps19MLt0IIe7vtpBo
Z1BKxOasQtXQ1S4qpp/oEubouQpLHLCtQkwpXOpciX4yEVQIVRMmfB05dABVUc2s7oSXJ41wwqQD
uEg7bq/Z+lF5zpeydwnLD05fTkIblmpm8EuMeL9LGkxwO1zNA0ZzhJp5KH9Em0BFR1ldmrjbVRrC
6inqX2OC4xWT+4EbcMjXBIEU8UQ7pqfPTuNG+5K1KTEyVXZXu29UNjggpUO36gnBcVqbW+4T0U2O
XR1D2Gzr+L4V0BU7Oh75UKQflzV86Mt+fBl2Vn5YL5FSu6iVISr5NBMBi9SXphyrKKhaubtY2Qih
xH+M+PSPqowR+3oO8a8k+xct8Ve7/GigW5LMeThlS0TH6efQQnWoeH7XOsoU7VWElIfhkFhFy1oI
YS98MtQDl7qD6Yz0rTGlcYoXLylkXynuyyh+JVUaDe5zJvufkI2T1j8GvF/es8oFLJnVURmngS2e
c+Re6h/ue/QJgiwEBggUDFlCUGHvsHr+kWU0ipCCj+j/17KGQLALIR7eeF0R2Jyfj0gYtDwusx4K
b+cx7oKGj5eQ4WlwPPBoh8ApVSdgmeTs29EWQcFTLr/cUuJ0NMtD2+JKAk0FYSh9cv/zmfLvB5p0
Tk3NPFQhXFCF0KdnMn5nr2w4RNuXUzOkwpTbzaY6QjgKcmu7dXa0jm6BTeDwzMVo2cjl7gwsqNuX
Wk35pgslsuPnR274zpIyxshyQsGbvjY9r3nh5ELiyErY+t/WWmBDVMBR9AC8aiW/PZJlsqrcj78i
h8NQahHOYMzeB32v73Mv2LJFeTnniVTh1AmWeap1ccHtb/1owi8YhxnVOuZjOxRKnf6xRL/0LC1F
ocGlixiw6UjQ65N1006SWNQrvmJNWuDVo9urFl48nTySiwXBDv8bfukP3UoyWaJB6wEBVxI/pnLr
3UGETmj98xCYcXd5eNaWb6ACMoYrLst3R6TcjAey5b2hRMnVi5Kx4eIah1KAUDECfIXeeRm9yOE5
Y7HgTmNuaoJVnsD8Mnq5KRoLN+GzFf6uAev2YKweJEyCAaAyLzmbtheNX1Aq4igOmxaC1poHNmOp
p6dvIJWlE4Zew7qF5nPI20XpiemffRBONse5eP+zDV1fUEDAkj/ArYgtx7x24R5eT2sPNqUpIZr4
0H7RWD3XjF/MYYKbi+okoMgtIyLSaf99mo90rS1msuaYeqgIEFtgrzQTPoTZcjXXzqUjYKGFFnL7
yWkk54W38macqgTPEmeuQJkuuOTgeMeHu4+ny6cYnMV/uFGUl+42klDTp5xl9/Q/ADW4N2R/oyz7
AsTmFeuUMRdkbOAAMP0lY1+IVestryrgxrvpfuCYi/NEGIP3CRuM36OBMUAI8cIsOZGKWa/FqC92
htqpiXFEavbpme71caGzIsMLsbeiccOVt6AXCRnRqw9AL0lfpF3ENDsTipc06Aw2mMMiJ1Se/gjK
yCiESanagJmzZo75TweBU+WQs9nkJSYXbqkmrJwGAT4de9OPGAMcXpACaf9ggWIfJf8OIARA+AjL
SvG2ynrxxT667SyLWdJ/gbK8VAtHLJqlpbWrxHIMCfhbe63AycTZdw+JBOl3UbjGAdgcA5ZpEcGL
ZOHSaRj9/wSYYglaiPnUxmvd+c+jJbLqRfFIpavF6MqhrqN7LPH1noB7Zmz9sQYfqr4uuZgB9ENE
58zrYG338+rL4FJ/nL50l83PjI6Gr6WctLfN4qlpxJf48MJTx6OpMCiOWY1FJ6/bhDtIB44Uf3bF
hwCp0FGgINFo7nKJgWKp/q4vUTZjD5vaaz/mBN+HERSGvWgHPhQVHIEZKaJ6RwrRrUJ2IyBwXPn7
BM/tNT6QxOMCq46gOLXDfwC2CZ61p5ZnQevyFB9YLASCIxvm3fn/wuafRbig+R68edVbfJPJ6y1f
h2CKaSaSb9R+xvkrsQUiAiEp2VbK9r/mGtzy3JZghL4WABntd0eCEwXLhOuypS4guRFnVButSmnl
Tv2nlbfiy3MbbgY0nBetBkFyKbkyV1ggAHvDcNxvnXuepQVYYyldRJwoXEBcIAKxYxn1lRJMfmRg
w55GhQAqjdLJc+Adw2HAEvqP7l3FWkeSLSP4uO47GzYi7xSJOHPqL+/1VRTbi7bHwi7gXCMWqelS
Do3bEvWHIAu5FWxtW1Q9vz9ABRN8yPfFj3b6bCErv4spXlGYX3I5t+isY0vZpIidPAaDMIetjjnX
XJdTo6JSYKqtaUp4lPS2rC12w5E9yWQCW2Q0wRt5KFBZY5Sqr48Xmqa2jabA/Xn4yQeNWddYn5S1
Bty3AStfv5doeb1/nwkKQIApNE9JxedZ/vDlWfaiZiz6kqHKzxfRsmcjtVIN4xBYzg89cfeJaeSE
DJ7RI4mCoRoaEKK1a/h81JfrXaFCHzPt7V+g+9eIDvlJpvKAGCHvc+WR1erdSqmhst2LxLxuIpsP
PMZcYVzsM8BEy1U9bhD/lGl4Zdew25ComoGWh4fd7cAqrLKVVryeftflpBMmXTEozYpAKrAgjdEg
JS1KVUiu9FVtsZWmFSVr3pjPwoVM+Cq7/8jjZpfRw/gwEOo5QruUwAIJ5O7YU3y0ZhciXqJoywpo
jL0FI1ZqX1/UI3c7b6NHtEh4y8hWivKadAfVpUegh5Q9RJUe2a51dNyNw0W303OxgScDLge7jane
e14vmNNwp0PD5IbJflAbIY5zWEdnWz7dqKYXbBWWCh3BjLeJUl+7GKEwN/0EsrCjQi/z0xfzbDen
UDf+089iZ4eUi1KT3LyvFc0GldQZL8f/r3hIuFYcuUIhkfbsLmIA1eKq34lvtgPdcnf6FGHsDAZZ
ymeQ5n3bLMcuPccTK2IFSDbRAijT4djO4oTFhJR+4X5/21GKJDi1RawGTr/TzguJh9Q35CVppiO3
Ulw+CGrsdwrRTOfUVC5j0kRCz9eVJf1zP/ZZdu7beUFgPFeSYF+oY2Ju++FB7oGVWQWabaBTs+/A
bQaJnBaR6xISqXG9eUgujBYbwt8n07guHGdJbXdcJr/L3cizB5br3T5Gvl6fjk1yr4v+Ad7/hnzn
L9Ok9c+38XfEkYW5SLyZbjlozsUdu5iByMGlMXeyQ3MK7N2n+fCdQ2r1ZripiZbaJgek5gcxtpZl
wZ2MlyY4vIYNVUwRxTcRvZpEpPUKAqYzv4/tEnKGfVkJHvkptdY47nBma9mGi1Ulj8nzrXIOdS8/
VTF7FRwVJFCIKRToZ0VEliKqbCe5rEicY0tpZZWMT3jFb06w0NN8jL4xpnP9tPKrjw7BngjpMBG/
go/tDFGY4Wpn84B6sTXFdNiblm6aw8TaRO/PSbn29OSD9rq+GJkadQee+ZOSCT0qKcncq2Lkj61v
I+kBLDqyBqx+8XmEO1Oq1U/oQxOA2F1JOieUZ5wcYYa7VL88Mb9pzmxnRgFdH0mI2qDlGwuZYtHm
xUYgf9RaJtFN4NzRmSRGUsIy9Sbo7h+SUPR6zz+ABnGQdhEb9E6tYBds90lnVR+eQa+W1IH+EmNj
jMJqIq+FU/0wU+11/bypG191411gApnqerd2DXe8syEEovNhqM6Qgfdz0BG1662cOEPuF0ICSeeq
OdwDRI3ToI1l2QHh+7KIiRUi9JQMKzE6fhiDhxEZcv7vyhwwtvaFmvDkkqStPMYIjTzpuMsHcwvp
819RcNp0DGFKgdD7Byuh0JAglDzJDdZT0vn7uHFwWbneB1NFBavkY4mMWOCWnhXSRE0ZORwdU9Wo
9FzH9P0eWO5xMaGUNLjckglsDZ8YdcMS9Z48tsG/b4FtdRvH/vyVSLbbR33nEQDvBRrH95A1ZARe
DqdB96nkhJ+2P3lOUkTXj2s4xxUtKL6GOz2fFWHGDCAk/HUTvd9n2nfh3d04Wo9HydlaBElshWML
8Sb1ZTz3eJ/nde2F0ZBW0XeD7vnJvAbcXJW/TR5pxzU2VNhRnCO4Pi/gZHRZELHHQ4Xsusm0fSQu
Ze2eyZHXix9ocDfds19OQF+TFb9FyKiaJ55/FHnFvg2nBOQQmvnz7Mes+HvNC1n807oZKqwI/btR
hqllQzrG9demo8N8PpjKy8cIzus0CBO1xRdR8p64C3Of5pfIhdCt9R2cf/5/X8mVhWP7BgfREP/x
Q+qaw+CK6cJ208nNVQHVGFKaRDLnmLvDBegxxZupUCdenf11iaRO+GwjF1SdyYQ5ux1bozpM0NAN
LTIsYm2Qnf2GOy1TEb1VFCwUUClLE3sxBKiFGfJQcO8j0uZMeJbpEVtWsASmkF1/SBiYVhGpB7tu
L6IVFHXEVO61VxewwIK+xz5NzU1W7PQgKPURqNnFOVd5e/1PyekhPqFZwmMPKkWuWZIx1pCYv3Gj
wX9+BY0kdF+qWJpJXmcO4bq+cHotOABN5XfGVvN49IdlDJyRRzgpfT3x29/w/4FpA+iwdE9HYfmo
Imk2WD1vSmJ9lb6HXbaI89LspRjF7/phzV4frl+koWPcxeKeVQJRFuFayAvLFolSZ5In14NRlaFg
I+PBIGdftqKVxRH5x4DrWTehvQW/3PrwIIX5w7D069Qbaf6po4xaz7r9JUJSLVINhUXxTgNEj4lb
QPGMBS9M+n7/VMBovvoSxGz8xNXHZwZ/nqORuKW3VZTqYAFMjtT06fdIGlxFNXZNBdjpDOmKpOAc
WQIQKrbNdtsnk7MaUlQylq/DQ7+Czb7888v9B4wx3WpTnvZSqvajBvHnY7+5onL+X6SPaQINKD4F
EPQESmXAh9NiJC+gKyMTeLsI7Ad/4GHM7A3nggwnE94RK8FunIqw5NZBq6GWgM2WoEHmt7JHwS36
MtupeTrY5reNkQV/a4ELuvlN9hwXabsC+03NHTDz9HtKacogvH5uWHSEn7ZyN8TG6FQ4cl6zEZt8
aKYnVSfAj0dRDhJDQBKu0xwhkaWzMUzhJo1hwkIce3fsIElCkYKX7quaXNUL122E21FQMd88dJNG
G2N1PjWas5GX42JOt+hljUAP+lv7SfcEI0iHecY/HDTU4k2am9ooFFMGeX32WjSjt3wqkHFjifyx
99xPW8wiqKklc/w/gixyK4iEenHg7FBa7AKFvAM2vYiFK2GpX7z0jai1XS/VfbfWf718fqHwNY9x
/4zS34YmWbl6Eed/6fQ3VTwgAFAg7KvgT/Fwt+uRddPofjl1PFVb83ZKFLy2tCkYnITM+k3d4Iuh
B/QhTW1euvrZwONFpGLH09y/uVaok+9L788V9yz3OHqtTNQ18QiuIO//oFDzn4K8hhU6+dm1GllB
lZtTeFjG/3EXsqtbMW1rCSSjIiZzHwj4MJX4kMZOwBOh50Jy7pWpR7SCHGG6pbhI3JM6IGzyLn0w
JW2gouM1bbYw2b9g87dkssEzpw4Ax+RnyHgG8oKEVhxEnW+59HC6G9qnvCTwxWY5QbIrXHZgmqni
VPZHputBSOz7m74E1vW14cM6RFxO5qOV1SrBhx8rW+4S4fES6J/12Z2zPoiinwNhSQekB05lLake
AbAzqBfV1g7uDLVwiXw4DgCCZi5YQ3EgjDxRmmbC5ESC1hlvmP2JH1/07esPrwx22NGImlQikrC3
Mb/Rp7mx7bLssAzbupBSgBBXjffZzFE/4gwlwrERTuJ2jvW1uK2o0aUw13iYYzDRe99MgVSznDcW
M8qNt2GNlCYRII0lPFA64q5DKZ4wpeDtu34cVIGlL0iZuSgjM4sVSY109ezzfgiPS8xZLbjTQnFy
WN+83ckaskm6XE+DsJwLgZXrdMeVyce0N+fpjiXfesdiSNM8dfpx0byWtucB82laOPj4axupey5i
qlJjqcYoGdnhAqYkhs2U4J5OYU7io6Olv2xOvJBtqtE0/VZm8X6DZnYjGwcOWyXLZIKsYz6N6zxt
RfpucdY6PoaYW8qhLBAJ1B2r0hgUjKo+7QSfzU/aGga1fBvS1Xw+eTefsMvQ3F5MiKyZGhW+VUe0
2jmoo5DQ0BzJWj4VlpKIp/cP3o1ZD52tgq7nE7dsX9uDj0Ks51+wZ+88nq+/CJIQGkgCX8+ecayK
DBDJ2ALavQmOw99HJRkeov2xFg4P9ONz/aKfm7Ok0O4Tl4kMpW6RHMI44qJnokWiBHGkKFYSB2KC
oROdQimr4657Jy7cd4jTKGs0bi73dpzxT8/ApCsMZ/7C58S7IuO4oUvy3wrWQdMM8FD0FX8/IPHd
WJnpvWJ4JEVy2NfrvhwBeyjYIUJRsbqjC6lOy45B2P66LWQptC5nWLEIf3X8dNzcFinirpRBTJrG
phiXXgDatrqej1yPD5n37LIOMnPJ+TQ7UT27qHKLvax1FTzUAXR7c7srQP7Zg1fboDJ75QuqgRB5
TmS56nPwIKV04u8qFdNnlyhYjiyFHblvFxsZBe2KdLC7KN0zmqhcWwN9Pfm1ki7wt5IfFkenFE2S
rOdTW8qaX5tpi2fJkLzVy1ZPs/We9ULfobnii8LCmOdOF8w/ChK9oAN0b2kOJE1kTcqtsE0wCW4U
EQzGJ941t4LQD4TlAL1O690Usws8agHskkLgIEgqZkHCpsSPqgcFsT4I+Y5UVnxPdFZCQU/0k8Tk
LapNk01jIKQ4sJT1Nk9Nv0Hh5PLHiVC8atJn0NhTH3y6PmDFAw/150ZKu8cI85BB7rtxyMyrebVi
2QMhDYH1cFIQa1H+K7XLqNIvapSXHncxbXAOEmiPeb7jr2jT2ryaOiNUGnXljCBFNIlgrbVEU/QD
1Xlxsh9uO3tt12BqEMEr2LCThpYGqo0b7BKpPtd2M8rE7uisZ76WMTA/pNn53snatE7cFqwAJC+1
tirudCetiwe4u1nCfg+L2fByx9M0MvzTO0fgUa35y4JiAjpiMqlAGP5J3RybHZhDyXEYuLdysIwN
nMfun4rpGjM+plYisBZOqnBWKUZXjBon8N8W4KfyxkCyrONQ74wYguYGMPxi0/MoaRUCN7LYf8ZS
VN5i3bvGuUMqBHez7gaapCbXcEnptAT1ZZ91zBORW8U/8gjnNYFW5id/RIQjKm8KrK8+tICEFKYF
OyXh5fgrixwnLtefVmCKgZqSciRz/IriZmz+qSGx56ti0pLKLb4PswOd19BGfiI21CddbUg4P8X2
oR0bEHYqVY4ZSUOTDecPLOJDBtd7tlubWU4ULGBZTKonhRJecAC2Qh9s9/ehIklBmAciUP7sjCzm
iEFDwC8kJV58Kj1dPHoVbsmyKlTdjNHeQjzQmOpM7OSt/KsZrt5aXj9vcHOaTDYQQoihGxVr0f9f
3tKxJXlWjnV/0EGDTZtbttBzrKWUzgiZFLsJjRn4uHA5HFRwHdq72lAtDGAnA/R0KAjWyCqx4CyL
cSkiQ8DJ14RujKdfredpAp+ENpnPx8PeqDjEd2bUlqkspuX/MxKY7OpZKlZdcyuK5nUzOewfJRSs
e+4jfI+M6Q2zknkiXA0KBaula90MSxVupSzs2Pb3MpH4Sq5CZzI7mt0H6USDcBcXHl9uLGzVavy7
8zrEUaXBPzbJGJkZgFbBvv//rz/aeunCZCNsq2FmQLrXEQArE7iM6BM2Gda7P6ENga3uDgXTG9/n
Zmd+YZ0SIiQ4KAdsMM8Dj78k40VNxhCpHylsVe1IOKq6l5eRW+Z8AtiRXHPXBBGnQ4xTUk6e5kdW
+lSHgqNgzuQw2zIHs1lEEzVE+n2/ZmdvfZoyToZdjC/RlznhjQ2gGRnNw4FWBdpGRp6IkTg640k7
rIcQuWAeN/da/i2WRqMIJJKC921FRYEcUbMVnjtA2o8gwi8tQbG8JrO8q8vrSSHLCQqgR8Tm3jSH
ZRXtrgAOKZtgjS3GbDAtYpvxanxHhMWbPSjU/PpuPMdKH93+QA+Y+g4fmAjDLJdN2J/j4VnZoEwM
od5RkIqy/1BUXkxGYq+0nP6+79nkKs0oVw8/XUqjsBlohcztqeNDJU7YF7bACC6E5c872jQOUQOA
Y7deoJqGWtyHUce2BFMW8oOZgU/AL7jeCWATgrok7Xz9aYBz8sErt2b9mNsp+jUWbmprSHymmFtF
AMpBMVbeLxLtdKDc3em0xm7PkwODqZo4dWW6QXqJVtoGzRUxi4OUM/UXYEqLj9mGnN49aBPmbnT8
23lhRyNdF8LysgDEg3+8Gs1aq1tuQPi633+QXTKxCSJMg+VzLzCYFU9fCACDW6Zac3bwjh6+Rz4a
Mr6dGdgwc2kAkjgn/UJ0CRSw6o63w95oC/l+ZygQAjAULw28Io0KlKYV9nPUxCKTFDQdIK25j/wZ
P1wx8t1GCed/XtyzBwpoFuKzaMbeYOlrnQVaBr73Wb9kl1EwZe6ts0kvJfNEBlE3HxWICPfC/4I3
J+eOIX98Cx/YgIDayqInqfEHLW94RHAYWdyIQWUXTcn1j2uBgkFNrULoKKddAvqFvIurGrMMpm33
etUuuG09uGmRsemydRbO8sYC5nQnz8qq5ytXXGeHYDCFT4/vNCYYeoEtKgyKWcCKGKjZL2AjpjR6
j082mrRYM7NKtsIwsWRaLU5tZMUezTqwCfDKXljOG0P4TBS392/e9QU5nzo4ovnUwUpW3cPHzbe6
LnVCXwdXGQBS4Fe1dRQ24SZrhVPDOhVPzK+xtUDZ9cXKdXoL156ZFTpBRqCLiKLCqVv29DHphsFE
mpuxx1BqtK7vqiuISlxFb2Qe0Hk577dyYSq/ZU8agllf/NeA1mW9QCN317iyHItzatAqsUlGTDg+
EIFSaMMsbN6Xf/AauIMUb7aRtxpHzNQk5z19kQGzBxeGQKj8uUO2LtTWWpNrNGm5EJCRgve8ZLrA
cDmuwVSgVGdn84A/wcyDQ7CYbwo2HGBwEwtgEuvrE8Mgna8xq18yEeON2VF7EoJB6He2Yo2pHD4i
Iue7REeo+GlGDjxTywDVginqbkbPMhyKWvf3RtgcI6r2mOr2AbeWrGvRNrFdw5yzWE/w9PT5zNGX
R+iARNiIPAlOa8If7rm1jd1D+rawxjGP4gUPGNPPkphYPRS0xPyWdxm5oWI7DqxH0zzsFCpoEqYS
nH+WVQDUo2ABzx2z+nUa6udtPuQi4F+HptOFd3ZfUOqljrc35FxQrKkWq0Vvoj+At8X8utV/7dC6
0ykh8ZrZ16S6xHS4NEicFaLbX+TFk8MXX+5vPQ/pbdlsAs8asdRBO0li2RgLM2QRK+l5Oq6q/Xhl
nIhxHpZ3/ZzmD9xMzLxRux31C0RKFCFgJCGQ6tzVz5nvePw6aCDH9dpHafY5DRUM4AMj142HJnZH
n45Nx4kAFugYeGkujN7AyD0mjKTTbml4pXrZMxIoRt1jFScEUcaiHGQViBBdM6qykwMXq/4ipmvC
AA/3WmGNJwHPNVrtJb/K8xqamfhNQ66X/MbmQVwR8Ks+YhBpcvkyiO/ltyPCoj0J5r0E+7qcS565
uq7efzafL8xLDZbQTjyID3Sizre4LaS6WjNERs0O6i/6Q+DU6MlH2hjrQZBdUB3A6QLaICAdOZMD
moehF6DNIw/K8gZFfvYmQCeLlU5ibYJyC8LkljWtOixuWl6YT5B0iM7gqNx8PRYeLLNqJNJMICX8
ov0jPbZdqpwlko7w7Nmj0CXF1Z095uy06M8szAj5YAP16W4zwj6N2zq6KjgQ3yhv/0DeVZcSDo7V
WJZSZzWOURnNiyg39mfelJmZo4yrnwKnwc23q0WcT4CZan4LBVvgAnzflPRTAfFTapoU5dGUO8Va
cgtX441oTxqf9L52kDarySPVgIUGV0dhNeXFQYLDGFItaOWfZqHwGMG8hfrv9Uhpjuz015Dx8+gh
EsCp4A6VvMsVhTMJj/sPrBuZCKMAwTVU5bXKA1sWR9Rc2tLNQkhqka/0VPoBB8QZY33wrEMyejAN
wSxVPxUWzcrdA8URdmVSdDpNVYBHBG1p4292XJesEJfSQAlarJXA+MoY8IpFu0KmmQXzVY1z9bo7
OStQ0N+yKZgZtq7BfZWhS+zKnR+6vrnRDxZ55NEmR4lYmg7EZ+9xSIQs3fy0EQQj1zO/TTWdQ4pJ
yV0bViqcYefFLRGJb+N4Z2Y7geCVf8Vp4xX6kLx7KCPo0bLP3hEEwFUpIWD4Gbps2KqAkiGWTnqr
GTfj2vD50tMK6/JW6pPHNuSkkWc+X8UuMDvhjwPqd2UYTn0lSKhSxD1Nc943UyEFDy3EWWlQRhVB
T3Qvb23Myfwfhugc+33IVoGI6AfTLSP0OI9NZ3kAS3HvHqZagp73PtqppXYyeZfCqLsAkr2n9xa2
bFMdFixDoAu8/hDBTxCp7/ih1U0YJ399FmePsinv0pTso5ukTvad6S5FfRxeB/TxoLjsqMPSxbTw
NKqNiVxVyAKq/PIgwetXFDRvP1zznuJCH10nZgDdn70XW1++XAV2wu8liFaZBExttQAmMplmVIHw
MAWRWrzlaR6mlO8UxHc9uwEPvda8jrwZIIHNpXvOoxti+e2I52TSn7IjSKS0Ucr+OXc4lB//j8ky
frKVsmbTXoxN/r4sGtJL0VpP+2dgGFFvuVZRgR7JVuPIqOluHjvK7Ljjfk3p3+biBhb7fnbFYwbG
SVM5ExZ+5/K5EGkFxhpYz8erCj4MVhHuapjWR6/XGZ08+pOYoAa1l9Ta4PrZnEjpgEMGaXNLOGym
L2OQehXcGS+7P02YpRO4qTk3snWaGZBsCbsa70q1L1BLVDP06ECHkSsspidgU6LnAx6pQeiCWfs6
plaZd8l3Y/75Bp/3nqt8jtDB/+v22upKwy/1GQDw4B2i/c8o1r+6EvqRd+nxjQgN2OPmhGl2579K
HrLJEMg4o44y1Ooq7Ous6SLv8NMb/oYyAz7ZafwEdEogOxZJpm8xkADeSs2R3Dppde5jaow9RX6A
sbDzhXA6hmn7D+7q+cSh1getqXxy8Vwy9rKxZ9lKITKN1cCLoIxA9gqnKUvaqIS2lCCsGQfeqk2Q
z3K5A5jJJcwBlw/4G1NQKETCqunVyvAY1ZWLPcrfYzDvS+2RgS7jXXKDRLe2hqWveuua4C7T71KE
4SHvp/loRQTlJlnM0+GjflWbtea0vdbVyftGq2lL1VsGrfoc3OpCkgWqIZarUxbIDCoWY/gR+iuB
ZnIUIHpxyeLUtGJn1h3R7wI1+E9XbT8zjYGekdZSeUaqlBPU45w2DuQz9+v2yQvmA+DTKSWD0tnY
KBgmoYlwFItDokUWusRCgrNCRafO+kGq+cKyfXiIoCon1yN5z8XEoeHY41Rjgo2XNN4ghI4vZa3L
uutH0ld92CpEUHdI8tpMU/DtHxcP2WztA+wx9X3QNqFzvnhOWkITjOAOxs62+PeFS02/qopGwVwC
+VtR3BzDheZWtkB3DMSnJnghCB/1aVc+0rUD6m6NHanmSvdK8DtJG6QfnmiyorBweE2H5aO6AoKO
bwv1h0ERdVr2/IZFEepXcpyzcAvJ0cxgnMQSGX8hJyMsVbXKfRELZPawyvW6XSVDxr+JLIBOw/SY
gzO7Y+9f2gbJeYbS1BnX5AfF9WNQ8/5pTsUJ1rh7P7i8Jr1Msp/exIgb2bQhiRUOFzuezYmEtxsL
zCZ5zHBZo0HyH0Lr/E6ZylhlNtaxhdq75+HRH1tMVYYF8TTB2afSEVeOHOVJP4un4Hf9zlPAFo+6
VVzwrkr3GNoK+EHvDi3GLoiv0ZDgeYS74c0HWEmQGiQiwTT9Vl8iduEUKb15auG/0TK+Dfx1/ejH
JnZGT5fmHT0e19aR+ZjbF02TTBwX9bALldfNLWMTZk1QBupbhIu3Ueqvevn5xs8ag9CDH+KAVpRJ
2CX79UGY3Y/R1MQy6rd5+PAJmQK5nmm2sbF2+r4a4LA4xFwHY6yitfn3OGUlMpGoDZ/onV12E2vf
LtmyAjHNBSdti0EXPtjbSYcm/krV+HgCuO4lY64nZq36xTM0B+GAi6kuhCqrqIlLiGcy4ZVh3Rpp
a5b1pkj3hB0gvjVe9YyPTPq/GrRkiVPBd+dVJH6NrO2RP70LbfIq8rN6A0BOYGnDzsysZJ+rRsf4
iWA/tcBoI4W3Kr4XnbQwyUjgxSIveb9K795Lx+8nHHGLEHmnEkCbH7cE5h+URudGwytqpEN3dLUn
2h8vxgqQwJ8AcjxGeDfpQYS9nBnt4owxYTjA1mgDpQv0tcTvyCYWpdfF9+P/3yhfcRwj2mjZzYxe
7JGwtt0aGL8y+GYVfbYu6VoAZya8ofBvMu5hcBWaECo/rSHtduV9mL2Dw4aGmv0br4rmn0+oTZ1W
iJBtPncVioIISQCzIwkbU45AADPbcBaBIkcumb55h/DNiTwPii6ciUdhk+hBp8dGzQNXz7JqADBZ
JIsOCkeo4GwaFa/lxSS+cpoT0xSDozKzeeYjY0VmJr/IavgzNR2J7UR7ht6PVS4PL2AKo0cjKDIJ
mM4Cjihi+J5YhvhURs/bFu1iNot1uqKmrJ02I4CSp00+f+eIDIDLHVljD8NRJEsHu6ggce1QtkeS
YgJzslDcFRBxWXtNry4qtZkZXC11jXk/Cmp0BfUZeUyRFwN7K40bbSUWBf7UKy4bLf8w4AZAe09P
tdukoSYNRzYbTIPQI131Sg9NkTXUD1cQI+KB5nFYKLeN21AOCP8TNN+FCUyc4fs8OE7wKQMsMGT8
RLnFvy0s4duwOeUTOwMGN8HY2urmG+qyof/P32p/N6oRkuyQktpGtSrSSsZN6v/nvwMzL9dkKyUa
nX/L+i6NLTJHguzf0ecfKHHr3FVLed+7GftHEIFLtLtjQPZw8X1+Iv0q8EdcqzWViSIc4n8wutPm
P5zIEv4a70pIf6wcSDyQFiWgbNeBBSHrj+7AQPtzHyTyL9XKicSTjXje31zML5N1sinScqnLnp85
EHsjsUkycllAZf9uA7YJwmkQkdyjiaPBplW2XMVeTQ03QpMz6E4se/lm9/Ka9ciPGB+MWSzrrefA
/ms5zXWA9jb/3NHTU3AMJxgwPsM55zH8tPGmUctsofsEmWPBbdA3hJYFJF5/sD+0QOMYWY/GSonW
lxmRpvv4QK5qt7ljTZvbBe2O2/EpVqSMjGscm85hYUscdnUy9KsAz5hpQRODSiF2DvGORWbC6i8p
BjmWK2keEkBYUxFRd2DjasWHTQobbJwx/qahaIyJS3UGFQU33ROGupifZ+hULcMyh1pRN7xJDFVT
saYkJQP9y5Ui4aq2KurMpkUlVhTWX/FlcmP3fIbcR7yJYU42epF/AEhCBfnJ55tGZLnECtoFcgZf
Y0SwPRgXFS31sOREHSYCGGrkAUierXUELJcWt/QMcMWWSa+5wAfrd3Xwvo8DZ2u86vzB90ZbzXxO
NYbDnXCEzVtqgow7M/+YSAGn4PQgcoRuwn0+D1GCYzoxatDiMI/KiEE72jQZtfl/ON7ya0JaJI0v
tXTEIUTvRVZZbkj1wtprU4DUvNH/A2F3RhRSPQyREa7fIZFd1TYXNsm8ws1XnSwd3rTOiRzNwl0H
eS5RRhE9FVMX/+WpZQMtbEgUsG4UVw9+XmxdlEytaGe/Hj1PFib+vSs2e51wIiWuVCCG8xwn4RU8
qO5nsOl3nVngxCQ0lh6B5C+K+iUMJlToYUtwZvsW3hI8sA4HNrQxrZCKKD4yCTvUATgx47kFm7MD
ldN/jUY/o9mJqxZT9eVZ5hov+JfkavjfH5A5y+38eyG6KJCy22cNSaUNDfdow4+5Ztrq5mwqNS67
zgxYR0eUeUTN4lE8n/w6nZ6/b7xeftLdmITyDsFpjI4WV9jg6GJeF0xKq8JccKxBfa78/JW5OyfJ
ddxf7SdDIqo+pQerlWr/uwleTvXdXuxj6aUgf6TaupKwNlimOuuvc4Pxi2erW0WwzcpZHzs/tGRU
QzvvJsiD6R/4bhbDEBC/+h2slyCIua7XsNaJcZEUVC1ljDa3WWLTriyDcW8KlQXE4qzgp8WdxQPe
nZM8k/tPkJssH3vf3CXOqBM6Uo+JHbRGrCzqUYDYsCeQHQtFcO9iwkLYWWUPl0olQgEAWGMBBA7U
vGc6OluTGgh+BRK20pZFr0Gal3WVsVb/rbX2vNQlNueKPV0PVwM+sYXY2KzqBl8+EcPm/Uo4m5I0
Ga8j4IzqE2NbQDdThev+UVzP/vmtlY6VV3YqmSNyhbgYwdwMjuFJk+0ma9UFnMpuu9zWedz3mBm3
+UZlkSkFB300opD+PAlYIZsWMppbLF+sCLxtVb9EG01aI8BD6kMzq3dbZ8hWdBk0vq7LUQ2FLpUA
GsYVgIjwj3DDGH53vAfqirSxF9Y63PlGISmWpp9DnFSE5eFN06MQo8gzctTZQgvScYhVVTavXdGn
uDNXvdI4Q/WyVW5JJQ2z7qYvpY7CTRDU+FO77kBMe45SLUVoNwl5lEBU6sDKulfA3ZI7PoMePITA
ZqtS+7yrlY5mwdk2EFmWowiFJNp1IkEQ0cMI0w8p5KxLaLL3iZufEFvtvGvfP7TOnlK+ggKfVomo
i9FalZAbvQn+P6geOL/AGrGyuCAD+4qG22fndKVBvSQ6PL1rFy1iGmTgkHtHBhfemI8+GcmYaQld
4OYHDsucL5YMMub6SrAldWTU0qK2vu3umX05LenOTq4/cvRhL9X7Uon1h1TK0Ld1UpJTk9JbdkTt
uvWFPFnSdHnn1z2BHyCXZKuBnoXwXnhbapUEG0VIovqak066T6OiNvZlNQPMyAj+qiWnrLDIthl8
x+7gxAFhjyXzDKFPIzQ1aTeu7+yTWTXKoWeShD1A7OJL3y4nx1ikC9R8gZGBCYdzRxTOypHgNSMv
fd943lQmK4jaWzrvZfW2rIGC7m+fZfDMxSk3SUbc/tkO0xIwx5kdjhkLhwDFV1H+WMmsma4x2hwz
Rk2zxkADr1HIKAjj7L7FC1eUOI0rJJwBq+KhRcTvsNuYJtNTHLa8f8x1hgZ8PcxswR/eryPrdniN
e6TqvGaKgZOJlZz3uY47wJwJXVo0cWigHYSas+66fPPnMbWcd2yCN5k2LSLjm20x9VgYVRbzwtq5
MPbL0+NQy96iBWQZKU7rzFMDCCuaSTSSYhkVh1kS00PmgRrcAo9801PjrEG+rNoM4s9VE9TGb0Ud
kr2VUSMZulfCcUrrrX52TeHl8r8H+0yYmWDqd1Ygmsu9GIWGtiEPMxbCTcvEInfA3aRUpIDhGLBw
eyAXLHtIucp+YCWAW8JwugbkLHjJOxTo4IYbB3DTv4sg83jhnT2UwRa5i+WllAPntaDp6s8vqAFk
mEQhxsJ/KEqvggGvluMy3SYPpB+YHwc1bZmvObbd4xzbkTPjb6DhiAb13D08V1G38tjKm91Y/K3I
UozWvBWsOIFKpCc2kqCQLvrP/J8zmdk1chOoceWlt29SCOcZYGWVCyyHM5Am3tVI8bOi6/8YtEQu
4TdDIJXMe1Wu2UycDnk2lEI89xMuhdECTVCFfw5phfu0qbmrITRQyVxpikV2KPIcpym3n2nHWZQO
/0YylFaxIpb7cWlh43QcKAefLnAhPn8tx40t0+LdxVUTotqoN/ysTf2QFEt9LkPw+xprOqnQPUh5
U7pugHtNJTq60DXXYu19N5bZI5//Ti15RSPMxXivoI1o0EGQf0LKnykgYfzYRElvI14SLTTHHdMD
LuFDqeut+BN0kyud8qYcuYdmrgb4z4OsldrjMd81tyFtJ4LIZrQDumDFFI1ExQHzuefpGIvgQ3Go
z9PbnsmS5Y6PzNTwqQ61by3gx762xTwQjy88rxqL9+C7ZULk5A5tbqXF/qUWelp/VZou11OQw/RF
BBU6Mw59Ue/UkAVUizy7QGwKF7DEwhsg77c6fuLHoE+OvhmtFW+i1c3sLMd/s/ClRk+uDKNWDNW1
5AH+cPzM3GwS9DL/uP/1NQ3r7zBgpJdp/1VhaWwMj3nCf0Xs5IDNxtPTC8egtppEKjCDjYMufdbP
EGjPY3zX9QZYy8NuRRx+p6cnbvAt2kqSBbclcKpXGe4nYj3JGPP/JqEueNnkjtZRQ4ysmA2/6O/l
cXyE/LmTSElldcd68BguVKqyMY+RUX5WGSVYcovP+xf35oydD36w2oMpaFOyQMqvYZOn6J+dfyNp
BcRQZuRJUt55mnyGImLGmrjfjtR7lVZOcVcrEM9iBwvv4p7GWDK4A5MHVr5AagToskbQMCQI+nJs
d3mv5areiKO/OtAic6rbYmFI3v+MWjWqiDGD2BuUck+aP2JPvuKF/bWz6vR0T0oMHYGLQSRK+C7p
EfZFH54XL/4qhe+/HjBRWWNTCWdcQzGrC0Z3lG6yMF6qoVMYGbLnYm1Q6D373AzZSl/4gIZ+xscA
0oIerVHGq3Y865ao4sD3IAe3VPErL0ZMXCL5Rk4hucKrKmfaXbXFaLD4jfBOfc47bqR6Uh80hznT
NbJkLmUEKUqeL6lKOTSn1ktro39Iwn4olWXMgxsiBANZXlOg7dAe5xTDVBnJ6dQrj4lKgyguMqOG
d2cREqFRNciGhfkPqB1qDh4mBXyLP+VuFXsriLff5aDfqP081TjHEoRkOUSRwo9DWM84SYQgudVH
wwlZx/w5pdrkHemmq+713GIjy38QCRf6IoBsWJu5s2PDyP+/l4AlI3DYkCaW2mAcg4gA/ILriBkr
/wycNsUn/w5zRLEvMsC/K0AoKwtNLj3x2WYm54U9TuDXzpQ542zgd/B5WX4A082V9QfPvEUeOHMu
8L0jHtyaTG1EbSl0zasdkbzTEVY5UaW6WyxRkUNOwJwdvXEYuABwPJxOhTycoWBc/+zsnfEpR3BG
IHLE3EhMgm2hrFLxljYhgpe+4vpyNHIwZQ2iu5rt2LZc8gh5SBEW9/UQ6cpYWxS8dQSgEoeqtAxc
92Hjy0DsZRsnPde1oFC+nBxRvUm+npe+3ThP/qhvlfKkQwL1SIp35pU0sqzPwtkDo1oQ9mjX+EUQ
3lS+m7BZaOJKnApj2TtLK+OqNdZzWIhI+r+Vw/VqrlyYyU2ZTGhtHVM0koUGARtkAofLnGcjKW4o
l4ufYL4AJksBPwNbigES3ilx5H0i9KhtUtDZKxU/v3pFbxeP9Aw26VPYc8ewFqQN0KYa5RW3plBW
qMhhQ2q45Esw8gl5Nb7I/XAs5mC/RTXwHq/uXECeh+EJbY08iQG+7lYAB3Dnabsq21Ohg7uKzQTt
D15F+Akwy/NJFGb0Z2rdRFDy3djvh6rnpDipkYpvaXHeou4AzaNjQulPy0nlNOK1R70on2ktYSbk
Y6KwzaGxJBzsLEr372dp9f0gybFSjUgQSOCRvBp6tnQX62I5V5aWbnNj2aO1TPjCtQzvvX9CQade
Zm4ewnwq7og6sGYNqaSg/o7wacjzdE/n78n+KxJR6Tlg3zQLONY9N435LshbA9yQgqBUYIWCZ+8Q
0QRsmD8WtjAGb3TEyjKWwAmcDvZ8yzGGkPDvj9o0LICRbS81lgrIWT4w8ZrwvYLkRbFwnTlKWJf9
4Z5h8XudJbdrOyVHjcSCKvxl0feuwzcXT98vF4/q0sGYsjItXww4oUf+L+l7YJZnvOvogdOZBI/q
nCTw1XKOcggRjUFGNzemtNoKuum1QvwYzvmTt2an4+mZIofPcIca5nS6t/u+swzCuvXeL0Qq3XvQ
JjLz6FbXr3FGLqXbgn3NtuoIkNJkEA42AYVSEb51V/BsVYNIabhUNvBUxTQ5fh9XhTNRkzarARaD
k1kx0LT7mBOhj8WquKffdls+aK0yfcXSc+hLD9P2b7uAXj/dW0H9nQjIdiu8CxUlylbfIitVHlus
SGMkbA5sKzo2sCLHnfwwWrU/NnRoLR3lFabvxhjwRm9C8Ra0vcL/r8wzRT2uh4aaJ+JAmcURSdM8
aK91FHAbs4dQByKf7xARc5lPvIflGMDaXrUuXr1DDBeQ2zlXODKaoWGKTmAHPwWCXv/jk9SFjaSn
2gbnQocZeI1Tv48met6NFUWqVpgF7KWNofgHX//e7w0yJv3NUd+RL9SBCoZthkZ1rrFzGQM0ZDSo
obJBUPFghhQXhtT/RMEGgPiHlllT4YM8ytL1heBrxo3dJEvARDodC8Arg+IXiuJdpMN1MF1OzGdS
YHyJ9bB9lwfM8lFl+4NYg5Y9DDPjN72agSgcpQJ+IOJR38T/cfLYNGwG/xi9HCvPt//mAYynuStd
qGqPaV09IsgTg1g1aCfP2GQmO44rScLARBJ4flUjpOoklFNPl76h4opd/kscMae4nl55j7qJikoT
eioDMGBKigVvTEaeOPsd99f5icrlm9YZ6Lj50C6o3woRUnk8v1pTA/wvenRuxuJRNCsyPNBnAjjm
t8pIRUQwvm/xVx8SZp4+eJOycRSJp32iklo68wzOgZpafn8IAy8l23GdAN9JIpPr1xGqG/CFZCXI
oMd9/FCNOxvDiBDJesZAvS1OTbSnNreMmmTdkNHK1UUZg3iRI7iu2WRNFli2TRamqM2vlN2cC3bA
+Aeu1dnE2nicFEW6Bt4wG5Ef5onR3U+RM/6cjUyHlQTXX7qPz9kkXuIxIhJhWFf8raU7gsFm1R+3
hDJpQpE0tKcmLmbx+fO5TxAmw205QbuAdknBNgEI5923O2uGCfNHO5dOFt7RMq5xbYLDiZB/oQPX
w0xJ/eYCZIR+72hE+esAcqNUiV/o3w7qB3skUOPEAbZha7mQNfnZoO3cvRkcleiUAjS1qEZyWx3O
LelG9BI75hJEY2evFfvzp+CFDKealFbrL/yyjxjx/XBpBjKJ9Z5QRR6geXHM0XWC7GJTQTzxGe6B
ux0jAE+wutIesVdwnVqxxMmKReEXBXlKRZ71xQxWLpG7waAEOufnA/eD3sKeYo5uMx2N8Epektus
bVvhUhwkyrsut5ZZbUKBaT8j/VL+bE5hhLmMRCaaWaztNw64CmMZz1pUPz7KBZO0QYgKfgxuQU3z
ZfzF7GMmaKO2eMa9zoowVOYFDKBbrzDQZTxyDu+I9BGc2n3i3b/yC+wbOaA+xizIG5I9kmz0TBCV
dhlr1PeWhwkv6q1lYsdFDpSByGYRnEj1cYaHDaOdbfbB/WtjnP+jeLflzRpDgeeEW0ghEoY408KO
S42nGTX50+Dca1BRC/HLHJGN5SuqSqyepnU6razFdfgp1tZGuYTy3w4Vca8cPWSOBF8jVH12eQUa
RWMI0hP2jyZRZyaL/+o88cKM1nU2nLdpS4uKTdDCzEg+IJ2YVsig6I9JOq2YgagK07Jsy4JbMRSr
G5AEo8TWjgQ9lZ/dM+em7ewUSIXZbhRbKhH0kmg2ISNDndGLAgTbZXZrdvf5hD3fPEflQlw4Gat5
obaIqhSUXOrMlGCszXOD6D1YWHZftaOGnGc+3WDvLs/AdLM+87tqqbgqS6ww9ybLD1T8dR75ddni
q/uJpkklsMEBNIHFzlf0npBFHYE8Z+QzEMkQxtMqZkdE354hLiKjK2Nma4mcS8cbkc/7LVvaIteY
2W5TJEgVtx7gIYIsZbW2P1VSVJY3etPmvXWk3GkLUFhP6Woq0UTgnhl0XmEjlSminz1/7mlcy9RS
kNVSAQSLZG+zxf25CLsPjji9KcY1TR1l/u+CjBidoPcGOZAbOthwEU7JSfShiFIdHDFtU6xjfDlP
obWB+K7rb7kCrlgo/teSjbVxnBAsQKl3ioITjU7DKQyDuqafDYSdjdBVMD1WWUlOF8/EJphXsYAu
3p64X8yASQTwb6AFOxwXA1yFLf8q9usUHtdbRPNtujRyHdts9pY7yjnNaj59A3+bssYZTn7cJDYP
bptGsL4jEG4WsAdFa+N35wb9sHHGelEZb72amXBv/DywxeyyEfC2eVfTXoq+zI17UwzrNltwwmoB
o5zPlbAmn2a/7DN2+CaGjUhllB6EyCyrSrfZOZj/SaQqlC638BvS29OcscZw7p+Y0sJBNiVl8o1i
M+BiIfsIg64EcmimKVITI+9tPzFf/n9n4U77p4WzVAqIJs7r8fWW8jQnpU+y8M91BDnRLjghMhwt
yA4QxsLzBmZSoD7/b1U/ic0tOISWT6GPqCjYz7ocgElTKiSKAPXtZV61FWjibosxxi1t87gh6Jt/
fUYJJZwXNjHYygMf+ztplA//9jRDI42yrGTQgx82UpYdjq1efDntiNhKCxVeMnM1N6JiUwup6AZc
cL69/W2n6T+5GiRzyPdKiQT0OslnUYDwV7pH54VAiCPI8vbt19BG8tk9PC99WhfDnxoo2mpBtWPl
LTBpuBsELkJdcrVzWm6QjnnrL9Kwp9SRAZ8WYW1G+9SELFbMhJvVv8hkUtvQA+kklAnYICVm2Zt0
7MXv6fD2MyWk3DweqHhY7vRE6VLA6hoFLbPaqgDYeKvFDs9VlqwCkYYj6uPITgx0mFIkGN7PEwvH
vuy+6QhSiVIyB/3od0LQG/H/6h/s+i7kndUtxT9c7VPvEpjqlKHO8oGcuCsddHd57eqWk0e7496y
COzH9wdD0uak73tBeTsgtvmz14L4jMCaJPYnhPMRQ9COR8V3snii1NFLMIQaYJ4LaHjmyoSxC6VH
F6CLfAn2HVd/K9RJBfKvYtR+0g219+3VjP7FW4mb+K0aycgpMUortpQ9vC/a+ygCj7qWyqmQCKwd
scPYtTDCttVLWtwAtEBdwpw0viBiX5MQliLqLAjo2l1PCt+J91zbaSS8jdFdXwLjzH8njEiq/yfv
jflL7x8Lhsqv9KY+CRRPvGOc2UkHfrNvQb8SeXwOQ6eSTmxHCReKJ0ddgnvf7xmqYT7h65r9MPBp
2dE3K2c9Hh7TepHultQ7SKaqfwF1nyRu5oGg6JiqnKzLd78Z5geo8dtMs0E6fa3Uf0tHV5GjxvKg
/wIRHMkAJRv2WDLzaBY7yG6AwDjtlxwz2T+MCTMo/blAHonai4BlJxK+41GKkaQdBlSrOa7RdlJP
xRSQCsaG++2zdo55eyB94I93uDro9wsZuJYcFJKVVc8QIA6f5+6RH5RKijym4wq5vADP9Brx63oh
A5p+1Y8x2XYXzWYuY9M3Kxza+V+smy+pe0Zsx2vopXZZUUX93Qagrd3Sls6bXD7zn67Ns2BU+jwk
3o1KRJ26heR3TEnsFDWNK0LmQ0KUAs5jVkSWg6NKES6+6Hp9v9bxVvzEe/4P1sSUT67HB2SfU7dI
tnK9r6VfvaEXBeIB4npj6jIFNDYyafhy6STsRWHysNrHyKt7a2CmxDEuYibjNlH8CgIN0BjPYHgK
OiMWv/NRVCrBC47aYo6nWei5QJZ9k3dXNUVyS2FKKsKpeNvoHvFM2J79gqXoq5ZrYSEGbaTUPfKx
Hg/WV+uvgqW/6diosfKH1LP3DP9Gs78w0OHZXZuJXrz5Gb9CyWIkjtVGKkO0h4/h5QXGp/Nq/Hk+
fA6+yXSGJQq4LnZqv3XVmzZn7WSHUvBLYxg13zBkupqOu9srSFY60ELe5rTsY2Q/O0HL17AypYjc
dl0IL5bWUPDsRmCNpTATtIAhbpdlDdnub2CCwRmcqhwQ47YSMl1fCZFN937c+Rd/hxdyJqyr9Bn+
Xv6y/cHcTyq05mzr5/s0hfVIfCGg4/WBH/hvgMVcp14i3Ok2Enlv1TjXb6iQphVVESyv0GPEm+RR
lj435w32lf04AzUa6SfEIWiyjV89MiA2vnW/wYvdeT0J79St/Le7o16fKdk0ftUga9JcjH/vZB62
yA/MwuvTotqjEP0RlPokRcZ55olgXo0vyumvR7pgVXMXKn4I0UwORyXG9SOn0nIg//xwOHIMu/Rt
278uQB1LpeGbZLGT3gvC+pQVnmSGE2jGN5vhOTOjtr8fHX6eVT0slQgRERGK/x+yzqHj2oXjKUSd
zPOvMxXOImoYdRqg8StDNgZOCfaIhUzz58H83phiYpLI7mnLnwQIJHbJi6mAuSEx0Qd3/pbszM7l
uih+htkRox6uCDNmesHwHmRCPo6FxcR8/Q5mWPdL58YOu5C3/YChpxJueEedVHM/utp2bXzh7eM3
HgUWHLYpfUcMjrUo93UtFq2f3O9Gu7Gk+enIRhc3mlkGQAiSZ8osyngjmGE7dcoHqNjWo2+eYhI3
IJ/afyLdL5ChsyQEB+vD8npfZ/sd1fXk5E82ajXmZ5fJi0qh+WFBbVHFniob4sRmKn7POwcCMhyV
Fk2t27ankrZdTMbOOqVdJarIeJOswauV4q0qPErVAbgimeVS+2TvunoUL0vQW5XXgVZASqS7MFlE
TWxXOqLg0wUDtu0p3xCetbtx5r8EMibxtvdc6eU0/T86v8vl5pu0w7+Ss8BWYEwU6SAVcg0N6H4j
dgNlI1GRXIBH3hAm26/t8o97Y+F3D075HBcraru9RdXkc0Vnjb5gnECWFwRX14ZKFfBnh6lc8VsA
5qXQZfMxs1piNfm+wDq3dzhgKy0XYTdfADtd63d84l5VBBUzCd1+R/XEZc5eu7YHH5TtdBG+R1Cw
YFdKU8LIhbtWNN0fvfJB5RxbvhQrsPT7KMfIF4KeIdXYNmrkzG5rMJKE4I+KLZBbUT3X1l58Jl4r
FGdNCm4t1ZhoMxNmn5g78NsTek4C79pIXZX//muJePuvaw2nWQHpolV4V85b45vpUzl8r14e6bXg
8X1BRyPHw16sXWd8epPhxh4W2tGNEKrsZ6/qJ0rdqy7tE3Cl6jQDuHAW/grAVyZ3B4b5XNVTjkgp
rsrwuExpIRONzdmqU4t9gfYvLqqgMKpUhQLwNBQ/L3NUF2IrNpawx8wT9U5uIkm++n8v5JO32Di4
3yaFs4A0SW3ZK9VyOspXb/n9mz+tm8ZVgw5NtJ7E0f+29rYzN8r9z2zC8Zw00Y05OpnZu2o/K28O
/Idb5tyb75zoE3sbd4407oT1NN4cObx01a3GY5LrYzpUuJv+QVEn6/ZG6XiL4s2aTQKltuldL4VZ
lX6R8cEluuEeiiv7gJSVUcJOaQoFL7YYff9p7ntiNd1o4zq9/iT9Xir3e8m/CXJubx0TeugGjRSV
Eazn3WAPDFXUZjUCoAv+3pe/isoqHKUc/qMcQUgckUvfG+fIP2XO2cr9y2l2TN4VitrcOEKdbvYz
++PFjm/O052jAQbIWo8LBJVtl/anQxn+VV9N0SHV6LPU2gWqcOryRSIHLaOvKnEUPjqRZ2TMPTS6
8TORwUX0MmV9luOomeNhwthXd6M6iYSbgJ/Q/kMeOelwGfJfCM0X2G3qS5HyBmUmKsVqW6Q4aeTr
1l/IniqRhPmVzOPVgwlm1x5aEQmJAnOKDrYX6bCx/v+jTvQ6X5kEPg1yEowgpvd6kiPafIHRW5TU
StbCAJknQ3NCvmAvSGfG7NdzktFXCimR5m2LRW5uCMEYnrqg93hHFYvdATPU2xK5ASai9an2acKX
XjwcFcD0L44FcO+sLo8bzIFMMgUA6P3lPhCeuF0ARwWx7bnUujwCgj2EFNAi8mVb6R8sPD2b75eD
/wNRllhh/pu/ku/ZilZKg7J+D9rHVaGn5Sfa+QVysaYoaD2DX2TTry9Pa8pXDUG1yIb4Oj7eDIdi
SolUT8sT5B1qGQ02dJduVBlrAM82O+HJ5TnU8KKoquNHz6nIh0actHcagzgkMiljSCmmA1kCm7n+
YFxCBZ42iuEAij1Zkgfk4VmAT3WdDtvFlwfJ8J3ICXOZWmwPnU5vaksCroFfXRSbKiJVP7woL+E9
a5ZzloJggpQAgSs8w0kJKtULbS8IlrwO0YLZW8bm1r6LlRKZ+xx8oTAO0xQ7DEchXaIiKJ/HRKhj
Q0WE/aer5fvYPE4WkgVfNuYQ1ajstPclE7N1hB+7L206nKcz4Zw3pTiB0fvxccXjZdkhQJigU3YB
yGZWvc0c8LqFHMtVFb97AS6JcQGSpHeseIM5T4ULRILFAfLSLtrDcfMaUrcjs1LZrNXHWnOpW2d4
F4YNK7BEyKouxlfDbW9/OerqRLGHXy7mUFjTBLg0iNu63RnaXvIVf/sCrVSGwsMC9kHKQqy4mSZu
DPJWFGQXz9brzJfnoTkSEDLQRNA0WJ7Mnsh/rgM+FFhNtjQRGe2U9Zl7W/X19cVPZaHJA85Qt2Tn
FNOtXjxlCR+9qT48laRHDW6RoSTEAQeCrJmAcULqxXiQzUnxz/5wFveXpqNKJmX/i/1BX+5OJELY
PGCGcrDnLhqziajHgDYt3WfSKTe7m/KYVOTkYLiabp23KtJisVagjSrtj7JwJP5Rf1TjhQKwWzIU
G9xWwbz2Wsr21hKM1vVbaDa0ZhUTv5BacuFgMWqc8aqTNs7WfSxYtLWNsmD5YzSLBOtj/I5LyfPf
X3N4puzd4VZHFDZt3XwdoVng71aF3/AIu/aFllTHzZwSiDTKi9AhuqtJyNxaWeg9y8xUdrSY9rVu
AHGFTDm0SydG1N3CooBD4pAkQwnuqvE2LEoibAFvQzHFg0X1j/fnKhI2TISyYMqOcJvN5M2Zm8FD
mCRZlkSQTEwwFOnj1qhfP4YMpvqoYaHy5raVkudeVk/PLz7W3Jm4Gmo4qr7zTPuKJPVG8avV+kcR
eL/eEznTgZpTtwP+o82N/4lnDQlxi0g0QwTKosPt0eyEsM8aySyBzK8J8jH9mW50lJAykw1lPahN
dCDms0uAUND1l/8yyj+m5qhen1P01i2gHX4fi5mQ8mE9z1EhI+l/qi9finV2jXlWbdHLtLdaw/YE
VMggso6QOJsF/Oe6Ja7LZxA1dRHF12/8yLiL6vd2YFJ20m57wJyY4M7wt8TKOxuKFY+ZjH9420FI
4QP46cQdu8Zzaobny/gBSO0XoKlE91UDHFwE0YqzEcUk8XePFiNoWLnqkR+puh0y3vo0mAAc8qWt
5PEBo8+hDDUyrXrlBcnNQpY6mm/8Uhf3oUx4z/ihrTCyTD27NuGhzJoFsElSuzNkEs/QO4gTSFNt
O/R5CVe2CQfiR6IrF01nNOcHFBj5yFdhaiFFOMrNLTLymTaG6DsDQMO//HTdA5DukzBF0Q82tEpl
p8qIKMe+jz3aggtcDXkqANrQkRF2gSp0wspqUo/tysvMWGtYHMQpnzPO31+fQq7JLk0nDpY7D8j1
2/i7DtpkJp7o+uUkjWz03ebaeJgvS2twgi+3s4Xc/si4DfDEDcHW7HbrsYSvkfeu3OE4fdQLtDy5
rpvL8H2pA2T/VDxsFL1yn4EQXINhk4JO2ZhTEMk9XyRyxcvG2AYStWY8/eRPXB1jevHZ6zq0oNut
TBZ3Xlk8UTz9d6tYMDQdJy7UdWzIBQwoV0SeT/1jbR0PItRFBD2ilnGfDDQlqK0/Y0m39hgEBUyV
OmIB6qu2ZhDeSjFMqGJIZhf6fzwbbG8V+i0m7+cEyKT2/5aN3Y6i6EtWQfVYBKN7Uf3VxI4Pis9O
NXEOBES1VeieFXXCibDqimrSchqauf39iuhq1XAbuIewkuAQSw+EhScwSsGoK/bkeCRtln7lI58W
WSk7hX70vj9zp0PniV7rsmNVE/PpFMNSa+2xZS4+m4oskxWansqZomnDYv6Ye7L/cuP/PTF5kMw5
2p3S8UpCedc1aVdAUVraZJ9Ph2AVNPzh4TG5Ko7q7nxz0MxFBAWP8E0d5B9sOiq+YCB3iG/kawTh
jYaR4JgQ9N+PKoDu6ENBsgn6j0vx/NoBoorKNuGlTEHgm08lWMRhKCqbk0VcRIugwVDF5nvMIq77
I1JPBGmQwJe16Ny3cTpWGCjfzPLOAYcP960SWXpb6FMZ3SMsrt3/KQRPWRImQu1gDQiCmXHyKd4X
3a+moEwa+u3L4N6bqR3VPWaqEzSArew6uLfDZ8Wys/Z8oTRRLoxMXl0I02W8nueKW8TQs3DLS5FD
IyFHI8G+ILVtytT9K8UObuerWbWppb2Mfoh/bPd3hRlUFJf003+cQ2eOxmRRqPiDO3PWjwcjY/Tu
6b1L2y1B/dquQbiKMpYjkmw789o1m0tQ8eaPglSDQr32a13ZkyQ2LE4ILyPcP9qY9lqJhXapRJkd
o+aoXLHE8Pgi5pFYKaKt8osMP077gwOm2gcXAAqOn1hs+sz0IMvVO0c7nY+BvKIih4r+nWWCDqmi
dlkL+KTy80UfcDU5dZxlHO/2lWc8vDDvCn7l2Otp/xaSPGJOtqcxblRhQHXCZ6MC1+SXjgFPmePL
eXLoKSvHHbaYyOA3S6x27VeCNZ6bl9UlXgPU4Ki69//f3X8mZf4uU7bHiulHeUiaF7n7KLrwejs2
GCktUAP7uPCtvkYp/Ng+BtfCg231YbcwYwjaoNP1WBjB/9DF1Ky0UEoUsgsL7tzOwqbYS33fDxBO
yYl/FKTpNIR5qNNiI7P6vt5V9eJXdK3MGuMZ/ncM/wrmntdBJ9xAvc9aK07Nuh5fFy3y5boUR5Om
Kv6xhCJshW692aUUEISkNM5F1PiMeHkO9SKYC+clwE6IMk9sG0mwTjize1fkx8cNLdtkZa/IwDxm
tiRYyMOc9+fErP+HpW1juq/ezcLTHfYQQ4sOG+fZTNXNif89OENrYkfsCgrDKmeudN4NntXUnLv5
7V6LHfZt98f8MVAP5r6/aVIycMz2nYfXkTYbQKKxDa9+bepkE/6WgfpjQeWJJ+Pah+TS/DlnO9y1
6JMmi73rZqHIAm53ShytmwnTzmaDVaDQkP22UIvYsSIsDZvDOiqZoUkpV0IkTihqLTwphPCkkXod
DKKbnyjuUm1SAdwD9LNygI+LlR0B4pXUwuuwHCIuLaFmgBEWEiJ1VOSmN4dyWQfQilhJ6WmsRJC7
/GBe/apTp+A+LPUocRv5XDpFHsKSd5OXliDf36M7ZebEs2JFjJP3IP/3B8qKKgB2uhFr/llzaOd0
qofmyxgI5h8+cZekqZflpiaXGLVHwCV4B0zuA868jZSVNLty+xSLJjdowLDjwsT/FAJRqbj/VBw3
cEofcbxgxiNFWNNyWees5mcThewqCx4tOxq6UjEOyayExNAiv3ixNKuozXjREB/fHLJN2kU+eWvu
Vz+ee+VZWYkob/viGVOGEB7BK/qQOjZf7Wgaat3ajoaq/Y/idvwdsQCnlQNI/pOuJpJ7spyiYmLM
DxQ6SbB5qgySmV7DujN1hZw2quR0QMrXK22sthBrMWIKK6G13F+MRKWz29Dnkxo5mFFHar3Fv8tB
TJoKQsL+k7Cly/WHmS+xmStZYgEMJwNGdkv3jGXMGMWpTd+L/+baJjNaqNw6b4Djzy5xKzYQJlOz
RBv0qLiPEt3ctZDIBx1Muof7rv42dsyDrqloftqUuuTKVV6hmXJSptMnylkCu0EVB7KHqPg18hx6
qHOzSGif01Az5FhXMMHpyguG/fE13REl/DRuesccGBrTAH7fhbmCxKDg9qLKtE4GHCi1bp8O//Yn
fpmuIbSHKdgv2P9vJgxY/TOEer61q+irR3pS6AvycZ7EAoBg0tK1wsnPCbMUMEPjLryT76rXSgVb
3VezmPdDUJXQkNIZ1JcL89Xeo3ObB4yQTP/LLaIAsx9XeZHUev2X865G96ZZKazwb1Z03D3dSO6X
prRV+38ZcFEeuvSdpAOhbIIBBtUiDMiwHXteECm/7oQCA61Z9r5IdOMp2Gozo1vUQbG8NH4cWU1a
a+EVcBxNpX54VoB9i8JIHjTCLxmARZCPlFZlJWl9J3zxCWgZq732PWAU/+GhZHfv1KHs5KYsV8u0
WrvsDoZGseeeIAdpiGvX63ialgBPvV287/de20ta3h04bwqaDZ3ZBvLROwHpbLO2ZKvByNrjNBfA
/i8x3Vv/7l2bbqwpzkUatZr2I7leIoATjLr3+VCE44utdMXOGhKNHTuVjexedE6yn+SSqUXDAbQ2
cL6eJ6yEPMm0ocBrXFx0ojiRX0JTtU5y+BjmY7ds1JDkvHfgNTQ1QKHZ5hO05lRV4y7dEiNM/dP6
lUqzXI9GPuhYmlDxP7JT+heb5CveGYkMxLriAzJQvVbcmy26tJM/4HDu2sxRWAqbNDMfaLGX9U9C
FkBG3EICDxo5G+Ly7E43lmDuLPrziVNKvz7VStBWtvxdZQ+KdVZ1GIWNLpU+IPlp9zQvvAune6UA
u/D35AGkMH55PegkDsEAn5xvWZ0dRuW7DvhwjRwe18tj3uGbNN8bmti0rOgHnlM7BdSGXTFStieA
PNGr4E6Dy65wzVXgJH+SWO87C/LtFR+qr2BU9f9hAAJWOT+SpZdoBj25tFY1YMbl0eMNijrxh9YQ
pF/izcBtGl5qHJCO/oWPA1HgbsUm+y4we+4+XRwtPC00UonKEY1tsd0m2WL/V0JGfn/f1QSBlz1u
Z3bcwSSLhpmpwyRR0LOft4frPG4bzXC1iBZHdywNCvgvJ4k8142cmnQ327qgycC7C2GnPOidRYjZ
xxp8QSu+YpLNazg8wxyjoe4re5K8kWPIASU7DSIBtbZ0H/0rrbeRblhzcWPreUdcOQI8AUWeuE+5
NLMMjnrdg7noXtTfmybLH8HFh1zb9DvBbZcfWekSh/QP96yfezuDV31WaKzseMPdNuuIPWZEANzj
MOeVBtfP7oemmcXevIWLtf4Dj/3kZasTZlNwj+S4x6DNEReb65nECW+6/bJq+yGoY02d/VtmCcWr
kdFtRIWaZdlpXB/sbRFpjapM7ZWyQhYNNwDJYpHaMXB2EoL3uMS/KKyUch13YCUWrgeg78VhP/B1
iN8yKizcroRYEjr0nHzSWi8UTIKLBkyqhk7ebd4iQI5d29UPFvQZBj3gXa6nXTr985Jc0a/CXKYl
6Mys7ezbNhxsgi7669qe+Rs61DUCnSzr+FYtwdZo689tCi5DBKmrduk1dQL4iZ1Y1WtvA/sIevxv
6c0KkQg91qKXAqtRvDVOxwzqnYNhsQSZHi9+Cw9hHqfZDx1SfNcscGC14MtMP3TmSPQWVxR1QrDp
at2c31ceBhfXnQTnVXEI0lBfglJCdsEhDOLo5JoOfzabNTN8NP+H3zYjKyescCYBmB4At+YTGnrV
bDTxEcvEmVv0KrKK99GyOtCRd21BeYJAhvdGXNKUMrUY3KgtgyxBvPL+ew8DIrXDeiwwcpK5GPxx
Epdg8/1ZKvGrs3Rgy24Cr1CMjpHsr1afXarS+E2OIuyn/W3KqU+oZ5LR8iq/qY9+DHCxVXWCyVdn
9cCPvmSgGjomSG4iOBI8kofOXMPmDi4eOJKK/axaHGiO3OwhiAHIi7uaHNoHzmvToxJJYwdnwEkG
kP1u7wwM+4K4skgU5ch1iM5UOoxEul3B3p3Db96irxJEGaRVk7EVopGeoTUVYdCgnEPQNho8aUbY
/JhOoF2/H+QtxMEbOYRP2uQV9AmnE72E4GMLfd++2WHgFPtoZYlCjYfhKrvrEb3/PgdT3Q/USfiX
Trz/6aHXPoCf+kInJev1ELCoHXWiP76K8ysoSntxbQdVwC50CNkw+P2akkCU+wYmjXRS/HrLx84N
YrbiCqRoNv3xncSK7G/zXEj4/8RUj3P/JMxdGzEspxjFL4yejPCvkci1cynF6Z2MDo1j35qFbHUI
bUAOVo7dH3hZTP3kNx8i54v6yRZSETTgvPz7oTRBKTZwi4Cljj6o9VYLlFEt6VjnDN/5exW2IDKT
hbu7ifxHrlaRblqldJuu3B+M5bUIlMUmNN8EvVyiPXsqFqI7C/16iDuixOdx05WvxaW/q/rMKqV8
nLYIfc1sZ/MU/6s5e5boNIe+5SBLg/Ho1JoobM4RInlhSJZiDtDthXoOLcl0U2oFwbyIyrtxVSQf
EI60+WlBVC6fi4Vvk/kmT+0fL5WCSPy0qUnHhphLIxsryWu4pylYIBg4UaSmpG1DlV8TYqE8R4Pq
NHlReG86OsLK0OPdT72uJvv4U2bovDUjY+HnpRAiQ5dTTc5KNeJRxhHuWa2bjJRjrWdUdqCSA8+K
EvXffchbu/ekLoHjfnd46f45CWCrl+eSR7KV0CDJAvz1hBBudRcOE6Vo8P/mevmJF59yGjoC6kCF
KwxGojju9W/cszitU5sN9z7m0YI+zYxcDNP/KE904pK5g4TbspEsS50ZzM9gwk1A8yjBiJ4IfMr5
ofs7bcG27/aFH9fHZUQgo2LfD2gGKB8XRMhK2nosAgijdNb/bBN76QA1GEdrds/HQizVJcup/pfK
K8mbr3lEAUdlxI7J49GWTI8OcZ1nVZ0hZvV2rg8vyAy1+lJi+nvzaoFShk3N0TTNE1rTBBPEUR6k
tA0acU+2vffeddvjEajW9tgAmE5zAw7f4pKqAjFhxdTox4EzszFr6XuIgyrUM4LtzDnnULeMXxCR
T07r+jjG2a6VQDa/3/l8u4dC9Y8xj577Ibkn5v/qDIzG28EPv7sBGSPzpw6td/jchwpJw9kejDrB
bBfjNI7Lbhs/oI6r8MqhxT1kZiEfckZuyjnE39IudAbdj/ZAHRRIjimdz7D+QibxQK4BB4C22ydi
nEJhspEs/x9/vbKtbFCxRleg3NT1D7yeq9J8RnmEgH4GFkiH9B3Xv9fOvujs4kfQnsqbAVuQn6Gp
0COKnvTXLg6hrOb9w8TGJGanwrIbNsjWUkbNz7uRnvhi5L6rRT3Li0yNTxeiyvV0182FQc+W7J/y
VNTj115+dtTqNVuzPE3ZExgVE3SrpDS7+hO5Qfj/r4AoPZVRhY2H+cCtUKPpwMB3Ya8krzInKkLh
VA5h4Us419FFR2IoDBUyPgJsmfq7EQnaFGjN1f3HMYs68hSDirRB70+3DfOHmXf3nOTg66cZIcjP
qZgUXtA5fyl8gLRfbGmlG6T/zJl/ycsPoZ53HBflJS/LLOggrakLFgrk2c4YoPB4qlMirFJ9Heon
cwsYpN+9hrFMIMxELPFRW/LxqdRz8h9tY3H2rWOQLzSDJHWhbWB6BYfhGi/AGSBeZrG/5GTbhGaR
2ngF1OM6YBDCsZRZw/s0WGquWo5rZw/svNCaC7kQUkCPC9V8xk2KX6cuTaFhZ/Db3Jj2WgEwOvfJ
cGcnf7OvqrSGeJyroh7e4ukLz8WjhVTEc9pNNd3EobuG65Dl4Mwo2KmlDPlv6B+DvNXep8hPsFP0
1U9vgk0HLNFI7JCN3uu2Wl/S1S/t+j0ghuQbI8hgB57/EyPt5yCJfydY1hdA4hpFYwaTW9PB1f+s
/Pp6/+dgD2SKZNMET3YPVjPGQfAR1HlX8VkKVutr4KKjXySPG7dX75gp+fa4IEQxDOL1O/U1ciaK
yxI1Hw02sZTkTqNzPBRDMRnh7p7dX/jxexq68bxDjQf/AUSaTnYP0UHrWhFIByqWPIt4LrVK9q/I
uVYWMMJzEj7jyk9fQVDvVZ7X91c0B9ljU4HTA39L+Ytg6v6sCnGMU1Sz765LONZtnA4/ktMVeGw0
Sx1G7Fe1DxYCbCfTKZQcsgrbTPJESlz84t4VHmvCKATsqA+tGCkMa3LMcD2ERncv5cpWqv9GDgU3
qgN51wW8Wm0Wmi1aARSZ4ica+1+vCkVdkjJK68ISp1cx9Fqv+2P20Iuci3htWSXOvSSdmGvlB3Oc
NgtltlyZVgh7J+DZOxl8ojpxwYQNKhRO2+tAjq2XDEs6qb79VojhwTT+OZHkgSy3PE8BNX3PiHBF
igjTdmTqxBfNTHQhEaHs/N4ZEE2FZQhcQTF2iR/S4aTLJqA37sCe24ePd4b2XuCFTmX2I+OuahTY
p/QOILvtB6R7Xwa1kgV+Hh3BV1VqvH0qOIHn4V+sJ6o3SGGx5RGI1VX+kScD80nVZGeoKLI5Pgzo
19OQAtKJyfStvWXlqv1+QxKDgw5NzvED1G18uYLJtz882xViEhZaxaYBNcAcdWx+MiCcjd5paIng
O9XgIg4rpLKXwpBovLYtvccSyIYsaPsspBqgIpLx0IamIPrKZH1IJ3/wYqne44+Z1lMNz/oD80rF
X+U/7tP1YezozdfbBi/+0/h22kzennnmmbnOq+NJNJW1taGT7Kp49Cn9sl4bDdy0h6xQWA5nT+Uf
uiYv78GTOnEuxlbKQ8SgDkTFAta17ohJXZseAYujkzHv857vmihfjfS2jhWupapQ51SV85IG4SN1
+VOEAOEJURXy4Bgs/22+qLLAND5SZ01TJe+bbwDAoZdDWL/r5kkDy+s0cRjTl78rR5C6bq8LYcSO
z9IFgBGyCDfQ9kFvYjMaQdd0ZISBZmzLDwdfcNlWgZovZws0NlvYQQEGKV4VKZf++SZcbDsA7KYS
AvlMQhoGTpWZ6DLvEFMmcLRd8NMku2CF3gK1fYkJauI8GX3un6vGfGN9WikaH2l4E5CtSeLcDizw
/Dq4KuIG9tKpcvl8DU6DmeP1i4rn76OVVdoPrSeTaWodzjsJIwECTotaI1QYM9FIrnegHCA696Ao
vghf7+R7AsmDF+9aV806kbx0rvhM8995XHVcPIhTUFOHcEHgyZnC3WDvzdHP4fM8KthGGHNwJa1N
ZkOr1zultBSdDTfbWCAodjbEByVgPsNJi+E+1KMYb/uC2eg1Awd+B2waoz6lK1E3o2eyRV8+2Xsg
3pOwEfRTmRfS7NTPEq31IrkC9whSY4qs2B1XgNT7u7yvOsg9yiMuyYs5BS6a0QX3fhm0NmqJA+kl
/1D21FYnNPvLQ3dFVR5qX6QIulooufWuedGsewH1IRF4MDmBSoif2EuJsM/DABYOvxPodsC7NaUw
ebXX2XSR4Bvr8zJahO3A3R6SOR9xaNt0VA1EMYYwqFvzJPTJiaU801/4PLTWE2OXZ8DGKHvRmpYn
W+Bs47BDPhWUn2VYIljYoHj75yKCivdxAEqg4coKV6vdppi62nCyiSZh2Jnria94cmrS0hm8bmg7
0tC6Ev0rYOn8bt4+aCrWslFHkWsj7vhbHIt6/TynjSFSmw3EvSD66gfOW15BPlNFs1CKgD+sCfKe
kSt1oprOz3/Z7r/LXBYO8NCc80MDTjEMQeLTHXRXu1qHb+hqZJLKGiBz9JM7eTaWs6y48tSyD0oX
aBcXooHCsdcc9FYwBF6vKf98nEhwipAup97gonIrLGgWCuXTDau5j2UEnIQOe38+oKyI2wWtn/+Y
RxA8XMSMumH0Gwi+TOANfl7iiXw0t2+6K8Gyg4Jv7N9Q34NtMD5cCsUFAKor++Yrb+J0WB+O3D/p
s+PM1x2kamE5dyldCZHJoIpzBhVNImXe3bQn6IL3h8LOEO86ZdWC0mXpnRl3fK6VHM67+QG3wp1I
ZDsZATzh5H0j92/feWdHJyB/C8G4CEpziLTENZYsHyHw2QC5Id5QZ/z5MnjtaRUOYALcFjlRnCHe
cKC4ETXhd1pKCdUi4A29B27ABTTw2iTUGvyLtalYU7snVeu1U4pJNYZDjVI5nR+XNK8StuT+zOAS
dDgucakHmQJGI8uF9bm5oMQLRwBhZYQHHw/2+35KX15DPdiXLHf6VGU9ZTEBgzXX+Ee/6fKdwiJS
OlJ6gw0y+KgGMhK/DYERRwMEHkYW7gjYz5l1ty8igSEHd9SlsDhJRn+WdOLrRAdgz2byPfr9sWm9
ZgPNI76DpWx0Z1TGGG5MvbK0pjLN42y+40sXg+QAKuiE/Vx+sjjXGgx9eulLM1wisgOnYVMUPpAP
+3dZRWk+oyIZUHHxB5qmvYT/5nkRfKTD7ZBJsLrrhMevSgdTQ5MEvoj522CAgcytyPqG7LuxdjFA
gAjOuutR0JQkYuHNrA2NaKPLrzW0Qhpxsn8MMNguyOcjIN99I6q7zjmMQvfrkDNTUAoQRMlIjaEZ
CO9d0DNczrnIBIXA6igkaNpcC4CnAhl1PJuVbO1GtTW+rFXI7Ti5nPKUJEC2C2iUvlYMW/HanB2f
bteZUPEg/QlWS1YB7wOF/Ox1O/FVT13H0p+pIbHp0eo5vex+l+Jvex5yl58VYpsh5VfVaanZpAKr
xe/COqnqbihpt9lVcLeoIwrzziY/rCgoxOoNxwQaBWzNB9eG4WU8ejvdwdKkuolzOOiJ6oYasih9
bD5KMqlMBLr1FhEc861tifxOmcCwpBypO4VUfA1lCmNmrIbp+YscMkmiw834Uchf5NZwMsA9wjUj
FYow38MLRn/eAyNc5PWbC3jj/yR0k1OebW0o6o46Ity2YVd4FnKCjPTijYvJ64UjPK80OyEmZ7Uj
MrHQGe9lBl94RymdWCX1mBKEt0A1f9p0dQzFyTlgOkdl09Y8Fgny52oTQTI1dEdJmYKSFpQhTBdm
J/c5Amrn+NLM5vHUzCjxyf5xqkS94k84uhytPsTdnzdOt0/AuF3D+iGwuCvCNkVON7Luf2ZraYb5
9VFpZdo5WRpM6ki2ggfl3H8aijpkYsMo3D8F0B9WnuNnflieDItw543Nfc+4P0kOTF2zxQ5Ii+o6
0N65zWTk2eCi+YqEUB8VaTfJ1KDPBCPQicI1yHtlqc5GTWvrUqeGqbcp7sueF4/KY2GRUg885EFm
tHoLSjtN2kMWtFiMVav4nUSK/Dd6qn4I41qAjmYHJLAKhW2b4UMeCuk/LzhaxkOHrsxYwUBftyNP
dqi6xpdu/XsUyRg6i44d2qo2UQ+me1BH1rhPLfAAdoNFvC0kCVHh8R8xUO0r5jTXuZcx748Jt3Ks
HaugB75PtqCsMO3fdkISnTC5pdKYz//EJXmVvvxV8PL2WhD7Ma1vqzGxIhWweFJ9OFnqQKnOIg5v
GfdnoneVSW3MO1faSngcBdB8GbsGkYFTMW1gaRkhsoXnB2T+7L9+WHFK7VOy2Wo4a+LhR6mlrRCR
1HIy84gmTuMl6uxzBnVEH2JsWaOrsB6SKmAokRseFgRawrT7gN7FPHdw/MXelmwNo/bvCaPwgqTh
gQMmM6Ox8MCrclqL6eHqYREpfgFMEyTGX5Q8drv44YRGQnOJuoI1tW6M/XlfNxWvfTSTIPvQK16I
qFjV5/NFnQV+U9Qdbsh2u1eFKfq7xGhhN3AAVS4SydcIWgBG3WcOixs9gz4uwLfxOfT4KFmiXjQf
bx5VWl4r/g+Soy1wlHy71grvGWgN9KjuTfkHcQsH1VKbaJFA8t+O5MQuP9aOFMDGorQzzGFhRK49
AYK2OkCSSbGtboo4CJqLpmruAkclk2lvTgX/knpbLxN4x9D3CUjLfNd2UJBzC61oR5EHvmW21vTX
B0smEQxJ6deUfwc6iIF6WpMsDxhUN2GxyB/Vys4K3/PGhM58hFuXC4FUOxm60QEpkGXHR6CzaYQ9
Wo35vWh/PpsH1PuNIvO6ERQUXhciiIUSwW0caYUhIPV8yKeU+B4+eUa1O+gP5icnHqz48sI31S6W
PjcJBSCaMGyeaNveAcm93ZoecFvICDIntB72EMaIwYuDwfjywoJuV0CDQi7xSpIEd/aKOiSBrTxM
ojkJ9QsI1ih/dF7YSPwWPis1BjgjXtOShdw3GuoGWlyNgIui9xQZMppaQ4NRlsclz0CRvTRIinZ5
4s1DN6sXoRn5oNrjqzMuqY3FZs01iFRTxbZS7/NkWdb9HuujOnHkZpY8hWfFmhEuJHLg7eOzuF23
/xszgJm1H2zL6o6TT4f55bheIH/Fy8Ntl/BbfE7JWlfuhvvgSMk9dG+buGRqbUpD7LHna5N6iqri
pXbeeH/pcO5mq+r99nn93pnunGz2AAgOKpsPH3rv9ECLKiav/30FYTsayibusdy1mQNrB/XfMW2H
+ZlJ7l2jGfVYl4Nh2xjL4rZZbjzowg5Skc3kBtJS9qY+NZX58sZEe+zcWfpQ3ub5p1XKYiG5NPUU
qaX4YTWn4kIxlJLXT0L+gyLNQd1gOM9OpZid5f9URwl2OnApC2fvoivak3ubbkY2YY7I+mKGeT96
HKnPSJ5VIBOMXDG+WI/kDTLO2LV54PBkCMlw1ri+DFsBYpXwj+APrPlW+2pB3wNB3budUlBDpyeX
4Gj5RdnGAOHwhCJRcvXQkrqafh6OGo3sy1iWcSBqoQQ0F9HAsdHkBVV7y4ndS5OI4pDl24QjMka8
ZYOy4D/wimRJqhm6DjF437VyM3YqZMofHXmPsfbMM/ecJmpGZLJNSMZr4P6Ar8Xa9lPnazSUCGyw
Uo3ORoK2rthtwgOvzrQiUmTaC9WZoh8ibfZv8YASvxSOxrwsD8jbhj0MIRdzTUrnCoYShYZ0xSlI
jZuc3E92UyXaDCyQz+AgCu/6JGZ5wQIenhCQj+J3bkyQ+wrMZS5nA4HpPl09z1lVbJ0IBwXGT3P0
YmkGYSNpKpyzcyf4uoF6OwQTuuH704V79MRwI+rXW6q7WVtCTdLAU4GLIEGQX2Oz4ctbqy9N6ZNz
gq2Vw1GWSEktXzX9BJqvhutMBVgn5USDWiRGc/N8ryLj1eVRJ4NWcBR5B8dIcQmr2dUAC7dml57D
Uv6/X5vSEz6cJOUbnQe17f6+wUWcxqDGHMyUD7hrXv3C+S6NC4v7EL9yax6CTfV//wqn7AF/jSQg
nyAPmxLunx0dCaRyB9/nhrYxOKoFhl1VE2/jODD7FIkGF4H2Q6nkco1iqmqcfijUCLQ4nChtzCUn
UAwx+6+b2Xy1o4oJE8Pvt6Lg6gegyLucnUn9S9RXmzvKteNzWg5mF14WaTSYeA9TqDMkCCRmuX2W
EHKugmhLvFMNvDSjERYKAIGKpYENrDPccV3C61beNkZnP+/JlSMo1qV6h1yvp3fRhDxIQiqOW1qh
QSpeb8Z1XPJrcMnMsbCsjTZwdFP4gicBn7AqvcSg9Y5ibkqFt4aj/jTQdtZ8Cbw8LEXdrK06qzp9
n66dex67x0vknnWbEJXDY56/Bma7eZuZ6CVCKxgmceYRyHruhh+h0ZkJ/3NjId8vKMOmVtxh++hF
aAbGrO+0Kt1YsnTEEq0s1zICeNSXI1rPlAmYPmDdfzWyIIufO8Fz1NCd9XFJiFK6vc8O8kDRsc4J
+30+vVtwvik+dnNWnLyaAJAF8w1yKTYmFWO2GPvgSHgTnONPPTlbN801p6z0vx/9BiMU6zziWYAS
rgSDSqRCRYgoSD9nOl25fqRDt+Cq8nRdOjfkPrWx6miWKNM6SkjSlcJvTI2Uphms/N7IVL2oZydR
W8H5bPonbGky8MaU2zEIV9kfvRsur7MagAszqAvaUDEzPMtP3txa//4AlgOuHn9cvvL+cwKgdoSN
VxUSUiL9Q72cTKN820jsM+TzYjd0LLx11R8pSHExbdkKDY1XBlG6U+yX24IrooS64nhTN62QqNzd
NWLVwQrxIzDlQHitRv8Sln5JLxWwuwHM5A7PnPIP70Xjk/S/k4IUg6E8W/BztG/1UbbTiQsP/clz
bUHDhdDtewp3GhI9vC4Av3d23EJtY2+FQsVvjn+xkAMURLheO+GGOJhOi3BxcI+yZMU8Q1AlQJev
Y8nF81fn15JTgBSik4gHpEMqleZ8rnY2FNWlHKk72a5v4ad6WB6s/ezY7RKIjQkflU1xZThLgtxE
fakOTOJT7/wty4Rg5gNcwHakCSS2KrlDlvMYD4hJsGa79nbnd8psi05LqpX3Um2OIN85mTEqmNDE
yE4nEgR5b1+8AwlNpDXqrc6vTakIZaTLQcrP5W53bax+eg+7Dt2XbYXW8qhCeX6Jmh3rfGrqgxct
HvyIp+5TxMTZoDBNaOmRo+Ko1lSYYEw7D5FHQHcO2QNjl6rNO9+ZD346mC4zcBB77ZfKOC9bxOO5
EAFmI4+fviQXUiMWwu64NGi3bpO5k1Xili7j1+04v2qEG2syxOchjXyuimOLomP1CDZ6e7eY9bUa
glZ8c2HCGYo7dltuNeQ6eU9A4fCVvcoTIBbtM2Zy+W5P6sMSKbSekgqML3XSjKWoTWm0t3pO4zvR
2uqgoA+XwEj9plu231I6qSV+8xYw3xtoOaFynwhU5VlGGC4PZpbbppi0BxgpgLe7SIuspL2ncih/
u4pgGoovPTxQzpo/m+T65SM2yMWhHXs/aAhHpS/nXlQ/m5i4rk9pY5H6T/G8nrLssrkTMOGl3mi/
JSpRoGsSevk/HmFnsRcadI1Krmz60rrQm4r2p8VVWyHUBJ2gNk1p3EUKMU447kiVVcdOJU4tvw6L
g8gLYn2+BUGVYT8ycBdBWJ1VNltPcFMiapzbQjxo7m5x9Y/kww4vg9OH7QJFKHVy06WwdI+af2Qt
S5mxeB0pshNgbzPqBpYra3RRe6WlBGtzm0o1xJc8eNwOqEllOoeMxWOzHpY1WyU8eEv52oBsuWeo
bep7SSy6SYWMzkWnnifsMrHKLf+mEUO9bO+vAoW+eJvAwl/GTq5D3yd4j8A//LTzMajcbAHH4LXJ
xwFDD7/+QWPg0j7gZTgzM8hPcwn+xLtJaynhFE70ZFKwBBWCDEC3aDbTOGI/cyQ+o5m/6Qs02mPQ
SgTs53UjlfN2T73kcrsWo2nfy6nL2lqz6ug9TMjJk6T4Dr/O/6HPAe5BqTgsqL1x8h3Yy0wPM2lL
Rsdv0MaDckGSlLz8QCDdWkolBjlP3qZdWwslkj/+N2UNFPYLJwvbHwkU9vWY8tksBZK2XOmO8sn5
ZzOqPIcUwMHs8MCTZLDcU8qFBxfbnoCSu0+FIXlsBkxTyfmEkuqCW8iUaWLl5NgybIl+2p9XVUPZ
2Mr9HMgUdNvA+ALJpqB8wXbJ3AdCrAs9acrIr6iWGsINoel78lGhZoccz9P9x+lX2Tg9KVKqraJt
jF8lwiCpXG5sX3bFnt3RsMFjH7kBG5nYU0Wmt5efQ0waQo614nEvQBItFl/8BRgGBlcLzKwLWCna
X1rP4KOZ97RRzXu4sLZUP6espH2mU8gULwzmKadGP5yDKk0Dk6rn6oE7drIDSQ3pFiuKvcQExq9U
yzPZ16c9xVStMJMgMxX6Nyyd+2kBfTCJzIAwUAwHLgR24rwDk5O8XAdCny718M7nio6ttw33N0w1
KPcV8zYuJEp6ano6HzW4/1hSfG5dp7IGgA5FDHRjKL9IP8p8iAvipRitnSZca0WWNc9ApDHqMJ3q
Cecb8eLez7eece4kHkcMl4jp6u2PjWahdIkA16PowrXRqB9OToiWCm8MCgVnMbeWfHGCJL5RDO35
lUtD+ml3wHGX4itEXVZMdMWw5Ar+gNssD5HWiHcIeWiqrOCVBw+bUE1HHhWBTlTcGoHSTGRrFUKv
xG/UL7GUF7zkb/Zw/+zd2OVYe30i5lbE/R76Mu61nf0CCHl7+6JdmZQlK3EMu+HPprUa+BZh/fjm
xEtQ8W2NbmsYX+MuNzIvd5P0YVuNyt0FQBGuglfImLPj7WbYGUSuTGiz8heNuXyk/9otRGiDAPax
cObbJmNNxcYgJapozUr7jj8agYVefz3sOmdFWTFTgjEcDlLyemFJtMVyJMaj8ahHUSRrmDJ9rLxs
pE+nJRxpIwAAM7YAeQpd2Gyn6FCmPg9JZDZHVWiRKrECghu/Rvouff1eaasKt8UpgeNkTIQsN2Os
llqY4tm+deMqlZ/QedNOtz7F2irv94aCurJP+YgK/zypE4j//7g4okhG7he24N21yxAuImNJRty1
Et1fC/G3Db9gg97WWBqudc4CPs+Cf8FCNdhqp7UiGHq2p4m4XB53Gb0GxD2Xxs9/CuBTPnghs8qm
7LCpb3kPfdvBpkCRCBJU6MLfXk0ZiujNETCUe47dLxuB+3ns7k7NZkNhw/gseYuccyV9hNw/D+OM
N4Gu04ooEBAiWnP9LagfAsfraY11+jY3DOaCGggOA7p3pJY6gYbx93iF6oMPNFQ9iMde7BPIl1KB
Sv/fUugKT0i/mCRQH+7JSxY4MQz+L0gSpD8YE1G9vo3F+n+trsTX6W8JWIeCWAkrd8pEa5y6QPJt
ohF/jefR0zGRWKU26c7dFHRrwbVAF2Da0V6zCg3I2xsXBHmXI2ETTmo1daIvMjENviiVGpfr6640
4ZXcnGUv14OvIX8MVwBmt5lRV7AIC1JRGaWmIPlgrM7gV9TjzMLRbKdiO+JASY/kKCpIUQPtf9jZ
M7zY00ZQzj0s2gVLEKIYsfMIpwKfohwu9wG71xkxaHiwNvZp+qwAcU+6jN4t6/YREkl7pUhnA0w8
ZumRYmZy9euE5KQAlnoqyP3Cwqa/TUUeFSl6oeeKKBr+2RlIQr0JFihxSQJUNPuIEcFa+N8kZHmd
hwt0nsnQaS9dkoLox81DQ+qSBsw2Eksh5hN9BPQ8B5OUvmo936WareWRjXhvBJFdlC6qcXlBgXh4
5qtxlMfduYiwrRS6wvimogr4K/bczVz6lVXadrzU42K8aosn7wG08mQikGVB9SusoRbG9EUABV74
Ml6984D/RvxRRx4y6NMpJZudpy+X6hnw3k1tY76pknkdlf3t5Ahc8Y3idWYPVg5DCsz6Ics6Ubyd
vwFusddC6PdldmWyflFIRHaBBRJqsAE8xJoV9SLM+bycaA4fWIBc4qU6FXXfk+9rCzqnyrTJ7MuU
QywTX/fl8l3t/vEBWHpGxGe9EUDY283QTkmt2mz345iIJtKC0DwrHRI7ZjdrKsROUZ4vTvsjV7yX
QwcnrKYPr+9lEU4jKmCwg3lTGxRFFsmNvSSBmOHb1u0s6rbzA0w1Uqgv2Vncx619mtHdh0+9vs5g
xovpE9lPD7ZhJ3LbI/MIcYRkCPhxGa+39qDJ4kiswWJpHSAsuC7zroe2d8WFurVP1enLA4qHlr5q
mxaY5VkyuiBdRzV+DP2jmeUUUl2PAZ5nVqu78VysfrZkPtyl+Utmm1WQnfuM6Qb8teyKbosWeWWh
kFSlZ3sik6OUBPOFfLe+H4U7PVlmuVkDltOmQkEJnYWGv9Lzgsiw2V5ErU94nEG0r7UrtM1kvSmM
rnBdsPnn66yXMYjEaPD2XxHDhsnpfulYTdAITZAsVptst/MsNICJ6TCl9TmnDtsLMBlFTRLKvHJa
Keny6HdzoYH3FP6mmRaf4iOSKf8w9f9PmN23iRTHMCAs38z5IakoPLWI5RcbHpTOr/9Z/InOoXgz
axuYnJEXejyjTBlUjSfMukK1UAHtsxi4jv8UcblecuVRN0P8rVoSVgLRHDCYdde8kvBGb3zJIUUu
LuUXKKKCpUteSNL8oDDzInpj2uUSJG5/zXFVkRvANhNNgxwPiPMd/tvFWfP0ytvkXMeiY7cn1VWK
tW2IiYEcMD0w2eNgP93cLsoaLAeXX8qBqIlsa1q5NEhI5uORmLUMmG758unm/nWvDJqBOei5e8Ta
L23geFfKy8nRNpIvX8KF7/42BYBA0iFOURuVfSzuKJrwv9oYlcDwWWZvT6nochIRDrH3AJ/7quda
7At2yVe3M3hkEEmoI7GH7b/Dd3m5LU5s+HVQtPftGWi+EHA466ydDlV0RAfStl2A1ICwbDgfnyQa
TkmBbLZwE91rMFTWxTHTnCMkGSjv8VQmYqimCSj/TYlqOJutVO8gAd4zIwRlwGWS7TmrrodTSYWH
c20KNjdN3pP//CRuWaf8HFYJ2rYpX2SD7ET9rDuyyaoOhNHM0/rbyfXWZdXJSPtwOcuHVwelU85l
tu+SGgwq6urOZyLZru1BGwiryowI+1oRz+1ExPU2FV+aMMRSdQOc0FgsFihUlXEqFD/JppxDFgt3
uVbBPTuxNhBK78gltgWE+trOCV/BwH7BPKvR6+mrIQqq0Qq+IH8cjiF7apW0AM8NQEq3Ba0jZuRP
FWMOUycjGle1541ryWCGehbneWV3a6H9wvgERqJD70hJHVsELws/8zp1+ELYKxy75qe2elh4bsEv
NJNYAEPaVwJ67hEns0jyQAKYxEBuzVPLZ4ks42Z9srkZM3dMmDLdmQ8Ey/avbngkMx/n4nrR6xtT
bS+pGqvwdI3IzG/IsQnEAc80lqxKlvI0YwqCROhqYJYEK+p+MKVTKCG3sSSJGZl2qY2LttGZDVke
Lmy1PF6+iB9Y0B8a6TqcaYO8uOdI1y9uUcvuqpXc0qofMLzlyPaWZ/nWewhmh/cV3Q3wFELurB66
qRs/dEdpd0Cama29bYsLWPQRv9ATKbZa9/PyAxZtqrZhz8rbT+FgIvWo1VbebAT7dtcxb8D2vlNP
B+RnOd+UlW0TtDQMlKtrhave4S6YDAtBV/BiwO78SwpMgtcRqGKU5P206APM3XsHa3qF1zK/mo9R
ZrOKQY1a7Qvd0vVnLPAD8e14Oc3cc3D5i5QiDj1m0/HR2iCB/DwPG3Y+SvolqaD8ngKlYKeXvgaJ
XmCEzY5mjf2FAnNGSFNa2ssLQJUAC5vgfgCR2ImGdFVe+Fgza94/6cCbCLljwzyodCR8VxAjsYeV
cyATqLJet2AyeWq2dM4gSJJRLvBA3S1DdwySy4NgwQT0M6IR6svlSzwp02vEbe6r7KPAAfy5MLY0
oqYRyxeUy97P0gehlc6ufPpHY1B4CIPv2n3/3b3mkOi7HZPLhzKEVdmPIV/mnl7QsH5Rg7FCUnLR
gEChqLdh4SU5A2MK//wkSakfXhjWDrXUAdNlf3YVCq5oz2wBZOsTdCcQe0Ci85au4KNL6OGbFayG
z0P/P9oJZWsuukBix20BhltNcBqqhqM48hFOUe90ty+rMtQxxfbmy3HND8O3lrej79Q5NM/GDCWN
gAQdvFtp6HBr9I6b9qYtJpM7rQ1CfS5x9ThL8rEBidHrGKheSsrcX5PswJQnaHoH9eoBrp7DV3Vz
r1kEEPXvXD0AwlzIo4P7FaC6/2dD76uvql+nXkYJF4Ts/E4blDL+QkSW3qe92oPeHV0TegyFwZ24
Gol+wsBk03OezTgjxBgs6xCApzCW8R3d9fQ396LfzICtlnnd/0njNoJH3s8XVcUvZz18w/rHYO9t
lb4HsPp8evYMYNhWNSn2ecYcPp8MEbVPooPCfgCsk+PBxHMsw0+OQ33n6cQcMCz0hM3TzGYxttza
rdQyCz7DMtQQR2ag/23IGPixhZ51YZaJa/I2m9uIqHcTOd44uypawOH889fmz92v9l9qZvyjLdPS
4+NQTfV+YKK85SYtnL4UJG12uxLFwM2cPpzE9GqSPdQuSyJT/Yct+5SBh3Eslb2roAZqxX5LUX22
VXcphCivRin/JF9iJ+9WFFLSBuiPKVxwZI9HZfYPssaieP79MfnW9iyaGPMTi9Fy9f9BCIHNK/x/
pphKkanQuVFqR9+QkQ9tecfAoyXmgoEwyjH9Rgmig9/QrTQFbwLfaCII2zlTrMzEn22Gu9WRt/hq
EuyeEm/SplIrtPDNan7XwVGBc+LbtIaIQFImqSmYHlCTtTwVDujtL6e0Ib3GIjtjVwELRV7imOin
+CgWMiuFzoOxiQ/SGXqGk7qPRyafYakzgQsSGiDS9FSYrLhuQZvIWMCbYrRjAdsBl+vfdEYheICd
1wKHtfpGySu/rZxQAjQT8Un/tSbQZL1Ype88EtIYujb/viiy7u9+lUpIIxJ+EaZqRFOiQp5+A4Nw
2Z9NbCiHYBIwT9rN3I4+xaT7F01I13Qx7vKep5dyN5nnDf2HBy5W/g4qwiYpOt0830uFiuQ5XUhm
3XP7GSgghLgkIVgv9KBUe76upzfS/Oc/suS2qXvubLhlnL96L96NxMPn2c/yDgYyLPF1FcIfEu6L
obo4fL6y71kvc1039ReZIP4raX9b/atMHEZ4P5EfWms0N6yA1oPs5MczUK7cVz6WvglZzbzdlxAa
hH7fqbMACzMx/ZF95nWcqlWaxjwoxo1n5TJK8pWWOAMV7vthb0YL3t2FF8fF/7OD3BeQrYpaVXZs
CqfyO4RgHczP3J4JjrCh0MufAFVR0tbEtEuihAY9SUG1Cptz82KPnaM1pg1834KYRvYlmRlBIIdl
u/VUwufqDIVO2/os7BDkD4X5aWeUE2EjZkX2ceJS6uBB16LZ6C9/Z+iNIlfclgYa0y2XmfvTUtwc
SynQjaTouAnGWu3ff4o6P9QZf4zue1cnwq94r/aM06DD0J/9jc/YqypS2+etCAs1Z7VKoS3UxP/T
3iXbhF8lEzr+1HJq9PrjD+N2KoZwePbz+UyXHYrSi0D7gbWhT93nXBTOJTsUHwGaH9KNvV8XsxQm
IVTLAQpn8vEXC0aN5Dk3cxRTz7hqpkNSl9Xm7wSe5fcl9reDt4P47Qp1Tb7y80iDR8UwjH2Bh48u
YyQSLciixizKIoCKTyFmbckCK3+G70gtAP6WazRy46iGRyv+k1niAp58+hHQw8EJsS+qfG6l8gGO
En8a7ZyiX+gNGcYqW1uACjl3yxxLJ+aJiNM9laqXwexI77MfH4rBeL94ui4R7qD2ViTfzZ+XE6Wf
utRsJrrUbgg/pqAAd3mDxNFZXwn2oaNuhmY9V1kHqDWFbmsi1YgQLASa8tkilFiL2OI1jnvQuiag
sTAD0e3WNjf2erkhOGAbyvxGyB/pQ2eRS0GpH7ILAArAzjoeUHjrt+ggJYHpXf7pbrRfllX9gdSk
QG9tBGYc2H8YAOuk8j2K3h6r8yWP9TWxkPpQZ69ouIah86Ta48SJKAWrmYPN/e6jeGGWJkZ+tLzo
yz7MXPH5QDNRnSN/1Ov5xihbLTGb7g2XCJYN2iaZNoHyKssAHINGd8glsGRYga38zmM3YT5vcSIA
i1P8uYXr4HBcO2ey7eTxXsxmifjnV9HiTCxUJe0ltCs3/BKajcm1I2nD4BR5R6oiCXXziZSnJ0Tz
hVBcl6cGje4/7ws+4UBCWCRsi2LaDphHAW0X/13t3vJ5+flmjwWYnpejEtIAxmdEuy+7SdPS+rvs
vcOmemhsivvkcZelnsKtJhQ9HDiy9Ch4J7HK2gnH3JkuTeTFssMxspH+eofR53FWIOmB/dJ8oMUl
MPmSdW//fmchLCyM3M9jZXQ+kj04bSPTGAil39qHlIuX6qMKZ4CBeX3DAJmJnTAe4F6uZhvZvrOt
QeGvU9koU8N6ia+7ksOFIEie5U5sXyIk4duLHCoWLC83kf0tEfjPmHLuBxsTI82tQIj+IDSvPcfe
IeWVTL6jd+EPvV42Na4nJWV71JQ7djO0qtoxB5CGrproT/ueQOIZ/N8eHu9A9/dUc4pzZBcwaRCJ
WsUsXr818Sd9pMbamL0PI8WlYgS8OGASbe8G1s0GvhkJDH8a3jGQ0syox1V5Fwoz1P1p/n6TEqzY
AsJIgiVFmGfXBWrUIXAYMhFqEfd0JbWk6UG4FQEa5ayrXo+RSbCRuI1mcKuwJXQv7h1KzDKwxxoK
1dcXsqXvJD5dcGceb/dG4LI3jXsQ3pGma4RBkY7RX2KDZHeMLFGS8314o5iHClpr7BOtWxBph9vq
OB0+mQmaeUXVurVMtiSJMyNlCMEsyytcvETc0EdrWwABRTJAvOSDdz8DJrKLBSG8kCicAAcaH69Q
g11ywOs12wmoRLFo+TFw5rHvOAe9kw3NLSAMUgyYDjvi8X4ImrNPOBrGq50Nj+5mbcjdnSfD7KeM
XnOI3z/P6qRyCnK0vdfRYaXrUwTivTsRY0cm6Qi7GbheOWgwD9pVbOMazsDVbL1/yh1MoYO9nr0R
zbg77QCMSqOt3Rd9erFDRwPbYRKDd1z/qB7Cv6OS8MB8Ll7vhGZd9+B2piIyggku9GzhE0JbRBLi
Xr/X7WVRWJM9TMO5rK0ZkGGWGtg+DBBWOygvaJfaXjqe1oWCDvDNQDqk/hOtEMSRtUkIPUA26TpD
BY8XH/jHEAMIVWJ8ipjh9y5XO3ZEdg6Hm7/124Cp7BDCs7AQs1///C5oWlb3IA6wuXoaelH5AszG
ZwjMG+7YDEMOLMSU04oGU2/QjjHnvMHVADfDxgO2/YvuMqY9olOJtR++2q6k/elUH4nGy7HdHi53
mJMmJmiCMVhUSD8Mm/mBVd4vAWT/LU/qDeE0pqW9jE7595mkefr7BHSP9uGyVe0y8tBwnvM55n2o
tngY93v6y/Ije00UxI5LfXA32w39HQ0tc2sqOssfVA3p5i53RjvOWWlS/IXAZdZ6dFgZFxrz+GGN
n4KCSCgpKwZFR1sHQJsVI+VsmR6ed/fal7x5FfQGbLhn/qXuCeAOUtQqwRYQN0aI/y3Yr4dneJo9
FJpYn4ojL7UBfvQommuop4jqXPS2ZvO+rOlqr+K6TcMqCp3hsFWyrqZwJbV42nfRd5jBXobFV+Vr
18HHZN6qn+aSfPSh5KxzDy92969iQJPy7h7eUf14Fvu93+QqzTQbqtZjCrlLvTx29i9uVqB3048C
eooCToF4fa3qhT/Y5z0mthLCp12EOzGnR+1w9D3oRVYdR7GowzJbaMvzlBwaaKjQblNySmQTwKGd
nQ0qDKK3tCO0Nkvi22UEjdIsf/K2d9llyZyFUd/wwG6sT1917wVFaLwGoNS4S/9o0VFX05TDJz5y
luG8i1QuD81+npLmJBdCMrerXFmRlnQCp2G7xcAH9t2PsNfUhvTMYAOaWgDgmWk0Xp8QqyAImyVj
21okn2iSj5iSaqTB6Gip0yKoGsHqgwxubrZKAtUhDchRVVXHMbBsxn4Ot0NNL1rd+L+eygFnmcro
Ym6LCgExrtViTvQxOGo5stCjf0Fu8GvptejAQIDAsUZ+LEUzm2YQZ/Su73weqFBoYCdlNLJ+rMSV
0mHVUrm7Gqq2FXquNGj8iTsOjJBT9xIaCIA1TpvrmpQC9Ds6MBsu21NPIJn4++6f9xyaB2vkl7aF
1y4csU5VvnAqx/2GGepHgKi/kIxmqA4WrTLknbsYcN2GOpPXJQ+sOyz83t8Q611Rq97bW0KCV2Ku
9xRtWaQ+N/diVVMJDk5ec7SSePGyH/iygUjMNPME38qVNdmBFp35gzOab3p3F9qMsqCWWNMxJUx9
51PFHZrsrDQlHKLgi13YQ02MlX0Si+Ko3y6zDnvKPAm1Fe7adNJJM1Ukft2MADSwlgTorOjAPS0d
h3x0oYLS+ViwpbFecW6vjb731QKxcC+qZhPrugSm2Bog76SZISg5paWYaygtR4LM4IosCRfk8Ria
rDsUF67zC8Gx7UrT96VeGQFp+HmJ2YqYA41g9L5emwhiQAcqu129trVipMUjEmztQRtnuEMOEQWU
PhwnEZ73AJPBy3qPbLhdcCxK0ZpaZnq9oN1eJEA6cYN+f1zn88WYVKuG1RGvK6JcShd2WciAtlRj
gq7D9/p938R9GDm7g3aWUqM8sg3k5JLGlOCtPgvR7kDt+A+X5oS6ztQv+Mi0G/lLrw9Qhc9etYLg
bm6fWaJy2Dtzrh0ghNDXPI/Mv628PUHO5mBgx9SSm0YMaSgN/nyA+S1H5NP7LeSKlMaQ5oy1D9c1
lAELLRnYvzHaOEYRzd6wbPGnpNS8F1DweJc+pRS6VpgzqsVk0yC/CCS6VGLypTwZinWIUvSwib7v
UJoO7ha2EBQCBWlkNDzZ6Y3/SHWmDxeUBsurBnH9G+UzhxP9k/r904A00i7CvIqyz+rK5TMlw5Ra
uQyOLMUNwbxo4sN5duxXEzDdJJhOniIHdz1riYDsOzLXR+42E/4wpBdkRxt9DbIbClUEWSPTBGoS
Kea8WgzPsYu2vamMsASLppluVjpQ2ZvOB1zpldERbnk+bv5Tgq3fclK87JFKw/RkJYCqZ2uRZv4N
bVKv2iRb5675GnTchKfznq+2n2G/z3pbGXnxH8j5sNkoWC/b0ftBVjG1l3CXseB1rPTxrJ8ydRi0
gavw0J9UsRT5cP5Y2o64xe84NYrP4y+1b191kuu5yZUmQ7iKU7Gh199vu4d6r2NZ39biLoB/YZB9
Pr1CLmeJ2GedfZ+EcS+MTwWx0Erptn7yXkh+206kfxhJhUrrLVO1KruZf2/xF6/3J1IvwEj/UfAV
VpozldYD1sxAoMCITItF5IADugkxseqSWtPysewOmNPWx6aA1y2nbAZcoe0DUxu9Jhb4CBWY7z6x
/Zk82IBv/v+lIuxNexNXbmVC8fnnp9m4NE2NU5XsclQ9cgXrquLqQ94/uplyjq/08KTs3zbSrwAm
E+OuTLNkuHk7nD0i1mpkvbgx/vxc1j7wcgERmQ1mBCRWi6UkBanJd4wMqdcxFv0ibpWjfp3WVI99
yMUY6/NCUJ8D/ZKLfV66IoQBztOSkakq+vaiKROQZ77FFoe2k2fxbdgEP8kt10/BzxEPXGpxDE78
UYM5AxmhFBfQa/2ElvE8xlJ+VO2MfyUr1wF6/wTKn62pGz2MKF3puXHbGDYWDXgQL4mRlkXQ7OUk
8zfgtpcYvSb8gW46DeTjCuYOZ2xbb24Ev2ykX1k+xg7vF5ZxlY2iL6m90tTTpXuPzDs65XpmmpIh
ATiEeQnJP7a3ndUvzaGhpAzRo9/wNjrCX0zdjGR31cXOV8X5l8Wowsz3d8U3vXiS0/x9020XEd7G
dFVtCdw6//uxQh4DgZPyIn4QTXLfTv75j5cV160Yy2BUiihaztayjI3RO+2F4TwMyu0MpQpGNSOX
RZId/zTKor6rui9YSQvfnKD3oUlKnDmGMPKm1tzQk4KdYvp4/WGREiggy7EJlF3BjIqS7Xl7s6uu
kbIYfaCbi36tj5+OVc8u07aamR2cTZu0LLo1g1t3jsx7fkHCqVICmy68RbXetmXHRUuVBlFOO8jT
UP3FKZbR7q8tVUwaEXuQ+Xc19zIl12QGmLQv0lJ6GyzKW9kZledyNVYrKoaJC2BeNz8q04+06vPD
ctxjAsD4RKv0YGNuktUT81mW8lcwTCPVCNmqig71uyQkorYoEXH+KHucR7zFDxHz8IrJzfonClgM
/mx7ZEGIVEuBYHLGKRRhRT5pooe4KIbcyFXm//eM96w6Y+y1DhTS41Tksp6zVVV4u49duRoax6zX
lj/EBQf7QQHoJezZs8uENs1+ufbDmjCU2l256MCSOsizPjppmQecM6GzDBwQ5YfGc89DgLBAQy1t
j2VrMZIWmFMNbqnC24r0yIs8H286hfDvcx2yIsGxjvcueeH4bKv/F2XmPRMVNhclp/YdYkFj7PNT
xOr340TW4vFiUNMljK/MtaSpWXE/xDO9Q202wSZ/Ug0Yfyovx4uij52aLGc1ALe6EOM8QoOcPKs6
s3Yj65+Gcgt/bYZgk1MwYGgnTn+kS72CPcxKqNnsGyhEPgGUPtlAEY3fHEvy1To0NS9vFhtVh9s7
DoCgDP4CVqJ4ZVL3XYHSfuMHT5CcQEfvcVVDrjaLVQXOjU4Io45FdHq8UA8hUH+KX+VK7f8cOPjc
WCudNsIHMiimCp1lnXRAA/xq0Y/bidLvvgrZgTpaeViJyxEqmhCxgpfKY9M0PcKxgocueX4Pvv75
wqgQ9K812Sb0wk2z+mYDm3MT39EMWf4Al2kvq4nntcNPU/gw35Mo8Z+8gQe0jSgOYJWTb0POX5zQ
bj5x/IW0AdK5/8vwrm8ZPk279QNPRuWpdswJuM51/zF6EQHy7nMOCewPHokIrtk6BF/8Hjm0joGs
xxvL3c8VIvPxuu6bmfYZRdPA7dY3/K7Hn8rm35jdM3PC3e76Ribiqr8Dc3xqofj1GThwL3+pzFyB
eF8/HdcGReVCB1LhqZpVUO7zRseYoYUC6VCi4lvVg09YVA9y3X9GM6eugPlDlJaxxCOwpVpQ+CfI
mWVIFHZVGCpZyxt0CqL4gV/Xbn3NvsbyDvYYsMhTrqM7tZo4bnu5kI07DbwOGLbM4PFLQZzEq1BG
2wPuZdjJGU1wDKm945nwUF6p91q1gK/sj6v/IgoWudH4f+LKkcdnVX0Bt1t7MxlIHOR8TYh72Bt0
5lfjqNKSmeO6Gea3cSx3m0pZcmGBUgS9EbAjRxJQGp+oLmPHEDLu7klxgIRMZQ+F5v4F3DT8/XU4
myduugdabp9qC2UNZCAxkGhLMwQtk00OgVC6TgK0k8E97y1uYW8wyxU4qpEqNHHZGb2H2VEBZXMZ
QT7pM7XdhIaG86E1v4oox4iaukkzsxOe6A2QylzDWwHsHCthCEO5+AAvat7nZoPQv2HSrL6H6dBU
d8N5e6NyLKtaEf7F9DgCZLDDxo/TgfjpgQFUDZNkedn/gAtsm/yAlOoeBeg+1JBi8xgvjnCbJx98
+jQb+PO28/gcApOam+GpthRQU3qcOfLXsGG6t9qiQG3OQhVHInG8Erjli3CG+oWxWBY7eSZJWJVo
D+O7rwnfH+Lm/X5MmFC/CiTaYqobWfN0gyLMJWI10wC1cQLFkzkLNcEwjCGMjUylwlA9CWu+RUHt
+c943Z2ul3KE1eWksh7UvZR/R8UlMO2cT11ULfnwtfcpXu74NoLd4jqKibqeayFxA4Ef02C29VXV
kW0xl/u4CfgyKgspglsdWqpOL2UHtLASu/aVlSU2D2pln329q7+Et8UKv3k/jRciSKXCIwid9h50
rJLzi1zdDNwbuGPeAlvzpq8a2JOQ7IPCqnInqWbJ5mvhSzsQlLCMJJSbJKP/IG7Y95R4RcxoC5YW
twF6+s173AWn8F7UkOFUxEf2d+Mtp1TRyLuo+TFEj7DWPeoHZUT86BRTE0FKaoKaZN4jskbV6YY8
Cqj7cMHanwJXgOuvgJY3llTkQMk5AQAW5j7M9T1lKHLW626w35picIyKqDcEd5KapXalRCSYb4gl
GAyh/a5AMHYJ6JThrx2pl/+Kqp9dg7nnuGV+teXHqVYB3f8AOJSPEIBZ5s/qx/gJEpN3PkWYYAb2
TlBtrcFICuq/0q7XEi+dc+LRkj8g6UnjkZgBjzFU/7YOtObZnvkmJMu8b80YyI8cERpDEyU67/sT
pKWMi6d+LqbpHe2+JkD0c9VEptUXBne+c5IL/R4QLD0L8TVzbS3/AxlBo/2J21YIIx421B00LDDO
ToCWwmm2my13bU/sYPwuoJLVAerVwIM9VT0jRMzYlVjtjCwUH+buqzeEW7kDTZJt4cQF7QTpxcA1
wpDcpel03b+DI3A+nMVSC7qkoMRPmBpmvkrqV7sTcaLr1nfrlfAzRhr+kZT2YVCiEEHibHRVaml6
2FTwHGFpXv8zlJWO3K5tc/qO7OsfOuOOI1j5zKzikWDGt/g2L9oDkC8twhItZagKRlhBwsgunZG4
X1O0O0N+2PepSc5A2Y9S1wbVXgQnbh/UOPd9VeBTuFoJa12B2RB593U1IY/GSRVuE5T74p6JbGto
z08yDvNeCguLg3W47ZBPsM7deUXrKEiqzS0Q4U0bSmeiN/L9eNQgt9o2dAVZgyOXoaElXYuyCbHy
ncpYHgzKe0r931k8PILra6hDl7z+4ccnc3zNNLG3JwSkmbC5baWYF4cCEO1aMCIVAi24tJRGMjbr
d/Nj5uSXNH1M4wGSCaMccIPv5bjBXdVFdOFVTP6Azhj22VkCIzFx16dDr3m0+LH9mbcB3W7U+L3z
opmgSTpE5m/3TjoAUt0Lf7Ofoij8whDHDiKMR8ncOCOmezfiOczQll/6G3doFIdl5cH7Xc47lPx2
BlrbGAbQ4MOSboYPs0epvnNG8bfv3cq+71U36THT5k0ozzDkLTwXhACxKkN8F6D6tBx0FLrEt2mP
mpcVlqcSrENgzAdUIfb+Pm/e8BsO+f7bySBvg7EwbRi/BIqa3CCEg0DoZJLGJsM+Xhw0t3Sjq+XY
JcOdSfnefjGNz2UCx5R/+ZgbMhdKKC2HL1VLqlJ3TsBr2HNd8ZOiCWN2utcMxFejJ0VMk9ZaIT8U
GQbRev4N+wyFl3A+xYSq8bfMAeC/qRpTx7/EzyqIc2013ROgkeJtYlxWVsfDCMrL2RbuATkNjYcK
d+3B38qvb44b9bxUpd8g2dTHQCE06nq9gFCK2778A9jbz055r+sW49LWsC35QdVBG+70NrtBukxx
sd21Vq5YTNnVt9FZ/GS1rytGY8uvoN/by/4UP42ki6HsF4DE/cSeRZAWSyaxgFprCGmQL5ku+bvB
LrVujwoMZq1DCRYHY0HzeeNe68PbrCwUuUJweCmFLRTd0vIJ2qCTEtUINEUjcBz3PxPWWaK6iIUe
WXm5L+KTSrFTlTFBKGmu9kmdgfguKhw9UEIPSLO1C6fzySKig/uw2D4MpEI/56Ye6odCuq+rquo0
qt4Pi3Whp+bxAZObd2qkZM+mtmZHZlZg+3wnts2aj3FxD4uIgSXFYhB6YB9AAe31pLshjSIRcyO1
Nf0eziYGJ5Dxs9BSMDo2IrmlMgOHezHz4vypLFHW3HbVXJVK1V18j1tVoGqanZ+G0QzY5D3dZ58x
NqTrb8HDUVzJohNUytfPFkpjJuC4ulzxxFjsozcHYXkIBGOnh2zLsaQW/72H2DDfppD4C2JN2xn2
qA9B9Wsss0g+Tvfxl/rPi6fxqTTEmcA4MfMfc96t+wzliuAjbmpVnfa0NPJGqAhs272mybIFBtbb
kCJWHTBf+nzXiZb9dTEPlYO3DkV4NoNZQVIZsP0RaYscaTT7AWXI4pQa9c4YxwaGhphnbAxy9MQt
z+1qly7ikW3nDFstnLnwCzt1vxWsPmvk/OKjlH+aNLZXlWvAngNYDFu3BoqGWZyHu266UWI3obl7
vsCcFK9x9Zbb7jdd9+AYsI5S1JE1/KJN9unC+nyAu3qGIrBPYvllTV4YlWu9dnHJcWBlcY1+CP8d
WKzXbcC616cqixJiJ5Ji1JQS7D/sCFK9j7p8G51uF1sXDmAwTH3PuspUyngzHzKlBBnoJT9KZYP2
2JSMtP6HDFR26vYw3zRNY8pIFiPJVqqIHV6WNCQLZTU1M8EeFnCs8IBTv+qr1fQdpv1MmgO9NZVN
qJMIp+32Rp22hxdSRQsKAiVpAjL8ZnT+F6IAdhjBzkGsF/6l/+v+iqbO5JgdnUDSr9eG5KJ3xDPH
0mkISONaLalLrqjsctd6pHcicbljojqh0UCofGjBigSIqhtIxWU9TeA4JH7ymRpjo6NoArOSPhwh
k2Tb231KxNwM2sn9RZS+Yor2gLrIxn5j7oZgmEWOoGTTdpYzknNfH8LIdHony17KcbJwdj5yHDNl
ocaMEzqXw7+nn0Y1li7mpO1gFgFJVd02lQGhf/KTNOf10d3939lKdk+R5tfCQZxwm75IiC4UaWKo
ecLeXNUXezr3IFkPEddXwnRblX5c1bJFzoNb+xOsL79lvl4qR52Qq+Cuk1Buxih0y9EIyoyvKBYc
1cx4nm2oDS/s1IeBl+DEoXrqz7B8BKUpHFlGViez5D21SzsZ5Z4pccO+iSZ89cvUJDPZyjuNNxgA
4JUjkuZo2K7ykPEH0ZJ9HQoEDbvjc+vH+jEK87hvfGckC2H53seALCvt6yMwOr/Q70XFZKH4qlll
fDrRVwJFFDLhjq4vcVRgYhsyhnhKnkxL7oi1lKOpcxZD4wUSfmF/E8dAvew81s++IKYn/n8Cj583
SgLKdXqrHM+DKxvXdrfzH9e+eFNJPjsUdMiZENPhA5R/p7zchAiuDqd4O+z7bzzdtB0hX0f5W7RI
1W2LY8KHp1c/9GhR7BKv+JWy7vkVXjdbWlDxuWO164PBWW7CLLSUeKXXX+ITbx2sduU7FaJb8126
j6dKJJtK7e6WRt1JdTE1CAl/XySILqA4MM++g3BlJihtsIrvlHLFv0z0AiaP0ewdgtNDmkLGwaA/
LrxOfgIwNVdfuMeXyFAvB1VMEEJWJrRcw5zlX9m9dURPeg1SJVLGGQbsC4G2mvFZ5mn0nrCoFAh8
HH3VEqGAqx/tblbg/+IAxC11pxvsArmMnsMrYZJnLE1jRT09YE/AXV8W5eAeMLLpys7dJq4hy7IQ
bz9clSxe4Iemm8F9YvdWmanUaBr8lxikIfLFE0nxQJKTP+LSVOcn8yVIyl9W0I6D7DA8U04dLQGp
8HCe4JoP7wCx/rC4Nj2WiljiBzIVf1BFtk8j+CDFfTfColPige9V1xqk95YOFAdDcJXJ/44XsLZT
DBQLJOXCGpsVQdAWRSSzHm410FW+j/r2xApqkqqa13zQGJLKagr3hUtecCmQfpfHiGha4kr7SSy0
WhFDOGPpS7uxh1wWIGAZxU2f71siiryniCBNrlWL1wL5Q6y16yK1nj4hJKL3mx9sFDXTNHR1jLdE
CWJbfAfdN26QXBba59FwqpbAHVEW2ZIQF3h2ePopkD62yW0YMuZNmAST3vrIcWAgW8voSINwKB69
RXCGHngnkrio6a3VIoNHF7VwYoVNqBVxC3P+lL74aFjCn8NdunIh/inwaK4ySutEqU5xgOQhO3kT
LAYF6BbbO4aBZxsN4jrZtVwy75LdjXsA47Wet87II+P2T57QmuhMwnF87vCLWqNKXgqCTR/4AZuk
ua/jKUUUv8ROSVTsEKTLkgutQkjY+IBtPria3yHQ8mbObL46vOBVRDLQSar2En4LZqmGC/pgog30
9psq+tqiktxFgYbXOb3cvi1ol3hHzXLOUGLq1nDnRP9Po7IUGxqpFQ/TYpzDJMGA0AYpJp9y02pc
Jo80k4arRWDlG2EbiB5+/ODZf/hIkBnM67ocVh3UD9kBA39XThcKw4sMvV2U9VU2yw3EIQd+39fJ
3lRK4/CVa1JCb+nEDw5nrhKoYp75tZdafIB8wXrnf80rkZMblFaOKc+E28l9UqZ21uCR6I9qLCkW
Yg5N5JagRlVWGJcI0b+H/JFs7+t6vpIKPECk1z35+TEiXnxUM9UO+sB1T36F6A60u/tRuOiXJSt0
eaBhElb3SfzWzqMeT+4jN7AMVBJEpGKAUVjfg5738YcO603l5qSpZAcRuv0ElGIcH0am9B9VW8js
WjcyRQWIl5cNndk/5FNq3QhTUPRjn8F4zwfFNBOYfVfq4YFISQLokrASIe8kdtaVyYX3p2ciQgNk
Cgk3e9ODGQXYm7fPa8m26RKpYvj3L90tFs0nInngqMvbzg5hF08VU0NXc1CEmCc9Fn8yue+hH+r5
Vevk/aN/poQxO11W4vqtc/0RZADvXS3XuYMxONqlwVXRDVw+JO7mxNEwBT+Kp1Pw6HiP0O+3fTSP
G2vpQcwEWmCrJflWYg61//N9/2TXJLlqcBfsZZRQzWqJ365DGXmCLlN6/zDa0sim3tWUjTUCrnpd
0TWz0Yity9qdE6Hoffb0Xmt5XLxN/cd8yFBeBhGU4PxRb25Bwn08EnzucMokVq19vUx7GKuUF+Qv
aud29cGUIC3ErpA/L8ccXNL32K/vJvxUEegGsKx5A4zmRHIA8ZSkVLZEWmvIhhpZlk5Alml/cBXJ
xwzusjJxaebIR/a8JHn0p723+Bi0JgvHcck0Y1FSaXP+6SKmbgw0EbGTYSuswKIPZu6jjhGlDNkx
gDtG6P0y0A0XQI53Y3aFPLHnVber2mJTdvw/d/hC+f+7R0EWheG3gElzPvbT641vJO/6UYu/TtiA
JGOr553gFdVhhB3kEKHvmPYcgc/kq0iy8eA6Y0+bvUiavLZEqfrkPztkFtwjpJqGd4fY1se0vztu
5lGVnMY0Y5qbq7wzro9TjBAx05Nu+8UPZKkavWfzZvW2FaTKQJSN9I6JWervej68m9qUwZExSHPP
wYpdAYsXTwNpUPEmaz2Ebg6guYVuctJOTw3tVSfqibc3Dnjabf913d6FCdNksVz1n5XaM23PyxNn
heWwuZLsGfwXObsZ9r9mA/a2uB5dTYI6QQBUXMDzog03HvmvjBhTsVxzcSj0qadBi5792+lpMVuT
Y3wm0AGV39Khu1jn7tsAIVdFiQBI0Noa85NAZrGpQKNFqdZLr2zZG4mms4OiQyIveJ1fEMn3WQqh
mYHHnhAEHftPi0TpClYpHU5Yo4HFaAfPGiFL8DlkqLAC7qXu0RuFitZIoqlQ87urj1qx4+c88Woz
vsnXg5GRszFfffTLPBNqaYwJm7UPr+xeRhlqmAk+L7SbFR1Iq+XUZntyTyVPW4QRhOdj8/KEAvX1
EwkRtzN/LzE+W5Ca4/QT8T3M7/lBfWS6nF6SP/g1ABHv5xJljphJu9W007e4GGJtgnTaq1aynOOn
KSJbAEmv4WDMZX4wjS6X9obCq3ERb22QLCbFlP6rER3IMcBJMFU8008U+Z5WVLUSbPNVN624BdnD
D+C0/sLuHr3eBunV6iQ9OuEVG4DH59/8cTrB3UYpt/V3aoWBuLILhpO7hsbpYWDnRgXkuFm7sm3q
A1AqAMhKFitkqO1okoYOIFLvFj+Iw0XpMzo0xPTcKtkBSLpsbSCdRMjFmSwqOqKbZYB/V8RR1TG+
u1GYGrmfRNRvgrnckVhV/sBhTqj91i+Rt963Tp5IvgI7sx5ZkkYVg7HXADuZH1e8FWZYQNgpjB/p
9NdVykZLZgHcvi7olKZgqba8RVC40Qm9hWUofzkijgGdAVkQ371Of3lcn36ryl6SR3GRl2/D9WPA
wU8fDRkAwTwubJ2u4lD2CoKSl6POfI0YvSQLbHY5MD4QA2lc8MlbdqrmFAbLLmHgCSY22OSlEDd3
/HjwpTJnNFoVaMpdzI+ixZzKnQzVE4LKzMf1pQoECsHuLIHUKWbHGgsLxZxSWnx9PV255dq4doyi
IA5k9hiBEajgPXSaKOqUZ4B6bfxu7iEsBc2JiZT07tiwEqFk7zaTVQLbFfSVa9K6SRFmccFdtY7j
SFzuUH8P2jYVo0e9No9MGKalt9pykpIgZBvkbvWlNgf6mSsQ60Gf+Wk26iBaokNMd0bDufoZIyyP
CC315TmR7ti2v+vM+nSBYdWTFphq8vD54xb4QxvW30see+DeY1GtJ/kQhDh7KazTZQfhU2X5xHS1
44qshTSgpLmuErD/xYPL+P6t6zQaRfnkEl2zr9RKlNAazuAX213OhHKK4YtOwy62zjwLMQ2+OUte
JutuAIs6mhAhwsGGPLrgW4TD8mllg6qm5DsCrjNBzsi/U7CA57dPvGSZGbvA/76gWf2RPhpviNM+
sSJ1FRFqhbzgS2mmh7qSXx01CDBe9usdZnlHQHNfqhTwgYWkXTdoAAFVe3lTTjMxiHPww3NZcrv+
gzo2oRojB3h8cnMD6DVFsFxC5WZDaZmcBu8sXcix4dPRyeh1yYtSrmmD+4sZQzR0QGsXC28Lz6zM
wsIh12r7xf8GMNl00kVtWJMkyVbepREPIdQ7Ch5hwjVcQrq204xU4DXUzX8r0n+LhZpHf/uvimFH
p/cTyZa3bekRVXVS9bu3ux11igSEQk2Xi2hLX2OP0yG8kPgy27Ajwcv0K7AtjRQip/4rlebrr+oh
ORzPNTzh9vEkJXGqty85oW4+/NU6WIue+1ct7loAQq3ESeizFDCmzOcIaYEQibcuL9uLmcrUDWZc
pWi9DGdbtfXjxcEhyYJV0w3KKH5NfpkAZGEcDulEUKKFU2Ib/l2ijzJwhFaju0cZoWBLDr4R6qAh
L9PnQ7g4/YqvHzA3oF1AdaUx/SDVZNs8VVJH/X9Ep+ifHAiiyn5jkjhw23cnx4dWtsJHr/+zRNf6
Zr7fHNnzUsMgbF11JR9BQHsiv5JFuEr5EbPyAyRgV4MtezdJH5jljaiEWq1JsPU7tBfl9wDDaQgZ
+B2JdpybhT/las30HyLK/Yuz0LeL6c6WNPzsjjIwKpS3eceucjiGdkwHjBwblLHgC5ATQ838rNaQ
CcSZT4tVK5KxgotjvMccn7gJVjw3lVNE9gaKYIL22IG0Kfstw9SJtucn4Jv9+vt1nz81Zm0CLCd0
hjmC84K/ofEFOo5FLrugs8Snavl30AQtVCjyzD7CYkUYET0KdfQIf/hTfZvX0NXceVAM5YZDTsPt
jMqJPrEhEKfnTBwcnsTHBXcIcXF7KexwU+mBRG/KNCuDYn1XG5C4hiJxBxTC8yEgdy+Mefyx0pTe
QzoCwp/5sq3af85gD6FfWO8WK6Ti6dYfq7t3vU1aye0qMQwSYAXyXuHKSFo9NAgqWZOL84k0a7GP
wMnc9pQ/x1RilmL1hErUlNeopySMUKsKKMjH/VANnB10zrFsDARBIBatcp+bNzq+9yPtEdcnYfXG
VEFEkcL8GSyTJpMSpKrLD2SgDLS13oC9AZmIFEskjs71bAlerCRSwjQJ/mTguxQR1uF6oVQxXGQg
kz9JCC27CnYVe9zz88mnvT3oq+ECoN0qhJOREOz6J5ul11QitGsR/EeZVFSREOSzwYNkzeEPZhJJ
QSgB3r0LJIn9ziGmZzj9WH2WTByG42b7A524aKcgwRthB43/YSS2/Mznv7uH58RScIYE0ujKec+O
RU4moJc1uGQfDVDKiE/TkSLNOSLASEIn+DQ2LIKFpB35Pvy+YynN6968qMNFdLG2lvhewO5XsA0o
BWoUVg4btqqgLKsS7jxAtWQg/Yn53x+oJmHuDBtZCptQT9yLX/ArfBATtjmY5MgBJcwmbKQjy1Xx
Z5RKpS6Gz+73x0bVB2+MLcgKN3ZemZ167a0MsspgLbfwRn+SmzUO/diWujbwyOFzOGcTF3y1bMBd
uDnXU/+Pihy6x87awqF1TlLHTHlj06Fa4hxLGsApi7bbuikb2eMSvn38Qh5hyQh9Uj2ozM3Bc1zk
eJvZFISHxdO/kdgp6HW0WX6SX4+4iFgj1WHv9b3mcdSgdaxEz4rAWYAhakW73nxA3JLvY91X7FL9
rZQha06BrnCXgX8C42opaDBlAV2zI1d1U65mGpA+TZWVqMZAPbmG2K5bHIX8nKu2REHCqrhv+OyQ
UO6O8xmlngHTAG2FvNcowefnOL+3DyvG1yvxi8cpvs3OEHVp/TcNpTfTuUvNutKB0YoREvSzlZFn
4imb2BSg8YHUd6xudYrDYFDeuKnlFcoj2DGd+GTKhLKFouSjDJK93Fc+zsqelXrY0G7prVePgaEK
Ugmr60fJibeMD35vHUStignEtwrNglf+SZajfE5ciOV8PL+DcMM4JcPol2yNT1+ZNln0Rv/Y+smt
AN/mGKDWym4t64KhW9UUadqHExPUL7RlBk26aZUSpPqOFhEEaJ4ylP02k+3ffXmoWmZSE0SsaALY
mDiVXoV53VQQJSqNkBqUsOEOU8N8oSlas2insDUexN4/G+JzLjm0EY7Ybl78P+nE9bIE2Vvopykv
Fd17uMjBxk3c7KV2w/xMa3a4KAn0za2LgnqrQc8sJhgXNUTaFLnDx1CMqxoww/kOJbSVs/WswxEb
3y7VmuoGfLPr4UAz25AwHP4nFxXd1pGTexm+mysNn7mAohKX+q/cY8KeHxiKY67YUvav6X3N3+C3
qPVtUiucA4Br+zvrKXQp7DP8v+lsGdSBgf0vQ+xr9asMJ/ZjWztiOJPVnvSV6VJAoVP3a+Lq2TKG
AufM0A3PLkOMiiontSfxRgGeJjszBwKPFN3QVcgtyobZXq/jUY8gzLuvqzsq6i1vlZCrS2f71XDY
8svYtThKWDNCvazCUD5bz3C67M40OtclYC21JMcRGygvhJHaYlyMLQHY7qyBjW9DhfFVhv1XHELq
kAokGH+3BrJ8b7cxe0vptkv9w+PTe+N8KoO5C0QFiBiwVgKbFyHfILGe2KJTnP2Ze5y3MekJmaXA
7eFEctnh9zSxQ8He3CmlkA5E7VEfFg3MRdZCbtgt3mOKJ1+0n/plpWW+prhKYxzSKDllkpX1mVVz
l/BU4pRTfWTVQ03Ce00t4E/I/9Dd713HqyWjMoQ1usBfvFOXoYQ/yvV9/vyiHiyC6F2pPIcb7D3X
LElsf+bJn6OgT69fnUM5IdfUm4Yj7xkXImHrULwMLXQ/rC/FBd739AbAGuvaOQVMxbR1l1v5ZXVM
DU0tIPupYskLPuZMdXDkfdPwFNuR5LLvPyn3gwl6o1hlwniJs8RYAvHuaLdyTUxqMeChUiDH7AdJ
s9N16v2iSjR4n9awkjQ5gAnnmJ6x6Nj2gmTHvDZVxZXzBIxSoq1h5PzTMlsnUWPYjl0UY5YLSVj1
Lq3jD/ZocjIhgC322sH3RyUo0grBj92H0h2QSCAcPIIjTXGxg7bx3gAXVizqJo2PPGGyVER0Extk
Is4e9m1HOdjmvrBkRwnBRfB0/abaeExwHk17SJcX+NrY2wY795oiAcMK7oXiAFR1j13VrVe4SJ4I
LLPe2DwlfcQaRwtoo9Yj+BIuWlSyWTEyivMVozw4oUKXjuADHUIkTaQkbsCT9obX6Y+keCBwgJ06
Lt6lEFmtogmNVvJUOHITiM/Pdm7CY2rng38xVAb9cA28jh6O4YXwVS9mIEI1fL644AEs8zoK+tjW
CylSE3NuqtsNQGsKao72D6vVgy5WwEkIluPKhaSCYD3T1IdEcNlGB3XP1o2h/tY3Vw7xAYIwoI6E
E2Vj9AJBmpFoYPSnbtjDtvFeqqcZuHyMkcHv2H8tS3AZPoPO+GbLhu0NtrNcLRtE0jP43i6ZJC32
fVgVwvE8TUe7U7AOhWE0cbxvOOlG65K8jb214UWunH4ZBsgymKuAb7d39IsSiOxC1vgcPN49zaWK
Hvb2acyAm7coOMIzw/sB/j3AdmVoHcCVi1zhO3iSGogBwg0qIheQiQQC5YkaqA5mfl8FuxfRRSUL
QL+9paMjl6SqbvrhhXul2mnIRpCrTmMOIg4ShSXQtqmwhqLgPjDW1UTy1t2LDMPfjpbNbGpUp+YI
moIAOlnlTuheLTPVEXWza/LQj2wTIOzBO6ru/gkmnO8Smo9Fjq7hjfThYcNuncFlScSnc8129KSQ
GDgPEsP3vC1tIkESh+beRRk3Oq9hmYl5locuXvdu69QY2mVF7VdmeyEbIr8Q0AOhrNHdxo84mvOW
SYFvy+mHmpplFlZO842F7gdoPJmM+oQuEBZR1rgo+8aa46WeGT4u4VADVCwEK0cKm3C+H4Uh9vcP
z3qP7/hl3TEdOymeJpmxsYG+bvumPrMLF10CF1TjYAR//Djjl6+2X/58poBBBOEiOvz8Xyt6lV9P
dhAhUkKSlvqvGvRfFjvN6z5EOBQh2fBrF0ZKAOHiLD347X3mTsVlwmo4p6XVf86dKiGfr7457bg3
1QTxK9ZOKF/bMenFeNuKoerFFzrorLbgDuUL3FaJ7IWeUiwM6rg1N6aSAt3rt0WHwHO+ZFX2zYx5
usAgQ1F/LmhP063hjPMbGbmmPizFib7jXb5TuI4gdl+3zLGp+XBgakep4d3j126qPhKVHMl3kmOy
ObQw1bCXiIud0k4EjW9pcqMKQoKXd7y0DSzAuEMxJIEUVjHSWqUipYAjvweWItyd88M3UfsVfonO
YsoakUf9iKt64DJyAjOuXLTjpLIxP8HmzhVNV4zvRCNaLRKr1oNW4LrI1Ai9w+1wrSIw313IEHx6
T2khHw6lG7RalA4jukTJ+B1JsyEs9tONzD92NZ/rC1DwJPKdqBvZXgj3HaDWFRKYWP4xad9jWnTW
FjEqSXr0P0xha5YyIgwzQNETjoyBEILz7YosqoFpfSca1xOyZCqJ8HONgnqJps4hZ/Kf2x/nftuU
IHoh7/IZD2m/CQ5kRBV5EVxj6lZv//3TOUKmu6gap9RPMzz5rvJ5iLSTS4tGhWY6NhMPgQTBYPiW
5NRqei7Hp6le+Z+bvekgQ86+RLj138SjS4R0Ta+mZSnp63Tm9CRPVdT8qFsT43gw/BjEkmS9hQ7J
Bka6D9Ulvf13MINWWQu6fwbRSvFFgVJ2RlB+8CcrMOGV996t0g6RSl5hQt/Rlm18QAzLZ/cI9Z/D
gwWdESP7WGC8vcYWYF9VWEPLUKkzoimU1iGusVx2DStr4pKUKxLOK/tTxm4hUl8S3yegimhiqIeM
VJiHcKj001z7KH+2JzPfeMY6wMYfGdkURtNGqSqHwd5BV2V+VS1YXRkU2+L4jGChOATe3Cmk69IC
IZAYTytDpXhNJf/tsNsfPLbn4Vvl/OAmm204AHoLPFJ9Q36rZfjCXmj/I8zQR1vVdImqPZsQTLMu
O72SijoIY2AZpUl9zoAEuv3ASwT5bxq1A3EHjUQa96qSeclLiXyUBoT+RdW/eopk+eViIHOi0aJo
8zYMdKEHCOGFxQg8oJO/X3AdEIWyOkWw/Alftq8F3TdqjAl35iIn1CQIRKyX6p9joLSKRtegKNjD
bGoju9TVmKbhlr9E35xzmfvdzDgMw88OTvJCGW+T6Xun33UyPjVpuBbzjHFlYR2hGoeEWsz1R1Yp
y56/s6BZKggrkDmZdoyxROMRuxCyJQN+sIC00mK5+8pVao526606Y3fQppf44g5Sy7BsuauS7TNW
QxMPF6Vr2YleaTktrcKgDxnKvWgDGecJTrOgQRP/we7g/M9rawJ/YLGOxEcEAh8udKlAAkCVRbcU
TUV5Sx6li3aAIP9a625hUUO+vW+i2WzHE+pVa8RekA7WR98/sF3fG184TvCoK8eOZZuVyCTSJaZ+
cUzN69g7oSwNkBZJa/fQOHkl7nIBvHmQ4EWzM57qMNMMK//a/FJcCrX76MqdoDJpBe3Us2F0Ezj7
zfOGt1r8YZP/ITXJwszJC3nZ32CoKk6yzXqzOudD7XBqgLVpjbuzhaziqoIicos71b2XWdmPQLgk
pSULIDuciNXpmUrUIBokXRmwwx+ZaoU1/JWiLX9mhZmSBrW7oVhLAwZx9pRGHlOhtt0B9pd6QaIf
vqD2k2Vf/kE9dxdb/7nf+y+Ia5NAegpJw//XxoOnkDjvyWDOHT9NiSU0NAfYlgfVKZk4pJpIkdFz
EhcpLHbKfxb9tWLmv1fO0UZcT2UurYbsLi4mQj5IkvbW0GlFbp3Aiu14QQccVhg02aojpA+HDK46
MUUPHtqm+9l8J6C0hrBL2rL+2o7vVPZnCLP0HS6Mg6DADH3q40GBX3h5yDbsng+YYcv7pEkdWz+8
fwnn+qHtV6sLQpHGkOXP3CQRjtiC4u02Bz80SA5UxM7kgcPghhEXxhkcq4LfOKUntKRNHwmm4NQF
c3yYBKk32b0e/EFF2/oxGdniURtLI1s9K+QZitjHho9EgElRZOu/MIo2h+3T2DjqWEvj4yRX8723
c84+v5+iHGoHeNS+RMgKWbtBmrF3S23UjRAFbfRtp7roqVs4xBXQVscMmBzY0fOijPWKlMaTXldN
MFDzFlHDUsPhq4mKOECuZn7AAS45RGQ8HHcgNl8tQk+0iiaVXhdCEqW+hHuXt2IjaZ8VKJN2FPBx
4hY8mN3XQ1n6a6WPFaPxcAZkRP1iwkguYSEIO2CsJN5XuazycWlfta69Nb4AV7DPUzCrF6A4CTmu
ftSgq0EARa+X0ieYecZtKohPqC704fRfCNnG1T+DfG3EzwcFUTCobdZxcPFSzjPc1d55BXy2AEn0
ES5swVO45M4slGWXRsHCkUQodxAzRCATjw5zLGdDf/x4lWEfTWVtYWKz4iHVAeKpbKk1piGmHAz5
GXruI7RBXCnOv/LTtkK/JiRnd+2DYcEqriX57vSELsxZ1QhTUOjzycbr7b/HL8oxPy0UCiW6bdyK
GxSDKNZFpDeBuSxTexw4NrNUI7sZAgoeyFz6lxYsXDhSSCnP0B5hKW3KqSDUNFT4n7IR+rrXr/hu
1J5gs/ioXLYtPb/BFYWFQnOFiVNqd9PNc8vcQp7SSj98DRtQ/rQsCvc3kbOcw8kNhjSGt9/4nrER
37lcANkl/Ku/ysJF44PKiBGuqJOLLhDQhMfa2BtCRLKWcasqaD7ZsSZs75+IVbmLqBN4rcz5ukBz
WzlWBSi9PoCTg/gue602mMBifWv6oBt502X+/Vi9rhDh5ZdPF/5Hpauy+Rkr9/xTaNkxtf/BOgtl
BgMA9woil2rv/Ymg3FXJ1/bfxHY022faFSyRTuLTlSqFYAXRgSfeDtH/7T9bx1Om/PnUynv51MdY
jqn5jYqPSiABhbXbZ2lT6Ybl/5+4A3qjdOyHykhzewk8em1YJZOOEp+kXhGimytmTq+cE0oD4bjP
SI2lEnjTtijx5qAvUNcmHD/Q7aBKJlm7TRweW5wDfA3c8UYPVW6AZgEUzbz6HMk0UUl0e1VLlYY0
3JN87b7GXeD/ulTpAyR7hQuC/7W0GBOaY9uftpV50uhxcy66eDyDCck6jj+e2qj4HW7FbGAAyLdv
sxyMuOX2Atrwb7VdvbsNGyxXKPga/urTmN9BMJxq777WBlRGDKdAlm3Q+OH0BeA6HqsLJ+lhzmck
8v7wtrsXwKrZuc1pBIOGm1AUtQiqSqNF1EbkWGkMYW7dv6EiHI85CnxYswkAovAD6Nh+NqyWdZXU
3aGjc8MBwU2XoL92SUWsxQAcOcPEeTC6v9npiNH9/59NfNowlsCc5p/ZXuShXGPfRVroQVzKujih
E4Pxrkw7vC+3H+a7mWyC5pZz0ktp5alZ+rHq+LdvGMyMBMs1ciOlOT2VcRaBNiaGW7Gqet/8Ugew
oTLqPtbXtSUoEJnt0sHQE1TDud2m4VUA1ooJb/DD1/HDxwddozbzlnKTwkAD5P7qpnBZdh66JR/K
fpyFF3nvSoD0+6YegAG8jMRZ9TMlrr6bWuLZLajfaCxCyjo+5JulZenFzUqSiYVFI3LDXkhyBvGt
sg/3qiS3xWvHAIUWrERVlTsaet1cVUSx1qjbXlLmgGi2HYvESbeP24/Q2bHM7/3bv1zXeVIxijgj
g6vRyGiTvy6RSzU+OyeIQzIfGh30AmTs8wIIDRdE40LcQaKhSPXcfjsF7cjd44WdIuqBF/Ii/Xcp
QB/b8YULc4qVGTgUtL4yK8hetiJCVD5oPXgm1FG2ROC26jlKz9MbeK/8QAoA0J5WCujvPLj0S6Fs
fsQTTp2bXmrgBpiOwVfKZBh/856VSdfpe7IdLoKgw9o2vHBKfUU4jJK3ougM8MHn+33WwI7j9QAy
gnl3Ejx9KRD9zPr44PNnnMv48bAtWC2Cbgo6XHgPsAQI75/sJvpZ9gterjkmoXIdv5Lm8fgu8yi6
ASqMLF5TrDo6q1fYLJDWyRvzHrHvAc8AdIE+ZBVBlnASvFLdgm0btbVmK3hEglCqu4lMoekK3YAh
OSbXtcINRsVi/8e9xtbrJaZo84T2DMr0ovM1DbxomOU6dY5LAbkkiLlllgTFwWoFBraVxxe2k1Gb
FJoL3omOp3oTHfQWKRle3pYLUGkN53G+3Fch5wshr46fQ2QIjaTIJ3WP8ebAaImYmsYkI5XY9CPF
jtnFWDcL9nGd83xobRxmectiIAAAKKvdKF++l14GYeBgGImr/Eo8lDvlRgjru7BXBh+YBDQ6TKwJ
jr85TbNkOX8N0kTKnHglJtNJl8fUAEhsCtF8lqgK2QPSDeUL/0XVuI19N0GLs4vFVw4gh9FH+lr5
tcAlmmA7MeOTrhohd/UFpcEcYVEc+2XibkNaUQXY8CibCkIAiID3ngqm4SV1hy3D6HO94slimEaZ
TZAErdR05NaK/MBUHaS9wtUWAks12R1NC6g4GaW8fT2DSdjBwCmO1VX8V0p5YNfrv7T086A+3xp/
uXtFGvFdl6AV6gB+T6Iqk26huzYmuWBHeD11I2TOtE4pgBxQpOLcevhSnHtXp9L97NHnnOutoFPi
ILpdByJt1vYlNn1bBXy9KeZ+RRLiVTWX+0eNmF4qqVa0x94LorXXUJJkcL6LCf9U+NrUwCEsi2vf
uvwEUkCclyEOh8vNXd6Z3otneEjcahyMA6SCSeV4lYXxN8dIggR5D42PKMP0EBEEpG662y8yT0IJ
uLuk5I7E1uIjh3zh2lqycEML45QwJxMyj7rViVtl7TXI0SFl7Vi8uaXm7cQx8AFiIB+vNiYdpSG1
4We4K6S9B1GdItWx2jfKBLNT1ypaagfEGu7kk/Au3ZYrpMYmoKrbmLxyQ1xuRe2MP9eejjt2Q9rj
F5UZWqejHzzAI40SnAFoKJZxLafLHHYSHZwJIbbf9HGNfftTHQAlxOhXixqOCyUVPD/fb6OVFFOu
wy+nuLiCRj89iISOZuI3Ws8JrGj/+l2e3AleTHeyppIwqUkyxZ4HSBZYzVXFqwaBTtABVAPRLoBb
q18pysXlNaK/5DjHRNj07ukt5mXzrUXBrODIOLP2Q2tLyumwuBUqPNIoLhyqaasHT/L4Jtjs3npt
D3CTEhN3y1bVwKid9gFO+jmmp6irsbnOolor8Ff7ba2LJNgQtE4G+rZmh8vOlgRXU3CcRE1qS4PB
hg77pMTR5SkWdKzQMKggPd2nleUgn9Mtr2Kmzdx8ie3Sd8B3pegL9WO4k8waHAr9/taLr4K0YlhJ
TGImE77wcb9dhRC/RU3Ckf64HgcUDibvo6OjIubZFoysF2+tjXnN/EMj4EgMpfj+fdhyNetwtpg2
gpIalEUM+BxjkO9mKdMCZ2SaasHQi/Bigc3Gn6Rb3CI2Opqmix/ZK/kzjuc6pC7It8dNvV1mBCpB
7FALed8uztPjpvNCRppY207LJdtF51uc3abhcZZIx3OrsQ9KBt3ILfjNxjEyie1KZ67qqt9nHDCU
p8HeLFGRnX+XrmcPXsbS3JwzkByHzR2b3xL0KbIeff7qG6BOEC77b+9fXWw6glF0KSpAjGKExChg
du6miHEwbjdpj+enszAQ/TbSzxlS0AwoMe9dV53EkNMmm4H5qM/uyWT+ionjbw6B14eXlQXaaCRb
Or7nLpcdeY5lFRm2i5C1F/STrWSfGXYihFdV6HFkCniv1k873mW2NSStg7WITnLlMSIjR6Yjoi6h
J7Zl2RcsgLdc7H716/BgnNtwzmXRY7oSqT7Fb+koU1aBSWSqawffipY50kQSRkVxh+HlusFtrlXZ
XQpwQN+uXTqh34vvWROcAk4znM1s6fve/3OIeR82SbXMKjKe1gb3d604cgJRAV1IypdKuZn5J2fY
ourycRd3dQfmA+cn8rThNxxmmvC2NQZ1xePVOPJ02GSO2+tyQJjopQF5GJa/Nykxdu2hNXGSwQ0a
izHiBsFua9R5E1hgCVYwPT0BnmrI8kgs9bcpDFW1qpZcu7xiF1HZ8q2JQCq7FU1AfrZi5ReODVp6
A69so6rkRcg+nNWFfCG6/OqpqOsiewo52f3DWghz78/S5rJxPsrOMnW4IzOJPaSIt5KjaC0kDRue
fUR5SO2B1qWVPYg1uqMPJkAYz85QBLePuqNmpTPhuka4tOeJBfobZl/Xtb77aMBGFH2ZDKQrxSBC
/GMJd0eoUGILutApx/UFfNFAgnwK+JI/D15SnRYsAdQ7OYe9JnxOceWB01bszojzwrfwS6d70bh7
OG9I3ghxN9NlGnvuhiDmNYHn3QbWoR7Bh43xujjPQZPlXLoQeGX3IYmsxmQTNPKpqaVTT3/UCNBN
QTtf11dah9VXQsuy1ksIbbtM9WWhY+t2FqwA4WY+cZCbL10n0UxHDSIcjGCwyeZR5AmxZUSL15Be
sB+AmwwDv2CUbJJiU4Hmp1JYbG5jWEspEioNicvCCG9vv6zfMjEUPAYJY47Br6xSeffDeZIQaEqR
6bCEprvp/eHitmRwJuZ68mZUNr1amuGaR0q4DuYXNg/teUqN9DQqFh4ZQCunXlDcODqN1/JDaeSr
W4W+xodRZiqcJGRwUtIShYCYrs9aiyM/vwb4TfQ2+LXKRLUd9LK5dIb1h+Jwfh/9OhhU98B5ow1i
yrFYlocx5JzVK8eL81zFxRDhAkXYEz3NiSg5mJb7siUVSA93dXN3mJP22R1Q4ofgUy2uk1o91ubU
Z1+MOSyfH8VuePNIkWVIPveu8jHHJAsePIxRiN7Fu8iO7m7tEDCEKh16hJGV29ekuQD3ZXu7maMe
5GFp4r6Tm40NVuDPSRS8tVFhCHEyHp80y/ACGWkXhI2RC6sHE+1NzqUDwE6/hbXwHpf7NuzxnnZ9
FFcOG64mm7mTGx96qo+RQNNmnZPqrAyzyynI9qUIzdHWiMeb1uDXt3Qbf1ug+jp/AHUbIXeB209K
2BCKhOxS687dCBsE/aj3ZUPrytHkV6+T2nGaQxK/0tZBxB2OH4ua7s3hP8dQjuGFCo4Z8sDIwB0V
7ONuIsXBtQz+9nR82y7SMQpISr9tpSdVJMpG4laFGnsW5iEFEtflTQK3Q2hhSWz8RmStJn4QyKY5
pGM4HU4scFKJouHSwxDkzH32Pu8acHnzUCuu7VY7bxn61wckUsuvVAWosbU8UiMzPQ6rKbsg7RfC
ul71AaKkSKMYoZfwL6pwrWzqUlg3evQhdCemBKkoCbUJenYGxiMCE0Pk+q6HGdyrU4y4ClaQ2LYv
CpPSFg0/WHmz39y+oGFZ4lRk82v095G8HIhIpab9Wh7AXMFJBSR2jUo1+hCbq4dFwcrl46wiuTlL
CQOQBY3W6z3h9WRSDf+38lKzLsHxwrsRc0wms/ueR0NTF92cuOUZxmbRSt0rkTazCEc8/Z4yPkT0
g236zTPVSKY00nseBSydzIwjmVe06iE0BSsQgyq9lpc2WGMVrBHhpSMhzQn4PKxegwCbmrM9Zb1S
wI0roQNQoT4vMLkawtR7JqL+L+Cf6A/iJY6QUV6onx2zogsNfjjiwE+RIZsGsStYKgGQgW07H6kw
cGJSc2r35sNdg63zxHP5gHmgMZykoXnQBKTTncG4v7cTE9sBBRKhHjx8/NhZThgEZ+B2n88TZbZH
ynt/VSu7KmAUAfjyG6ZriIDr4lFb55pE3jwD6ugWX9M1UZJhqO5fU1ZO/WgRTummViT13kW/Tegc
4CRlbpWyV1sGPsWnP4vPt3lVZ6uhwXT6zK1brQgZWDthGCOB4OH6a5bSTRa7K182VUr1a/Yqh3R/
P03yMH6BJPuyUPFhtYX95XsamHKtyZZSPfC3+2WnR0RnWtgF3EKz+/nwuYeSdLyLlIjvuWp0IQlr
cig6JtX7g1QVGNVMe/EBeg1ZxSkrKS4j0Z/RBoXo8Eb40JRBTvGCiGqJKOcMoobxIQLcuNoA7UFF
kCdO9hoeAQQlolAQEZFr+k4DADjOBZLlQ1X1Df9U5lytlWssAI41N2CPXeHrnCyIQhXE5ulaf8KO
NaRVK/RgZpY1HmTI8VwaoV2j+dt9UxUCzsJR2X0akBetFYJTmQ8Ghda1SpardaLY/a8CbIiYkzEC
uGsD5mdP6gvPI6VdTCZdXb4uC8e0oAKW9B38ULCUPN0c0bf8c6apIKPtilP6vWoSPCTfHEsSsyNp
jCQawK5p/HpP9O9alSMbUdex9DDi8ojtuZo3VdB0Nh6jP4jgN7c+6xfdHMficY7wKBbUvuu0cFO1
SvClGjK5BkcjkvbL0okTpk0bMfiwWeM3JG/SvZzdXhFAAp6GisR1s8ddaa9LVNTory111D3a8fHF
2FCqGFqgZxnutndKY9gelxzxjZIDBusiaaIn/yUfyedVmMrIq9CjOXTq9jehFqVwgQDPotMoM65z
NfigjnFJytZBhzkr5FrsFv1AnVpt9FG2M8jqv8LiL+wgOgVj26ESeA9z7+iov4ElJt9tgQNgiy/Y
bx3lUmH1L4UN86ezaoIWzhIjq2VOWKUCuJqT1UvFnwy6yErEKERWMU1EVBG3u5uN2IIsfWZjO1bF
JHcODL8fxX1dUeoD/M1j5jpzpddY76PSsHCEvfsFOiJt07/bBJOQioS6i7y/ty5EpBzkoWA3vnGe
U5w6uJ/4JH6lWvtrQ9j6CTy8sPYdIuFtI2TweuAS3g7ZABAkLHY2Qlew90C3KDkaX+svmShfGtt/
eUb+eZ13+8gOtOsw0yDXwNj1+mXPnbZKZI4Z9RJF7LAMME+Ul0ZzSFBpr5pNz+LxeI5LsUmMtxwz
jeHfkOWujO/yLHEL9EyWf02t5uKn8/tCoemB/YBlFlhCmYqeGEfAnhw+FS5nnaE5cP3/Lvpj0D5Z
SxCX50GNSzOArvsIbdETB2Caw8SIgU1nH6UPnudCdf6rh9Sr3Mz+sCE/dgUP7e2/yvY02uFGyLoL
Lyf/FazxbdEAjGUT7XIOvk3p5qRiQUHt4m1JiP0jt0JOaEsI/npycAB+DEfcg1tg8/m3Yk/s26CP
nFE4dZinJKOXMjpjpisQcmOJQDMltebR59AnH80AXXzwxd6pcOyho63xG42tp9+gwlc5SfimW7hi
6gt5wWzw5LWQ/DBMZGg9XYdlrO9Dx4h05RwrnDNNImLa5lSsupFzkiznVU5uNdbB5L/BZYAf79K1
C3rKSTDPvq/X51CPa1xCnLdyG6PgTmVpgqZ43Lsqh6ima4JuglOTLZ4gwEOiOotG7PpGTcFL+/DT
vsYPMD++idX99bTMAXeo7KHpZP/OUjQTCMy9N9+/4MmhBDsJ3DSauMEjdeV66E2TBgyJxA46ENwS
A6+qhxSR94CG+xhUc99kDsPs3zYEveVjev/6sahpZGRvcc9bV9CCPOoLeX2yW38AwBOX1z2YggE6
Vyae0vmNxA/hh93/7PpbnGpNFMIP2xxFzgMy3ocz/JYpj6tLAbuMR7vib6n+1u8Lr/imySOFEy8j
tkqIrh+TYo6857/+CKEIZxDS9PKdtlvUymXTbOR8aTuBik6zxoKTwNOcDFYvwYonMDOVXkw4Tc5m
pwISaOrAYRwLinimIgvlBGLAl/CsOtYlsFiAfwgqrpdZE4bN5DuHlvxPlgS4HPxQSo+y08Grtg8r
Jmu/Wfd6+PfkzqUVYeMWWzK0wyDM4CzXzllkFcCzIoeeUmTSDmPFzuvFRjqtU9VbHu60V1qXHJ/0
ddcWJYYucMNNz4aQM79HEOR1CzB/f93iaHZgjkKJLqD+a+KID6T5i1ux7HRi/BIpHyG+PkEr3Kph
DXwwsdntfUIBcX4UIoE+DnMCpAV+TrfwjtiG46bFPH05AacEZl5sBSVCUo27o+mWpmYF+KYm8Pli
OL/ZVZGQ7/tgG6o7iq/9D27MRb4nk8oHLXp1l/C1leA8j4sh3XhE1fZqO29/3Cf5ODNihC4+SO3T
S4+V0HGu54NRwcuHDJTHSYc70ZMDh8HtOWUpfbH35WJUR2mWKI8pRhyx87L8dGzLMGhs/75PIF/4
nubFEhqJ/hm7Q4FvNDbBTFTOJlxC7Q/jneeKcJ4iiwpWhxcyc4VZSFghyW2pIhK19LxbxDnhgVMv
wwImPz5DR7hTF8/59Hez36te91PegmVbZ3bXgi5bmOyxd81Qm5ZPlIdb7BZW0A89auJ8J5Es/K9T
LzOCLZdjJpaVVtEhLVuiSj6rbeS32EUC/0Am4AQafjfHfgW05JmCML0cAWqng6+4jYmb2OsqLcxO
M5owOnl2O5zqbH6QRsMtL4a9Y6zTsyVuCx2oRA9Pwq8KBt0u7dO4IUOfXnQ6ZYf0zoV08yTsyM9O
68UH9r1tojYw9Agvxl4hVrNaOiExDAqexykeAs+Wj2T4RelDoNT9tlwmvZLHoWY0RWf8oKg9hF69
ZcCQVMcITZK/52pF6g3Fr7zEMzSBEyeEq2OcZr5OGHDO7R3U8z8OpK4t42YhK0TSEYjssZzAkmWU
231ifoKXjkNJJK8fjyOpqRQjaO28Rhl+vWz5jhqxSFiUL6yzcf5pDNMLFZobbXYhfWarMZhW6rQW
nffGxDs4sJeZZGL+iGCdTtJzJ5VWY6KtgAjvZFCmv4XYGl3+qo4ZmiUnwzIc9hYa5drxpKtwlj7P
0sC8v0u9FbiiQ5KKORHAL2jZn5fL/KkgFqCOTiIdFhVS4UVV9hycJG7WOolFETxNjdB9GsN2R3Kx
5BGgMshRGJxF1pUdHHoaHu3T10hyC3qbn8wP+1IW9dkKQpBRrDxyxdhxbvFlnv8VJMykEIHuGKAt
mSoe//z3vo1Wqo1F77Hc57ByY4NVxEaZcyyz8Z/wWaN517KlPOqC+dIIdWgFYcP0lGAk4YnIGusa
M1f9qRHe54sO60LIaqCygQpUNI3lGyuU7kTUO3AH6AZoesp/zkPd4npoawn5nUZBOzswdExy8iwO
DsuCdlCTao8xUG9FotnUghLxJ12sLu+xBqI/INCCyssjRIT9jUVOs7T2r05cruiwuKfGjwq4iskt
9NHYR8c9e4GJWVkU8feN6ILxucqmguRRlUjIexlgdH1NXIvex8rCLaa638W73H8EoOfZfi2jagw5
OozpR52gPxS9wz7dYV9UtqAUNy1tM6A2LcaLIjpLQg2zmeqTC2EroOg0Wv+7PyXfG0DkyWW/vZQL
XahiAqYnK/p4EPdroo39Mxo3eARt6mZrv88+i9RK2BC2J7/URBuSrmq0cCffaDHRoV5pNoUv/yEy
I8pFSIQ+JL7O8m2pklVoKm/ije1W0f99DYvPFo8xPhkucWWkqkP/Yo8FjChsbMSUJK3kpC01Tiqf
lQDSH3+s8+KWHjgiHhpTbxpRQBrIXJgDM8Pk4hMZXg2VWXfgrOlXaJ+zuhJHusr2wFrsZiM95/0H
yj1GTIWRSBjvtsOIlB0I8sLuPUk5La0pAcVhe9965Ls2DH8ZnFsVVI9rPybEx7xHDQnUO6EN8T1A
iTOy+XhtERscF3QoVjGv7vskf9sYBlzYlVwO5SPYwQAHVaXW3967q0/TiPlaW08+L5TyExzgXxyL
Xq8FrrGVPQ9j9vjjvMzu6NDuKxqw1Z4fJ63E0NqntCsP+z2bUypko4tqCXbzPR1fx0+1mwQs068H
oHeGV7pX0bAFRbmG64wNV0j63ZxnJ6WaC2T2Y6Dwv5f7xg6u/8R3Uwt8PIQtRBPuXILKgYezn8Wg
jilzngzKp1nEfUtH+qWLGorhbSerawDdC3p5D/er4hJYZlu7M9H2VPaFDHTTU2eluhIbJ65b/cBa
XShRnG73aXrt2jSvZE3ikqI1j/AE7bB6lD3Oceg1GXbd/mulQ+sJNyEicMkmbY1OWT+wKqZr+IEt
8PMckCMYTP1AO7RZdJgbjhzfiNNJuIodv82jl5h2CRFFH6LYA/K9U0RXPr/3hTUGH4Fbyd6mxOzM
dPLIdvyF81Pe5BIYO6AshWszpuLPRJow/1C/BpDU8mIkMp6ssvPzjENpJTEqYvQhk3t6wMzzr5Lt
4WSq33YiIJWRw+RauHTSZ10+BmT/uInJH2ez5Dh62uAdl4zi7Fh4ZzGd5U9AhnsjiPfSwvR6DUR2
j2YV0MU6cWNG1yBqYS1Ow4axoKbCLmJPFLSQi2+5i9giMtPe8yQrQRlB/ROByFlMUWQLtxSgbLw+
FD2mw+SWhwJSXK82g+m4sWc9t8MFBMh8ySMOolscmQvkxlrz+9P/b7DJKziV8Up1cLODrFkfi9T/
HC85HvZxxqBn8aqySBD0ZktivTcWbAJN61V2kxHhTS45Fq5fN1LxN1KNrxdJRTbTQLu5bN5YuV2r
Qa4PgguuK2YLpjq56VQ9F9HHZbohQLPe5NQiI4ldc1cc1IckCj7H3iRTFWxp1bzTZdwQwKzkAGVN
SN65ddxKHw/VSDJF/uuXEpLkkuS2zQuj1D/Kk1b9MxRvWLJtIVVTQ0qrfcTtRHdAWixVH0LPhJRP
Sb5jx0FohPQsYejMHWSfv1UbdWE46G8Sn/5WzKgenJQ4AB7XV9ksXqkhiHtYt3nAo2OQuj0SlcyL
zWznPYDV2csKCKg/Pfe0bKXPvlNkPexNo/RgraLkxf3qa6sIRb/4BPJ9Op2LIe8rbK5ssGch7CtY
XuiA4Faw4KgPJogAVisH7ZdcOP2B88DgP9uy6l7VsAQy9QCqf3PNsjYhWhtG3SQ4T3hc4TZI5/FS
YIG8d48sPVmLwBwPH4ChFm/q/Nun5bWxqO1D3LImrFtPIMCgBfftkCoKH8g6u4qQDKcA1+Wl1nVV
VsMxCakoUX+TR5als3XC3UqP7Gd7FfOm7f8z7TKwKx15ufFop+vMmCD0brX+DgtXlrubahGs6PmD
4jZTdkx/c89wGu2oukRbEISbfMjxZhBkMelH42s58EmvmCbxcnlcod86Csz9QOzU20ewDhCZJKR2
WoOJWgHfgoya4logCjCWVPKiD7MDZ25JeGA0bpvSTPXhDh+jwUZUHeLEnnivEDXn1qHLNUtl3Pyn
AmHmGMW1nH8ZWHaUfzyTf53MnmyvOAGuQ9NaUem2uTv2xiUfo5CWlfxdNDk78V1p+QeSMt+sgb3p
t1wO2w7O511d/kU/7ooMy59Vl7byam3REBIyxuDR6ZG3ksAoRhTnaIv3ZciuNMlaaLWDp32XlUoe
aTsO4ozcphglNdkIMF4PyxyjjdzJG4hGbVElmkTjrxnk19nIZPP9d1jPmm4B4l7NNOY8WlOrgNMf
OhyhGMQHJ2jtuTVIRxOTfpzi1dBJVciuvx8Cin7p5lhmdzMZQo0F5N76Fr9qCv2M3p+mi5EohLu5
mdj+m+rhOJpGscBvJjNvykR4qJkv2k3sxnejInrI51ajyUK8Z34bITjo0CB0eVnjzXin4GanFNiL
ganB64g9TAhP+gLC5ywFtaj/VrZ9g8bJ+n96mpRAfFoHpAcuKE/QOS2PF/T1XKOGgwXTp9nBWQhR
swlk1S3ZfGdOxloXXsnKzkfV2X23Wz/W6u4HKXQCRzm5t+yvLps0ynGra0STXK5kF6BSGpLSc9H3
xXZxUX98qcAf1rb1a/ouNxyRFKYp/sU+l/9b2EYEyGznJ8ZsQkfiIl6eXHcFz5KcXxmN9cinXb53
sqz1WSkPzlzLmYr+hY4VeVP/Nuaqjr2NrO5VQnquRSw8mIDedExp7eslzAjCCjlERfqrfyQv0RNs
6fuKvRVotn6pc9HFei5XUqq5WehrYL1FuOpXf94IyuuTwMYYriqxV/zcLrI6XCXQlE2iizSvSTpR
juc292bFstKuAMAR6cPi9SkQwbMI7A2buctRFYc47siIXajTsstZCs66m4UQxQ1H3R/4r27gUo3K
8UGFV51A3c/dLKhsrxcb0gYoyoRIOAMZh6OopU+7J03Sy2qsC1qHswzlbMwJ/4jlATQzswDDDsa5
9vNN5hB3snor/DRSixbQwM7eNsNRepKAIdNZ1D0Dcj1Plxb6yKnj0kGFKLg7I0CF87X/RUF1gRou
T1LzuzgSwRjYPgZpq+s8QXEDH2H5vkf+Ecs0+jdUixcX6AtQpJPYfjC50ZScfkeaMDYXkHt/etuO
OciAPU2ui4eolfzUubc10HnlX82nDgp6kre3pVMWT2RYEhh10mGF2fGff97uvSqaiwqXDAkUaFpz
4GGEGklfYwekmEZkH6gyvFilYRd0B1RETz9l71xs0UToxLhwJVB6N5xhkegXrsVoZxlZxtjGAt8c
bXV182zSgzG4LHiuoLZ1mKouA053OwIrNLHjp+t5vTr+8Tytdm4d2o+WU7qqYEUsIh04EX9Cziyu
mqwSt8xkYs6R4X2FrMkUExuP9B/r63j2qGGNdZfbdYEeYTzrn0876nVP4ARl1yCx8Xr00MJQZkmy
jWL1v0oVLRG5HwYDJhcjZVa+z9FTATxpYB3mWBj3TrTogZosK+dxS0SSBZpuUKNi68HX8KZLjQRW
JySMnCtWoGFBixRNTLrKsGJ0ioZOUxqxH7KioGpVxH/09U8DwWJEWfRJTYHJg3G0qN/3xgbXQl7V
n4sbT4ECuJXvbF4K4RT8a/z1NkXbk0t7T86wiLvswUU3UjII3FY7o4x1jUhFuIaj6Zjo5eWZdLFm
/ooyuLS/Kcm8b9Fz7H04/pgEf3ShYUF5oM52C5kkpQyxPaiu61kLUOpVNz8H5Rtw+lcWHMzYeVLb
gLISqyt7ZFKnMSjme45XspX8RZNeVfhL9fAPHswQOprSYcycuqUFPzwVAnWZzdXrF1H6KD3gpjwo
EzHXvcNrpl5mUkNZpX+fMxNJUTBOw/tTbHkIhzG687EByMKH5OpdckxSbjWvU7eYiWbI8U2kQjFC
KiVQIU5uI5EaC4IeffQn3N9vw2qPShWFwTLsSFysUhAOThhd6WJE+FvfcwqEFG3qevdr5XTxiVpC
+KiMXIcGPcbMjXG6JpWszg69oApuDJCMxYtwonSCQb1m4qPNh/0+bj2jZs4urQm8dGluaRmtIeqs
YgfgnvQDW5YbGwtBhcJAvv4Yn5DQMo+ob+Rv/eYkK1N8zLX6LV4c7TJFty1V0v78Ig/ZU6LmKeMr
oRmpwVT7RIsGCzq/+q9nReiIe5Wj5QVa00ZMPkbXuMNtyb64RI8ULigF5wSpNju8ALIaeQmZV6as
i2XCidyK9VIjdTbnIU+2bs7pk5EUYy4IpKlM8Yq95SgX2BcbuyTUN+QwOZ+OTzzrUpA4LOo7+WfL
G13GenICtUi1VsRB8Zt02Js7PxXEx6ImIr12sIwg1rvIXULIoNRPn+Na/OzmvSJ73RYpR2a+LoHk
AF+D5aPvofWAOnERIZ307bHLZMF8niprqh/6sdNx0EwaQWjYlxNw89orx8Rcpss9sTYhJzZvvbKi
upeNkPbTaHs0FDoeMyg6xW4TYlNakaXlIR8KL7h4qp5t9pFxbeLg55LdLEmNHl4kz80zee7e7boh
I7iJIoCBvaXIXVNuJvygYXmlvVUPIMW2C5LjFDUfYVgjR2uI+oZx8qCQ6USuPsB+iWs+6K6an8TB
dr9u+gGUYW5EWWoH4XKEvbCII2N8nUUSALIUgL/Q/3kIQnaM3yn/HRfcL92xbhaJVqnIyBF5erkN
KWeG2BPcRd8aRlkaT+2zC2U+ZpfrM8Dil5rFxmBQHDcZWz9N0cgIJT3E0DsJJQHew/E2lDP5s7R6
WlEhFtcpVe9jpgYfRPCLa6+DTq/0UMeW8gAQ/BvsrfELm4xdL83gNhmfQTcZURmC0mqm5DSa5fOc
/AW1ZS1BROQ52ocALtGVh4/aO5LP76J14wDECIcOxsXVrGH02zn2ALVCsb7nLZc/qhDg7cBs1Eev
fUAhyHQZQ7O87rvsOCQJb3BCzXN7YN6kV+EBZKq/u88laKx0B30FRex2PhSvLiWSC46yxK3jowqD
nzG+Kw6leSKDy5H/yBhvZAUaotRPXPKL2YxUBx3TtWBinsZoAXIqaxK/nt327mSKo5XU9cXfRIKU
x0GqirIfYvhjMkOW8G/JMUt9WsXcmagy2NWXK3FzuKnvLFDiNNMWdRUkrGPZtkkC7CeuvxfB02ib
H/pFTfmPXWTyb5kJqACtwR6pnPmN6m8RouDovIvyQZOzMP06qI+yrvtvCQeX+3IUzje6AB3I3lmr
cZngS5O77nvZK5iMzfgzMBCLYkD9THy5DojGzQjZ1Tb6iTZuvnCAI3mvGuwzwMYHBIDeZG9mxlTF
mN5E6IkabxytEtqFOqvL4o/Fag7CKTImcW8Mxh1Kl3YFagwbqMZIcoCYp+xaX8BS+qIYfkJk6lqM
HJSOyTbsLHvQsK1hcG4bF/5csBvbA8KbyWNH0xxYnlvkWdiK8i8BrzRTxFS0Wzkry4mOQlJNkLhL
5umqjTtZwtR03aROBbXNQ0HW/jkk6kYKtuo2TGSNMVJayyyOVQkXZaFnnnPcV9Z2K4UKtAdxhUoX
gwu/R0OUGNgj5LbsmLaNkrDyWYMdGjNdhTMPsRqqyrdJ35LY6zNg+wWKGGET7rWMxFKUPIbDu4k0
JD2karUzsjs0iUXzt93xeUlvb5d3WA/jPAtQOvyFc7U4tFH3qKrgfTnIm3pqDcwarPOfBSN93GOf
1oduSzeAtW36VgP3bnfKqmME8kyW0npluQK7silpELzhAe94EDY324Em8tGAYNnsbX4b32NGQ+A5
g1aSU2E50m2BcXyPoDdja6t7Nk94tkPRz8fGgMZxfhRm4S1eOgOPUNGPRxoWqVlHqLIypQkwAfu7
kztcihD6nHEgeigXw6XIfC6xtb437fElIJuETxXcBsAipurUY2sNl0XAPCXgqsiEPbKhkffCrLCl
CeiqZ1zn/Yk3HcYCmF5k9Qh9KheLp37qZ88xXsrM2GZ9fLqzF5XTh0q/QGpl4WFlv1cgXouxtHhD
Gx+grXH1GfE0EjNxe3b7D0Emg6aEN7UnVRdOsaN0PFJ/PlxtOnMspcWZbJrR74iqKwkfgAOMGYFk
lL8nmi481KS610cn/SfWyIm/73N2a1jHZNfOWrs58CRuwPpWok4Bx70FT41IWG2GjSoDlvCxPqo9
lCkV70D7bALNaXeo/5FY15zxXjwo0RcBso0/b4zOwjIzOAt4he17eygwA/9uw7kLpjS/0vlc/ekm
jzFh5TE+ip6bJPEDVLKBObNt3+APp1IglKivP0CKYOv/pPLSmrZxj9BaDgfFxPjo7yyRWi4XW6Vi
uBDw6WpivBXZImqMBo5MHrTnbqjh2au92lWRFaWb2FEkjdRaRCAJ+e8EVAbpncpO35dQ3VXTFpdH
rOaHW+a4Z28nRaso9bit9sIB0hdKxAHWbZDsB9ycSKveGe2tS25MRKMsnXDNuDe7WnCcOjqQy5mF
DISk+NvfLRo5RGmr5lENFjQLeajHtGIXPTyXR0GJvsTIjjPDvqpV26kA8Rj8cP1KtK2C0gTdrDCR
cozkvC3PR9V2sqQ3B+n4hV68W4aqJNglF1iOkKDHKjqFaKNu5HdCBqvC1p+UUEI/80LxHyM2gh1W
7spg+o5gV3X4v0Vg+EHGLRdmCYkbbWsENC+Uh6qzGZ4CAkMSJp2RtdZBbbYXhnc5uNjUsWMoOvkx
LEszQVtP6BUuZyKt4vjteeY32Ae6NHqC+HZRfmxz8MfnIiHGapR+AyLTEfRL74GnNYmhwzsBPJtU
j7i7BqTLau0il6pKekVwd3eSWtdCzdrPrgUrquvIoY5XsAh1QKKv2YTV2SxpPbfMKk5BjdECGEqG
0zCLeSp6J1hcFLPoHsevuFB6dSwOWbX5+rj9R25MuAluv5PTndQLsnjwtWgijcOC8boODUc+PKXI
1xJsQvHVuCS38IqYw5sJ9SUhUM23L+Y+asS2X5ZSbotGljx87dRGxQ3udP4tgZ8Z8bPdlRB6LPdu
8X92sPLZJlmdc1d2sZtUTBBcI1FvmlCZwZdfFSkQwEsXpvOYf7yZK2jCcDgIexIS/p+Z2G6XqkR5
aAWBVYHTvGPz82DjFDNG8tJpo90s20zorl4zWa7XP7lRd9zBWTVSP9Gy/6ln3HaqzXLYC61M7OXn
Bes/AoLuqgCFYHQSguksW+TxtmiGNx/rIhNYes1UiqbXJtwpmG4PqNdWv6CXN9375kuJ/RGHG3sB
uOJ5JTmehrJCBGAzq27XTfU+HLOQNdaOc14W5sGD4Ok1ra9fwolC0v0N9lgCz3uFOM5X3h0aSpI+
6ny5d5qcg5T0aCWQidIv3k0eS3wfmjD8DZhrE2HPt3yiUzSIdgQLJ0QdkJCR0J0G+j98u01luBdu
FKvcHaGUQSZtdk1VPtT4sf3af7Z/8pKZq5cVh7BtLSEI+gxbdJYGS5H7Jl7tSl7gy6CPEcx1nVYQ
sDXZqDZyBI+HjNjhNTpzAzP+q2ZdWZdy4GWqzV0fuc8N896AazfqkgfyLwKGTvK3OUk9L35uVgpy
qzGrEDTGxLJUhNV2nzphMWmRGHzffrvYz5Pkl0j7kaGobpFFsX0KkjQ6F7rwntL96uCc1rU9uZOe
PgaKtKO6Pf8kNcJK/OCfPV2XwN2a/SN36L9WL+z0iOm+ADkyUDO+9aClfV1g/7muFADlsoU2+m05
wNkveR4GLuAYtjBqWrrIOcU2kMAuD6Q+OJ5U/Hdd3rGQ3Xbyrvu27tLMrmP58yUGP4xLOhDaxU8P
x+8JkMML00GjqTApkduNgsMM+2Etb4TheMPVnhuv7/NWq1xu9mU6R6Tx07HzHF43V8yx6x0UKuST
qJvQ5Vr5PuqcelJqV+c9xNtLk4YW3QOvrT14CljtTb9AJM7PQVYhcqFlLMtYqXrz1A90BaIWp3Fn
bT81bYuumyAf99J7ukZpXXriAjpgZmyW5Ol/CKgAFj13b3TDK7ntwznGlrMWRSc9QiLc1kzzZFY3
eOD1M1xvFSbD2uRC0qM3o215SVtS5ir95LbD4AGrYNoGv3gt4qIK22Ypn0D/zFIJvAVICSE//xBd
qrZC1KC6P3Eag+drCc5Ka9ML6vvwknAjHKtyDNwqEDLoGmEAOq0ozxjbxlcyXDeOTsHVq4hjJDXs
AWaR6wm2uz5Spl44/MV2mOiI8J9WMoX+HkSLEHZ8++4+vN9A8XUpjgM8dMZAs/j8oBjTFC1aa53T
Yp2Ez6QJftBsNNckUif+wo1Cthw/hEp+4ZSM2oExX8OH9x2JedhYz5jXPsUHXa2bGm4qycWnEAM/
cfe9vy/wAxmbEKTCFF/xFeK5ra5XSKmt2N6ti/h2gHl9Dk8Hxmu33iKfJNcwntgNeuDnS3N9cZKp
dVhjofH4wGnuTV6GXQZkqg7F1RCJGatX3uOOcSBb9lnRuX70iCs0dj0N5ydUqZHbPcK++k+0Iv7T
kMs93OxUXgKo770LCbsXSRvub19e1MslfuEMndO30bFz9yOjL7bRiS0rJbgX5sa9FViKAsxBlmxe
XycI0H6Xm/OqwmmrhehV9rEaiIMj5EhiCMffNIzsX2ZC8EArUh/yNIzQPdutinpnHy8eyoKeKMvF
G5aLXzzpcIOVs4BtnuLU/G4feMZoj5KbgN5aE+8BAUC32xyTo2K9//2DbnjpwMp5LH9I9fHG+z56
487x7oZESfRZAHREgdMeqbHxhcYJ4UPNKib/ro6NXAZgTSHPnLZG9We/jbDjobITiTdNcej4EU7m
yFZkhabpcCpehe7NEdd3IFfsCcSY/zEz8j1WBN2cwWy6csHrCV85mqCDxQwLyBlYN0Gln9/oSWba
dG7sX4vGQ8sY0qO5xLzydiq4AGpcpkahhcU+2pK6ICZyMiYDUSnL7wHTnlGi2B7CYJPa8CcHfaCh
JUbPJ1Mf8w/YhXgSAd9FSzTe0Mv+ShxvmkpDzwQszYLccjdaen0AeP/06iQhY9hnc2Kl7ECVWFbp
JcAxKegC5XkdrMYEhs6Ie1FhUeoGCUFDZDPn07cR3MYqfFnOla//L+JtVTPhV3enPvUSImg67dzq
iZ93qo3L7ejRioIu/FbBEY/IqPpjmUwyPtc92ry19/iqr8D1rgohbBeHlZqKyS1i0UBFeChtH8sO
d/qYfvLSf9MZkdsupoSYuajDs3Bs73WgIlBVSZ2V8xS27Yo6CdIV42xbaBZnpdHvqHprq4BzIl6e
bCCmGbulnFpZtXni7hulfqqOucpiNWk0H07KjcQB5oyjtPHe4WOVQQrF4KLHrd+hKiMsVOAhj04h
G06dcwvxVbkYyBXdgEZSJ7z1dBo9OD4hQVCEoDuXjSGNVWJXrFYGP8n6LKU5pbXKYbodV1HksApz
CHsZTPQt2u3ZyfDnydpyPYTtEOs+JFyhBq5tEEnjct4UttYavGd1jUBnKCaycWbBZ0uvZXxcTx1i
Yi2uAQvg61alT9StzQ2+UkJIkFW7qbC8NkC8nU6YOZU8fxRvaz1fXOSLRPTMA/uCwKeGTS2aCgxO
Uwl3M+Vc7zQbBxqcI2AqlR154oqGfKvxcvlRBQoHjTswG/LxXze59bYkSu4CJKEIDHjLLLOs2nAK
3HTP7M0a+Rh1ficu4Rwrz0cit5loBtsb0IlOEaewBEk0TjW2at5tzExY/VzC0EUEZjf2W091Uiyw
574yzFNFKOVp9z9q/zdbTFZceX42MGBUuAsQn2BVwj9zxd6LNRRnB0AmJfRCyGrIdRzxq978fRlA
uDEKhiPzgoybaZ5/rDe3FRB3g9WeSno81M67shGUjAo53xV2flgShSlUrcoAFiwqQBOcNATiKSPB
IG04RnoUZiX5tpsyD+7kmjE0eAWZrBICxT/Rj857iw6x0r2KcTN7Rmk80Cdd/qEB8a18N2KBVz/b
JM2Bg0qB7J3bPo1kywShVbYsZS956FmdMALTySbl4nvoa9msMTl2cmPcKw+Cn+zhtOnKN9SxNdIT
2vVYN1fEngm8YLXb11PLZjgepsveCX2TiHeWDY/dw7Fpg4cd/bMdpMe4SzihL1aRBlWQ+O/hCgq0
p/x2m6Hw5+0e516u+q3cjhQ5J8OD2CM7ZHxkR1Ind+D6ZOg+X1KDfMQQDkLPOimLhmfVWdI/H6+h
I33usdBn9/U2XAl1PyGtev05vLjheLcuLKfS2UUhX0+YsZ/HNMdQ6U0vvF9c1wdJut1njeqZt4Ra
U84nhgmvEwS6HHaqp3wMV3CadlEmIQKjEeMA1viX1ig+9CMQsrFa5gODk9m52YFawuRN9HSZNI7o
ewhzarfDaR02QIYN1B7z88Z6CThGO/SJY8Iy0hMzrcVVYgSWesIVh5m27cGc1AGJbTgqO+gvEeTC
sQU5Y80DUQ45dw7G1UeINgZLz3q6nWO+OsDX1ytjIttbNX8oFkzb/2ifLg0nVv5skqvJkTErMrNR
reIZDvvDig4i+DIJL7xASqw2awLGPHBGAxb4qEXwKOplPlZxrd7kHfLBBbNI3ivYYGmMesrrz3jd
7tyzCm09bokmMlYmqvwEbONNxXZbPUh/GtuOJxmz0e+v4jxeRdU91EvAEHEXFhWcU5Gi5VXuaGZ3
706F/b59+6/hJ5lGcFPjgzAoF2MWH3V1VCHInk17f7j6ACINIirtn1r9NqMMIeqGX8GIDFXL3fWT
kFov5eQy+3g8+DXJKSfJ6fdLNgkZPBnGi7RFh32GoniTq2t+XgCtw+sPJKUgZBdWF5ISLeq7hjwj
wWHuCplxsaOngXeVTRxSyOScu5K6QyPNoWEoYm4yGk6XhKEch1VlQMBEptXVDMRs8NRdd9w0/lep
lgIIUeENrKwKnTMcnqoeYPcCrxtdGTsLJ5MobWwEuVrJ2mL8DNLehjeTPAswgQTjj/KJxgHinWX9
yih8NW2pLtO3qBdRLSgfBJGCu65kXCQQyymKo14gA3xIe5K6LWWFFwLYP0xj1MHhwWK0kQUpMoP5
xxlU/3lIE8eW0jUL3KQk6SiAkSDz8FR5jN6q9LDF3EDThFsKbLBm3IvS3KwegfD+JlLiz6WKvSQK
8cRs8eCRFeCDE1k4pF5jJ890+cK/EQ8kAajsIdJ0ra7WcZ/pfTtARdUU7vtycgmi45sWtlNXjJlz
BhF9xv+SuF0nKG5BUodQvWk20FAkFHNls9WL/cO9lmSBRq/tynjOpf3rKnQPmwW2r8XTKqgQtpO7
szk3TzQj1DGf1p1xOhawMXAQREOoQg+KgNxfH7+Qxfnhi/qQNQ3eTbUhBfH+CBllbGtX6QVsJ/qH
V+o8Ap0PWMq12bvbeblLBQpe3Nr+QWRbGIWGPfNMde8Qlr/DiFDZFStnArw6/5Yd+/pbGyN/pAdx
QaeJXcPxP3KL3cHYS0hJuFBFYa6vIISXtSSCwj3SZfE6++Dk0aqbJ1t7v7XLq7XbEy0G06lBTcWf
F2krlGnBqicvxSbi9tGMXApL8vloazvDOdMuA6ZPVTci1b3ligCvizV0l0tcferKzgA2dG47M4Oc
no6LnIkeAeFphcnQZ2GQ+e8mCA8B5NiWob3lxG2BpkRGoPzj2uivxW5Ewsr+2XW52oWdgrsEh087
UKwDZv+fCM0CHFjWDzH7XGnaq+tqAyJtjX2cW34FVPDYIbvln/77EAG5y7Qy1jCfy+WTI28RghSs
rvTKMkJchem7POqtqX7xDav4hlBXFflOQ6VIYHHMc50dBtF4y042FZft6PifLfzzAT42zVL6kR2M
0fquUwFzoD2bHdlKieB7se8bcECbdtLGsM+LBf1E2nqydXodl16dheFdnH1MXwcfbnkvqNjWAFTT
v54qKSePdpRy9ZPYhtS2hha05mMDeAGRiFWNCqUFXKSgsIZn7rTftvdnILk9MuFJKu/i9wLPRciR
K9FfRsL0w0YMXaVKAL1ACzpRW0JWXQYfkqn5ve8TjUngEW6R7nwlmPKVcyXSVdUb7JJFSV7gyt3d
L7/zdAR1i2Jt0/4EZEHQCdZjPQ2aaQoyo6TkuJ3sWCWzCOKgTVkehW3Ze01ZzZ1vAPvCu7OwdwmY
hvYvfJn85zNu+PwGmjkfdebKQfWcex4+MDdpQRGap3tow1lx2FJXBLZsv+zkDce9NzrwMNF1aTnQ
wnFM70ZZuxFeTypDJ8Awr7TX2bcAZ3YquIQmGYE2nQBDeSFo5LC0U68R3r59uitUgfRJ7A4BtuaA
HjXVA/nCNM/uY1N5S6NUiRc4/NkAfZny78g0hMjr+9zr+O2p65lxXrXaQgxd87MoByYZrLj3U8Eq
2l9txLpheFCCy/Ejwmul6YFXD68gupq9DjX7r2plJjEX+jC6bgiNbpL3fjal0hXiEmr9ntLe93uy
LxssW/0D2/NudtCWNvzLTCqf7D67c59EMNNf2uMubDr+c+HkdJXadR7URFCRrn+cOadbzV1xvkDY
ekp10y76Xo7mQ2wSC/0LsbkNAsG1h9Ak5wtE2l3otVGV5c+72Qk3ktE5PdY0KoVjWXN8agzchVvz
z7PwkZd6HB9en9M8qJ11758j3/yRJk/nVm6DL40LUF8EtVUeqH7WMJStAoohUUctIsZroMwxXLGA
wRSPk9vt1KdRc/XhVE6Qmr0VHUVp5SM5fBeVoAQvVvi4QqIgYrjD8GV64weBZhLKcwZ7zsyBZNRb
/ADA2HkBhxjqxIBhg2YQi7s89Dcb301PgWaF5OeT+vOncYqlaukXNJwm7uDZLECo+xrfh49IgfFX
7LRo3392k0czWCkY1J53iF/LXzvSaH7+SsFUIVymA5LDgYc4vFOptOsOWzC3n8fVFOB+sXDiIt/X
h2KZZ71oWu3JGahuld62B/ikRE2D1MyebE+529d1GH3bhobI7f+0mzIPMHlrZgfBplcMQxBDpCsB
L1gtp/71NJxpC5cajTgDiJ8dlusvvpAlXnm5FcmpwuFABtHEQjX99K48XdpwFZRhQK4TcLWkiLV9
Cw+d7Q8B7osT9KYeUZu9PDYz/oY5nOzaMqdh56DR1ysqVttvqbFRgy4UdrBXj9ARIhZUlAzHCjwn
81uT2m0GRVlPJecXs5+KSCvXgLipQouBqjCfzGBLhzVOMz9j9CizF5fUuaCsksB/XzLsXVTeS6HI
iVNBPC0UE/bZsa0s3sb5aBizSCXbrKOp0CwBpWTPG4eekHS2NxX0l59lM//dTLE89ZTYaQtYqvGb
gpTTkH6tjYzIGwLbcdcRHbUOLCMouWa1SCRXYZs5dzKoVBsPNARfoLKLg4/IVan+BIIvfqMpLwfu
mk3Iku5fOF8IjYT+6GsL24qUHnilNQV9GRw+Qt2rB86Pn8fVZDNgukw9hYfZVU5LygNFvUiJ/c+b
6NZeY3TCqE8XD27Aja4jFL3BFdSXRF6kQHaqWDz6D34YUMA1DwFIUuJm1kNtfB66iXJP3Hd4yhwR
S7Y775hAuBDGgjev/2m1jHvkiMD4AbltCyCc0fFV5iVFIPBYoMcTCuXbpKr5enRdIRfR6Ob2LFrw
HUIGTm4nStxVzsCpBRrkiQkcyCGSyiWtuQW39UazwJrkLPXza2de9CwAHYLCOk0qZUyLgxSE90Zb
yc4EdXnuTe1hmj7AhACN3WkodVZlMHj0nwjoylha3EOj0HdgGgN3e4/Sxh+73g9biv/DDy0Dglu0
dN7LIRmy+EHfDjfyajYYKbcCy07pWIsa8gqLtTT+DWJFbUFIVIE8JlJ2f5JEPZ40I+153myS4qoi
294WOWSGrZHSxNtetd/XUlLvSr1S583WLijfJ0JS1US/oyGAE+VcleIqaYgLo1NThjSpIaLf/UyW
XC8SWRgx3PYvL0e+GZXYTNINIErwTz0CNaTtqSJZUpW4MN7i3z2hC+MbiTU0EggdWWVmCnHaeZUe
ynkEqEVpdGNDoWzESxXCNBgfjtTXSOyZ402Ix5NpqsPNrtIKjV5Cnd51nSTAhjGdpOz4TyAB2/vf
9tQoLPQBKciqxNG4SxshCp+VO6GsBPIjKoh/daP9THtUUzAerW4obVIJmM+HL/zTFoI63e/wDK7v
jyB8hwQdH6x//uRkNSia90AipEGrV+01NCzW7FkB91dCDBvl78CHSPBrKJR4AWhaMcQgULSMvrud
NvrcPbxm29Ncu1TQ3N8Ssbq58MkCKWJHjY6guMoCQi9NPKMnIWnD/1LWKM5HlAJmFl2ZdxfY2/LG
HKAlBlbDkLk4Kzvevo+5x4Azq9grZywMJsqMeBGffmhxzVTfY4Dt65Auj3eT9A8z3wEnaMgvgyyE
n9m0MXzTmGFrwZDaZy4bWb/8IZ3MSSAkQfNCJHzM0b1Zu/EIdkK9AeAsOp6chHJtERKmMeNisRx/
L6pMY2MWfRafSOLSsi8muIafHBc6eytYjm+6DwV+S89E4lPZPYonNED0kPoCtQdj+LMa19hg71bp
E8oHnqz2hURuaWw/H0U3/eHL9/wOYRVWxTe/4LrsmMm5w2RElTwGc+Fe20Ho+K9mOm+3Ld7x7V3I
mJrvQJ+wxXzPb/uEUjMgG6SD9mDilYGcAw0W1a/EzznI951pK0Smns6G4fzQfAWAnZRob6zT/MZ8
4I62YwDDWBkLEGytqz2viwTA3OYEMsyuU1/NB/ui/dmXdgzBTFq4F0U8E4RkKL37QEtYAz7UJqRF
94YqdIKROhsoJXNYx6pkodB3i5ic7F6O3hhxkdneo6WZdLI+cCoMshQjWCt0rH+P20Fc5VsMMdIh
iT8wxWxPm9rp8Qxn/sXhfCOGegifqSlpVaSH+RqFGcqt2z+kmjrg9is7PSnH2OMSqcfJR5DUpVQ0
+vnXLmYW4NzXoebo81ecGwYlwIjy5OQ7igwSUagGm2uIvvWUan4bmFZqGHilj3TarOher6r0hD/L
Vk3/lY6e6w4cER7S6wN4OZxvKVyawFHjpjQYpXw7u6FxvXQoZBRU0NqpplQG6KofrX5HBM0lGpyT
6NeAtJKtSJi3qdWA7WRgr4OZ6ReYsYwqdo9qVAJ97mQYiTH9/ZR8l8m43aIQ2QC0xAszwActZc2T
gfxMWBtR1cNIP0iQTwmq/mjQlV9kkB8fZwsBPeCid8b4zZW7ULKAqXl+GhR3rDFf//zH2OoBLSZU
ODPbpZlCA6TpKIMjZzjL31feDGgNllNzFKYANy0Bh0H4WQsatgA0mDiL0kqn3EZqn2lKDmh6jVqP
FmoMFXSAlrqoX4//ABS88RoMqlgsNaS4yQthJG0nH4Y4cR12/1lqhMnhqpxQ5N59WPl22DEm4LAV
LObRliL0YdOVdb7lQW1ED8mm8OxIn2Ur1XXttEOFcnscGE+9dxZvJgVcWB3BWlCaK/BdevidE8VB
MXkMs1mCcsnMsxhEWBi8qVb5iRLxNB+K3gjExD/iwhop369oxIYWWP60zVlmycy469NLuX45Jr96
g0JdIh29u/eHnedXbvKp9d2mNQhBfehrEgg+CvbGWrUJJ2KiOC708CXy7ze2xH7K8HoTIMuLsT8T
gCtGkpTRkYQOGNNYdSNf/UKtd6ouPE+rcih0QAz9s8eET2/rY+95L466sD9bdDNO6voMIz4lfoI2
9lZ8fTq4mov0/zSsktRcCCYF/HtCj850+pzITVfO2MlwSSahI0h/989mgA+7T1MSa3/miXFpRcQ2
G8/tOOOZ/eCdSn8Lg/P1DHijDsustKcRs1ToGQ0TlJ1kY7ym7sHKKEwvG8mHmU8XikQdqOjFNr8n
kxlhh1Fe7yysbNMmahizsmFwkcEV7/D5Ez6WiXEOHceOLgwA5ASf0i7SaCM4nGW0Wj22yq8Vcdw3
QofNmwE1JfD4/hVN89aAybFEcUlX23oX0XI+xM0y6GhsBtxi8L0HElI96voDnctXqPtCjTBcsWjy
f9sDXTzpir47BL56mlPAM9QyHUUTWjRlImrX/7aqNSODuJH2GKIzfjVPYVO4VNk+9LPEfjCuKBcC
/XsWDwnwQUFE9KAiSSfO/QSQf+DAWr2pZ6XyZoPIfdgCezBA5+yINjou/WlXSlnfC8I6v0uKAGqV
KsXBH7uSO6KJjeirjqNoJtDZe88VKkpAbBgOBgvPRej2hJDcsLBSYQ8h23YGQ/8WeZKamAx+vkGL
WZzPT1CSvjC7M/xUqjgjVEioQOeeDqSjaBNF9Jwe+T6NifsiCce8HvQ1ErsAUJbUTTnnBG39DVDg
/hPOIVEyT8oqG+dvIJBQmFO7Oe8s60c9kVLgF4rMhwbfwVwr+90yDAYx7d3UmwDjk2aHKsfIYm8z
HTZGZaGXj9xrDAtz/7nLqDv9eU5AmNU+es1/SBB1YjT7pbGrRCyTyc0GXg9ednwyRYK1nVWHTWGn
5NScubp5SFyytgkv9sKO8PleobOrkzBDbSTZ2EW2WTCr9nsZpZlL5cxmzjlZuFhuevHrCBpNSw99
CLVevMNfstonabF3jx3VZlU0dWiOFCf61mNA/vH3wTsK3Jgynqur6LxdOPxNe0jhcgHzXOgjQeUK
1/BWjbSYITnjfuMhMOtOfiS2t+Tke+5xBoPUOmEs2tiZ8t/P2AIsngEstarccI2qVSP9sftw4cQD
irZXMor7Fa7qgoD+Gh2SaFB5EpIaWITu/opkJAB0cxUDlxlKokJDWj7DbTTbg6eyIbISTjDTP3Va
/D8P9pL92DrK+fpA27JDoZbQjMdJgP8AgTIvCx+CD3CdItOlP8nXSE3s39YeBep6JaGK4x8oZXsC
ONF8l84JIC1Ea/uySk0U7xClmka5mSD4ahffPfUlbEhlM887GV3P8+1thS+mW+N20fBa1bcn2nZ2
X0PLDjc7O8zgwDqA7m/Umljnln9ohu0BM5edXYr3LfcgpybS4zccvfLT2BFaPqq3nOyjbNVisZoD
2FH8cLoc/d//y3uEhH1jP1IRAEtLws/Fep5cr4JJ0XZsKy85INCgu7Rf1hTPigyayG3IyVwn0iAV
pOM2WF4dRB8HIFQohWl3oOHG3pngZ04n1rEchNByS+Sq+dn1uiMXD5yT2Vh/jocq4IzbjzDEspIi
bKMoTHaxIijtC1RQbsRp5ro5hcBe8sLq8tJqTTUR4a+tufKRQMZLpJJv65BeTKGImxGi+rBiEl+8
67X69Q6Sad3Rp8W/+X/Ti+afkmfnzU2cNJeyQwyynBpBW9PUiKgdmZOuhO3ME7hWH4Gyj0/PkSGs
hUvqA4YyqjX2s1LPli3qnz7Vfsxn0PZq5xZL3YxSTpfdzxGzq8eVbCqHZqZWTo0S0lsEXASEM4ej
OSYqDBnnr3oPiykn8REYHoiILESDp2GnT9RGzDvJ9RirnPfm7BFl0Pjre+JhZLI1NdeQzMedpIlQ
icR1IKjn6icmW9nmFiog/zLrg/kaJ4ub0SCQl7uTQqonR2oRg6sWejDbGESBxmOuDAmq0GeasiTe
hEmMxVcnfL1bXBwJjqaIlvOAQehaMXn8QAY6KxUiNJcwfJDo4TZ5nEKOxQ77Ef4aSQuDnZ95uTbi
J4wqvmnvWYLrPuyP9tnZzKZQHUFQkDjY0I1tEFBvxSXa5M5CiMAmjuL9ZA9KqJJbXl1HqlJKNCvI
ubyJgOqIdqZVX66JO43JuwA+u1Vr6YsgzNV+SuCMWTH3lUJ8b02AOUYV1mnWOjlrHjYocZo7Mgo5
Vh2AExmTPSdz2Z0pFhUt7MWvbPCYAneRyrckna5jhdfeS4cAc6gE7bOjxMy2DWAnoKh7d1RZzNlL
wJC8o7m3uY3ZjIdgomK6BSnj+JwT6zQPDcHHsy8JT7BJ5CeuLSjO4gqboUgkJtHqu69s4pWw8La2
dUoHnqdCRXFv7yudc6q+IqZLve79V2GNxDUofWcoGqxkSzOnOvid7C8TMtmJOnnD5fuetoJdCY58
weUQEOPjpFNZKu0UPS1lInNttdG2gYmCN/IBYbDvILE/d0LAHJ4AgkWpa0PQw3/EdfmjJ7GxdbWA
d6EnaVCdZ/us9xNa6XPiqKrZcoKKhebj4dReW71tdKckuiocnW1iLRhnirmVwb5yZxD1D8i0Uu38
SSBUxl2J7oNu64gA6czd+rZOHxY6E477QYq3u5+wNbl3vyS7xqdDACvcsmO44L56U6D8o3+NuPSl
WiIK3/yBBpDLziq6t5EVhwqg7FLk8ld4ltkkf4rEu1qdX4C6+3sG4nxqhSokLsV8TGXiMdJ0GXvp
QG/01beT48d2tTI/6E0FkUoFGVaXwMJowrz+U0HzNxRgPmoB9ERoo0xSCxUDcLyhkc2vxt72zN7f
TcKXCJEM+DD4SN/I84RshwRj1ApAxwoCAFwt1uq/WoVM8TDaFODJKr19k52MXVN4OnuNl06VXFkJ
6nreprk4KCoCHDZ096DurYNTzGW1FatzfDthR37pXvTNQrqCARnWljDMVP4Ugc9K0eZe+MqoYSUY
+0jWc5GUrJ7zHvrwhjzEyUQzTeNl9emVPUVHaB/wEuTASlxmpUMQUOAicfZgZkKdDfgvyCfP8Unr
hrxBfYRzH0IxuEMpxcV52DNPi52aubXZY72Ij3d23tbLyIiXmKX69CdDTJ2F+s1aG7je1GBaDMuC
AUWoW6R7JJwWmO1dx2g3aETG/NLL6753Wb+2TYuhvJhEpn5B+4nJ+Smf9UqKaXPDSTberPu3gDi6
k3R+PNl7IK4LHh3vW9pY0rb0+0TuWSvOlo2cpRzQn3Ne2T+n2FpjAFmhfS0liOl4EtR2e83U3fOg
ZbwQvBbUqASihyF5vyciSWVB6xV0Y7fpa7E6/Gxrkv+8LXwhZMN2WnzMuUMsKII/pLpuzxuVtlVk
uES2FXHNPGQY3Bdye0yDt31UXx32Cdb7lwLS/BRdOtLrNnVidLP2KPcq4+kkNJz/dFIylZg1LJKc
CbYBDhdLL6MntXB0SpTxmQYmU5whaZj2oNwiJpokzL/dbXSqs8WHJamAH6ITbeMyECUvoI/65CWq
+5Yp3lVKH42A6c4y7Elq8WHzEGtIafNprftr7MVQEK/k/m6kx36yvwqOAYVv/7TIi8VR2+ctqR+I
zJWUPqwt+yj6bcpFkyER09rdwNrgTUDNJPg7RkTXs3n91+qtLbDxqUnyGj56JHb+TnYhGuAgZHCW
Ni3pC8DmK3/mFT7GgEkWHRiVLzRwUU5CL7KQOvDERq2L+Euc1yjj5i+yn0bzbAOUvMsx7sRZwFSi
BNH+WoUOGZAJhQ7D0ADTbffCktAl/uthAt8dDt5EYBz/hzU4NgthaOaQ0o/fVw+V97ZgNXhaY9Eb
++d/9kO7tnWAaBXSkCXqHMSStkmbo3VsBCKZGjcViYLzXil3bQyuUMpoK2fQ52vaI4SRRunvJF16
Fw+PrbFbWShWy8BJgJF2NXjuvKMEjOlQSy5m6+sdbIM3hg+6M6/KnPcnrRjXHJbjwlvK2t8O8Bxf
Iq/oNwV/bvTYKhKiWFePus8fALrADkIsn38x9rSCY2D7ZCfXmnohNaoqZ1EEztsRUDhrRGsUgMP0
80LzunRFG5/xtz9EYKqpxoZbhFOqnw8p7Gjs+hoQKyMfWQXTBGfBH4F/inMmMTjVvEoZcRBTmZyu
OHnCPd3kvNMPAeHozM8LdhipbwC9YqnXGnbKos6UwbwjAWM+YcoA2+dmEP69XVSiPvi0yAmh8Vuv
hA3yEFAgYLipfIvYzLpLZ7NLCSXHa8T/I1o6jgTuygjK2czHlMN142wJAqiH8OU1WcV3A9tm3lYa
lmaYSWUxB7PVj1O4lN6t0O51F+QkHnpU1YsX3GxQ4F3b/87BylcTkSlNO2VrSltbJ/WhgUEBJHMr
O3rYQS2czrvI2tHZVcawxC92VBoEQQbAqv8wNaj1DWECg1bSEPilStLnO7+zL2K3NaDAlH/wpbbB
+M8N+QDyzTFRdyzYz0aEZBclZH8x6DRqDj6ZX+3xwAan0tlv++bJKLqbuZqgHb+tITe5UfFMMDb0
fFUKt1n5mYy79hT86BEucgo0Pu6yyVmuLCg6EXJx4XYMRaLwwPlfxiwipXwOlDL2u6ISIdOptBWD
P2hKWCo8ezi/QOyE096UAGVEkdegjbxowciKe6gkSJ5y8xN8F2ySzOmkitnRU/p09ViGp2NE1Hmq
LXaN7Q8Y3xsZ8eg4D29B0Cn8icoCe88OILIkep+GMlpPG/6F3Ar5EJ83W9Aig5qtYwgdKRWEmY9/
bu+x9u0IPw7wthdDwXsO9q1iTUTZ67e8OdtFHWaH6qIhCUTINun5YGy1Zk0/6uk+pRR2kStofZxz
RvV57UGlQapTriACIBCRqnv8NRiJjNDVNDjoJV3pwMARouVujHL7EJGvzcCcHiZ09IKSlYPg3eUb
c3No3ouCpNXPr7pFb3onlck0BUzjz4CiBjQDPqpf7gT49+N1x1CFJAxbXGCg0TiJmvKbEKaItEPI
PlHcSY2ObP9JwkJNI7qpsBETpyM6rjmsYYG8Kx7AGoZeqYAOPwWNIuHcmc4zwqOPXvxjb4NzxrKh
ZtBKSNdP0iYHrHnoCaP4WGcr9tgt7DFtJztrRMC4bw+BBnyyFFGpjPswbRcGxSlg/biaiwGE8jUP
ZtoNUU1uo8Z6MmndpL5TF61btgieXGMUM9xOqnmHdeZqPwGKspBZQ1jHJIDLIYjd3Wfx9dI98Y0U
Ea5fQBGVYUTci7CMxzlmzryeNoiM/AfAPtB8I6ag3/uUm3Nso2FvIv3nUmxplFGFo5G8z+vplcGR
DpDIjG5MAuVOUKvPEOCjrWQqb2basxD5YTzdc87Dk30ALMWPZExnQjBaGVCjmrDXrh9WeIDPmeUc
lprKuosOpWAL/FedZIPvZFrVjXvglE9GnzGSKC3TXGQ2jZeeYTaclj/71WO2QaYvty4NPmkwb0Ua
wzZytpyzxnUp+eiRlpwi8sUzswl6s3G1KwNuWAo15i0XbQf8OitXy1tSmwSq9wGs1vChsgQ2swti
rxOQDykb4EDh713shC6LD8Ft8Tq948HHUmR3elb9NGGkojsrw/wqy8iYwj7YjgF7J/XOaWQ5cYpF
zo7OPhxcHpInAqiGe1DjtKVaYrFWiISsj6FuzgFvnjCKKUs5RwGVb6dAB3e6SqePkX3lLVtZthXt
YzNNBghfZY7fAtzueAVQ67vRyfI2bCr+/aui785/4a0kRi3JwYd2xG3LPe2xV55ip5uYTarJ5Cqu
SdAbOPN7k+NUb78VYkTbg7rvi4ewTFJLGhEMockHBSojJBJXm4F67eIi7cWGWnbbI/ecIx4U8mKB
IO+aHUfBEXGQjf7mF7pBd2zEzx4ht4FbquMjGpEGDD2Yt1I58RVfPOSuM/TsZDay223WRug7c82f
9HnhK3ajwPrIrbXzFW5UHPdSX+MHsj4wKW+wiHxxTQvnTV5X3Pww5488F9sAIIbZ9L4AXPIfwhS9
d+b0ILxEuJp2OUMy/LvWCEtsUYcLxHIaimGgVZ0KJB6lMxf6PDYPLreVsWSC8SolUWvm6SXg6ROA
iiwcCJHeBtSA1GI2UN3pV34zPt4dbFH1WfarzEuFePdzksaP/WxwY2VB95ZCyrMgcv55d19Z+spv
Oj5O+BagfHk4znt5t/ZqXviopM9Xb9XbbOwFqlhyt8kZKVgg+E27FZ6br//MJhDU0Cuq74iz4CGZ
DxSoH6nZzsYLB4mOlOs0oYptv8MHVtNzsJF/R9fppY8PjR2D7DVTV6r+AIyQNps0aMx6R11QddIV
DnaljcoVxG3imrsb0z8A7oS0HOW8p1hE3+5gycfI83s2SsrZSdmegyx7EFHGZRGHHdcmsB7cgm0x
aUM4VBjJ/VxdjE5wGdH6AV48UsF3hws0XQlf2tNuwLR6f1iHqJ3fhuMIbnq1cG+u0kSfK+bAlDh1
KVIUX6uz0Zn+QlGHcAVbrmjziR8Nujtsv3Y1oNA1SG3iau07lncNjw9UzcY6XWgQG9750R+4JiiX
kZA7LrAASMpT7BNIaOHZkHTzWD2JoCs4xGNwPCCuKRynfDN3PLUJdZmtUo7LTOpvTgrco69QiEqg
vRPVS/e04mhplDm79Ww0zns5qzHqnit/r1G9z9c2pGc2Lw3o5h4Q3qu9SrKRkfUmWNypSzLbY7B2
t0pg5uz1iGwn3IW3FgZTfIj5BD+pqgQJ6WnnPTRvs5+6sUK6lzY5nfxrZ4mGSrggUSGvN+anIdc2
FeOLzlXqD7/W6jN4lQFsEpQ8G4WAU4MJ7yH9MyFZOSByVfZ+vQXihmAolEaP8Y9UXKknP9dv2NUP
w3BTe4m+Ch51qZKQBP7vz5r3xIRPkooRnTZpUZ0T4pgWGvmNsl7zlDP053Zvg6d9TQRSDGLcwo3A
q0ShsjGfUw3iZz24bdwTSodZASFAUXVZqdxXdQ3kcFl50aaN5vyavxYSIpHtPl5DMrT0U/Z/r1iM
cBaHr7Ipak4fkzxDT/sLRWISni2msd4pdxyiCflh/7XcsYx3nYvM4SGK+2sM+eT+GADK/hhYIR9r
FiqnhASt0KDSatjmkm5L9DMRhx/WNep2L6W6XX2dkljNtf0cZDPHhR2HPGu3jHbi3Nf4Ewh6NfgV
65FlTKjZAatsn/rzRFJ6cKTVutAePCUglHACTFekrDnF1/Fgks42/jpqIA9uittwcsuxaAMquBqg
Fi7Xv2ogXTI/8s5dDr1z51rqE5NU+GFgUOWyhuA5FXHPOQHPzkEUYYBdAfFR3kKSbCdlHYVtaZP3
bBUwlxzYwnTHkYJor0geSSzMtjq7haWSbinAAwV9ECB7VMjdIGjA8rWVVnp6DuHPhuaSVUwuPuPt
euyGn5SxqC+JZQEVsnPMgP2E17CvrTQ3ZD3kFj1Iyv931xSCLxdpvDL+WTdPoA0D+tdx6+Oml+0g
KWUr3A8mysl1APf80srfOWGz/vTPfcf404BXu7oKsVDQmEzqNv8BQdTC5NoG6lzPnzrAAD+d04GZ
T8LxhxWmC08UQ3PnZ04B4rCRJCWNOWQ6VBNotoxAX73HTqsvPy4N84CE91FB/GTVq+qF9t9qf3JT
VivWqIS34+1RSWQIiAhVBhx9LruRV3EDtopDASAQFPtHtdnnsrRJpxRPPmYvv1ls4bbrF0HWf6/F
e9K6vVyZr2lMj56oCIKQP8V401ZQQqYtutoYtHeFbxM3OT7iQr7G8h+H/G6tqaa3LlUDNi2k78Q1
Py+3nw3v66XTpUVzzOXJE/ImlKQMc1RK9dNahsHLF+t6Ghw5XPSFPiVXAs+moYRzltPIAZEgAEa8
vJwO59cKDxLt0EX4oRhrnzOjiV6DAaZsdlQwipVxL6szC7tphDnWmPp5y7t26H87iCdD/iOLNe38
asyHdM5oKT55g8xq0XJ6sensrvO5Tw4zmu/Fh+0ojJzdYaFMeSbFEpsMH7F+GXLCE6snVgTOurV6
9Ruy45Nqx+fP2u81BZCGx6XhkD7liB5G6mXDODPjB44szbWBD89tmiduYXkphoNuIIzOtKXZTzDp
oTC3UO6iQUNHULQ5hQUPm4YVuOdxyG5vPCmKT8Oew5KOWzNtYR5ShGwtYLpAdIebfN2eO70wIydX
r/mPCBDO0VnZJ4FAXksghkzrFNNkEFVVN+tZ9TwmlLnc54NLD6QIXE1bwTclpoTJATBP3thAt0ag
DVHYNpjG8DcEftM6JrEmYODGdBS3nWOTbXhVYZlmOOGrQ3VroSRT6AmGZyeBxeJWnDVu1nsxcHEc
2HhvKJStbgY+Wn8rvXzvVttG25nEG71KvWj5K51XjnSod57qYnHnGTRPOhaSN8/LaO5TbPiwxS5T
RhCRHCAVj/Dn92/Y/Ff2emDdgOxDU4fkPNPKVlfue2NR6Nup5ehLrfExKrbO64frX41784BQZNhg
Zq1inHg33VutObTZPEggMg6LGHLacXnH8d4TYKk3cfGOi6+2CJRbEn5ABqb0/lfRYDVJRbjfWl3M
RhQdzEm+bedFhZZAgSs5HPaRbGgGI28SNLxgllTf1OaGTle0mfKlpCSppxDxHRXB6Tntw5/hVC4x
AmtptQT8nZffByEJi+xiG556z4lNL6lOy2N2633RcIcjQrmqiqrTzdaxRAwEQ12FjeSao50MZ6Y3
It4kjHTZCh2f001D4Hq0U5UPtIOktkZSsXwLlEOwokFxD92M1vnzc55owvEA+U2A7wFoAEe1l3Us
KyHhTnf6gNFZEoqv2SJWCWgK14PEJEy1DvWgetHmaXh8hIay6eL9376hN0156qe4Lnk7MpO2Bo6O
ZaudKBWf8QwrgpfG4Ul0GnaJZy4+NIXfNrAHMPT4RGemakbfFmy46sbIUhIR9p6glIiW7G3iLKQI
u+Y2G4y999V2lUcUUaMvXQfxaSI2v9X6tTgPz6vn0cJ2PIOfKADrPNMr6Hv54L0enNRidK9TP+ox
Xx9yCKrvkwgDg2LmykST/wXEg1g7UXiMUC+LBtpc06zTJjoH3zrbzDQdMKam0a+1KeehWsb7f2ij
PYVfjGuDQ1+5KftGM2VW8EEykLwJpHdyPsEJihdZsoBy1JEjVJbUfw03orINJIJRG7NB5FGcvm5a
ERnJMeQ/g8eyuT6kj3xWPNh/IkrLoM3q0MhNxOZkTgEPPJulLlze/5ib4BkSxx8xbO/ZWE75sjKW
z0eyHiqMIXGgo5l3FXKI6JN9UXtIsBlfab2ci6NnZwquKDlDRBzQd3nu5dXFfmo0CVGRbV+wmgve
YMHYA8R0B3l/QA61hO/u9KJYvsV7Q4HGLKIJUyZV9cSR785Oin5+qvLBM7RcqZEHT3AmkgxQEF+N
u3tAYkvmTG4WSxdkGyM0ljVYWo288X/dRnFy2oBkzk8QOsGoU7FS6+ycacJHlx01YYwLZvK/WcVm
Wka5K/KKjVC1w+1rBj1qGEiWPrJZ0QHS4y9WQ7gguFcZSqnY1cfcG7SgJyuqsT5BBlqdHj2CaQSS
4jSpDvCnLhrOMWyfYASLrQ4cwo6QHRURSv8UvOViELaAlPR+cFM8z+byy8jCRktshDU4RvNp03t+
1mdkzmX3KmS05eifqJ0y+HSRkxyGaxhlY4oU6d9cZRTwgSNM0GBZIMYLwrrM4+YSK7JRs/bxPDWc
FkapX7iFZCgobmfLzAadx8lIU5180U6mCNnurjqS4xecTF2Er8kb3Refy6LTtpNqDvVBnjBHsdvB
OiCtAsJBpzwyUc0iYH5Q3iWGrESqpKdek7Y6M3kA8uRlUeJfZTwjdTklmf1aY91pLxPrTU6bLXQv
TppMFPDvPF3xPB9KA6Ycl9+FgkLPCpdnspavT+9ElmCfXohXlP05ryA3WWX6GFqYFVrZD3zz6+n5
CKa5ofYGtZxDNsgICaJTreMut0mQeBEddnGImW1Xuvf9jkGykf/aTQFKtRNBw2pq+4tCrgGY6zCX
PZrBwOtseWQ/fjxkrbOq0kkzu6Mfo2j4Hg3McmC3E8sgB5/kkeOnmOR9M4v282z7IhfNzrxuFfmr
SsQu4SlVKJCRQnQdXzz6qdTTjshGCcYzCDwBSx7TmxKD+zoDBsB26RXUesoRl9c9h7Qq2dSwxTRB
atfIoFJSxncKFspqZGyo+xiS7jtA77rYCvZndA2BfxC0k7EKs/Oq4jBw+83uC3p6JGIN/0hl67l2
rOmnFcwAzv32krZ+F+JHO2QFZ3Yrp0e17q5EfLevqauANnTECnh7EM73diu+N6QlFYobRCI/5vYu
BVsCgtfpLpVHW0l+V/j8rlJzLlyJ/B+30Xv0M7c277Ca5Dax4qYsqQjj1a4RL2yWKR/VrCFpOM3q
aXBkiP/wUM1QEnM0Emq7hrpPrPM348Pn6EI2oCcFNUkcsDHgAJYddHWk4hXUQTUz22BU6LTMuR4c
3HWRxBc+Hlsv/dFxwCerSgAo2wgqtCofBVb5yCvLKrcQ+x6BO0KjuxSNuxdgWdPAoXRzAbbPKOHQ
/1d5ZHMNNKTny6vFovzAvRfeNbpNwIs0DfC6rxrgD0YrDPsslDS9uXwtPpu9I/Koo1hszATM1Kh+
7n6kilN+UhluSzN8A14QC3q3WC5w8vKWDGJ99Gamq6ZvrKIDcMJ8E7qTKM0hO3wckwLIcB60EaV7
oP2dcgRc0shCJOc1b51bMZ2+kDizyHCXW3js6f48k4Hxjr//iue413goB9m2CeGSxH2YxgfjPiEk
71BgNKu/NPmcmqSTeVVfcVPctuLh/gpGal4Vqr/7d3p9w5+MLbGpH8pACt+aY8QnMyEnXvkjPtyd
CAWPHEv4ruqqhitJ0+11sp40sWNcykhVREzU0OfY+8IlPMlNZsyXzvcIrqDsbTao9u3t3qMf0aM1
WUKLKh0oGwC/5ZGxS+ebsDvboFJ6dPtc1puKBvbW70rZslv3qSyjEIAsCET5YrwKdXb0BfeFSqEP
j+mf7shnZ/Y+zq45Em2CPgTLanKxmLaS3mWqErlKfn7FKBjZYjx1F1I66ptC0kJnOHX0vmd2K/Ty
kLOo0mj+sqEbjFpJ83rbjghpR8jBJTdTxJxARbuQ5zoyz80/fC/zNOrhpUpq2PV3I85N1R2vQ4yf
yGAk7U+3k1+t7tFmQmiKhLF3tGInpzj5PnhrW5C20X7U3tcTrI5DLUFCfcwMWXU4XUjaJmvNetfE
VfQRem2TAKvWhfrdDsRMa5rR0DJRlPU4qf0WTrkuJiylv9W+SMjYNb5MAcdfrNopwJba+OlThELa
n/bipPPJnwzCHaIq5p737/NQBIIyN8cmza88mZ9MLsaFITeAJqREkh1Z22AXnmQOYHiIM+M3OdQE
Tf2/4aicRyLpwKGzPIfAeMiMl2JmKEcdVvtfknFPUCMgDZV+Y3hAHfrgUwgZ2BYWFFjP1ksckqt/
aQEbLtIRuylXr7DL1pIYNbvR9Dezrckx2NGuONqHOJGMLwvpkyVm0LxkC0uMHSs9HQoHltYVK2rI
g0i1E7lHXj0eADuAXEnE2FJklvKxoUyIwxj+FhPG3d/UCypG6k5HkA7rs1AMct4giMl1o9vJi7tb
Bwi+5cOVeo/IwJ2U/lTVyO4cNU1TfbrtfiRdt7/bVCHonw7nhaNyXpsiXe8FpevEvWqWGqHmJhqT
iXdajNG0G6oHOfcWXO8m6K8eKRIJYxr8sk2dBHxgvpGnqEd2ijVSLOfnDJvqdsroCCfYk15SFXaw
+ePe+MfCMEKQgtpTuCRdVVYbNx4h1Y2VRcTYq1RMTg+wQnRVenOkJPVNGuGorSaH9FKstIzFWMfC
T5SbS9ZRLXPxccS8uLRH4dUqlQIQgo3Q/d2RTNKKQyLWaqkEav0fmkFw8ho5wEQG3tGDXBd86zhm
2Kvk8T0QxxmfIluZKaQxmCDbRD7FZSvCcx3FBIsQr1iPmFKvbYhHgunIrt8P1TGS8bYmIEODnY5O
PFQVHLbjP/OQoZOgjfyz+xaRG//U60TcBu2wvM1tmKE1EgSDN3w9gesxUX5pe6W4YmyFOK6AO6Uf
t6D4lLjBk4Sqa3Jr8Vin6rDVmoIis8DyXm6oRHWm5XcDl9+b9qd2qgCvFtVhhts4wNJPqDBzTB0E
+j5L2PNty+PnKuhXJ3WkjYLgaH8IlMlg3kihTS4W2tKcGIyTQ6/nGuRgBf0HMDM5yHdbVO7KgrHK
r5HhMYALwnsHCPkFgXEK/n5p2ubmOrKYl8zSeH1FKcvgX8luj7+VRR1QeO6PSCLZAHHPi3fQEbsH
gFTUn/oinxocKH7KeI4ehEPj5dxGA33x5+JwYwdqZbYJxMkwtqQhX7W79T4Phygh6frNoSVIWqrV
i3dHGdu/e1/QAhLGIlRLvjcG8TrH7TXhG853J/oazZC/g9zzMezkIhp9uOdIWfiT1gb+ct4MsIf1
yUX+sOaWqx7NXbPkT+8uLZB/ZWhjQ/LwaxjBQreEM7zRI6SDaUhAo0vqUtsa2Z3qe1qCJDDPUfIF
+s8Q3vm2kH5XEBWOkaie2B2IrTZmrlCX9hOanbJYIqtsYX5d/TI6lZR3AFQ5rMLtt29BssbuRmdZ
Bhceh4ZlHUqONM7gr5ym7Dk7T+yqF9V2s102zauesCwhBKKuOLbnxmFnvjjaPxbqOm6zejntJs7u
6kUy8Y3c9sSVDpJKi8WpCOSQjIrbKwwii83BJKqplXOzJcXRivaFOJm2kIy9x5LIgVaMwH13Mcok
LX1BgXFezu1gpIui1n+HNQz9vlqv1e/v9ZBEldLj5FLpI2/WRaaJY8aeVsIVlH1eyizN8RXz3TE9
7PtMhMFboQ5tVp3hWz6nrYk535MdHLrHWaEct3la6hamp22AHwXQHZHzU1sdmjr187/l4HOzMNF8
UBbc5CsL78Ww7EirNYRm3Yjq4YPUJdhuZIAccjo9DWdAYV/1+s1RNP5jcchBZ49L65jZ/iEfdPqP
P3IP6kLHn3Kak9m8uTvcX/3O+vuOyLvHvFmkJ6C0Si3e9fI5RJ4cQNR2/UogCoB/J+b2ZcxRLOh1
9cwLVedxzWIqiQhGvmZaW6aUfNl6rvSSHrEfCkz6Ll8lj9Mly0bWPNBJfQxerCK1egtilBw2ldnz
KMIpDvcsl1B78N9lzAY1++/Hl8j0t7xL62tQG22z70DgZHuzDQFftuTRyyeIjRz1c2CdvJjDYwC0
kljl3oZts4W1UOzYEZblhh1si6X4W6YbTvOA8Hk1OfenNo6qegwIyQ3i4Q9egPy30H1+K0t6i4A5
7qcX4DoAtRF8j7WAaVHlg6sKK+NRkDrol/ErW2abBE1xjqdjRv3HPW4t0+CbDju5sQ59yIB0qH07
ywh5SPhEq9kK1wq/8UxvJk8jcDJv2vXCQ8/jidM8cuDYJLcY5eUIyTR7sIyFD2dUChCufHFKWbC/
aE+g8P8d3oCo/+hCIV+XTxe3MyH83ashPqZ1ytD+2xDqfBhHLLrLWa3J+dLfhtm34VUUY+NWz1cX
Xfse9q1jukq6ABxIzu/kWMs+Xyi02rLjjKIoV8kDsPIVSOf6mLnGLFUgwNxqSXyI/x/y9W7OlGLJ
EcAUdZPbYpGwwmMOes3uyhhnWtB5hgXhOiIooT/jc1UUvrYbsvpl/MO7yxxhRd2x7STsc2ipYce3
niECo/SFxykfG0kv/lW2JowCZA39h23Nm9mWQ5G7VJPnLudyyFGLKz5GwX2+QnD9RETdJKldwnSt
+uGl9WCEK6SMVmatgZFaqoPhbijnFojPnjdIR7P2t+BJz1dERjrqwlfJLXNBQon1Wzgfdl4MVqJi
soG55CmgWkRZ1lpmUEb7ue2qU9aqFKbobAqLCL3B1lD/GXt10q4c2P7jMIlg48t7AVE44KpxdE6M
al8d4Ce5huUpddk2RtN6qyjegzgijZRKJNpAz/t7qzHqF3bMesE2hRP+cfXj7eo9gVVuHQoldRxt
Gby7/J8hPhovA7LIY3TLKQ+V5SNygcWg3eUPbj2H5ndVhBM23/yG0gnkE2KBJmIHvKqqHeRfgp86
D0YXbd5W7LQndq+C5mZrAyMpblFinBp1IpQM3ctkVdrRisvDUbjmHtVbwYbmBn/EGMIL0dAIzAiO
k+Khz+6EkOSp9qQIdfPBdH4E94OSgJwqBqxhGVyn/cFiXij1Yd3BJNL+qxPMQRFMdJuz1N58XguP
lm4OZ2twFQuzg6dA0NQcdMhjcvkVktLvZiixyVb28EhX1qaYhEfc1cm3rJAj2yYqf7JqLn+7YAcl
tVKembAH2tzBcCojcY4wiygJJ/E4yKq/bRTg99DgpvMB4/xGcdBXyhleyWbQ4Fd5Wzk4tacjv7YS
mzTdKKQ46YxXHgL7f7lm0fxxy1YrtbfSjezLof7aMBLokMLVkfY6vHB+4uc65AWLOzYOCV0D1dc5
BX7TAEH4nKxx2ptZF6gPBJx2waYSV43PykKmZjZS7C6kDAuMlr3efj/xuov36VtAPzc/5l0HmbtA
Z1BBuyV5MJT65FQ2+YOH5pnsllj+nJZsUapUxZ4/rCaZ7abf+V7dOcnZaNuTPfO0PBXI2nHopIk9
0M1momi+B4F9SACufFFGbw3bC7JhDTeHkoFVtlXnqHYyPAsLLE3AlpzG3Hqo5hwJndhPvslWQD/e
cCAINYTxyBcFX9B2nkgKCyCNoIyJ2cuGXEvzoVVr8pFDgsiTf5LRmsIzXwhJY0hlgc7a2zssNJnC
0/L5iIhxyH3VoOdwH//GhtqaqzjzVsSAh1bFoVXmb0jo1l483ZNsIRie2wRzGmgVMYOWnvXqx8+K
qXVk+WBsSoNVFuUc4NUNEHqKSFAYNplq3NZiEnt9CIEgqAgvsZnd0sJ+UnNyvWDePnT6fItGBbuT
DNRf6swejn3AcdOz5TbUgaTohgidgrKksVXx1TCpB5xt/vL+/H7l+WjvOs8JPlmCbo/IE6O7jDVo
Di7B2qkivCT8+ZrGQGylnI3DtIOBhdJfzg4Q8P28czEMjCCt9KFx4cbuafDv/QAVZPFeqSpDwozh
Src+bwVmVn6ZOGoz7jEsfEwtzU2oxuKKqOUXhlXUJdN32nTgcfQy3GhU8ou9+7U2o7eRoWM6Msj5
JF+C8VImqpOCtTx1C9vDj/nlPVpETIxw28aiqaYv+x+m7NRB4d+E4XM647WKV8ocv2l2iAtocwHF
Umbct5MCSiI7MrkkRwSBnP4NQNX5M8zroDnHwcsJExfNfq6GMGDE3QjBSoRGJF7Pj/oIgoSibLNO
Insi7uXk8PYZREs+YeLRwIe+zrSyDxxvLNnBe2jSbgTFtmboHd97PFBfYbYyuLn2DH7pRNc8+iYF
zD/rKWQocD0QY4BgD/dynIx32u5naLbzSyLE5LkPjVOWA+ZKZvgaQvhgwneaVePGy0kU39/NxgIO
VCtxfh9XfQGZsg430gGnXz/dL6pM95hTtDq2E2Kkqg6ErYDZAIm9QAMN/R76JnwOQcBnXmMrK3FL
FfqyIZxVtft398WFk2llA6xAN+IMtvizQrrw/qO0I2LoAU3sdUfhYoubGFrW9LdLOiFa26wxgc8C
tkiH2K2mC6pZ/RkgJSM5O3+vZI7CscjUcD/2OcEJzP2IJxyBYvHqxZu86OYyQ6e1/76jCZN7q75N
K//kLpIlNBm0YCMCv+IOrW6qb/cOMOTVuOLBOi+8ims2CglmdXWlPJKumAZTYQH5So1x/X9fkRFp
FBluiOzGgnCScuiz2fDLt8VPky0q9dC0XyfW9jH8wO4v/NPLsCE1EHRolLMt3mM7rGAOHT580BRy
QuQJ/+cGzMHc1LvBA+SGKxd2Pruo5bZ/fDyRFq9Lx7iN/CEpdVeYHADae2IV5AzhdLj5F6ZaIHKf
yBW2XtRmUOEG39dZT31HUioj1xlikvoWjWCNyCW7eX7Erc6McXHAXWjVTV9eRXTxI9WYuU7H6aF+
xHWf9JKYQSdPhOzqZqaqCSRI79qhe4RI6RP/NyMCXZ1PXFyHnmQFnC7+fkJkQumrGEM8il9mwFLj
gIIDSVK1LoPd9j3oqclWihfD91FFM3G87IL1k09mDvxlL18f6W51Tv9TNVGtf9KHtn8XLKyZOUzx
B2rYIj6+WlPjlGC+pPJfgUEC6IZSj9i6i7OQozKselwNj836v0QWku7ZUY0WuRUbRP8DoepKwg3Q
NxomTtJGv2/fgMAXqZMrWaW1OA4zHQDy6ies1JKLIYU8PKYvYw+m/UW3jQp9MTdSY/1GmVJqkLfS
X9fgF2Ugb8TW5WOGFluedMD2nlRmIw9xVy/BCuu3FM1J5vMcS8iufX7r+XhLV0Lnh3V9GfCKJYhx
U3KxafQtaLVvo1WKROfP6CD6h17M6bVF0tJC+StbezTUjpRBaGFFJnO/xLX02MQfrHR/3GgQFP2d
m7RwBl98ZLIHvpPg3DCOy1+KOiSE6Ak3S5SqTu8LIDphrUw909aLoWLMcOBXJp//BbKsjiy1vZXF
RzdVkL/9dWvTbLHBue/+6Dr7LZmzJwFa5rFteNifOKyM2kMxSZYym46TLmkXrPPXngchOmXbaoG7
l6N+bmJRNddyFrIWh//yfPTOLt1LvafTyGkwu1dxmK7M61MjDQaLQtv/y8gbRYNn3Ckw+d0PMs9/
YNwtA0Es6zvC924CAa1ufyw5m5eIaQfjvX/dq5MLG1eeLIsxOdu4R5iDIxjhuGZFAeNAB31WoB13
8B+MlTbTkxFkEbywcQXNJnT4eh951966kGIQGtfMKTtGbLLfGYstn4r/4dP2urbWa/8X79TZNqoi
fXMeH6Fq9xpKh7jH5n25KYcl5LEpM7lbEdVY9Pm3X95ocWfg7/0a4vRNHlInIUeaMsgM7YpsJmgW
ZFj6NqBLuO4lSHZdIuKwnc0VhqXYxsd+xU2utzpARhdgIWMqRNXIYt8HeF9cnVlQOBhe+htJK7RG
/i+mws5BrwSqKBJK0vNSOHrh+6JRJHJgO5M9nhCSqQX+z1PcDuI1Nf4ZWLoqnC/+/IjfoInbtlu2
27HvekwSXBRtRhKHbnwGSLBU5TB1tbK29WBi5FfFFz/wgPIRZaT9PfcdOZlKmOzWfhb6qpL0RuDy
qgSL+M6lT7ZJOqcMNAJl2Vh1alu2u5B5ypWiD/QqlCsFcDevH0KQEcGr6ssJjJqKplkJxrrF6+wY
utf/jYUb35Wp9pUrcy3hFY/Cw3EWtSLdA9HNKkw8/9ktAZ8wkz0w8bBerSpq5G7ij4vRK4wjfewu
3S7Df5iULLvLN1fCgNrPlwgMXf8rXTW/Zj3Y5k+WJFYnmjOPHLfh4Hkp2RrYY1cbZfRHePsxS5Yi
sNGUcAT5ObFPHky95MbpYT77AlcusmZtrQbIFRUKb6UafZCwIZ2wzx/2EJItw6iC1QxYc3rIZAVu
YmrH/ehhg1dgI0GCTKTGJGUg/QObucAJ+927rAGVk56m6+GNIj52ye5cqB4EtIPQwveWsrMZNPJK
eEYbCN9A4fRDt7DdyCT1L0wrEqirDg8pwcNq/seTWw6j6kB5APWICgWknjj8LV0NYQZQhg9nWeb4
za7fwqp5bOAv8bOvztptT4HbJ8aWfz2J3FqWsOcpZhAc1o+ic2b7q/YLLuydNoz04UYTm/0ozDCZ
MUzLYdgz+dbAbeOJdL2HabQwuV15Hdh0DDruTeyigp4Erb7MVn6hpKXXGau5aDs/IU2/KGZ+b7H0
qVxInJbpLC5ORIfqwYdrgiebMFBavdsp0m1N9btOwbztrbGkaibz6k+evCcTscaewN9tG96eKRiR
Q3ZUVZXDUOl3nWD+YoFLz0vbFN3pAa3Bh7/aEVkikTc7RpswyTeejunpxBv7EBCcy4/Mje/dhR7k
Dr1KBcvifbYGiWcrwd8/BL0d+t+EGsmtiHWebgTNuverf+M9pGef3Brld5w1saPt8wO58Fa/r8HZ
FRQdpywtrp7YshMYdBX/0a0Nq8Git8rrCPsqKqfilhJ2swTQY1oLyeXXf5g2k7JkcMG3b3+YrF+1
G987Z43Mx7RgwjhrOB2z6o/1kFAxUHrgEAOOfx2H2H2EEXCWKUV0+bYsVRLbxrgDT2CiezPXCeCO
e5PG0/hbFDM8o6+vUD8//xmckgLFDc4jTBhn6T+gmhst+Ar/QkdvF1CXY2tQT9XmUKowsuakKdUk
JVR8k3/oVp/3/D9yXtnEAdeiq7e8/G4N5Dg75C7Kg35X/xYG1uCClM12RtzORbD4T37g8YqR+gFv
4a5l90W4NSKyaE5vBR1ccnRXbYiIeHM4nqYtzNLzPFPB1fFO4SEc6v49PVNU2OrM6AQKNNqQ+T5U
pERjCrWSoV8fOquz33myprtzRAxekZWXMaRhNCjT4gIqZg0bVj5fwT+s6LLlRg8zsWB7GHfORF94
MmSSzLIY8XBAFLhJkID1x88cp5Q+DJ84l/6FG5mbAtmardgbq/Foj7VAj+ZJrDMHoZHa0Yi9Vedr
ttsBQOEw1xC69qFWwkwcMOdfUh6Lhf3r+8Q/TWLi0INN77+x9W/YOYUSkDcIU2Yd7vz2dsCe+l8u
dlww5lXTGSjRtXqjZCVaNurSq1vQXzhleWqtTLo9G0nTimax7BnfXuneO9hLZCrMz4sI87TpDE5Z
pFYI7VOH5oIINA5Ns1MSe5tmQ/C1q22UJdBDLu8o8EGJEQ30vmPaU6XagiuH5lorfR0v5DYf1zpi
JxOEJmV/ldzvJ9PULVXCkj/+y8BdI17/OPxAcw0M4L7Gqgw2bC+Mti88GVY8HxqniVCoZM5ndHA9
t8W92vQjS/PJUOOOvBekE76p/FME+sy/l8F1hM6HXd6gpqZD+lR7TlRtIG8O6bKHj5YID4zMrEfY
nbsfpwUpRTAf6kyy5aSxpEVZ8zGM0XLKrFkbGrguzXFRo1aQwMfmMEM7dV4NT3UxjAWWQIjX6ZQq
phOH4ToL2Y4Qfsv7UWigZ/h1agtT+j5btEsORB3m58dKte0mC/wLzNa3FZG+/0GsFQEBSTOS35rp
E9bOGlX2Vq3F4s/pIE64cI1Of+HmIkk1cWCmARCXss36qH//x06o79dOuiJCw1VnJwxgUBNaRDhm
KH5eRCzBx/50Cd9DMY96RX2gUlJinmscR9ojBXS7qDUsEn/VYKgQAaZ7WBKK0KitkSct/UrHj6vM
1iZ7kCJB6giZbQKx2A4vwjX0Ek1ZFmaOT/P616ePe/ZZLgroNOeZSPIFtXEYsP/u1LaLEqzVCVHE
r9U7cEHRmAf/UmeYyUxbaM4APiuf6OkSF150FrrjpsPmoFU3wBD3HWMnK8RunVUBxVf8Nb7Vsh/B
ArwuIDeuEG79lSQs1751QHZhAO1UdPI+RlyahuHAAFWhcnsfDrJR+NgMxWBtveTZeosD6rQTrLDc
vGj2VVvgWoSnr6GFA3UQ1THcIfitBwQd7mJ09LAH/Fhv45diavKNczxrUdxPVufrjHpFfQ4SdJSx
HYa3RtXt3qVkbzIIA/4waHCmPc8bAhniT1rq7LNObUyEyvOEWs8FG1lgxvl8SoS/QtWMaD90ezPA
6NeBfQYHpDxVTXBnc+JnSGGyTba4CkZ8CcQDCbajqUtAd04yJcCYjvm+MghxiSYroyfrUGZFnjpB
/mywumyKFoJeVrdyTfcq/xqjjIR5RvK1mJLBItxMXruQeRt5oDXnz1eGiqQupCysjQM0hMa2LAOY
hwiat/MxuxWlb8kEwP4WsvezRs5Is+yT2h1PKJeSqMx9xHEITaRaK3iqaBWlB5Iv6ZUAVRvv2FTG
SdUq/+EeJkuK+T3ZzfNnyr9wWe9/iMoF19FCnqBib2XFegFlp+FKn+NWNFjGFD4KAbbw6TvZ/SRO
Dpb48WSB6gomkx66ji6/YRrk+wJyIfT1KpOZ8oNuW2irQAQOUTRFpCZo2bo2/pB8cbHce+dvWFp4
yfh4HMjQHAwDTonE6MaU4HJbekMdXTtH3ya7Gr0K4L52w3tXm7m+l5992MxXhdqUpWtYa/sUaQj5
4KegOFO/uIlzeOeK0fGCO7zSHxlFE+qgCGFmtrP065l4XCga1bO9V7AHp0J8cBEZ4A+Q03YY/d6v
MDcxgiaGg0Y8RWRPUPoduvojo3ZGhBtYy4L1pFjuI0Gnymo0gJobZvQm7PPvw/2U7YF/uUcwin6u
W1gDtbIT+OeUNSj4GONibezPlv/qufOJAU2TQnaN9iNQt9y3HprgvQSLaKc+0MLreJWAhza0hrX9
ywagOGouaeo=
`protect end_protected

