

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UTmxs0OkmJURXBOVdUGR7t0vPgcBU0oVnrXWTlGh9ogLy+aZVadnSNImcgn+4jLE3/0AXAxZXQ82
Xbw5u5ikwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NDHq9z13OnSHCjB5ixLI6v+O9siiJNJuJRP5KO7VWFUgsdEdfLm2msHdSHMZWHSOwKZ3fpyDnmNx
BgNrMCYycBeI/rO2pKL2N4HQAMnhKOZtiPFF9n2RUplezsx3A1KtfrZPlHnD/UnZMT1dsl6klarx
WHWoOj2BdFWF78jqP/k=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pd1c/MzUc/ohRsjBZ9c2FYMEVEx0/T+c02CO5nj1hjCkjBTD1iExW4b2fGAqq2hXvApptvjN3kao
diEYImrFYF0oK+4fJDQ0NDCFSHEPkV9IuYgpAy5fNfC1Dx9rVAZAI1tVIUXAIZsy7oaGc/ReA3s3
/Ev1+YSM6X62ouq0EXc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ds2lszdMaBUWm49P9ovDqEJCNyznNiiJV1s10TsqQV85Goa2s6Y0q2oK0nkUurPC2r1U/lFQ6UkY
FyQj83Ie6eOpnawKkK55JF60SUgc/KJzJ7bDwIpaZjrpb+XlrqrzZU73J8jBBHKLoF1/Njgvn5Ad
h9N2MGH8gaas+uT9uDuZCA+ii46LQ3K2yd1YWXKK4uzoENDnOnWVcV9omYQiZt2WoMmuDtnHiiD6
BU9fNvTDJc2E+yqoRZLq/i7Vp6O2raEB1EabQzrK+1rVqoRBidd5D+df98jf+SVXW4uK81yOCvMA
LOV3/ZU0qCRQoJbwjKLC39h49ly0sWjEpfW/gQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
df0vCAvcFSWs5BffbtXlfaFIBd83+wey54D1uX3YAx267SlsUp8LU636/ulbSzkGShRGyHAsajTQ
lak4/g7ql/uNS4cPDTprvz1MsadnxOACDABIUOl7lg4w0zjMlnHliJydcn6lPMrRHgqJ6QJh1Ypj
8in4rFzqjprqSxw1d/10YsZZxkQoba/tmtftne+6yGg56W2Fvkku/OTLhJ4+2k81Et3P6Hl8rQs8
H3zDC5jgcWutFMz9ATChQpuoW1Bt6ol0u96wp5xiZl1ORv7DkneMNq66FiXR7uQAikRnfSIiT6/5
QAjuFDJ9beaONJ/7PX0YKv+VUGzRFq0ZFYEUEQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nCZ8D9A90hmHjnYoY13nJu1ipj+rg1ZVc4+qcqLwK/I4sVkFzYXzOHfQZXQ7YKW8qcQwr7Ja8l+y
rmS/aej2Bl+/GBm2e8OPwXjYQfJZAcWrX3bukYUhs960X48k+oy8IM2fpLqIO5UjCHWUKDAmMH8s
veeZjDOkDvXS6zx4x9hZL9OB3MW0oK6L//tk4UtxPcVZEJmBR7mpHfQdetJlD12R2NEAOMEs9GYi
egJoRgy2DcxVo/qhMUxikMoNK8DRbPimHxnf/gi8Ss6Awc1pw8Haokg7dho4WvcGQs5jULvRh435
wbmLZ1FnvnxhHSbLJwY8aBTSiBsD5Jozey23DQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504800)
`protect data_block
bfQPtBYpr/T2HHZpq/M+5JlfAt5urBOX8ih75n2IZjT2OOXX8TH4MrYacgzFuYrzqDqPysbKpUAA
hh4K5MjHizmYQEgjJBA4DKw7id1j12BWS6jpU76e/Vz259wf3/RpQaV3X8AbY0GzwWWXshHOdYjB
kI7jnNeOy0CQ+1RGe/e1CN9ZRQ6zdCZ3YBYkqS0e3KHZ9L/oYC3uHVBT0dcqk5tA/2sP5bYbh/2F
B8B3h4PTzs5kO/LcfnA8bEw7SJyNgYOA05R7QZSAJPRL3EGgEJtsSHSo1hYJLgjvke7vySACrpXp
bCzb+scbCyNFx4bYxnE02BMafClv6c29nR1t9CG0C2SpcT/CfXM/WQZfX7Y5HMHXRwKDxsad6dBf
kMgQKN92A5eylZeaW7DqyKv9Ib4t8Kz2B7bdRHIMf8JyqvFQ9dZ3leDO3mqAmbRq3C4dzfxREtUU
B5ljt7UXdXlWSGbVcsyhBq/r0CIbq1050XxqHJlnOhviJyeN1e093EYtWWbPQtV009zY1Dh89aKu
8w/36m8mKzAY+2yDZvYuVMZ6XEKFeMiIFFo9SI787WE5hWnGu0C2Ibni69eq6p9tA+kiI0IWSyaR
91iarhlEH1Lvfb5AAFKPghlwpF89fXyGVeaXiQmYYVU08ztxFvEU7LxrDwRSb/1t/LUB4YbNuTTa
EP9Jz2e3UVz6lujSaJd9e+lDXYfD9eYSJ3JpvxKjJy5RIbWu+yXjZdua/aRacOk+Od9ZzyH9DfNZ
UOu4T/JOA3B+bk1ly/sZYffpWJhKIKMlIYVCOcRETVfGhQNUwIvF+LLOapkNiZrtBeUcTr5ZEAZO
rP2llneJkHivZRD/ho9Gik10pjE0FD2jKAb5ldyXKjRQyi7apLDzgDIsnA45JFLaOmbiJZ+8cymA
65H3cou8phlbLfO3Wh9YKWdecldQXCS/2TOVsU1hQcmUa+ZZe4+Rel6h2p4hLnx9XF30pyLAuvrs
JS6hA35685iYWtDButqAzWiDSgnhPXEDtCeRDMX88/ZzgzO4IWnLzoYpMU/iUmpSMkvoJLLfuBzU
kH84cyigtCRCZP1EjPMKeWt5caGIv+P055l0X7zgajj5Vume2gTfj3P7dIJK282OJzjT1zyntPcn
XHp2x9008B/1rzN9Nq4x3emlZsPe6XmoJ3hJNY5XM+nToYWDTLJMmKvmK6AhNs9ikYbb31Xv8sYO
EBmexxFeewVotExUr2vIZC18VnbPOay8INup/Fq4W7+onwrMj9jSRq4cjNOucQ+FQxarvrosr4bQ
SV8jxohGbTnZXFx4N3S05PiLRiXR6lwdXY5cjSE028hkcQwVEMFLBcTAuwCaWo4rT094LSeebYHP
8bMzv7ENCZDQi1Wy8sz/IJSmgN0jQihjT9D8Roy/KaO1dxcY9zJal4ySdjca+JmYmGdhg8jBibph
ONvFAF5GWQtFow7ywMrA1XCWpAkM5kVr8Wsc47oNrIoagnaZsYA8wr6/jru3VGEpfbY/VIUhT1D9
9O8wkSer50YwQw+PVRaJGLtYZ8mvV9JyoGY2TSv41sZK4g2wUbSkfPKkHEXS4SeixWIhs3QvaBxG
9nfPnx5xnHi+T1jyv3iYsu8fY3J56m218cH7rJrd9zy/jYxNfw4V8guM2b6ZoYx3QF+RvOZPbn9E
l60y9+BflV2xQA9yKkqshWnTmdJzMv7rb+czi4nDFXwrhaYs9vV31zt3kAfeojHLEocp9WwuUczt
xguNtX0B0MuQAViOyYFeun8kvas+h8sPGkKKJ2IQW8lJr1dikphUJWg5aKIMG0qvaxGAJQsighjZ
lTeAK4imykSp7YqA78PvuA6MK8WyhLMxu8zqqMvibEk0d/KxsEiaKX++u3VaUAFLHjnIxNhqzbuf
COSlSkEo0JIzdxXknNRj9NaAfeVYy/zHulYKqQ2D6l3qZN/J4Op92eOkJw7oNf1tOOPueyqtf5vv
OEs1QkIP7BxDz/b3Eg7KVOMBn4o7H3xEAxUOxSljHTq/z5Nx7FFuQIK8j7jSWorgOJi9t2Oy07XC
mXMYSC3h2iZzUq+cssQ5rrvggXudHI/J2XtWTsUYA0lDekcMGcsKsMbVVNfkzbHe+K8qJay+810A
PsKiNMjx0GbxWY+QcaAF3pyNmUzzN1riHU72qiolmijsBFsbLfAqM1q1Kpz78djjLIGBWAchk9Qn
2bjtl+CPByJewy8FiiVbtvf3Gmvb2aHA1abyK+CyoN0YCtZYTLnKYomYiM8nkvs6sR0Vt9mfStwd
tKpaL1Zt8d6IV/f1AzA1cW7hp4sG0Yh4Sc9A0SPY11AykVVjZFP1mbNl3Q7SfNbgiqL0cflEwZQ3
q2i4VPeE3AIYdbQdSoZiB4umnhwuT0n80wzPzcAHzhkYiqm2zOT84Fr35Yj7tBRJzhIXvfFDjk2/
96mfGb46S4CBoiEctTQUc7hksZUYHAUVkOAftqG44y9f1gkuPSUsDnrdSWM+CZn48oFrPL6iZLJV
CuB+TdPJBBTDJHNTXwGpaKeehR10LZSlQOE8aj1lKoGpWybgZY6SejQqBJg837+NoiVIE5/ahlWI
AIKajIR19BqUn/7uUt0sW246tG4ffmD+A9LeJus2UmzdsjBJlbxwSBiLc+kiBvKt9b/1hr4oM1IR
sBiuJKyjp8AkUT2fMis3pv6uPvuz0r0fVuDB4vTZLk7VqlZsoMxH/bTL+XINFtTcO/Qcrz60nOPs
HMtEozUoi4KiOL+E4yHqs1GCvwXErz2SzsUy3kgjgpBjs+cDy6KoGb69Eetn5WnzCuYKwTKMk2VT
gwU/XDqQ+kmlR7Ct1VRcoNraFJQ57q059aOx8uetIkUtF1h5I1TUzSIB8RFmr7WuLzpXre3uGFWH
BhArmYoXu0MYZ+4WDNjxeOJHsMtP7wtVSMHXGvvgJ6okD5op2E5w7SW5Lx9mmLJh04IOCbi1x0H5
ngjGA1GKCkz14xfzEHWX17p8nAXvGpBw1MnXOYgsiKGN1hrFB1ubn20oDoOdtuJyzSSftoW91wJo
4cm0ZTSmcPy1bQgs/n3oRQbYRy2JgVDrjopjopdl4nQ8k5gEYRRESPEmeEGdx0UKhy6OTqZK9OMD
V33P/yBduxNBu9bqlUBmlkGGQ9y8z/97SJk+uPZaQN7GJB1vIajmMKChlLkNwz1jxYhRbsmxO3Us
tE88TaNSclqysGjD4NgbAbv9Tk53UWvmzvhNyrDuR4UrbSVK+byfWesqk/2XcTjg55SVCGh03syI
XP2rQdVege+6PkYIAnx6avjH/k7e+QBBRWAcrdvnQjm5B4NWTNOHsO5PfmOw4OymojroXuSzpHS7
Uo7K6ixsAhnA647ClFQH/VCGQCSqeqJJ0cFI1GEbIpec7D90vaFs2rfY2En3F7y6+0ZOz5195+YH
HFkeXuflzZqpCZw8RUb+GcslcSr1a4yJxzZFmjX6TG4QSKqSyKnrh2oiNLYbdeZKv5rmBdU9U4s5
ekXrmMryAaxHZ71cIfSAnUvu2jDkHbYldgqjYTUPLygYri2ceEMzW9x11eiX5Xi832znlOEgRIxl
L9AMUQ+KuYn8QA2m8u0wI8s9gBykeZZrogBB35VvIG0SEHHvzlMau3X58e9MHJBATrUDhwJkq+uh
LJcDPDF9i+tRZrryoq6YXXXLkSj78KkCvTllDhA80exEQYwYfqUkArXaV+r3C/u+ywsDimPiLrT2
y4+XqDSLAmQsGZ5Xq8oIzupJrix+NjGgHHJKYS3bgNpadHrXxUbS+yda17+mdqJ7nACIHrBlAPvo
SQc+hSBzG8Vnei32g8mRPPXw9vxk1x/ZYgfPpHTCCLXFumZHqyOBZyBAv6U4nxiuHEC+icngWNzq
G2ysSc+C3DbrAbeHiXHMdBYZe4wCtBzJ+FCa//vWYO/GWhCWH4Rpw3MVv+tI+cP22cH1+PWAOo0g
fGdlS8mwzs07F1qItLhIIIyhqDPyjBNqhvp17V1+BLgj8aFI4MEb15QWBMRhlbcCz5mOQg6QPtzi
FPvEEzgfuU/e0BdcrCKEv+xJUi4wSwXfHs2Y5cH/b0AehI77MHReeuV84E6eHVGaUIUZD5ZbWhpm
5gsEObXhlNsyNtlII2PUN63CQwOsgdg3H1QJCvvlheAMsyhOg7ks8YGKRbV8aOsUSjHd/41Gv6vr
2M5x1YC5synMFw5zenF0bsjrJZ3fFuBYRY3eiO+eCbk9rgMu0i9/oZFzkOahj7FIO6Mt/RniCGB/
hZk0gUcQQeMVstxTZYlHmRfWmIATZchBRfAthqp+WrlhJ5RLAzf7yH5Yz3JG05kayaWdU9hdYSBQ
IpOLFhzDoOs3bizNSbBc1nEAxiCNEusRlEYgzQ98+Sz7b4N8Va9D/NEGg0JxyOT9nCNxz7ViDUG7
13T4SFSk6OEuce7Kz6eL50W2rJIDfQrGl9tThyUGHKKz7OpC2KeWIhcMoz3qYwehxbQx/5epGkSf
4NRoSvJ5AJJdo31VF7vYAKsraJt+tkcNLg4T9j2snt5v16L0i6k1FmjQddN/NQvXhGFxPZDyj3o5
RhxPd6FLQbitqjKuS+n0sAZTEQbB30/oirolA6lKp1frwAMnXOWJDDgUhA8nUuNzo2NHQ+RSEjeH
IYiRR/aDyuYwfGVPGkw8wEQbgKYPbjbN0Wrjy2Cn8HlaZQ8NjKHXMZCa3YjcveHTQYJQj/Zackav
BMSRIszrSO2ZegjRPUMillP0kTW6mIaO6bEm+oAFIGCcjF4pWw4TUqpDmfz7xwl4R9Lak5mhIGQG
kqIsAPYEepn9q4sgvNOqZ5q8yDg+UqC/unm9va+3Oj2aKmVfnxNypvUvlNw1gsH0pI+blAv9Rud4
4IHIQrZFndM8fsyQiurcBf4WefVZdgdyZmzZRWjc37nOPSRgaaWFZtHPpQ2Lt2+cJFGthOcldGeT
SDKIj1rS+QJgkT6AMSnzA3EMsvJ48uBhLXhP7JdEG/7ceBSrWQ7yAzaHE9sL6cAEFf3rbSnUyaVK
YkMHcaayF/4hWJGaBewFFvbpzQYsn6bkMYXkwUhtkBiMAF+OghQlfWfEpY3ZNckOyvYfzKKv6xol
UaPq3eOQV5M4e1yL4R1vcD3kRE2qcJHlWnkCXrMrnXvt8oWUh+hWd5EANCNivQQtPNdhB8TrOGaW
drDy1bsqrBFVRrCNHaSGSU4iWEyR+bo/0wZgw2jCzGluX1AJ7Y71PZ7FmRcpOomakQF+/htxbGX6
Jmj2TtVTYqaN45Vm+tLakx0ge2TjixVamFb7gj33lSDgF7D6qKSVZNKs0UNI5C0LBP6JWSlx5P4e
5gZxmDgvqKRWp5asZ2xsA8v1CkwdNwpzPGXK7M8dXvZbuGgYa6RZ4oukqMtkjPVvcMggy3zrSehu
SWedkOL4MLJQTVvF1LOlGDsv3T7zRg34KXPje+WGKTDGoXWyh+HNQgMk2yZk2r7JFfy89kfIjHgk
YnojKSaNDz3hSMlEgWjb+r++qxUoi99L+2uhD867RDv3ZT9GYoz3kMxTdsw03UvRennZE+ZdTnyu
OMzt3SZwS83GJzCrv1vI8g+jX55GMo/xAkPdFp1wG1xnPlWNyN568M18wZxFwruVBApCP+5JIChe
sxbNTX8fFuUTrYFgOgFzNdsvh8STQvTYKxNVEY/i7J4Zv5zqybbkFSwFMNxD7D1chn89dLk3zn6+
75bxDUkx5szDLkZFBfsSy7dWmpT1oapnk7ueVoltODyUUm4ONELbSUXxili1w3eesbfVX+8evBec
PIcyx/DewaQgaq4RgryRhcgpE8lZ/ZAEJN9GBBkMCwC18CLlCPbza20AhHjpHztLg0BY3f0I4xBK
Sylgsf4rHPnfBDesG0AppAfFXato1SwTQJyjNtZ9HphK3RykkYQur5r5UNA67Ytcd1HG2V6jpmGs
seQsyIFMurttMQ/2A0yTQ3f0R+suBXlvuP2uUaNNa6VtXB5um/4RHmqM+Ghd/W7LfB02mhipL9NF
pRpmqrvu2UgqSgtymgIN2xvVAultB6rvCq0UVnjWICaJogguZGtLk7zkYRuRAaR6/NBIyd06xF81
79SSrJgjf2G577dTgnhsTiCTlLaHtJ8LUrxbPFM9AaBIj9f+DKe9TeE3CEePwGOmPAD9oUh8FYEN
bGVHDdyj73pEvB9bkDCMQgfo1hPSMfyv6jKww0MOYFwFuRFiKOeHkIU54BOcI6BJG0+bQt3tEdL+
m8G2ii7rFdpyVDC2WNXnt0d9lxz4RqknzCkjo9YmpvaN5sV89mBCuzEoIgNNcJZqkibkqnBSeZpg
mDK19Dt87jTw1kQIiil1GDEsp6aW8tWBOHGAypCR9/yPPEYy5jEC9KivB4Hxb9u4ObnHhY3twzlM
phXnrhT/eR/oQQmYlk2EO0x3a6GO0rSSRVMZ/Xj3tu9yDeUa9qYDv+eC2miRBFM5x+3MnBeKUVW6
1myvDU9b7BfI8bCVHRP9FDv6WSf31nY4cbdPM2CNb9yxj87DfZ1ODY61TRb5r3SdrXAyMyW7AgtK
FZW65BvQOb0m3CoEmKUmduZxcNbGZSMrma+zjR9FiKP6NK7itUZJINIVJH6yD+RRYOIuqpylhqsM
1s4QYGE/bUBH/lfvu79a/FHjv5fFe/ae4Kzo85Uu8HLV9N2ctLsJNr0QMF6LpWf2zpQSUVxmZZZm
oxdmSP5zhEZe4U0PvTaEhALQwwZOI0EwNZR8Nu8bvMChRI87zv03Ky8JqHH6xigJIu2uOnE+7W2A
kue777iHuwk8n6nSDM2ymaT+DKXKV/iPoTiOLBxEVM7AkiGur/u+PsW/yzxDfU3GTEtqNAFC4R4Z
0WRzlNUM5VzKmRJ9U1LwBztAE+lxqd5KuJ/wkaMdoH9J5QvunbGQDQivlLMbBHW5gqc6kwVNpX4R
IGWuNV2jI085fe0kmhJBlAlyUKXwCEIk5VakmwGffHqyTbqWVdt9qMfBs1BSOf09MhK6+6+z7PF0
Vp6k5ucc1XwdhOYMKyXgSRXaZQxy865w2w3JrflgdAXcYOgYir1SqjuI9sfxrDp3oq8l1gD2wKhr
hGcyg/L9YCSxPUPnkosSr+oz+qx7PzOd3VoKmkskdgsUTGPdd6g5VqtJnDEyKLwnho7sEFZq392R
Uh86AwiVj4timdP2mHy0QnfcEXveVRibeZ1WPRPTorhfa+TCVjDUIl/UzaFd0poXW8I0OXGo5K4S
SsCy0tIJVzVSyK4r0sXFo4VJMFff0Yhjv/0sx+JcOKtrfja+9MEEV9blmITuTO1ZKZLSfzp3b9ft
4gX+jWFGi+HoKGGR8cXzfUTBYRvP9WYqTjFUeanODwkUGA4YynECS8h2m4H+sD0oYTweEtPhQmdk
aafiwN0vekCH6bQcipmRuGZTWyL/pMhc+Xs2sap/RwLWerQeMjZBs+dewSP7YR12OHa6IF1CDo3P
zEdwH+w3g8de2gMblNVs4HVR4nQFll2mmps2b6hT0Xx3/vg+hg73nNKp6fty4FC4QV80Un6c5mmV
oc9J8bw2/OmJMPXl9VS6WaYvbQW6OnDd07ujuxDPygqwkY4d9cuYgYEMDB3bJiZw/yOQyGgVylPG
f9c75lPBCzBUlCXzJIXfeiJ/ZIq/rW/1lkigU8UUEnFqmZoUMtXxSwC+Roz1sLhin25y3UH6grRT
B+rojgWeEJ5vQ7Lb2BB1EQuTgM5+o5Wxs8b0IBg5EM8O87e4I/9ANKRiAqD5QpPE1yvYLJQly8TJ
zxYGHgtFCxTA3VuxnFK3FqlLr81uFHC+oLBP3mLNYE0cFcPTFc/snxhxHnUceOosIWocIJUrALKz
uU693IUULOgbxEWuwuy8S6gwFQGuqGg/79WPv2Ef4FGZ4zdmCiCPb9FWK5SdCBXr4yBzXZ3OSGnV
1zoSz/jOUzeA9TTDuGjLcHbani82+JXTCY/uQVKW1TVgxvyL4YdnOWB1ZXN45IzcM+d4TqKx9Ftj
Qbk8a3aJpY3XTosgmx6C35qDbhpntOCZal5zE9qaK9WCg6UFL6a+OXGr9BHHaOlixzIQ+4rFMRLZ
e1fhlmI50hx7F0IaANkgHqzIh98QyFz9f9L7xsn7veIxby9k7iDXZ7wWRJRAasDK0YDquEOgltG7
SKIsC1dU04TZFggG1zTQuz1P3/t29sp72VOzpj7ibvue4nt5j2QLlmF486sEce29T5FlUexhde3i
nN7MpCh9//Q5HJrnZAg3tG5qlyRbcvYVL01i5yLgkAq0mjdHqiPHMIPot4bsjmFCKkD5x/O7ZbbH
jbrL+vS3GWGfhL1mKdlDgh6aoeA6IHyk7bAaqHP+jM6Zi1RwIWDi+sMZlelcIrlAQzmTelWhsxRr
U4U7w9uAxbirYqfvBw3Kjzp3iuwiu3i5D9MXUeZhdhUs1SIqpkk1gUThxD8+pH89NGJrcUvSP54l
0keC3FACq3ZuULqnpY+Fewo/LlMQZW7VxTtT1nv9tFgkWM5fLlkiEXrwG3lhqez1eLIp9C3XTIi2
O++ANrF5rDHkFoAHMsUqSuviT+0Y61yLVDb5UnojQRVzQ7XV5PlOIlVpDPaCIy9+gfcZ5YBDpNax
+32J9GPfS/3ST/FPKPxHlV5acH6oTWaIJcKG0q3rDhzMB7bCnMAtiiMk279W7AL0GFrhONqgiRib
MR9nSaGUMMh+aDDGYvWokvMQMiaCnqKwHKDw3mWsh8KJqem5vRN2P8ltnWtLp1juk+L7Htd/hTze
OCcPf9ZaOcqIw/zaw54rBdEeaFF8LNwu2R6qMwBFHmAF3KgszE71mg5esdAOJAyiLyivvZSMaitx
xFskOg9iCz2+lkvUDtpI+DGYiYJs7MesnVGKnDNakkcodihL4twtXKe3iw/dBZwCEZyKbr1mZu0g
ihGzQShYBHfUdHudDlzDNKDECXKoDMjaZk2ljA77cfoVEEM+5SGoacXwY08ENJc9D+SOCdxOGC5D
UJl3Bbys3XsI1mf9NII6pS1n6wiB6rv6kg/U0TEWx09e5Y9cdPh56eGmrDlfRAw7UxQad9ATZ923
FDz088165hw6isL+p3ZgrKU0N0MXUWrrVMcJHQtBD1qm05dPayusZ4CxT94WmDnwmdaPoG75BYT3
w7THQRweAepx/M4u3tBq9+AvcwZAig3+K7bQd8pEG9y+1bDZ5TNOBK6PgEsOoWjRtJNKVsBHT0ME
MHJCKHQDomAB1aCxLf1bhwGfEM1S6xJJE6z7yy2VV25te2b2/3blYOKxT4Drwkz3q7/NhaQh6EyK
m9PY8jbbW9m+Z2MBR2UJxiS1oJ89cGC+elGy6aMCvQLWjVlyb7aCWyzPBIAiXEzqUIMUkKyHnvqT
8bzzp4LIIhmV1WqsT1sWE/AAJ9SE6fUkajbUdDiL4skyxypQ9swylVmArS6ndjRXjWYCJjNrpxEJ
LbSezGgahfFrEmxl1TEy5xeqPWWh/6GdU/03xeJGcoA/b6D3WzRlylMrTXSF1VYLzyWmxkEvasNH
RKrQOUFEkOn5cbiqrUPlgUVzYZVzXtdHjO4pJVMInyajklPmLuToepIeGUcHNRaRBWpQiRQw2TLU
ZtQBSgNmNsFaD+KjyK6fDMYYyy7itCfWWnRWkou8t8Hb3uqsNpXOqXve7HMTXAcicoOlbIyqcoPa
mbSpVIgS9cffG+brVXt7p9SF8NSibYZJbCG0dL/qbAYkO+sKJhrHHnQY6NAHP/4CR3NYnx3MB2Rr
6vFZo4iWjw5wps8lRJ/GBaSByb+C6ExBUX8EDtefjIlXYj87aOnkreW797QHBcOnEPjXawUeOBVO
4N8o5UxJLkLCcpuTL5BB9/2W4+D460G1ioECGWwILvrqgdRp/C1QigMFUEHgzYRcvcVceRPczJTg
rC+Yn/0v+vZyFZkKuoIcVJR8nsWHAqEZ81OKR58Vki1y82Jfr4kORKtlQxsdSCPIz1bp/D5fciyy
nxM81ZbIZaoISYYyGAzToK01sE0iushQBE82CLEZsaTOTQeE4WwZgWASaaB5521P+ElGK22AAZZk
xQvfCr7a33K7D3jWXDGw4+xdLePC4b8nAlliElNFV5RiMfksvzYP8+yCSkCsmcpNhhx+v1mjW9Hk
HUYn6cLmyXNWdlAoSAcHXF95ijEQX04ewKJepNZBrlTP9T3AXdkSKosKhX3oT/GXhQI0X3tNn2gL
zeNOtMP5ANLESSzuypbfQ+mLM0JUhBX/meHv2yArQGY6vxMuMLhlAks023nRjhv2VZVybUnLEWSu
hiPfrwN304io7IGA2a2Ly2zejDIFrFKC6yG7gXO4fTg54Werwx/OtvZ2HItWUReaxuYUvwSQrD09
Fckg0JICNAEBuBabXVk4aPZz8zWZhLM9EdoFTwAMNR3oy6eV0YSGiuahmjIXvhQ4uYiWKC0Xq4E6
34HfDAdp8pDc9nUPgdXOvh7VmXeT4gdclEJhNVcQ9GDeO3hNqOK0On8NWEAKDhR6ZktnTQARkLuu
2AfYSyXFMtx/O7A3yuOVBAbjovghzC3LocR/WWLru25iSU8xjguzhmlvL3QNrixUsAt0HQL1dOce
C97hAJ1qfiHp3cwKjqzWiz1k+lwZjET6UvYllgC0lB8yPaL4WA839l3LcoN2wDxfbOAhruBX6AZN
nUznHXBXuoVEVKr3ALrkQSqJBn3bxYIjrIg9iD8EGr+A26EAVV76ISUJS4DiUTk0aBkMWIZr9WuC
7CwezjXWBY27Yu8ClRpvil8f2wEYOvHwUFpxOsQSbyY4xINl/anxNbbaGLi762epjkm6vFpvhLdb
lBxZ02mdLnzGCeoPYcIZX69LJHfIo1oaJ2joZUtZXtzGorn1+knmyPAG3i8GnGUCLycGKL9FQvv6
yOXJSzVxLahM+H93fnLqthSo5kRunPgMyHgyvWRNr8qTNwM8ctN0dOZ3BtIYRtqLHnYlXTQTyRX/
4YN+wf9Wn99lWADSGnb8kmJGOUFX7hazz2yyOtWO0nVYhxsxZIzGKyQDJ2apl2vs03mrcTRucIW5
N73P3ORDJK6aRnta0LJUZ3wFbII1b7IRyPMPWpVmftchAQjoU1pvpk82wcMrYzH7b7XtMVBpQPxb
uBf9iRKSePBFqkYeveftdvKIuqM+XdhbhQ937PXanM3Pl1t1rT11PJOy4VvkR+JWk9VM7qImzGQl
TEtpcpTFGIWqYttZ1yZGqg8lrD5PHFRemYzuqkLn5ghcqJeMhWQjdO8m+4EUzfG9hjRqQD5eVIPU
cZsMAPMzqOS0LsJVTNc9Ud9Y3OZ5kSuXkXTUbtc+GsNE5/CtMmjw4Hk0QrwHOGRrBNXyGbFvAXgI
6mlemkGYWpCIo5BmcbpQKa2jvaDLPNXSAY9wJo8toJ7LWm/ur6NcSFk2bf5STYVt79/1JZu793qi
tc4BWzMxILTm9U35kVQIzk7gFpNYSZLo87sIhMjV4V4Al2+LR295Rs1lTTl1n7/07BDpLcNByN0L
h0+nSAuSjvi2qh8zOTWQIajjh2EKfuLko3xhEwxz36Xr3Ljx1MX/YgkeogIgdAvzGcneRzzXOVqY
sjVU6bMl+dV6pC7CS/QKzwuyfxjc16CSP9eB5dP89YVo4KbFzyZpRdJi9FghcWeYaxHkj1Z67ZPt
BAdXkkkEj+G7wRLywBSctjA5rkQb4FfeWcQ/L12g2yB+bab2S9s/YtmlHFd9AOaZOrHwyW955wYa
JoJ+EzuPLGn3ka6vhFlN1d+TOhqD/H42NMzczuDMGIsSkTKwMIqFamfCunKN5cXqV3OupPvuAago
II6SQA/zy5hl+x+YP6bXRK1/kb4KWAwd0sPaMbI7akVBUZgMt5ZbT43bINKkmizPPfLGudIpOXho
i5jzwg2fs+7xgq8FmHQmx0gbezn7FnphkrTfvYva3K494cv9xk0k8gUJGr2SAIBfp790XQI9kKXD
OxQgOi/y8Hd2gn5wQBx1+KEJp9O13y9uKkYVB8AyElwTGEfX2bFmlRM5LRlPxAko4jSQJLpeHPd7
FfuKjMwQIivAZQqkG8poeC2m+dJNYpfrV3qI/HrHMvv6NvlcjxVTr6ZmiQNE453pBf8DQvMdUn/g
mhg6RBi8n0ssPafQyRbntj7qajWdcHdwCatxK0rqmMXsOdTGuCu+AG+8gFUe7OLBXTBn5oEsNVE6
uGSL9ND+PNoeFCozDjZTax5SkZ+D0tCnTc7MxKJRaVJve0YWdBWnsaybmxDYNBXdBQ0fvJjrfYIe
lo3wYew/iYSGlxWMIqqQXNqIOdWFTmDR5FsOpNVtRgcAsxG+OrMX5pQgC9poubzg/vkJe2IHvDzg
LP+74h28PWEwIa/8ci+K05KfIZ3FGgerP3lTTfMA5th6ugBkazly2CiSRbHtgzkx1x8qvTwxY3XN
rXNa90blXPqPJeyCQtJr/Z4zuDd30nXEShS5eaximVMJ4Sil/7UbCi6M5o6cnai3yRBf/j1u5Ojq
VVyoT/ZcyHlCV4rrbQ6qyZruGQ68i3OlfAmVvQofiX+q6gt+UBK849jevYjpz8s9V1Rq3xAdjnFT
5g8tKCCekVZtJrie763mI7UN3QLKs7QNBTt3+IKRX+8/xEKArzQ/s4D4qWM3JgVoeahslwllQGFn
EbW02QVAVoqWhVu0emg9K3Kpw4grP0Zrt/P8bL31UTRM7rnoOuK0x/QT+X0wng2jGdC6PFkbpLkL
DjxgMSRVwe90rsU3hGnaLLRNdmfP7Rwogv8VLewI9qMHHnxCylmNIMQF8YK2tOTC8MbeqGIZcjol
6/nDudKJUIVp4ogpLq2InXkIpeqC13cuzXMA2v8sGRTNjnhw0i3b7ZEswr7MI9Gc+OcirZ/7qI0q
fOtZnyYyKDP5wbzJMipCVQc6eS6YyjQ0tRTXLcSAFBQWm+wO3OIxgCdlvvrIwiZu3MxCk8dJ0jqV
qGsrKR5CAREjftzMHzTDg7wcvgViqVcHT7wSEyLTfv+F9pMEpwNJ9aejIYXkO0Gj/9ovRRM60A5c
czL3QL7VUHjYtsqJBj96O7lm4kICo0C7a9w5eGOKr8wLm0ad2/tD3/S24CPyEEx++zBKktcBS+h0
XJd+s3bY2WyCcIEB4TTmFZg4wTYp09NHT1wPRkfC8ZwQsjK1/jgxe0qg/6VWfSD77gk9oXAyJRnG
ZwlFLtVq1N7g1XnItpDcBajGcn+LiwErApu2GSTy48oUNeYDi0l8DZsn0x4ZvBep+tzv5jmJ12tC
zPdE+HlsXosKO2IkGY7dBzPxq4MQsD/C7cpBZbYoAEGJy3syTWJBNJ+UElE/mB7WsRGxCfCD3cg0
bkjgXGM4Fn/hQ/nBZMJPpdNMBwHor7xpSG5Cb+rBCxZRidZoGCjstQCp7P7qGw3qV+/kvIVhsSep
mjwPvTvi71R0ANs03yU6m/MqYAmysu3RkzQRSVbIck3J7sYtrNA9xxfjk5ccoi/pH+Xghg58FSc0
C0i8Wy/LIJwSubyIsa2yBSsGbpakygzIIQbdUh9GM+g1D9863Lltcg9dMtl238XP2tqUucxMEyM8
S1xp7qoKzHg3EPxhaSt141UeU/Gm1Zv35qeI02zrxVCiL04ylrEK0qLe6dBMjw+Gwbz+OI3NnTmw
s2qrt25ZbKjCPSg/1ofemyCcLEWZ0/5xZElIHghZxSIfmIlzbBCU6DuhcF7ggqzPOeg0FY7s01lY
+cqVCkp9I+UhOpwUzLntB4mTUlIOCckUfzXGmh2w5YrFhOAdO9poZ28t55R5IvNJrUcIOqC3woGo
GVmBicOMGV6TwEIfAAa76lBqnI75KuUNGmoSuDOkK95slHQs+wrk0cX9NsQ2PHWYnLMC+0TP6rvw
HWxj/u+DEphONPgoyY4Msb4bLZH4rkjVYzeFf7EBnTFqC1fvmXSO4fOdD2za0IS2sDip0qqEnaNn
DAN2WeLXYK0ICP0zp4pLkVMpfK9Fw8FRNLWQjJldaHA0Jn0nQvOC/yuKl/+X7oQG4SeZLm0s/VRZ
NiF1jWnWtMR1zJ0huxPM5NMHjLitpf4cEJAVA/S4u+z36hd+6kVaC585HUlUDbTTwzAn2S+9Pk7/
neE6cjDC7eBWqtNf8W4LPvaUYvs20dQux2/UqLkSZoACClY2AQ4Mmn4ToGi/yUHPJ74TrUOE0PSx
eCHlE6YxwdkHYKY8KREOyVTtE4x3y974Ne+6eugsbqnnjybMyIPgP0Ixcjcq+lmX4AzEEb7rlPEk
wJRZeF7z/Dq5UnRX1gQfJSYEr8tMy3dQxbwtvljh+kPS1Gzsu7CbUrf2wNcvm0s20KaQVRQNYc8U
L8D0z6ZMigiklCZRgiBWb1QSq8OgR2qznJMkONr6hbXMa0J5IywlpOhkXr2f1F97pBF/qaCG+yvs
PwaKSA8SNT33bJoO2zp8ObsuTmFEsG5OREnaa7ZxoF8nPUzeQ3ZUDhFjiSV8W9UukL/vewzuYRNY
dRCNENRbnH1dWM5dUGr/1dL1lIz0Lodtkvqo9o+rhI+6qxel4a2o51RcdK8VNrPz61hiNfBCdCKR
Zh2XRu5yNakmXVO026zTLlnt8Kuti04ozCyar1XJ1Ra1xuGbT1lGHys7Sfc8iUBR56ttFBcIwgmS
vdkgG+RbI9NWIADwAmnRE2PNCJd7+muASl7oDz+9yQNI8Z6Pc47tZk4SMg+w0XZMlcVOXhMuSZXh
QLQqfTSTW5erOC7yjimTXwZDCnhwyctuBmfDB/WZ6slG1dUSny+0rRIS6OVBRDDGPyVDLbarhq5N
B7fmtc4TgkG9pnGen8aPdzzeESPaH//emd3HkW6mU24z7JSMy0xHhUFm/z/payaMjsd+rJ6+HPx0
jxSSfKHINbXxFpB0fAbno/M+eQLcWj31kdOJQZQ4AxkAXxe+Om6WZWpcbwIUBzNfY3f4cTGXZYk1
pRT2z7dyzOwrHxc/CsLzBjL2V+BrjIoFBiTFwLNJzU2MPpPiRYmFDXZ9px5NydBBwjM98XNmEiYO
OkxztrMRMlL5DMK/DfQhql9+bHxzyWmZX0qNU1nnTkTj6FpA6nYlPZ8tTdGss+/ltKGDOMcB9wgi
0NXFMqqA+xJw53IGMoPiOSTbEdDevmGFaANvUxggQo0NiYXAXr1hrfg3sMw3a7DWf9DMxI/UINxs
VFxk6QrBkYXwMdEhJ8hbYWOGA213Gm/77DHYNAWjXHriywEgfgWyfjf3I5JEl44EzLONBNQ2G30B
Fi79SeaTKhHe2SvtaUdC8sLCZcY6dwRcY0bNDPf6587nY+39kCf4j0rkCzGyuar4giRNMNTcCzhI
M6KMgZ4wlEPd3xwois/TFAiTlNcCacIFF8GKoYVi2U6lmDeAP0CeJxEbOdVk0m4DhLiKBUH2tw2G
74f9MIJJMKWlSB6N78ePXTjU0zVCl5ab4KSdjA2y4/2uZWlcVpkcclqieVcu02mpdzRsvD1W9iuo
PEM+lASpUdqK1iv4vsi/5kvwq1ayoVblNonjKF2HHTukYtH31jMVD5AdvT2gmojzu/vuUCv4QYmP
83SZxGIFDC4lSKDfZepNboewt6LzDSwuNXGUEdnUDtdLCQnWCJr6MjTTCv1ovraf7s5R2XjtrJqx
GwiA3Zb6JN+dX3kQeVysMAF/e01bRSDSxFfA3l170590b2bA1UL3pgs65VnYEoHCFsQwIL0MnhL2
oZLbnTVR7OvJn4XokIkMpadYwbyiELZF4bI2QqpJ3RB7vz/luVRmZjpaKNVde0chgWbLtk80534t
OJI+qCP9U5W6xu1ZPh0hc0d89oSvEkCbq1e2fjv4aJep3JlOlndwXLlZE2WjhP4QfhGNusTWIFIT
IU4ysngOayh9znH7beB5qBESgr/wWVh6lO4uquW3iJ/CDr1ufZvoLgoLEiWNJ9v5ZWfJfm2UxBGo
V2UxqxZ9hNCiI1l0v/Es7hRU/8pW+bKnXVXkB4OHiSI29r4lUuh3dxwcOvLujoVVr2N1uXRAho8A
cakUxM6QHMXB0oy7jotPdHFpmB9bOAPtdvQLaILcrjM7+YVMBekX0vfxxFRJMDsmS06xwdieePrC
puCo9b4XCiDDlKAArv/xNZ6jsd9UdFrDaFmMqhTZIuRI8KfSEX/Je4xoK7faDBYhb5rr1JPtrDX7
X5T0RsnWSug9fJot8of0VRIk164zQV2Unyjn6kMGf4Kl2z3yiNOaOgHeV6x7j2qH7Q/ho5ZVJv5v
3qC4/z2sbmCCWkGSH5zkiJJD6MertV3eJFWzoLzo9woyKjkneCV80v6BxB2P8I8slQBqDP0eCGWX
GJJXSWhBVLmBpuE0vgzkQFUE4p2w/duknk6XnxS9vzaVYToFDlfoKWlvtl5pXL5Mu8MRC+t0TkDd
ais4Gk6x3VXYXLrFm7YwWIHUWI4j8Rxr2mb9sAyJhsVoqhCXoluykuVgIYUt0x82qPK1odADZSa8
tmi9D80Hz1Vk83lLv6MXW0KlC2bTFPiyxl4GZEoUNnRWJDJaZzYgot9k+yrzzZIY23cOe68ErpuI
T5nA5eqtHF0NzYPfi7ekf6KlN02OwDpe9+wdEGEao7H7np5DTpBhWkLm6Zb6hVLBFbHnhZLwGmhh
TpBVF9rx98gsWHL8ETDFnp7rNj4W1hejtD7F8M7DmbP+A4Sj+rAyMQ/JkqHTGAaeu9kiqxvUbWSf
UbMC6fa0+vGfBAg943/UrxTVFODgWt5jJNrvOi36w2EwKMlvFlgfM0f4fBKaVhd2+39mrJvUEK1y
Ik9XiuXJI3Sz4E65JXc7w7xp30SqAyZ+rtf30iWMtVNHof/O2ou7duM+UVph0cQ/Qsl+XnyBbPHS
IaoUtQJd313fie8KHLWcsQFNuPwJ9CDGHPZJtc08aBPFWl8iwBlZQOxRk3VptnDCzWtbyaE3flFn
7s95fBeuF1/yNFsFzdkMzc3pQplXJaH/9Kl/sy/nBABhpAjLiRU0ixlvpQfl2O11NyK/IAdE3cLT
DS4r0KGt+Oyx7E70Kr92gyTz97CBKUSt/ErL7wQ9ZUQQKzv7TvzGTWNQtctGwiMlOaibzCSvgEXx
rMZliN7gKWxI4ieeZ7UWdCJflag3SBefz+HJjhLjDixA2GiK8Ciy0rPWq9Q594YQ9Or1slMkbwjj
nB/VAsEmXh0+ewTeP10Ao30QuiyU+juS5LOMW48zngRLihk+uMhvYX9bhBBzw0Rk7X+2F9d4BMKc
SQIppQsCl5CQRwqGw9JFf+j/+X2tbNbi6IRFlE8miN/G1N3mt8bWv1GZpZ+pPNMZzY6oB0ovb1NZ
ovcMIJrvX3UYROfuZO2vU7G9NdaFixAhXreEvt4RRSDGSdAXzSX7nVsk1LFSNaEx+5bRnjaa4mg/
n0T9zIki/FQEq9lc/WODSeUgmxAKLTRdl6TziMW047GMaX/VECBaUGen0wQS4/ldFNw9164NEt1d
QkxfvVRgnns3r4Ky4SbbS2Efdi27g6EkbJEiA8iHFKyjEDbSkX+FVZzKt+7LcxNxoy1XH4xObNc4
krVmFsUGcfnJotwPyCJdTzfZEEiXTyHTBacZy0A2CdoB0e7382P2qAW6uASjFf1Tq5UjoCEKKD1y
JB8wBz0+oaiUXKqt2ql2UNd3tT5hpl6CpL8fxKTg2j8ICik1b5IMlbTzvPtgKPzeMM9JM6nQgscz
uxwMOwDs4BD/m/yL6RLdnwzM0eNRW/iYRr2uKFZgcJYz3copu8aQ5aVh8arAoKQDUBqTjDAvoQK5
49o23U5XWDIGwQ96K21fWu8X2Z1aT+r45ooTsd+MOGkoGgIthDsbQS1NFJRdxGhcKo7NEB2cEyh6
HSv3bG+h7LrcnY20sDqAOY/SOShiEGZsQSIpIPqvTgQQRhPKysjO3/xaqXcxHTKzfXUg6nItTa14
QvifMOfhclb/HqLaO4tkwiee/q7iTeMf9aCCfHNCHi5OY9Pci/HRw0Pz/V1duHJdOrQUcvDW28J1
JGxJGF11gOKdW/ExihUeIyVPvwODl7LP67r7JfEccfasu9FCgenfNvyeHl4Yrr772eyzEDE4c/QE
9NFQEtZ/blytQpQw49E9UIcO+AUW7heODDIEy9ZqFOfmC5l9CRhqdJLv4/PACv8dg9vAFyWeSZOg
3dRv8qU4ochFVAvpxktzk2CvRQcziGTzUjd0lQzifl+aWEeTfnFHwjIaiFeAAzHngmzVYBrETOl8
90wepBpsC1QZ0m0qg42kvWP/Xy6PsBesfzqo+OLSi4UDGXQ9rzAK0Av9njD5LxIKgIjyREkwfmZ7
iaIycHZme4aFBjxwxnUyTsoFuCoW1dzGchQVop9zdc5PlUUxr7MKbbJ+F0r6gQha39YR57sgQLTC
HY2DJQsKRxtKncxL3+gqHslLG/Zxg+hRMyUqiZC2uPOy36yzOU2y6GmgqHPG+XVadhMNTkc9f91b
sI6Ua/SG8NKmtbuKGHroFwmRXpF0K9ClVGuw45oRXgVVBo/7BVIO4t3VjBkdZgyWTeRSrnDCPy57
PAT1i4X9Allwyv3nRO4SrUo04YJ0xmlRXKJUsQqOo4PV+O5ebD7Lw3m8haKD/rnqsaJ9egxWCM8D
e5W+zkMSGpNDSHG5qVBn/oqkm6HXKpebfS2adPP2dDFJ7k6VBTuoHu+J8QRfy0Nk0/nlgiKuWBJ1
jagtfod2JNvLlvO/+8JfDiE3BsZ1szIpftSdYHK9zXlAgy/Sry/SmzUHMIhGIeDHXRiRN2vctMLG
vUOooFbxxTASj7p6WP/jFzY8jJg+3FFbig47XxpmomnbSzo0dEaEMw5BnYwsl7lRhYyRm98e4wpq
GG9uV1AFBHk2kVeLAF7ubkQKLk3PINcHgkvnP4TNbw2CZof+XNmAlrTmdvRLWYMPInmkj10PAe/V
G8JFZ81zH1sJhR6r0uoRE0uyKSwb18b2z/uYb5Np1WRZeZ5iYikwTKZkNU8KrqQ1kBZZmrnLUUku
WWLp7y9PM0/afCzo8c1Vo+sHlaa7IuN73mI1vnlewWiKQGKPc+tcU0gchlxpVOFGgs+DRVVHUvFG
PVgAp266gzdcLmQB7mGRzQFgurOgHbVx0hLQOQaeRWhWLkgh0yqKEl1SzHpph6EC8sVTT84t4/l7
ygBr5jAAsVOKe9K0r0Pb5purPzJMLctxT833MXWKikKGcVrU+3GIXFU4C1HUdcQxC0C998qltNsC
5iS8fqFK4FHSPtZCdJ38Pdv/7RihZKP4nYnc7jzq/4I5SeguoPSsseCrsbvkmW0k8Ca3OPllLUTc
hMNPEbftFNEtzFTcymVYeBhwqkMKcB6rOl9ENMMTxdJZ+Z3U8x15s1WxA5XUhtS/ytCMukt2AYjh
B2oNai9e0KLMlwaQqwNcj5bELDC6oBDH26lqjMaDqSxkIpwAn7dQWYcDzn2YwKuqChBaB89SLeYx
hT/L+u+Ye9TNuQs8aWd+qQhMY63yPKyMM1I2odgiOBmP1wKs9XCW1IN2batGzqG88sYVSPdrXD/Y
NRZaaBD4OG7FriZ/RtyAkkkylRzA7Wp0YxEXiJxV6vLLOB8uS79Q9AeCygbq8B+u1Vl3wYOXGh62
AfkthtZX7+3Pufx71fe/npHKOq2vb3NL1681sZSviAIUGtjbVsqENMZgFTw3s7mJl+aupnkwr9++
zFNLr1iuFxolbxHNApaKqMLvr5ZXZM6b1tyWEgBsYiQomMuVacpLqSrr7uuy52RNycxY/OW4CMVP
9ISntPsF0MYFYkALJrVQX3myXI7N1Qz0ofMHDWkZ2PRT+xRnpWFw0ly4xOleJNhquUXj/PcWgolP
G2LUngxTYq0wDyZgOlbEewLtTdXwQoaXNxsSgIlGgt2y8SkVlqyF5Ihffsmk+uJvYetAPj4vfP6e
9I/pBccWgfvL8ihlUXEc0FgVLcVMhoOsiHb4zG/z6RCNl2TLV29C6CA+Klj8AR/tObAfilgKGT+I
7hgGxLbqDp7LssVuENu5AP9+msoVMKQJ+hyOhpiv2NFptXBqONJeYTTJiGndELSy4k9fr5mX1tx8
H8XQNTEZejFK2DIXxfKx5vMKc+YxAoWRV0h312VnhMHau//kqZ8gRWlzvt8sq6nAZpNu3+sihwZY
nhcovF0lvvKIJDHALTIR++gvdV9c0cktua4PreOAq+bgXbcd/IlRB0fmP0QWRVcEGqCPa12luN6u
Hnf30aRyvdz9DGmW45riHWIcxl9J1cMKASri3R/7H4bmU7fxirJQMxiLzIhNbpGCmrtADZQ/FHuG
wrRd/Mg/+ItmQrwY491jJozeMfbC4vglWBfHcDbykcPX9XF4mJE9t8vubwrEg/QM9vEWnbKQea5Y
m1AR/UuOJjy2DpXqSbonVBBFMIIwmO5DROa/ATjwH8u9lquEWzCLt6jFBVySHpDFFthQMla7xgZG
uQ7MaeTjqkxXVS1HjcMKRtdZ+Grac8dVV+hGJ7EbT6XOFTGhUPHvM0K72pCa1T8zqArEnkqxRIkx
81rtFThd/3f9xPeIsSvvBz4/WgY8gza0G4Dmws1Bko52rSQz875beJMoAyGgVYiOxnrTeTTdz91x
fvkQVTMTXh8Koi2oXbDGvq+V3N+HAupc5tQJDs9IxPqqew5OWTIILjcDhab5Ui08pNmn/bljyFmf
ZM3lhlMxUBsyHP5YEZJ5XZjLSNl5978+YP4L1X5NK53uy6QI2PB58XE6s4V9Yq4Het37R1PWsFPs
fPitTOgPgYrVPID2ZZhLjFDoTtFLN9DYmaC1YFFF61/e9HeQdx7InXR4tG1oH0cGrs1NnonI7xDs
mjDjwOHpmzDLJHR+K+hTuWTnWEvsDjg+k75aHR/AG3nTHIEQnlE5gCBQlLx+o/FDp4DwtTA0SgRI
H8m8S3hMhT532+MtILOTWYTKFimSlJjTE7oGrV4Eozf7yiEsTDH3umrqZsGUPC58BgAxzvaQDblm
kXSJBi+WicOevfhr1OG/SCihDcI+XGJfRFaDMU+5G6mwza6KVXOGsGSsQWlN7JIrsdt3sbuLelyw
c9Wlej689gxARLeRHCR4nlJj4OAE+Fr5iFF/I209EyWDZIvDIWhRvQFZeWACtAzKIWAFuXAY1zJ3
E/PoPlUnTmFlk4LvVhPtewvAUoQU+cRhx90tPe4WhMcMXe8UzFxHcFHrGKkFDJ36RFHp0m2gIDoT
lOCzB2KxqFvdOv9T1aDxoBUEQpoLhy/QyCtjn84Bmp18DRcFFGP7DBR1SQxfgVxRAxcUpsk7vEah
e9d8EAMClmluDa3WNxcAvPYLkkybkJvBdMaDVBAXtYCZVleohutWcA/HzSpcUTF0qoUBm+JgpI9Y
fpAbq2qYuFMre7Wx1mdpomvZp1e2FbT2erXPFRp4V4L8pHtq1D15B1ZRx1VbeC6cB//f0ClT/cPo
6qhOLt5V6QVmyMdkktRIH5O9F38Aetmxeie6LAHacXm408k0xvhNH7UfHhbgzfuy4R1NVOart76f
7RalS9Nq3FOYrtF35XCSZugnAQqEVHs1oubvn2dOn/KVdurz3GLqVx6XNeM1uxA+92t3ABnKYwdb
qnAe0tLSmbKP7gE+y/C9kbLYuk8CGg4wU+UmuNhoisyl2+cLs9mgFzV+LYuho8iAGZ3ms7Wptcst
q/Jle2tWPPkZ1udnU2UIEMfFkxEFYKrqaTssq+l4N5vM4mUwF6CsyhoCUhB/DbfRlfq8uXqMtekV
cRu4fErYU8Mphob6IfJPwjZq2AJWMDU8jChfFMrmFE8OAZs0u/1KeII2nzDyVScHWX2z8kOUQsZs
0VxRNpKR3KINTFJ1JMyjLFY9GS9x8C1DSHcStLszkIYEtkM/YLMainbJqinzfP4QRStgHEZRGD1Z
Zv5LNnE+vHLPr3LOTMEtB240zN59NoCwLD0Skb9vAhK54R8vs5cHE7GfULZzMt6n+k6bnX2P6ZOs
5LWBpRXyh9QVnHxu17XYs8jsD+G2Fd9gONBt4EBn8Q/guSBWKb3XMUGbPaXEBbGPX3zcnQMmwuGg
RFeLIoqHy9H81y5LyrOFTXQanZ1CSPLkcmdszQfugj07bWPrIe1M0frGvQsCLbZGNxa0YSmCN2RO
Epfqk1r0h/iwP3dHxipG/IcKOJYjoYz/FuEQUE2rRmDrPnLrmPvSTT85c8oH06I2DZ5kw4SaB4S8
nMG4yILGR4dV2vDNckD/e+M2kuy8mxEgDdB2wEhBc/ju/sxyCJbdiGy9b2M49KBnzTpWv6YFkCga
VUzz4ACCfoqR54ujyxjwpWLO2FYrb51eK5Te2EzM7gb6Y0KpusM7T/p1Pe1LG+VKnIS5utGGDyEP
a1KJN5a1em5E487ZM7ZguJ1ErCtxFFdZiZAhXh6w8qoYtEqE0/PtlZDMxMWgwDTrpzgSqkaIufsb
XlYd04zTCWZbLfqtCfHnqOp8ZpRcGDJgbTuQ9OdKUHMqTqkC7HC7nwAoOhybFZTxisGQgCWBprer
PpHSPlXxoCKiX/wF70SkuvJF9sw3BzD5RstzI240XNO4uTQfqQVtrX53sFjCe8amCV3Jl66F6JPG
GhHT/fjaDHqLGal6+UU2f2KrpqDsq3U6BkIct8Dbh7VANthvYvFRzBXf4nEZtMG26qdvyqomi4IP
1YWH5s8Mft66CQk0Pd4os9qspDxtP7bI2fydYKujMJZ32tE2eAOXjFdTNn3YTC7Rysn7w8xKPFYo
E92sFIXsqe4suQG1pVgT7QW/eQSLXjqX+vK0WpkpT9dK38r94O85YECvjrCLMZhZBnpH9QQyLv1A
xQo0id+KueNo+psGW+h9TGY7f3IxpMzQMJplhFkvLDtVRgLSYjxsjIkU+oGMHMxIjFG+Tk0lerDv
3AMxV9SCI5eJgHqZlmEgqM4S+sVw9dKgiTIWTHwtPw/KHCkvzdVHrlG6vA6Mro2zZxGzyRdhnms8
fR5fOoK6jxZ6MZzVHfxaGJlaBnV7tIpDw1cC/mTXcvn5cqbuKDpPqSlrq25JKi3wYALl0qJwYkky
m6KMzpQpQLvqfYNIolwPlECU2CreDXcRILJrF7tNXS2dLWx4vU6xV7Swx1BY+Alxh8ZXmUQiU7Z6
F+JLxvgA7JnsCrlqAQavElm/35EjCkDRB3x44Vm5o1aXckIKKtoRyuaCSITNVx23SnDj8O2By9ru
OZKgCZN7Ys8eZlSmYDDi4TCjknypjo/QxVJRIQeTFCqo4uW7SdZaQtcQh99iB8du3xOvydDrt5VK
/dMTXRuK0R16NMjSr0Sd+N+wYC076/XI0WXuAnIw98i/FSk5yl7AtMEHTCyo0+vuF+UCo+SLJfWQ
j2/uQd/65wIDYiznOvCQGQdG/GEGFo+dNLvLiFWkVKYZ9upauwUuCZreupcAI90ntVBDpya+IRI1
OZpT9EagzyEzQW3VodqDUOAJl9q9LI86fwIKlqWy2YW7VE9o1m2zcz6606GqZWMTSscCzyzGw+kc
4coV9Su3ULgF0+jf5ZqBmwx6w1+gYiE99IlZukWcj1Z7wXsFUB67t5oaE5Sjhd2n3nKXh4/gR668
RPF6VtSQA7bBSf20/rt0FsoqNvTi/Hc5w9D7bXVMcuvUmidbEUdwzoVrXs2jek6sD7AAOSlG2bU9
eOnVRcqzIMdVNtO5ZDCOgqrSJ0z3Bwr8flLa1GX1h2hkAfD886+DDBq+XEknjzdsJ+2XZ48FB46x
rs+z5xMyTB1SuQe4cOwTSruMfryNTnKOVbAmwSbLWLZIX4BEm+n1/tEIeSEaufDa2yeXCAmJmWea
qqZk60TmK4tJMnCu4aJwnBGvGtmRrIji32vqvFBRO07GwGWSHXsSNJEcL6Suwxc7D4ds+r894hjN
Y1GOy2my3urCBXcrx34yWLD5m7NJWo+YYzCq+1og8F8ilLok7pDMnPXi7GjOAXoMqtqCUeY2FD3+
JFSUYy6O0aw36ek62ik6DVtbZgfLwDErU2y4XUA9P/35LMwCHtCQOwD9vCekWEMUeBRgFdjpDcDG
95eJfjfvpaWO2jP6ogJFQ796bbKERU825HfcusXhxax43lVCwWVXDUat7+884Cf72ekoj9ZKzAZ1
gzLxBUNITwPt3TnQsY0K+e9lAMmOp8f842yDKvjihpPZR6hKUr5HVDUKx2Ut/SmRfElNqfJZQsyJ
MZqhXFgmQJrn1QdwWcZMvsBM1TFCvgJ9N6F78Qsd0xmnlZfOtHk7ja1mTj3BIJCuMBhDch3/UCdA
Hah3oWzVo9vyIIVp0yDB0sZw2Q1Ksj4ls4VUEBv8btnR97RNYVPGAwHKrHhU2Qaad7dAw4hd8WHw
FBZ7oHD3W0CPQ/iCjDdcDhrUmpJF9JP1OKkISHtwryNEm2sOz+GU0vv5c1JLz69RKTrBppJWvgUS
d1A0K8CG4IMdsPrg2x++IaxqEPdpfbCQh4+FM5of3FA7nfmRHjnXWBpEHZXRAM5tEWwNdyw1HLVF
ceRw9LLPz8osUqbJ2fgVeGq4ftbypgx2BMQ/RkOhEIrwPrSffSwS+DNoGuzY0afXaQyY+hdNmM2T
vRDXYjzgpBvsNEiNYlxcBNnSjeVgcuaBlizqiDw4PhW03hvu3nWMfG9BYgytZxIkUpZLTnQz3nPW
CM1jVwuD0+cnt7ZbLKPzFcTr2tbaQqATSl8uynDkjHuHQzmbgG70MssEsxfT7zomt6VPegvoNm/c
wwZ/UDrOVRFVKFpD2B/+Dn6KQKCNRkTwyKImdF/97EfUf20uSsyR35Zue/eqvQOBCLhxl0bs6JOr
61K4/DgAMucAB95fDGvvkoThioDVfO9ZZAZyyE1XZWEfU0WSW5lLAhYj96YaFFP6FnYZCJwKsB1E
NXLwbFsCnA/Y1Y3FmvXOZqdULbEXsn/iGAVt+OD4KXZnYEDsiyhoI9VTDces6ipvRYj2ss+xuPoN
nAU01UBd+us/OPSB0LN+/CM1k1r94zUtH0MsWgeN/9aTqd9+Hx2koUBCUckQpHkxo5EwjzjzcLex
uynn2D2VZgrs8796v5GTd7emVOKm7d1GjdSfmDzfaMU6kj+JbcY+0+KThpWIvxHvSX9J4XNzxSKX
zsaBCuM5HX5gmRRaPKUWPiiDbwwFRmNmUlNVfCAAjr7jp5SW37jt2nKdAMJzOqaUdOLzEakyLODq
XMKOIBKY+HkQzBtX47q0H9TPJvbFzcA5L94dWP1oGq6HfpSRhyE3mtja7ZcPngDVyOwV1qeXMzlW
1niGWaJn1FwY9SLa5fx21ZdW2cfqE1l5nf/kKXHGBO1PVgvqBzauQw5PsZfpsvJ/tdP41AP2Qjao
WKGvo4spXjo2ryxxNpQEv+nkBFDUXrdpL0kKY2JzEf4mvMSivo7NgKRqxAy/268t0EEYqXzqLWSN
LEDP3I8AFO6LZnOkRhkciK7XZWlYSCtyWpQWhq+dcxFAMG+egayS3xnvUflzE1P/pnHB4yJbieyY
Whp63dzhLfaocv9JfZnADed8AnNF1LJIXSw8UH4G3XuA9MRxhMQZoxt+0jCjR0HeO5f3JGyBOnb8
LcO0ZE51HKD1unpMBUsV72GsQXYpJZ3NjwHxpjluzX9B1FwZYKvk9Xw4y/yogZytJI14RreKEWID
DyzxSWT0IM6tS/S9X5zByq4NsMwy/xq+KMUtwakgiGyBNRPgNHyXkH8b0fOQXtzmtxWpiYlHScU7
LlJ8f+erdK0ZM9e7sFVoOhK2bedeRnk+ZpGdPEDlMJcU2IYp7js9jWOYiCzh21Fp9G+aORLZ1KTW
2tbtnj+FuAX1g3kLV4aov817Nt3OMB+7qp/yEcmTTll8+TlDwVG4Ym4MHev1Sh8DhdQMM/R0psNq
RDDamCE2xuISBoGyPTqOhPNooRyGucXoYwH2nspbNc+z51l6sV8FjU1Xrzu/y2x+TMVZ2PtsF2Pc
G3pbvH8kEwpeZDSOB2ZhUvAlGkM1d5P3QkiYE0oyb9aJ+XFMsrCaDzgdghw+Akx7qPDGUKn4voEL
KtueGvf3msNyBW2gvHr3pyhsQVL3hOhytBBkdL6xsBkZgwd8ApP1viDfeL9it+nwPetlLeE1ybN+
sOsCLlwFREi5rkg9j/cS5URadVPRuV/t5QbJZgh+RbPMKJ9az7udbqZvnDghTdBMqp6x4cm22mFh
veoPENozPvnUS4KZzfovk5H8A6AUE+YjuFnCxa20S7fYp3IRT07SQ3U/Fk+q46K5F/1sYS+/CJ9X
aVtf/i52CoGLtpuOmzeWIt9XuS+3c5L/OMuSC2MWfcCe1qB5UJmUUmyVcig4qUwtdfx0eek8m7Qz
BpX/IZPu9mdDN8DYc8DY4SPyATbBin3ia4z4/YVoJ20Yw9zq62z3yW25N3KcGKUF1JCO96m7OFTK
r16ZoUzIVQWM//0diqs3SSD81/XaXiS5RUuqKY50PlmiUWviGtl5ZhYugpZtvHSe7CsblmkSVBoi
NbtW1K3W0po/u8MJ92LT4sm7RzZljXNH16a0EenmYZoEEJ4bR8N/epWBZhBE+1gCMKSolnRHqxkT
La+ax1C4zegvfxm75W310EDwlfgP2t5AhXDZ114/Nv166vUuuXDUSUnCAxEtg8BCx/+PY/uwp0Jr
eBuPmkOEJLSeeXcAf/ZJpFAXS1a+gy5X8pZ5S8tk1pTGDHRVf85gf6E4C5WH0sS9sFcCZrt86sKp
akfhww7UdR1fqoE26qDoayQgCGkFMmVhwpnaEbovpkosWxfHqQ8LfXWGl00Ny6nh5oyLjtEAxWNR
yetcDGLB6FF3ZxJs1KV6nxckWf1eLsxMvEqsinlTWANv8YYwaW4L4a2f7sapbLXC6KziaH4EnWax
f0w99xbU1Wvud3Tp4nnMgVqMb2bhnVR/q/bTAZyfUI8JlE5iJWoV9aGTHFO5O2bGrq7m0KpATbcz
GlzkRsK6ZgN2B1INgj0YNZcLUxF/7qVuWo98TYRpouoAI0OA4yEQOuhmk4OOLFMayZm4Ls+yjOcj
jEgwVdo+kNkpYAXnJ4+X1fXndB5zARLcs/hJQ5rfMfNJTmFcaXjNWZ7tsiR2IYM60FFxhtTkhG3b
r5CamxZzHqoqmyzzgDcC07PeEFLJh7JV0QKMQ2rjsOxt5byJwEOYQoN9BdXdmkNgUgEeC3JioalG
AoO/px3sVNbn5xbYsjpF6ifHtN6Cm/uKBsPc8VO3LLZ4oujMh/XTsCA1nkG0ypq+XVkmPeJYCixf
lSL0ZXZph0npr4+11OWJDnHh/tMW3ECxBQnl+oiMDY6EYguVAnuojEQxDCLxtoYybEyMw56lLslL
MhB78MqLHKEbZRdTzRVMyF3D1/K0UMBtCMxe0fRslsct52bUFXF3IZRZE+6iq3FanDHp+it8sM5N
xZnlcVQJIgLV+65Szafhpi7DPQBKu74cD7FmsJtYGFzKKEHB5959IaWPoUwAcZc07fSSZRQ5OKsN
amm9lVKcOaztwPF7rLa90HHLbY0ErAvepLW8JmrioPvSaRy8u/VJlG4gmvqrOY671zeLdPNBPhGr
G86PRBArmd7e8I6l8aMA26+tPWqORfabZnkfLCSr10TWugwAosqOzRE5dymXApgGWfqwApJ0RVFk
xJ4n+jZfWvCfQcKc899vLCoEyns/bxmVtO73gO9C1vdm0VAjuUX24bTiFKa6M4xOu7I8u8bJX+U/
VvvH+MgT37ufVK3A2qaq6mp9c9Cgz88IC3uEJlvWz5zCHAC5YOqc9sxgZN6l0EXIqQhyHhA7yUkd
RWxz0wsaQhW0zjFms66/Prjt6ka6M9jVhciU5MNiP/JchKykzuK7K6IrnvAg41zAyoaNCXzgYDsi
0WqHPbo7hDXl6Nqd7Tgp1HHCxGmM7ph4ZX4UdVPYBdU8IeRSR9xvkuG4O0U+RSxU3qdf4TQpqkaS
sDihTYt57DcZTna0ftwNFbsHPqqUEG5dZ2dlwX9xnUoq+Lp5h1nQGQY78VG5tqzm+zQlhqvzJfpq
1n3GvxjgDsQcx2KdBNCXAzqckUkaRjvUDRF7dvGX0FhHTb5xyBwEB3EhdUSlwOYCbZnHEMVrok5/
coSx1XP8HoiIdb1CHOMxQYQropwHISnQF+LS6gsR9oXH6k9PlYQPgMohTX9IuRG0abFHGKuAYw8g
ahuvmX5MPW4eR+nMb+vhwJ3siLnMm0quyoARu7L6Qmc+Xdobr0HQHc80y3WlgH4b7teqsihyIkO6
6nE0QyhbA3PEwpZ/Ea8ZIUF/MrH/xzaY/BAaLanpvbzlELMcbSP7IALAGiRhxl+RSTfxjvrVbyYf
tprJtZDaOKi92CaTiGGdeHvtMoQ1mhKMVbD0AzKFdfgAbi9/IqzY6koSjH1VURqiKUmyT9zzWLHC
JQ+9q4vpKW5Y4qa9pmK1vU20+U0JXevHMrieZN7KOqPJptXg3XEJbyBXn84oxjkbXkEMI4UYm3Lp
KRdBqC/gntlCXhK8J9KMY7dHFajkVVlTZ7D+dA6dHbehhqo4B5m77v7S8eBwD6BAOMbwy3O3Gu6r
l0C/QsFhPm5goct2DVCXTPJhsH5BZWGj+GGVCLoSe/2WM8dpj5D4PJFVlmC+8KNZa29Kf9RrFmtg
0j3PdPqc/GLTGL0NEROUWupf2KrfaiU9Aktc28vyJxyTR9VrREEMdt+W5YHKzKOztA9TnmcxkSHz
fKW9Y0MkyuSk4li4AZRz9dRHUdFyZxdtkNOU77tOygkcqoHBXfIlVg6kFlMXf2jU9JJm1vwMjppG
xlNWj0IoaKVM72ncZvxvBVOAhIKXSEowgNocGFbXWzEhOVPfmwyblrbfvbNBx22RuaXuhyxRRTXo
titUpkprHk9TkTSXk2UBTvSdR1qv1VEBv1bmyf96AVVCReBSibnOqby5h5ZUSpL8yd8S7qv1WY4A
TvevO+hR4K7lN8pxwFZ2we8Vpb14+t2iWm8wI3bXv+jxcP0ztw15/q/bilAErQ4uXrIjRP1yzb0N
Cj0l5ayfpZfKeq5SCD1mCX/aat5kex+p9rj82iMllzyO3v3g69j44fpoci+fX4kx/p46Fb4SGO79
bSVfPnjm1dtKCZeGfgVLEG4P6NikQfSdLckineq9WfjnXSMOuGqpwMeq82NSXMntRrZRDyzPLHNQ
p41L5qGXwc1NW1ezzWLSSLEC6WuPPxbL5QamGIFBLNMCZSKTTg5MLCb0HFpeIcIRVgTeO4gkci7c
+l462tqohXI9AlLq3dST6z7AcT9w9AqOcO73DFydmQtlr7ZcW6fEFK2Slh5G6jGScGJR3xC54DQk
0JWu91Md0sogjRR8CuUVOJQ2WGpwlF+Roebi4HsPMR6RBxLAGvWBJONkoy1UqJzpP1DoCDDxp39F
QoIMsYHSvxSYEcjbm4+8x3oVSdByB9Yzk+lQX3VEvA7rYB6eN1Zd/qqyWd1QfSWmm4kHcV4SYFU3
RUstxCsLb8jW5iaYEOFR3r8hd9mp7+EgzBmxO6T7C9l+7l3OJISsDURYXnl3M1we+6R6ZP9qRioC
J2+5Qxh7a9ft03nrApihkO09DD0vbNRFyj5URX2sRBdiq6lppL28CaAXa6ykTyjKvzZo/Yil4TJB
oTGnlyrsHtYPRIvYggIwNsUUXParPya8Zkp2oidLXeRsgdlD871TQxzeBDH1WD2SXiNzlS0BgRN3
x+9yKbVzkp0Y5ryahkHTet3ulYwumTW8Vcu8LIv8y028GVtqlD7e5VOd+aT4k5EsXGs/4KP8kAYm
CuZvGqsDBArtO0hbSFuzOeCdkYarbQcQyEB2vFX8oPMw6rVVddJwoTKzkqjPlOZEJEVcW3+t68ld
R2KpEoocqsJYne2OlgwTVb9SX9BcfKO9tGAfRdOqd41IUCJePwEQFliQVaAJt50LgjiatWIBuU9m
jxHtunC9SdHe3lAFUvetwpMyz5dA3rxPUqH5UpNXMyOnFA4Kt3KYuL3NgIJ2Q+y8EUaMKcCjdgx2
hfpbEPemLbMcHzBKPaNBe6u4TmgyJ0ldskk4xTIJoXHcN4CeraQpSzHQfqozO74YOpaHdf3CWPSo
SShyOgKrAkEFd7LnfPtyAfO6zSIn3yGo5J2zEY6oWljrBZ/AcI5v2IbKy0QF+AP7ukWJkpibRsrl
wPPav0uWLT+0fVnsKSzjNmca4AJtgJJDFNH7kPaoFgqc2cbx2R8NW3tGs/r1UcKeR4i+KRFftax8
AqYhr9bQVga2bFu056mxHdFrhc2hFfy92oyvCkYVMv2K8UYZGXWQge/tXj2ie1LoIjUb0YoMrtGK
ouaHmyRjHe1F8xsqtBnv4dlRL1b0E9p1HLwlikigfQo3r7wbmP2FbEvGnAwngreNh8PjgSUOX077
l8CZtma0VXa0ziht6Kcb8Y3BJB1o1XuhUcGdtJ6o8zwbQumxhMSwf42wktfxB9Jmmgklrv1P6jUS
qy2+kEPWviMXoCrTgkMnLq7dBZ9V1IEdgEQsgRcOMhKp3F6qVOHXL0OTw1HB7G7bgWZEwyb/fLqW
2w/4x/SwNL0J8NTLdcJ5Et9q1OVciCr2hfpzKwnLZMMouOK4HdDBDWHG4D7UhOPTUBwTy9Q2Adqi
KKzO7Qa5GaFy2YEtiIba+ZARFTU+sdz4j10qkl4qDXlx6WkeYANEYl88548CNuVYvhJAci30jhjT
Dy+6K3ZnVi2uOLzLL69bTSwuxnP/BrAhs7o2S5ydOCJQknnNrSvpf0hudShK/oJWW44+i7LH8v7w
5x+8WGfFLDaVw9KOMs4//Ew2pWayG5kOQQZ548VnSo7KpZNRU57W6lgTpw7FS+LPiqIf/dUjzk6e
3/KtVkmOuXdOkMSgqhhmrN8lI6El10pt1LuW8ftC4Swv3Ax5zWD1hNqA2fOee/oFeKtNoA4Lb5Yg
vDM7j//IzIQ7BxkjPbpEQSzFONwR52AccszVjIITvj1keAplsXrV4eHjRMo8LIw74BbRvxa45Xeg
QfOm2DauVXmSiALiA2m0gABpN9Dhq+uPgCbit0SvVmiwc9sPyErZclgfklZGlNnxYVCllOBCT4KN
+21M7qqqL8mvlBKO/ESHoTQdtb/S+oKjtV5KHczR/aDIEU5wO+PgcV2zooT4061pirbaARLZ+Glx
Y6xwCueOGnkf6Ky3txHVlaNZdG7tSDxDV73g9HhmEiJGfgCbTP8YQX4FSsyFTIKedkhKPZMNmxGR
Er0L2vOfeFejOBY1sGx2QleLx5H2iQLxbd2gyrhx+zlMWp96dLvqCJa9E/pD0P1UMXbsn4oj6nBM
7qVh0WOGY52nbPAcLwKfG0toBJqbOmjIxzpgO02Ku+c45dggPQ8E51Om3wfqHTXcvPbkmRXZ7zjx
5WTU/DS3TvDBcF9t3P3hWjSe4QKMLkzDPMxlkcNH/U8coh7RHFUvrLJjdS2u10GbuEwsZFeuO2IG
aAP4tnRLBEdHFJ61jTEI79VBVEQxGX3e/xe9EHg56xi/+XqQiwGdFB9gXNZovcVXrOY9cNBGaNX1
boRRovdW1wHTVSmRbwJOe/Okzt2+F4Du+AJg33DCkArBkdDExX+L3jzn8Gul7p9u8SwP9yt8DHk+
3cmSIkwBlQGNtNJTlHw6Npfg3UrKJ77LhG3mVTCx7ex2ulE/tIrcT4BenAiVJmbr2cYhjtmxmEOM
c4iQ4cPhAy+Tn2CpeX8UDFyKBY0XlkswHH2XWS99TdrFUPTgoQOc/MmXLhS8Me6VuyDge6YCV4I+
umKRk8Rw1SaMMq1IsiG/cAr+Fa+mA9+RJj1zfwkbvi5QNapsKOrSvbIMObTwbv2LR9yghptrNNoO
5dty6ZlVYiDgC9M+kcv8cYTiRZwmEIVjryg+qIXmFZc9Cci8Pdcm4Y01Q2LlkotIDzYi+oFJIog6
8Yqr3XfPQkHXF7ZcM76NdJI6DXOMBU4hFbAvAgVggGW2WfEOwcxYqrVBxU/HeNr7kqUqV7nSrd8C
DGBTvnZnStKzR8mYVc7F59BNuG7ru+CkvKfI6ZKGJ/0GPM5oD33Ia/VhTWMYiLqlHXRvQiraPtOI
/ANbPJSokgJAn8UlRguJEF3KC8Rk/hBs7Zaz4iG0tvqPPwZ7GrNzLBTth03NIV44XgleuJ5LOyXb
PXppt+D+ntIxuo7mkbXj5Q5/lvYZ7ilFgyn2m2sKLTR+B/Tjo4n3cXECigTKbO8rtWkMuAALpNLx
LiHsI4rcRXM5j0pq3t6CZSDtAzBoIPYv75WRtfCca0UN+0qS8ppvyCe0CkYQ4MD9uXuXy6zfr9Tk
cGMdYs7/509JN0+30CfxFt/mgIEmqWYWuNIgTMEQfAVhk8MSwOWc4x+uxGgxFDrRKD66uQLRcRfC
Z/2cMZPvX1w8SGUIe4B7QnAQTDcgx37CyfUeGoevj9CD1xKUrHCq2NbfxflCgn5ANxmOEpWKdvww
NDXslkHYDmlwZzXPkzooR+HKAcasFPEmciiAeAS6BiwvB+GmNgG2Y9ILRtJ0/SHtFCyA9cbD3Pqa
SA2ifQTFCTp7cRINykLD7cXJ6j63JR/ArGBTdbgQSJs9h8Qk8OcAw08YWPkR57vQ0xbT9APVpclf
fJWYGgRKRS8345MwCNRUaB/9sU38CfY3UcB/8ZXcCRnWTgdGTudTGMrgvzGPuEn2tKuukl7/RD82
JWDseo2quDENlG+m73Hv+OJys6C/T/EXuWCirrzgVBSr/ENtSssYDaFTFsSa+xAYOZmB22uQ9JwM
/jbpTwekBpVCgO1jv1bvVxvbCRJSXWiv3ye/Xil0uAyS4GCjqJ5Xs114186etDU27ble0swJhnxH
zg1xnTz/Vbz6G/QQN9JjdzJ4fo1A0NXoEQ4Zgk8z9T/qirrzwwSlJ7l2HXX5pXmbRNu26RlQSyG4
9yWUZRVxunVgdbC36sLXxxc/bxJYt/PWdayofH86qvo/oLDAkrBRH3AAqRB/fefF0FzP1KyP8mhP
xuvNmv60G8AyOZREDObxghNvRk1Jv+CZPrEmiLxWT3C+A1VEgJwdkq0df+07R+vaY8b0qhGnCPxI
zrEZHxe2YZ8t35rExaRahs60r68IC836OJ8LkRL5+ChopR2yIsqDoPD84RRD94QRYxrVClsxTZ5C
Qm0n6SRchnlW8V0vFzmRfkWQHYkpFJ9bP2CqXjdsgH0/guVUWB4zKLkcI6OObQWA4uTFnRxxQxV3
uGNWo7GOKm8jZe8DTR6x6ZC6CrD90U1EGZ+MY+Ey1z3JIaKSrqgZkZoXMKV/EOA/H9Sc9dX9jQmv
KP5LtwfhXfLWy2fUBhOFVMCc2yV1Wtda1xJUXzNcKyHh88xFL9iQeoDLpApCWw8ke4oR0gVjnRLA
nAAl7X5g/rR/zaPxSPspECcS5cm/7/vMaj3u/0bpnqmJTGH/pOMmbyVTug/LjXJm0SkIhEWFUGdt
U3iNQtygyCXpuDcEtBoxapwjADEeuHX0CxMrZk9wA9VC4JvTIR02wyWK786vx+JgGoXOegwACFFw
4KkmN2aJHyHpcdUMfezoEMXPTDjl6YM8gLD68gIlLYASXceE+OIVNBfZVw97ZOtihp8gTQFQPIkH
sJIWwAvUv2MshmkrFwygJJMPx+5YJRJTdOmqvikJVpQlP7OjCchZFD5aw71DGnmNCgdYaFKHnitW
Vv456His2D7DQ1WoE3AolrRd8L1CjUYJQYhkcqh599ZNxNWoiOJlZ6EtRs5BJx2Za1uFpb+vsicR
G/5tCiZGtILk1xBhqkdd4N7/J4Wp0aqxc9qkbinlcFpclqa2vNQxIW5Tf56Jx/tn0atKZNK6grOH
//LjRfoKMz7Rt1w7yIlhq6zG1+iDsh0I+DZ4YSQ1E0GsGQNHaD/5WUqTLYdVstBl9SMtIED8v19D
iLZ/BI/88f8L+jKSqLXzqboDQKL1ULLF3+tK79K8bXtLiRQCGkyy2NxopdYjBLVwbYBXklwU0IK7
s/mdENA4Nct2WunH+DGFHBc6uiOgLscPW59k7SlAn0Dg9O2NPB3VUGajXIAFVu0TGkxGfJFgQ/to
Tv5n/93iktYFcdb522mJWer1Ml5by+FU+tHlLlpm8z+EBG8SE35Z2GaBLtN21YsfB+CCK2kKGx9e
JchncfghwtVSUxPMfvGw3UngzrhfYgR+6XsEDzoVrVTETHSvQ6i9EIw+Bb0ZdnTdeDZsHJwphHcZ
kA69Jf23YRT+B5l+13nyvCsnldlvvyYlE+HZpUeg/l5vs0PZvTuhM/xbKDxsfYlaWp94JalE/Wz1
+zvj+UuWwbfwOe3gEUQDzjx8i36k6DaATloc5lMOdRdA9RLPO98SfrWrTT28hjy1D0UrNORkp8Ot
ZPUvvN1PgrNGXkPoPkodpUscmQgQwbLamPhdNOJLGULhW9AfdAXAOvkk3hp7PctTXDZw4LCPCNGn
vP0VkXesSJkGE2tYcABP9gVGSrCstusU3aeJrbBjs68rl3m1X3CtjngCuqbon6YT1KalCGG4NW9J
k4hqUKTO65GiYkO0y5OOloxd6MVq9Jbr+Oe+c17X6JumIl+MuWeNzvxUisg83dK1VDcloVxRGwGp
i8OCNuG3aIIxG7NHjTEFcCpXetVX0zJ8KirTzO9TpjZL4EaMWBHPQbV3M1kj4WUa/hx/rWfR3zuX
Q6dUPpTVkRndpz2Xu/VtRF8sSJdrAy696PKp7bvn+KQL35/05dBQ0HUsek7Ca1otb8D1DbNtAFBd
AVJ62oy1S+B2UHxFnRjue5eGxXNpw95y8E3wo2zRJuDDrfAJH8K0T4Fnke99KgLlJSWZsnqlLOKG
/MiPKSBrTLwfEtfzeAM5ZGnasRM2n1aqyYpjbYwkdrd/HXkb7HPQsBAB8WGktGEmgz+fSKpo0/kY
mbovwLtbrCadtOOCUJIIBABglU+ntMlSQV0Mps81el+/+hJGEUIXRjmmhDpVngxvTpJdSmzyD7RQ
oKoMkrVqblbg12LzBiArIit7ZpBbl0uX0lRT1bz68gMY3nHr9iYXsBkMJRdkvPqURNkMM5qjINXr
S0A17oCFWJL6ZuZxo0OAciCsGlvwVGolkfw6zC2pMIP4oND5duuXFC02e7ofy23qeWOhscetFZIT
wojwdXcx4q06r1AglLH6c3IWrPmcIOCAUD6gjBYnqhBql3sdx0al2qr/q9khziHNc8ELvSaCnJxR
8uJ9yt9CbUzfxhuXHuUWQwMqUGefzdyuDHBNVQL8xuu3fgwvguDbJf4BZJEhPxW1UJ8UaMfNYQVs
LCbHP7kecj4SQhtR+XnlFIy+edKxHylGrToytdeChbtk+tcuUeI59MZWO3HNp689SRBbo4YWcpmQ
uCql6hJGm4s35tKpUPhZzi9ysOUqgHzp5rLaSfXlSbg7+6wo1Qgf7TGy4KSbzkiiLePfTNkQ6mXu
fW9L8EnB33wBHqZpFheNYDOgiHGcgCSVhFC9zZCIShtfrcJIBQwn9KiawPPMcFKR6VfC7m7tMcYt
OZJ9yVCi6gYNH25yVkfaYyRHiPaX4GiToD3UTBdrxKzwcIpK4fK2MTTplYZOIoyCnEHHGxSTkfTc
jtdgguR7BTGDlZ3o9MTREGFQEihPjRopOGgoOoje249QH5RLStN0Nv605nTqseOR159eln0ZKBRS
uDaGY2yprpr4cIpcp0QLFnTrkyjVEoAekXo2yZUALkUpw+/cbuDlyOM4nYCGuhEiS0bEcHOfbcRE
C/KfzpszISMhAyqCroFrdnZIi/pH71yjujN9FtsYhgLgc1cQbeZ5FZgQGaIG9/ndkTtqOZblTIl1
T2n7kiS2oywh7/qoUxi6sm/oXZ6C1owkcz75iOfetiEdySk/8JZ5Qr+k3zw12rxX2vFA2xH2XXF2
/l30lmNqAalhMdyZam70toPt86lXYhuoPJSn53JpAHXac6Saar2+bWfAxapANv8uOnucP/b2fIt+
R+1khZXXQR9YO7tiBDLcyc93+8EBt40BP04t3gFNAf4KbxLpwl5pYTmWewKCuacQw9rmBNTSyzDQ
NOTxhK/D1DdCIXqW7RPYInprBmDQekFuBZ10ZDLq+SBmQoI8GGMx3IfKV8NI7HW7Yiw95mrlCZQu
GAcKif7ptJTGPZ/jdFZEANHfGEpvlInlylc6ikrLwV30ohRIZhhTN4uZl+gVmbzOzukktH6oN7qi
Zp3YR7lsuELH9SYY4tCRY8G4z86YhFBSW50j50AbtYeAocP5cFBDUfEy/H2+QXlvVc6RrHWWklY1
nMcUBB12e3hv/CHuPUaqtWoY/jxgUuaXmKsA03aJgGpkMbk1NBjO1kV7a71lLq9EONbIQEALKPJM
Jerf6+PeHrBbTrUe3JBr+r1+y235eqe2BFeHKs74Wt9cvkRWmLq4l/TV6BHWXbN0mO0mIe6RNPhw
EESlq9qiGJinnXypKK2VIPrzBQVVfEDaXdGl5tCiYBXa1MFh48Q3lfuh3NEBDQoylh8jLScZYvcG
dE8fDx2w1U51tf5B0KbeS8vNMuGsoTCQ2ffQxISpK0w+YN58+ykwNfCKyQfYQmHo4KeU+w2Vh+9i
KxWLusxSUMcjJa1kHsHmkN5bqByhxZc0NcTMyltPNoAP01HD8F91VLi/8YOuaaedq8KGoDTJLMpo
towCjoCQ0vt6IXQ85p0WXXlOG9MQXeurO4kNtfubshkIBZae5dcOAA0MoW+JmEXziGMN1HhF3/m1
C85nLEB9U4X9Uvja+q0TxkIcPdJxxEeNWzEK7kHb+DTID18m2vIMIQPX680rvbIk1k323CQO4F9J
FUfuVy0XvRbImFSBT/VUrxSTlrN8NCOAKOHdh1Mr3FM4l2Cv/n3gtce8XsdGL5f8Oru6vnaBI5g/
a9cbuO6Z1+N25t8H7E/dz+MIe2qoRB/9U6/o9FJK/MrJ90eXu+YE5liZ6l65f1ei3/eIS/KOkb5z
2sOZF2SY4YhvlLIFrCDmo6g97MZuGP+cUXwHTkpdQvVzmZD9noFecWspjabvzcsfQeHJZhl51aJt
8Gl2B0ae3mwdMORprH8JNZikP7S7fHf9ton9nv1oe1WMilFJqFzlTWttjSChpKb5EzD5Xf8ak1fK
SZQRHl6jyUjzMzC6aSZdb3zaPVMiOLoD4etpYJa11ANyWnk3B9ES3KuvSBU8NGY5FYaqt4YoC2Di
WGiqty+cX6tuOSj2v6LDvPn+pf29fVdgQlMC5DyHsarjEP/hoCdytFQCjd40UI1gBxXgj+Wvx2SM
Qjj/Xx5lm+WYZkCmeJ2HpQVWE9lDtBXvMrDKsy0zsDK6DU/3goWDMWlBlJdYOQsIHzQnIaRJhIVK
BVZ+aLHj8kHgTeHysgV+1Y7/ddLq3GkkgEvRAEoIHJ+Gjocv+roZpn5I8U9pWWu2verlnj4OXxQr
ulQ5HxK9NvBbpFRk0OKoiRITHASkFJmS/yj9v58k6CtENQmES2ze+koBlS3U+6JoBtzmDI7EyHNA
7/YhSV5SGag6C1FygAvJL2IrT0856bu+2ICKobVqdCcUm8EmTt30AfamvvuIEsK9STw4liRCNmbs
dyi4KYak4IahjTkPcDDyxVDPHx2FlUiiLf7xGQGjtTWjvRo19qnC8+ZHctx3a1LBfsL6nyMhynTm
5GT9ymx+Fy6iej5oPYio9CHItIo8ZIYqE4u+QAzEROVRmPZtad5SPm0gdcF04pybmeULSnJYJbid
nQl5WR1ZKJx/n1DumSHSbRWXqQKQ3QM2JJ+tfb8giTbSaM2XLktImpmOjSJPlmSxRn3CTZulnsYL
AQoaDl0+v7R88upMUbS2+r/mODwlEN64qVsZzsKeHCGzp1JFe5Nmiu0m++nWrW56DEcP7+26SANG
Jr9MwZpNocTtxHVyEZbxnSP66yKW+ibkhdcy4iUjvN/EBJJiEtpmuVOXKK/e1apUnQB9gbkQ5c4B
qCNFSQE1eTvbxAyRMDxwkcbDGwzsCYFtdfL8AcU3gdkDX2MWHydJ4Q0jqnt3YLVpolfjP1QENlTx
M2l3IrSgOr47O/hzOTgZtirSW2YLlNXxaMmTLvtWhjdo40qgfzg1uFu7t794chtVAJNa8NtWg8ek
ccwm+aZyF+87inAzqd+l/NPGgKmabRxSSbePcpKXTlxT6LnaTlbJ5RTy6kMSgvB06sv3qvhqYviz
fho8kwl69baIyHCmcl1l+LdPZBVkIE7VZUCixbgZkoZQwxFoVVypul/Eloa3S5CX2qWlKw4koTCL
2VSNHeun38TDGv4hw9JabfQrL2CmhgVU4+qpo5QbxBXtsoW7hhxW1cfpJ+aPpn4N+XGevNwuRotj
6RLrK8U4mYv38Yz70oc4tX4n7cEu03iShvpnM9Xqp4p+5ZWxQnPFd4ijmkCCLr0KERHLnL8JCs0b
9fql/gQqgQ3Bi5VJfd4aGqf6CvomLZlZFm+ppZTTYn6nZ1TLG/p9BiHyo5p/rJfS39U1QbRXF1Lc
zgvlsGKXFeTlJPXSRf2dcp2ELrObIWOr3vB+5eVovOaOZX169d66dKtrNaieNSz6isHBklTvf5J2
4Krs43lcLaJojQVgZOUhT0Q9zQCyucKofuPAEcAFvk5AuqmwkOU1hRJ89SnjdMSfV252/FsLz29t
ttdWfReDszf6UTOaHdP8odvgKm4yaNaPXG2ONfCGAVwLtFmtA7Qx4vuwOFPwMIDnFqJ7dR1TJkXi
Ktfd7nBh7+Zx7qkQdUyXsAoHM+APVUowLba+fETjv2nEnkAYY7Fn/SmJgMwHnAMLP6MryY9e7ov8
yvBfR9ISQ+bFN4F2VkW8IgjPd2x/PmNzRAGIS3t1FfE7VshF0iegGW1vtfSxW9VJSqNRhW7TPfg7
ejxe3APal75Utbj1DGA5bCrmaS3dpuVs6T+2ZtMZxIuTwPmaBsipCMPMuCjIlkaomSi/CIVhK8GL
gEHz9gTelg0B89mUrQKiezcxu4rC9UYUyVv3y/wl0eXEfgHTu47xcsdB55ZGJh9m3rFn+XLRxSca
V2umKwnzcGUIgEBuGQ2GeZ52MZNdFHXdVZMYAX1ZR7RaBVy7Dssge7GyJCaGV3yi6fOocnT3onHR
SXoFVzv7jBejLWMwtkJOTa0sUK+jTCiIC3lxILvCtP8ZL/EtV8bwGMtKWKjew0om5V3mFOW7FymW
cgXoyJWW+6tE8TkM0d5I7HYbsXE21KN4liixeX10zJ6V2CAYYQA/ELLabF0We62CjrilDBM3dOMQ
Oy/4kZ7VHpHl6sTu2NuUrDTyQ3ajkv4rsLQsEKY58H8sRPf+GSNz6Vt8qWePpTAS6Ot+S3Vg/2ZI
u0PXCsgUKybetNN6vkWmJY9V+j8q583qECzFyj9pquh0rGGOdBSFN9Ba+ZLqgX0KPDNoytBoLL08
g6H2AH4Zu9rjouxxmBV3NBdslaS8+E0WcEAc4SV+Wl4qcaegeCV+xQwpqgu4wCmSp3iof1TYXAC8
vvwfgEyaYEDi1qdRtcO9lfw48C2aglqTcRpXPLDafnA7coaRpveT/hvq4zzH08hTck2n5N4WsHGe
AZKqaLNHPT8E2dOMXWHSq2vBu2SLAjofcmyRdEnriFuXIUhRM8p0dNzRmIlppB815abvWDCKvs5k
gX014t/Uk1nX+9L8icIex44uJMo51yilw6Ihgy3owVTbZe0ozFFVKQz+aIRq7s36SKiNAwGjm4Nl
6Rtet2MlJOl0p8V7J6iWPJqUVVVNAUqp7IhRRxu192DeyfYzocpsc3Ltij2SSz6AoD8hcrHQEQga
iLMqSB0qosiigqu17GXqk/bb412q6c3DR1Ugp91u1NCby37e6IgRGq8wnrLAfbq4f5VBxKIyIqEh
RETldJiZtGlVrZJJJg00PChPIkTVYo7zcNiMHsx95l5nMywyYUicEMmQz20ZqJeHygBKgbsmdnmB
rj0EbUiX8AM97Xm193JKlvDYzk5XSfC/t5+H62CmpD+UXSk1xLMnCE4s4XncUSRP7b1yPXaMk6MG
p1oH+S+dMVAy1D/xiitd/U/BbeFId7GH+DNGGwCh2Iu1GEwblZr3X62j/Qdz35JDZAFO/hyj5OvF
tyNOP7YGvEahdExHnouiFRs5KCSQBH7qPYIEJovsXlQJx1A2TScGadyS/9WAQkjbfWRhpgh8upBd
0x8YC6EU4Am7RULu6xvVFPQXUJOdldCXBVmOcYqjuRYgpc845OYnXxjRz88lwgCQ15xeYVGPLu+o
ezHy1j4X4RgYeYAQvQEksMV1HuOw5f+YIMlS8Y68ax4yNN75YJj/g0YhPcNiBTy1nncIUn3f14SB
AdSAGKvqQiKI3o6MI9rjzuMWNX20GwGgSBd4NasGJW7uZ0Vn2Ik23kGDuGCu1hIrbGYLQkpkJ819
TWn+nrNfxGBQEQnBQM9kzycvw6XHEOaeEY52HRfI9OvKhXWCGyMVc65ytFIlUA/b4xy4pwpjrSMJ
AifSmoU7EaPq23e1gwelk02V+DUkkik32Rb45fDbAFB4jgt0n5N91wbl/LmRQ5in8f7xfSoL8zeV
ZPIHV5k17dn+BaYRL5t6RFzAXqyUiklG4cnAgEYvXDSDZCmf0tZy3gKU7i51jIpZvJuW4f1Fuu4O
XD75Ie1zhIXqe6Q4sXhwwzLF0mptj1eONQ1Fjuv9mHeoC0v7XP9077NrYxMWU9fujn4MaTK3Bk0S
kmmb/Op4Ocvq946yO2wSO8/pxbrYMnT4DXKo/l1e5r3dqy7axLwbiCaBGGsX1NJJtBKziYuBcOzT
GSsk/15yanPITuWwud7mo06ofm57k6AAXjNHRoesMOwnaXyPkYJy3Zk4ujOCcCAEEtHJx/qOVoeY
iEu3OySGdFEO7DKoJHm1b1VlJsQuQM6ouZHqK82hlE3pfYJWL/68d7DhPmhninhgITu4ZNT1433E
seH7ejqzO4NJy7krflZYhTLHYsBjNLHIHON8scFid8PpTN8JrvjSh0rIBhz2Wfn6Xh0UfVDEYji2
ttTUe0eycD5+MI4IssswBXJjZV5DGjuXdKFyzJQJWF8jh8adHL30osWMkU6X40D5liCN2VtqOr/K
149i5Pgl3xR8tbXnwCQHyRiggSNr9M4IBoUfoItDJJixHrMsvXHuEhGLG3LDjiqFl+ubdiMP2xIi
08oSR15FIzJYWDveIHpwZqWv6Vntk49dgmgvAVFw6sD3+COKvg7lQHZfVTAsnsbx5jxpYE6hgmvI
/qZVnA0taRt/U5mzOesdt/UcfsdgpLq1UPGv3K3+ZF9aJm54yBYPF2iMoFRPmYmZGGIpjT0PVFDp
b6kXJb5qKNfvgt2QhxKrQlRHLz9DE4SsbMb6BqVHpWl5HS0L/RnSM8ZN0y+i3+/LIZPdie+ALTdj
ZIXgABoeqWxbUNChca45LL3rYxUR4EGf5t8UXMQwiN1nlfBssu3lXlWiw9QmTlmOTEumB5R4KURa
p/iudQwTbt1U5xjFvsXb9QhOd5s1g0XzPLgMT6RbmPd4kHyRt/7ozhroJE6+Jb2jcBzRTtl0B2zf
ryX77ayTDl4BJ7V/YZDnHKkjSmhwsuR0vzZoa5QyPMzXmNVKW4qQS3lxezql4NNhz3fq0qMk+UF7
1mPBs1Z4hpjtfms3qxII7V5S3gmE98iBYNRe4GLj5QCyWtzMB4oZvwQ8kQFNCImz0AdR38M3FvNE
xuo9qdgG/rHwxz8DvoHYruD72eivT3JJNC9THVsrZ6MmRjjQXqSsbmJSXF7Bsnv02Uj9psqRZSBr
DwCCG4JyBCA21zrKr1177gGwnNNcAcNTdItqTslyXcmPvdFc4QhrCwqoI+LLR1UIU6Lo+MN/SkRh
dRmhcK4oi+zKO4ypYsDQq91DE98Q/PS5vCeZLF94fViK/qoHnB6QDk9kXrF9d/lu693n/DuUnQLS
XEfM2GZjrmq/1En/8pgBhBdkVzg8IkCndtPg/dIHo09mgENOCRl2gEVMp9D63q5KQ4dG6+FBryGS
l8EhWMTTWdaVXB3mE/4PpQoKHWJcz5+Z/PO7pOQdkbd1h7gsX3ns+P01qLjX38zWwNbDaaFmDqC3
h/KD+GJZX+6cmNkfJQuHwQ5Mwl0B4dZ8xeC/lSC+GWVevrTZg6qhMDN7MkIiJE/oQ1xERZEaFDML
hh08M3N+Ld+bj35k+USIfCRrb6XoAgm55Xa2F2d44fQesReITzBQKttJ3BGU5IfDfIkcuwTsf06S
9mM1KjiMlgECzG4o1IJ9MqUyCej1BeR1vip5Uf4SKnyae0fLm4Y9GrRmnuMhF/lBZbqAInZMJ36f
0H78jFZvjL5R9j+RF39LKlY1UOvn2mR2SzmwE1g2cHqVFcryw7k2EIsIfW7ahPyE+Sva56L8AZ/X
klJQrVN1UyFcSlItnnax/zpsEu9194A9Zns/DCVUe+71+4Nb45dI3MoZkUl4AFogytSdsxCWeifR
i1YuS2CIBfsyYvpZFX2nu54IEC092vrwjC0BJXmciYrKZ8W0OARX0ZHnRd7s9U7+GAWr6DbWwLTE
pQppvCy8lqbPeY/Dr+cgESGiw5ql1m+esJUR2CT4u+SyuB4tliBeEzqTsSRZdoklr7glyCfT1vAP
22y42SP0q6ERiq+M4PEX7UtQ6vSJKndsg43ArXSbv9gCg41Y6n/QP0fYkkbdNTvEI97L9871+sIE
PMMtxyRZqZZEjf23zleqTJTH2yJGGQU3+qss8fR4NC/WAZ7IjWRfUWb14gtELmfjikf33MWE/y/H
qgrcsDvmQZ4U0uGQhKRVVUKusSshoHVFdWB5Z4XILs9Z9e1qpN+IVa8bqgozzTPS7yq9qNDU5MCp
eodRaW2LpE8qpTi+CQUIsLbIzvPKTTDZrYn2qjm8jTsSIfG4kD3zb6fQ015ZFJV0x96+LiKpFHkf
vaOHyogenfhOS2stJ5LvicJNwmRqmUFh6ejeIMNVib/9m2Dc6XlYGKiMBnJB1pRPIUhZrpdeaXV2
YOpi7zlroaHxpalg/QEKA3K6L97vzaIr8E8R9nfBs+tgc9zsgOvuAZ7esBl7GeJ/Yl2nlzuTbeUp
iLOuyOYYfT6x4UnM8MSuXayqgLWgenlRAds7Mk+YTc+Qse6pdEQEKHvI5eBxLmXv22PPvLcmQLnF
jub5YEcCp5Kc6iMIWP2AWqTWUpKwbHb+vyk3KsbGDkDQnAx1buDuUmjj4/Zt3/ehEcuiQoimNUPe
5CGW7aGgqM/7nQ2FpFRxPEvo87NBmFCwwMhop1mdifAGt/WTjuDpQrCwnhdJxNyvyfrgRnskZKZ8
A3ID5NP85ja9zoCabw9lRN8fa1sZ4cYWKQUk5C46cI43+mMnpAjyE5RQG0+IiJ++QRHDOTdhoyFd
1OjzCD4I+JU8IzJCcFhMJxBRbtH7/sH4MplXg6IWEiGPFX7+OCAo1mwohlFPg01f/Br1qLOYTn+t
xbaL8H/nc+sZnD1MdzvcbOBdtZ3gfDf4yDtU0UBRGZLZLmS0Ewy1XFpi6moNDdg6nBnle/N9RXao
0DEPTkkxt6Pdw9/vaC1l0B+vUQw8g6HeLguWlPj6qe+Tn2jiLwKgiD3ED4dx9pJylqQy8CsQoejE
yqmK1Fjh+MDVSOu1GcBLAjrzRni736Yh/jSVbz7okLY0Nyr8qgvM6anG/0Vj3O0fRVP78BXYW7u0
fCwhW0Q0A6kChWJqUL/voUTRw6hX9CBONjPImAC/sDnHD4qVmovKteKNnnR9Xqfr8Hp9jnPmq8a9
CObMoUwH9LuRBsb3kmvolwfcpCZMfMbVMV0SMkJCImsD8NbtTMLfxq1q1sinxBRN0OPWbE0s2UnL
2S1G6mETOTaB+aqvEBn6VwEZIQn4m3qcUmVFQUQyB+IWHBvsuGEhXxSH9K+wiKrtOkSarfrESOYI
VTgK8VZhjldEqGpJ/urWkn1rFmvn29I6z7LCeKjyHCZvUGkJEY/drpn06aep3WTNYYs5UQYWC67h
vLdlOLGgCVld337YNXXKQBIzFMohzC6IKGH0tumEGzc12nzGOG4kndOjghSIQPy6gQ6JhhJxjmBb
BBmYjCCmbIm5f65L2Ml1CgkUsa7MBV6zJksL8YXqrB1B7ZzcloN28dlMy+cH93uiiy810gMgKW81
60VDKC6Ahw51eAOaG1KSA46XtFt+ffJQxBc4FSd54lOD9AaAtFMTAZEjoL9hTGblrxG6TAduTdVF
JAWoDr+cqoJ1za41jU8RNs6OMkWdneHDPuSLd8koLsdFeDTljyPNVqOCumHFXM/pe4XVCs8MyxYP
GIP79fe7D5gzmzu3XwkBaaax1xlngY05BCXF3OmNQwjXrYdHkCOjwbrz1hy2gZ6j9UTgWYENSzoe
yiBINMmNaH02cis2XoFgZJ8wp2gXss9RlhgD0E0OoEga6qcTGS6LvV0rY5tiDnC/WPTv+b1wa8nI
BRZToZg55huUq93VqU4LZkF74gV42JY5+1wtxt4v3q5wERxyUQS8+/muwm9pYTmF6QSCRj2W2eXI
wwrt+F29BhLAreV4paEwXfGeF5rUPbeNhguZGsRcAxbIDb6jqYRMsW2WJPVsOM+HecvSdZEGTgvI
Y0ak/jNDKTSb7KMDt1GqDba8I6F+u5pfw9aTEbBmkGiIdvNasivLm2PoP+cJiLJw7CHb7L8+ao5l
+/Kvdd2dWcg/uR7vn9hy2bIwxfyycIyEBCzmgjglI58wIx9ue2KKdFiek7EKT4CPRszKA/xzVJsD
+wVMqkWGF4WyXsYZysx8U/oefdcCFwglkEqO7BPBu2L1ANV9dCSEJ0sVCFjwdp9IuVmc5kereZbs
i+o3+TQke3uKv5IGgd879XSRqQJLcNHgX2RbseA5ZTf8ygt9DS1Rv5l+zEE5o9tSg//QkX5/gpCk
dJFndcX0crLn8HJ9NIHtBI+9tvHkFYQhiWb5zbzSoRLMkYllYSQ/sZ9AkvEfvtlGz7IPiZbdgBti
HXRmljhHN1VEBgG8mO+VA1cpzcKbX+ip8sEAfAkXDWBtaZGPnWJeFmHlr/qALk8hbG/AdZxNGttt
m5CB1ZzC+/U9RhirEU99dF2OoaWUy7uCmkCC33zpV1p4lh+bV5hP3ugxvZ63OfGiKSJ58o2uRzDS
Awq3IEigPoALR6cty4LVzdkPEwAmy70GZb/KxS0cNOp+T0Asq5Jz3E9CYzS3O/NMWb9bzH5UuJuN
z8qMb6HpzGZNdBvObj2yFgxrxJ5jQFxX3EM1Pegj3hM1lWBW6S7IFSxrBapppj5e4YdnTpH7cOXw
vT/f/KePx5e5jwUvRiG7yIy0eLzYC7XjuA1yANPZry/nJF94MPUfeMCYN5W11puUphYypYci+bCr
XHMk3QBqeOlGDWehL8Bq9QrkRFt8t8K6tvErN5+/4DW4wt8r31X+Y+IqYPllQUBtkIhVVvkaYqgE
XXtdeFPOly1O0WoqFxmfLO+UEBv4O1Qp2nrG2Cnk2E3q75r1kPaWfQf05kWWVdEPqg8YV8zKobI6
TIdSgjQkRcE+qWP5UrQtMGaFHBjb2imM0oj/xFIsJNFzKe5xkERi5FvlGMFgxECsTTp+DDK6wJf0
rZYK8/zqZPrW2qAWRcXBLKzQU1OUfxFTd5cx6Njavj0tdf99/uY/Sp/v48XNkeAZfMb0sDH2FM72
GfD9jIbUkHGROUeHMXVbVU1tyKrBx9KrvKeJYGH+3eYGD3jJHPwaVYKXEx5s+Hr1ZyF7CQIT2wq8
U4RWqpfmWDieXCffMgSqxxnOD7YMNZKKqY2OMM88FPHrE/0da8S8OXihwXyvekwtw2cNcGMa0CwV
mxyqphp+A2UPlq2NV+EmfmgEZjIm2B/sGGeamDEBCgPQTyA057OPVOylsCp8bMB9xwfTPb6rq/+X
K1K+t5Dkx1N2/qV/svP3yazQHAF4+g1INrtrid8D4RnKAEPR/2cGBHxqByK0JZmDznodUT+cnsQh
UTx1OXOsIgiVBQIP4MaAAJ0+BvBWe4n05pq6gyq0S7mUMCvD5Ki7etUsLCoUzvhO3JkZNGpjpvGI
TyvYSygdTAhILZcqCjn6dPkDfBFXs/TgZgBilFTn+gMZ1EJtjdj+kfm+IUadpBRc6LiMILoz8suV
tqlFZJmWmbICaTjuwX3J3JRks+zKr2FYfw7FCmtz/f6kJ0Uru/DKdWIt3dSng9R2xNNgmMjYfi5u
c57NJ95Ho+xkbyLLBZtEWVUUfrxLnpck1JSh+v9jfhYVbtBHbiwZlBflMVuRxOo+OhSR+CyECbaL
HBAm/OnAl2EdlfvWKsekUwyHq/TVL8W9D8aaKpVXHxfdaAYNr0L3hiru33MpNriz9xkG5RxE9Vqg
JL3vLItaymz6zONAuYcFPIVcIVlF4FUkFzlP4Te26Bsx8iKQZRUH02hFy7s7pWiehyKNTQw4YNxY
xpuJ7cuba4ibKDS5WXy36AmtVMhdLIAhaX2Sr9e9CqiIUn0xSEd4zvrQdaaGYksf/hR6vtopVF+H
KSr0uDDjwBQ40BkQ8BxWNdawEFj/wTTebXab8hJpKDABvd3fXoXKmlAfWi3XzU1QzifGx42qnkP8
0CjQWqvxZ0ru8l4utrnKxKLYXe4gM9QQFsR+KHf4BV4O9HVtdVGzWw7seMubB4t47+IARuOGS/TZ
vYtuUIxPsYaW+WeoJUcch4ETqI68sOEQzMWMxRWexcb0e2TA5VQSPzgBtUPOybuKguD1zxLEmIXZ
S0YausF8yGczfz7+UJiyavJdPiaPFMM/0NDp+Dq6tyygbLvCz35ZYsj/DGPhUklPq7uGaObTs6uh
QQ7cXUztBmdpb4wRsfnK67PZbSbhkWl32LvQtuxwTDUDnqMgUhjOnvMcgwsjBzn7Zz+7tzsN7lpF
Rgx5HCW7DS3G4hpsDB/6MF+KTbuVFDNw4/yO9Z35EfZsIWTS2Gq4scOiwgQt9LHuiIhdoFPiJIeG
CMJOpFpHN3xlBDNUl7LyXbpiymyEVMmJJGU/sBGKO9EhE+Mm3bAbbJHuIyn3w2wSjom1Hvh7KCZN
BPd8G05xst6YE4qcVzz2FCwmttK/TyGOz7mmEMq8L674+R+G/W/dGuZF4ergCOAucKDc/92JvEw9
8W9OYmzSgb1C/qT932lGaETXqUFYife6Gl69P7Pmh2W9GvGMpac0g82jYuT3NrDyLwgrcvVLu+fp
EMLT00pNhcA2ycTc9/NB8sRUEHsDwc4aCMNERmvh7PI2P2gyiftb5Ex1dGTs0Uav79qkAZAkp11e
/vIP1sanSsqik0/kUjsmfPfqzlacLsaq9e7qlRj84ecgxZuehNDT7pu/ycayQCkFdOiQUZOgdpq6
fOZ2eXumFwCVYXDI5LCfFhyjnQhaL7BYXtZVBDwIR9KP7XSiTfTdN41tDXAX8+1ZSw5SsKB8EpQH
dMCoA83rShHrKWGEmBrI4gJwMs3pDwAELAZCmRiFct8tLhzEncP2bXSV7cfLokzxkCacwFD0Lzo0
DdKSXEvhUgbbDS1BKmzf6QD2uEEhzgrxVxzHNahA6vnOJspddxqmWACldx1z2bosJ5NDQ4U9iqPT
Lrb1QRMPRGiw0tLFsPTvx8uisnDJG11ara3PTlJrSQfcasLC92A5OcTHW5TxITqbCd7lbf1CvPOH
KbHLko9bDReoaD25EzPsgs+F7LYFEshkaQ+oo9zgfS8H/3ve9eYL+g2nNmwWc/TRYwyMrVZhNsOK
3dJCEDEfcKyX4bLiwY766Ndg2j+gtFkcSmgTcRRT7A+HD1vdmsF4X6Fm4YMkuXJ5/42kX8aNzitg
i26Gnj7Vt7NL7EfxSM/5IQEEervHdrmFfcdEEQSVqsBUfxYfyoJcych2+7HjoMIcNaGR125VYUCv
TzbpfibCG7PJ+KS8HGXeEPwWD6IyyVu/7Yp6H4/AiJZvOm8wcxh2VCJo+jqHSIpRljIfc53DgIqY
ayApxGqD7Gvr3XwvoxEuJdOExvz2JDhu/nI+uGUHw/4sw1lLShStjEiSPNmK3AUSDQuWTcZfhIBH
ANr/KzblIdNTDz3LwIWGRrcb6N2+8GKDQqFBvWdoHH31NXeZqoizlbzBpZLV2OOuAyaPJUlmCl4v
LoNAB+/yU0fRjGLb5uVXopXTa7QhbNaW/xD3ryavTiVB4kfIpftm6NSWG2y4IJinMSPRmjQ3KbLS
DUKXSyiwQJoOQTeCV8MDjm0dtCmaFwo1d/nyuynEIDhdUMc3PV7OcMsHp53p+DNhxUZRIkAj5LO9
T7mdGf+eYloaoLF4K3/YmZdGNrW097eh3+8ryPMRSTB4493Txw0MBZrQ79+QVUoBzLWZW6gnrOOT
MlY6nPQIKu7MhUEdy8i6Y4azbaQopZGd6liStMCUMhArZ20FWD6v62ajcR8xXGncCDt2caQ6xW1R
dLW3AAdhqYrPMxkcDi19n7OsLhgEQLbxgucBQtUOyG222Q7/Vw1ZNG4mW+OnvKOoS9/JYDCByKi8
ANaMmJKOjW1a0SP9cK2Nth/oFLXXIqaKIEKc7j4qPYKkwHbuIgPUrZkLPtfD5Rb9PDFAyi9V7ZRh
uFM82fxoIv8hzQM5S+gdC3z3l483XQeAIMdEMsLEYNSEMYxU9fyJZhqCkWPrLW/bl8ZoGG7ydX0g
6NKVALiD3zqkfyQp0kkm1lf8ytLh52hT4G359vYDScE8sr8KBf5Yeqw4bp2zOGcfbBxjNl6TBigJ
PeHUm9nlC5n6h3yCJbWsnbuExueJVvlDTwHUUgatrDU1/VjtdMC63CAL6GrxQIV7Hjr9eQby1l23
0/GB+mWOdz1l8U0jhAdegQ3gfTvyREDM2Vrn2sDMiVb9dMDe+UrpxtPuHHure+wLue/Ntnj7vN6D
vorFEb97i3l/IiIiC/gjz6XAVmbGnx1SP1rKvv4h5LRKoDmVUj2cBuRfCbN3YJ26Tp/W4Qw/bRwM
HmgDidTCSZnU002SI+fImHG8pAWMtSAnevVc8AaWGgG/vvfKFI9OkPvF6+Y8HVajzXb+Pkpl3eC5
PXyyX7hsIIK9CS6TqWK0gkYXJNN5kH9aQtCEsjgMR9uSobjZzqqfnms9lJdXEWePpgwcn1wQ2LgA
xZ2ARVPWZouJ9rLx36hp10LbkagQBGJX4wSOWQ9N0A6yLO0SeeytNwikJrWpHypJhkd6deNR3r6s
x4s74VFSjAaYXQsfXBTqW6rFuKMRMPg3Lwi43YV+dMkbG4uCvBxo9reM2wvXidBcuFCPgXIP2bFM
mXd58M6U0d2GMDoPGqSvDzyMDBLnR3NAbvWEVigDFmpBVNJOSk73d8ynZ1mi5DzBnQB3uanGZlgE
GJkLxZnchbAEAHbjby3hDZIklJW8WbCSCiVr4anNJaGW9Ol8AZUjIQP9ntndX9zYQNAeu1jW5DBx
40AruGNf43aebWf3iCD2FIg37Zwt7A9XvZDIfWJSaX6CPOKZwwmZTyEbcIlmiGlBmqIAigh+48Rj
MkfSpoI+8w6kXNTRG5fyUZqDW+LmhL7XPeY8c4JhebXClo45q2QL+QBvy4atQkZ4wVtJALBF1RZW
ORL9gGv6GSn065CjIt6wLIdPcQfQGClPY2Ya7WkZLL51CvW4sQP5EXT9z3fj7vKztgnaeOLj1CkV
fWV8Y+vGPFAmPWSEDIVXh+y5DKA3Ek9lM0Fl0p3ZxhGXz0g6JBebOqwI1f17DjAyLLmZktiP59Cx
oY56SS1mLoMmLeL06FY85DO8u5zN71BeiDekEaRKQiLPCoNmLGJrUnP77kWL2bq8zlcjwlZFy9+0
lCWVg5YGl8VBY29ZWmOZ6nXZUtuxS2Rfkmf+eZd9KmQE799ZaKvun29RcHRZPaUQY+aCeSxJ+5nT
yIyfW7WUf315B7Ec4xOVzY89382KVj/N91k7REKmiNksUTqFVitoshtXVrNLeS9m7tFhC7agcLft
XelbV4eIThwflHXY3om7PNPBqljn3Yh/e+qP5HYPUqbFXlHbh7XGygYEceTFtCjf/mNWZ+V0yijv
JdiCtVNHqUHiP7fTFkdCreW+rJ53TqRKszPrq/tVd+QkTk519fxI5wtbQYQ+GMc9qNisRX0f2bhV
kpTZzLvz10uRxaWJIHn7JZyoJscx/4ShtrJW5n3rHQMpB6XcEZeLTHas3H49N7y51Ab3B0rPckzU
vw4V6X6ugJeOo0K58BgAiBi0s6tHpN+eYWgt95yys+IuReRkqG214LEN9F7zQIvGZhlG7aI26Cx1
k8K48Dp65xpZMfNxLcu3FRJbQgmfOI+GofmdO7uxqCDyK4+BjqLWVOBveyCya1gId7y7n0QBgGiU
IOR99VD2RAsfOGoRg9BQNCnXklJKU4Af6LzbykUJm9uCeCNYcA4A1X4yHL80XpEcJ/G5KypJyb0S
Nbgs3EMe1ecDQxswJQMO1H8gu8kp5zELFNvnsTuq21w1lBC2bGWQWI09A3X5FQSUmgaB91P6zlCG
srRLudh34m8swHZ3agdTyUN8Vxekl0QA62Rfg+wMC2W1LgrSjBKkU5HfophEpK4YDPMNd2zBVnzc
gpuwfzBqBkrrfVASSux+/J20CJwA+3atCAlqdmSDaKKIZw1V2hlg9MYULJQ/ZIuvhJ3dBGSXZbb4
3WAwUAxMODb/DIBvBIISNkteFyTc4YQGnfbRhIgAHGxXBhmo+h3lJKhmY9tLT848C1e1fqbR4RiU
JzNJHMcuNRIa+IpCXk/zIH8u22GxCRFzXMQM5bRY0of4vcq1Oikyn3k9XNm6ElXVGsHTOvmxwQXR
TldVdfBCyJkNLwwldflqDODvTFMEWX2ffGT6y+6m4zeYoXy+Z+Sto/Z/0WGaY4r7Ap/K5wY3SAKW
Rm17In7N9DsqjWML1ARkMszKXrsrmCWiyTwQx0gmD9Tx0maEQwRONoIKXc8ptzbXZjp80XfD8Avq
/kF9X4TT40iHt0M/eu6kCYmBNXg9L55f3feUgjx9yFLxp36oV+Gk0oG0ZkIvFM0Agwkwg54IT+FD
GR8b7srlB8v4NR3sWSkm8buVj8wzt64Uv7MWv7xqzhbQ8CEirIrEhaRanFRFiBzjC90xaoiAIeo6
HNCVgZMB4V7dygrRch+OZlNfVmNO38IX0S+Rzt1q9d2a/szpyX1afOgIZaIrlksrh9vGn4bWNo9M
aUaJEV5pY345Ykqq3BL+5QL0i2h0clSOZDt2ezTpUTAKTeBQSZ8mr+EPhBgotQTouNwwm0PElS4K
DNb7HJRLopchozsAnOE9shNisKs124cWAv6p4qfux+nHpnGz2VU1dkrFpLhA++XcrmzYxvR07atw
VViGh8EJDyK1Pz0qvRC8CTTh6GpPf0GC9ty+vLhb0uLTt0SEm810AwkHkzHXI7PpHqxDqrbyBjd2
6YEIIHFEF0mNT+f2mdCEF7lf2zevkUTVd+aVCUR51Ah9RuLHuo4lgEnCEnA6+Gnv9wdg2k//PIsg
FhAwOuS2PK2qQdYBKt2GDk3WVhaDSFCwaCQjWmQ6nYEzPskykvMw4W+4VTxRxagulijg/hUSqRlu
DKooftpvq1PwqNmgdwkmL0FYReUItE76G71LsVM0qTGiJrEmYVqwnBm67T1uvF50F37UM1+9vWG5
pJSRp9IWbedVcq0pov0DoHpacOehsEUQxMSXWGAX+wr4tZf6hCqhY8+brK2ucSRfOSvZjg+wM2fA
3sn/Z5jqGBOsh9sBvSe+G5kExnq3FL/3H6GuHj9d8p+Xicbb2z+hBez9J1BMDhOrC9vOtQ4h+5vs
MSvEYTa8+Cl/ESZVMnVqTWkGPL6E1ZTEMg8vItqat9FGkXb7ist4aeyE8bClNLIxjtCjzaVYaRSI
DvtQFsd8QiLzAFTAFsw6h31aSmiZh95rbmB9GjPP8DVPyrjmE64t3Uww+9/4npfxG2IvnNa7B1/p
FYWSaMS41SC+gbVhf+P7mvlPcG37oEtXRLN/26vkrPxZK5a87wGXPZlxDwgbkNQfiijDQeMI2Mza
pp7lFlbVSOg9AebhYvR3jWuIVRPWxEsKpbs3Sw8WYUitUO9DT9Vc3CCSkXPccHu+dOpgVyFvdP0q
wf8oVl6cQhfzfd8YWKC7CNGdpFfIiaHfjzvMNOVqJCq92QDofkcqaNCIF1QoY3lFnEwhUNCDGsNo
o31tWBcRv+ueM19SNF/yaa7x+URJkbHyRznvv6kBoJMAtoJtLXyH6z+HUN1Ko2W1tpQPJF2mqkBf
SQ6CDf2lLEMM+xzMDk+qF1dU362++uMv58jdkzhgP9OYMVYYfzhli6UIIuhFNvPS6U9ZnlyewnjS
wyxhg0SNgPPemZ+jcqXeH4RxQzxtYmyWO0ihiCEEQ2RhuSLalwhxqi6z1AouS0oxTboE45azHA2L
ihOQv84M4Z8bTsb1o69iuQgoMiq3bgu+MncxT4Qp12VPquTX+H73Iifxoth91vdylNCzIu5fua94
tReLBliGvP+EKFo2+nrU0sb3iur7oZEyGT5U0StIBBlBJh3pB0y6WsqutLvAVJ/lX/MF1gDKidF4
TYIZdR77TSGKVUwFSrn857HrFNFGLZ89qA4plgAqCBZAUuZfW5V1oLm1Gcr4e2/7TwXQtNauBxuc
rrcb0RRadzr8wdOS2JiM5XNwa3rGV0j5EYwdGiN4fQys48ubhPH9khwWo60JIwYflO+L7jzqsSyi
Bu14txOd/EoMX8VUkhfko2LiuKoYNh7n4vzPHloarXs5YNGbA75z1eFoVSBMfXJgPXW30972gx8Q
4JaGNoSUEZxlsqU+aWd6NSEIKDfEnrLvhFCMPZ7uAvqNBolpKfTZ7LMPHYHrnh9gQNpuExuTJUH9
j49bmmOUZ2Dhu0elGzmgA9OOvh7/YiAxuZ+k9IgTu8MXhMtJvp8hmbV3/YWOuwqfB/QFiDDaxK27
/RJQsRDBMQLTjXnNOZm3yZt7P96IqWQSP56Stbw8neSMYgErDgZ20H9S1TQfk8i42HIV4NZt9+tR
YvH2mDjGNjfOUxDD1o/8AcsesmyP+572eTE01XZd522Z/kY6djq7amAG4tLQoc48Sp4Kuyo5wdGQ
iENok+tKsRE/cq1LFI/xeWSaSlbgm3p92e/LT/6EctgYHntZ+RqF2cPnPM+OSzTsGynmwWGuHHdy
WDNx10NwvAfTEGZEoUfkgIT/7+rDuXQwaP/LLtqYUFrsHoXs6ilVO7GjS0mCbF1BZkP21HRdkhXp
u8hB1Mk+j+XSNq73luN//2ftDC4ETc4eIhJtLsjpYq7NyR8qzi653tRQPliE6l0RoeJXDJGk/Fjz
5bjjtGWSchEp65J5dlCetDqIyMrogDFrGrNLW5HXqpnSFlt00XRxP4Z7dvMqo7uZaiJ82ApaWW3k
axI0iVCgM1rnS3vA0e7u9Z+NqrVUR8K6DmUM7qXbpnlzxygISLLvtB9ViouI5RhkgSzZcEmiM7eU
ibPlNq+RnvYyRKlERSnukPnyFHDEHckjEYi23aFlOTJrzq1wgPL95qUoJKjlRyi7/0V+TAhh7Yqy
lzH8HtsiqBLJ/h1h4YNq+Wa4CJSBu3T1tAHYoX9vjolLuDgQT5Brw6Mkmkzrc643nipGZ+P6ACGD
UOrQPBeQU+gakcSmD99TGd+2sriev3Y8G+RoA4Uh92SeJWgVVUf7FWQDyrBr1YgXF/hMLDl2iQhW
b1YEC/oJlXf0aPhs1qBmr8Poeayv2BFwyGXfoKouhGtqZ+1vB/uejliyQcxHWqhbbFqVmHGIyo6H
pApLz516xrC4Adc5tKzAG5eWrqBh9C8CG9SkevMxoMuy2nEeQjqCPaGuhcXWAjj+/Ksr+vUCiq1G
kdHm+WsNdIaXATuArd6VkBfY2UBEecjfTnzmeCgIJU91IUT1KU67voWzJuAWzeTT6ZQFmNvZO85+
O6h7j2tbBnQHB2My0dK8mJqg+8bv8L3ql0e/j83fGSVOFJMCTup+by1JB4W2sFc7syeu6wHIt7Zz
EbN0U2K1cRdrV8H7hnfrLssT8JenkmPg3oUjwmMop5r/phpvMteqr25L5/d2ekzJPrbpGJ3iGlMf
77ks30Xah5bItW8hkUsRPEe5XlZYZwNP3kltXjoH+qWM55GYMjnOETmS0L6hVFnpkKCbiGmBCM6b
jvAgCLilKuFEbAOUIR299X9uKtVmmoePcurbeJ3OX1OCveMLumNusBIwmOYBjTpN8S0tGhEu+0dz
pq9VkTP0d74gepZdSEqavlaZFOd0vKTFzlTZEQPPa5GooBoWwvhT/RRTmgYahYPx8Icg1Tm7gWH8
usG6+xmKmwXK5GLde//8LL6wBkUk+grYlcQGxBWeGiEMhgk6jZM/x4G+ULzQPhQfYHmtb8JMdl8J
mfpCdbUMpVARd2jzVEJmyFcoaJvVqE+fyxnJTdEB26bY6k64OTuYQzCvrek+ddjGZgqZzjftmEyS
ZAeW9SHD11xNxctNFrtUVOJh4C8KpHgXf1RFs/78Glub2fJ5XESBaOoLTQh7LQZxD8BGl7j2i0DF
qbZJKlSFBVyfQBU5rLbeKp5oQnhnJNzO6hlHrqwNXjNjs5DXfNkHJpuKqNGB/Mju3tRMHcKpr15o
+YqesF7qxSIci92hcMA4DGf+5ZNFsEdDyZXBuNqSoiii8c6+MkxON3vvwNp4uZ0iikPR/spFS0s3
KpmQFkcqb9R/yYjP/iB3Tw6qpSVSyp/mjGToKLnDyPRjhqzfkPk1wfLdTLfKqVwY5O5vdxZ5ovxK
4MO/TTj1ONy1df9i9KimmorxuZKC8JAlii9hcQ6p5CTs0gGoT/3YJV7qfJBQZr8vGWlKTd8Rt33l
NGuNVpT73sBFjExXb31gma4TEl7T/MKQ1ucP7QrrVAN5P9pwEErQDtxq+dX4WChOgJoV7q9z7uH/
AXUQbzJy4HeYKmyoF5dKxn+n5rinfEkMLlpmJz3/zjmVcYwmh80TK4tN7PP0sPPKwzk9QYdCHrom
/Uudo5N7Jxl5WzH4aoVmv+5x+csi0Ghg2F+xFlrOrJRGPhzc1+TQJMf0ZAKYcp3xt/lX5tes4g53
3F+09uGwhqAk4J0H8XgELuLOyGVMOiY0uNKHSpIoSnU4f4evaaYopkE2IbABijmyv+cH4JHbdmR9
3/lFVqqVlNCyCuMDNfvFwWmuc9eYjHqLO6LOFAAx7icwOxeLzoceG6f61lO6YA3hs7aWzVDCIU/l
yuUmBCCnRpVheJcQlCyxz31E7+TRi0qewpkWcT32E3qlk6cjEUpv88YX62Y0t0ALXFtkZFyAAj4G
bE8xE8DPbEBnP6GEAJQPOgZyDRV5g8Y/yZmqZoZkaCpMD/aMQXvkNmno4hgqU/9Q39zyYaQy4Ueg
gQ0Q7ivXTJFX5Pgo5esdQMeJtgJILsd7jPyfjILmGzXuT13uOHdR9P0vhoONoohH+8NCxWBR2HNa
BkywndfnPb/6Sa/5qCubPr1AkGuhOQuUoeTIzFGgKMKuLLNOjGW6/fl1SGz5fsk14XVmJA4rajqc
ldsWxe2xHwZv2moeWbolZcTxnawZ+om8BbbHbHcgvzh005GsHVPATOOxGntfVv3DuCSumhpVSCNf
1SjDaAOxexQwJIurZxhZJ7xuQuDPSioAA6ivi9R1SAxB+AFRADlrMLah4rJqaFLdNO7C0HEqPKeD
jaEaCP5eyEY2rJnP9CvaC9pOOcG/7y4Lpvw2dsnz/rhsk/vowG5ujTFmO/EiocKXPQeW7bvmJOXE
H5dCOEbMMCnnPV65+ONt/aouu/rZbKEkZ0hbOdbi0nQ/0KJ2izPu9pqPfbRXneYlrKStUuA7zo6a
UlF1fE3Yv8ph4sQY7NRmJUj3AOeaJyuweTy6MfVoO/x6VedodnXZtQpXaN453c5s/CeaUmVZI3yZ
apZQnH1TBtnhHBFjYt3unFai03xPuKeD372rFQ9a4GpVUmH693I71cbHxi6FQc6U6EcuEkjWNkTv
N8pJZJAdtb9tEXgyIav5IHTBoImpVsK+VBTg4nP5ezi/YvPpeGPAp/tD/hLFv2JlqAwPDJRQ0bhU
9iKIHCYlMuyZ7U1dwN/02DW//+Mwlv8MSk2yZFhD4Bwt7QpgUcJXo1stMtWAqXQe9fTY58e0HFCz
2gdUoYsG5A856Irkryv79QXOTblFOqbKqxog7FgAHhSDrr0y2AGFuoJFD53glvdV4JSBrxVhnwLS
FK3BK5OrFGppPiPpU2RW++cs/LZmK2qGrT1WZMI2cp9YLckTywaaFB5mBvSKunbRb8Z7DfVgVYBR
hI6dFnzlI3meFA8iV2yUOG2lGs7dIPkhIpcZ489Jup51sp43UeoR0icXubo7T9rf1/gY9sUa/3bu
LWUIaSJ931cGInU3Enww884YwXAoB+O60zfLhIqx694Uzd7+5+r+khtpkhFNZy2kCi/AJWxqkwR2
QAFx698KjoJz4eaOPtVx4V8RGEZdzZLGBXNWJF6fndNBHAwi5M6lX9tIfO4KUwzUopKwCe/LMmCF
xyA2g3MnXdZPbuhUAzsLnyrc9jmDQYxJe1AsetZhCE8TFcqursWiO4LAORvuCpc4FEHSgS+JpbFD
lSGg0GBv15OMoUGCtOBz6jDVw3A0bB2NFQUiEdMorunnq57cNmIg0a9bo0Y4OmCkssez3/yals+c
Ubd0GUXEAHYr6cUn1p2GFrCST7rHPFOSiSH53JtNsyFEyzqpOy+hkGlvdt/axKqB9wRcexGB3xPe
5hulC+zi6XN8PTZ0jrq+ZWQf0xaXhWht2ppgx6srnw+15W7W5s4jCD6bhNOWcZ+6O7I14/+0RlHK
DrH9doX5GkwfahukalhuFBywJ/iED+OkW6QmV8EBqxpwumtGqEdmaVI0DbDtZmzeWymS5cOxAT7G
uSQYSg7AyJoUC5cUWrebHRnj6bx34w4AMNZYz7hxQr65plD9vbL5oYUwGU8V9sjdht3pnIPj3njO
1ALQO82F7wiBKhWwUacF3LExGLyfTK+FnYPI9I+uB4g79FKTWwDU3adT+i0jr38yrjJIugqHt90L
mgGXu2ZSzslVO5HOtkzeIocCKCMBgSY2Go5MZIC88xmc5GLUM/f0rOYlqI/68OuXJDS7GSup06i9
SgCEnPxa9aMfLNMcO2L5cEXzlz86/7U1K2CtRSSRzt1BX504EkyCPgCvmvZThw2yPjsdv+KJh6ub
t9tSz8cgiHRH6syME4EjuvecEHV8H1tOcj8S0FxgPQHPyFFCaWdR1Fmx1+5TmOeS92/4RYWqeq1B
TUcux1eVPNiwOULJ5oa+1Aqwp3xL+LXvIEWExlAZA7nIelv/6+USNb2ESoH9aVHyOF+x+uBdurWV
WkyocJdq+5KvoGHRkfOxzgP9B3ZZ2ZywNV1kltr7KYhixhjWGdKNoGOESDe+oKIuEUjy5NMq/wai
5woXH2nKUrQOHV/T66QenyLpmBvLbFBoeZZbqX6bK3A9uUzGiSUZehOFvNUkOcHB9ggbthP+K1Ti
Wjt3zqq+RiLlf+4/CJLMgFxMmzdx0C0iNcPoOwLforfaZyzySI/az7kohkYkJ1TNEub+I6z5nua2
8O9G3umCsm2aMev/965jV7pn8vDb7OLEtPwYJTa6IM0/z8h60tIk6qBzpGC5kReRzvllBuzdiGyD
DL0qMYGfBDIfv2+uucnydZRLjKhcVpKaeZiDbY4EDjkwx5hksv4PXVZHZz68sWw+35vtogW8ZCqP
+k05rTt+YoSuIWyZuEsY80TR0D29EOCJpaI17eWjrJBf+wEveJYzzLT90zOFv7UFBkwFW8H9oIwP
coIyrCSuUNK1CCASrs5MhPdloleYqq86jry8m24I0wCPHXGXfkqAD0P2Am6tcyDHdq3RSmz/BaLe
s15g+nufCa+2yK3ilBXm5LNomYMJXuBDeYOcgEzP7tI2W8nTLU2QGc00eReDPHiELmAiWLAXXrGx
D86w1aSOYYc2uDysDkWA79nw+Un/P22jOUtbDBzWDfI/spjVRjt2dgzW1r8TehJwaIF7LwtbYTQM
aJll6IFG93shfFlpJDUILKhJXmw2bBJnOFs6s3gLrZmzMfi+8Cma7qbY5lhPuO2a/Cf/g819/ZR4
ZQkgEBA5SjGZfK4DsLPmdNduZcxAW8cNpJF+b9XEWXBlv45nGkfM05h9F2u1l4eMer7tzuPVcbrW
fP8JTURpLX0sTtmG5IiTyo2WeqesrmspZrk4SgzlGsdJwG/ynKNJdzW35jjBp/JNGRdZL0Zlvd5n
8xu5Z8a8+wCNRBgbYHvASwqjvOP19ko7aKE2FSPfOvpfAYSdX4A2OhZ0iCd8m2Ue/agXFlKJsFsN
QlUJIxIIp4Ml5QDbSiG3W4QIIIPr9gYR1cn/L/jHZlPIk9PhKludnDcmmLUcFw6w4fPzi0q1sFzk
YwSIe0oTDQ/ZH627nGvlI38cGkjQ9Txz0AYLXFksJKHLxiHHgRJ45HRS4jKCjrqmdBCG+atOtjUT
CbgFpKoZz+khaADGB6XYqPkOuLlibTvtME77YTnBz9Sh/3z2HH1IRUCwh3+0EvrQP+uMfUrZzifU
pkQzHXvD6st2sSZ6eSBQWP61IqddpMqyeIu2gA8yQsTcLOmYwTEzH2HJvIaz3iRCyiA+D4yv5ZeV
0sIZmmfGUZAhmu1Xj5JkxOJ8FQsERUhes6lMp1uzewGBvNMelFXjOCISrGvqVneDvTg1gtoDhQJf
+bhAXAStbr8Xxp6/OGDVJ0weBoeImSVQR/KYB4U41/GTgbbN4s48v3n6dVXYYPGG9qTyzrJosmJr
R2byATpCvDpYTAkBguF2DKM1EM6OW/moN7z2Jo4L6c3Q/q5/Qyoh9RVUZb7Ym1WvAAabCYuj1sNd
ycMPDdhJ+48hmj42Mq7QFZym2MvqezxuwFRU5Kg+gyazxMygYbVCswVD+tacpmhZCsdcxS7j5Uaq
Yh4E5n8POqKNLe52eJIGGUpTQAzTcR+//t5BiOIjm2rAF9KyL7omUEXukB/9nbwsAw8sBOhCmw0Q
O+EtVKbk2dC+dy0SEmhnR7wamuJ/t+rmuVYvwuouzObW21DHVlg1SvoLMrKCu4mbrOVqLMRmbd/F
ZpGO4WPefe8AfgtzFkzKnboASDft/1sPrbroRDTgROV5vvn1Bpi52ZM5QSe1mQ9mGthLUGgHPo7G
NFSg42FVm8salT+lD5oisRta7+o6PfTaPMvAFDxgPjkuAzhUqFWZ/7Gyn4icRjeSB0hC6KsFBpLL
2CpcOVYSBAjdk4M2qNBvQxtj25dz3vlUOdIxSq4pOyT3z1UWcpnBHZ3GzzFq0Qt8PdzGK1dZEqIM
EFHiuzzZ00TYmPKLK4Cfy8n1X9y9BStxjoGfWzepBjWljFyvTMVHtakGo0Prphf8LgWSNcp6P8ab
plkyYtm7cwlKcpiQd8wCeC6bDsaHQNgVIxJesZabUaMwNZ/9Ly0pXpIoKXHGIUX0xiKfYiGbBF9C
qM9TBrDbSb4C33c7DSz87a8Ml1vPO5zRkjQXczbs80QeISQOYtdkfZTnwSE6O1PpZXkBh+Jwza1w
bLDy3UB982fssrXJ4slbkZmyYBBfPtig9KJonF1AYywX22Iy6Ex63VAVcRBR+rdzq4i7XPA1OuNf
zWlGudUzpFSRauLg2W4rby5a/6L3RtRjLAh6T6QtvQo1qKPE89suGTznCf7oQ03/7wfQN+UeFbi4
G4imPjWb44jyjOr4NU5vkJipBkIihX9Z507PtJc9yQCniKpM75SLvU9aYiSCseMHcy2REhywBtTd
6+IXRZwtqxaj+TLX4xM5F1RbKnV8lN4CtOtjNVWskX42L9jzcuuQLNXbGbSUHk2uZ0sF0n38e0eL
uNQOlCn5WZqB1jEZMBtR+Wucr9IVafcjLvV+RMi6f6oOTuIKMjO+FQaptKtcOWPDRVzFFAoTEPjN
tIaVasXOoCY1vd0s351jCVgRGoRlj7QFlzKriw9MaabWHRMupCvdCxfpIXF8XMybmdFrvth+HTxR
+yQg5ids9z8pVNIDIND5dryLIcFVwSO1ipMmWDgLxlTqsBXbmQlbWge6MLoMq5qScZXBh8mUumEm
rCz7xszLpawg9Lipp4Vo+7ImA/P2BPR7FU3lajFqkMnM+81tpSNrxxFyObA5gdgYjVNusPCC7eNn
GPFBu5fnbBMMM0cq1ZLGd4c5FgRLNbcxIg1AadhRMXomNRZuHNEVGO572udFHh9YC1eZW1jUARIr
7ZmmAQiMyqX6XyGGFNR12SDVDM2TVDTf1iDiiCGDTRKGn44dkhkEKZumLh2Ba79BdWCXnRo7jAYo
CA4aEJMEAVnkBa61V8fwzy6DlDXH+TP+2EqHw6mDCAjUeDG5BjdKQgL1zZ89nHShNrlvp52pveB2
nCv2HMlNPxHXGn8JHcccrDHE7ZcO/BYvvsY9K+IgpwWDeFIpnWobF3D8MZjqwkQNgyRFk+wJBuQS
qIt5ktHGLK9c6YR8nQZd8jl2u/taD+g6cLq0TJGBocqzr6VF1DLRyIaozhzNc0LdTMMBxm0g7O8B
mpIv6Kb2flU5tFRDEEpEQnW2SP0S3NDg/YoiH5pGYRX6upDJKv+Dsquq0h7XHI8yaJuPAteVHxM3
T0r+FK23YLS5CKdmWko2W5PeFb4xvspP4Jb5pS3PkVDpOxoToEb1lDoB40Lmu2xujYIUcfhRz9ZS
Y2icUQ2p1Vo0Lw5V1bkqYeC8CPgrUIR6xaNFs3KohUqq2kTCQ9gqCK400j1o01mI1ML1O0/D4Jow
bQc7jE9Qf2wTRU0MZNAs/5DN6GPhZUx81MwTptdsF0VnBkpK08LYctv9EgIr+nEKwodHVrJNJiRq
NjITCOdoQCdUP5jFk36vL9XJb7Jz6eddjBOzoa+R+9IUKVynbEOE9f/hFhf96EWGm2t+SlOpjItY
bW0RcjG4pMqxxtb79OsAdnecwvku280L+r1uzh1m3aXfs6ylxB15G4cdRnFqcw0Fqp8Jik9EbCRX
1c9FtK5eN5H0Z/wKl/RZ3zGgE0amnA03x4F2Y1Su9FaMZiDIpIgGIZlAsi/OAsfS1ozd3LUik0gw
oMOqs89QBEcuBbCOCXAXXSlrMFslnLF1ToHWZQCmtUI8xIGCFvTCgiyAfN7h1/jN0NYP9LhBjLOS
3O3D6+MHNVR7vn/AEdwcK5g5WhTz5lqsMUkoYAYAADyzNNZzCLMz50e/SNCmjoAA2+xFc8zI62SR
6J8/Rj4soVWP2s2x3i8plgmWnw8Qq6EQjUQOO/Nq+hYPwjlSUPF38+tMY6wiefS3uJVo0NAEEueN
it67TZLivV3KtBdT9JqYJWKun6bN9E8XiseLZFgV7QX75nXma0Af+qbPjgXEra3ReptlszAblq2l
/7xMJpltBBcEgHfAAaLe0WmO0XTmKMI8tDbyH9e/axJKpgwq8fPI2nxtduXlyAuuhHjltjnhxCKI
DbyWo99YqJPMMJtVgwxzfQ/ZP/kwWOwIA8n0mQApEPFbmfuIDDxWwLH0r1sfxvgX9m9T1a7rlrSM
1MsR01HcRTrIdsjGDrfCwwlMY8kIQIGvFkOgK3Ex4SK9CKV8gi05ZIPnhZlZeWymbnVsA4J4Plrh
peM62hXOGYwlq3UN0pX7NBj0PlpMwOqLzELFdMs+3UHiScieL1FESxeGNp5ao35mTLsWB9ZoDMDA
3kCxovj+SjCsqeC5yAfaPytViZT9pxzEC9HWtZ/aqo0Ye/8W36pkN899XRldYFwK83PcDHALETEQ
k3UrKXgZZUOtfybDwo64vGfD8Ui090wo7QWZny7IjEfpwrNscqwdAr3Vm8t+yk/wfSLMc30QQiMi
zhxHKLuK+mTuA9CcS5aMq74U4jUICO6SDbX9GFNKVS274zgJV/TEUKFFiXWyHlD1f75JEBSggN7z
HRNYjocSfwpw8qlcb7fu3Jf3jo67dH5CmAweKacc3KWuS4ILi1Dzv+DlGL2Zxk94Z6v4bkt/V9d7
1yYBVsXnCZMdec57J16WSVMOzm4YEqUyAQeu4xjTfPZY5fAP2gAE/zmAnYjQp9gd4qi53afRfZPe
Ql1uWRTSWlH5zgo8Os8q2haZ4oOihirHjp0ZI2P55OLN3Z6BfIpZ/p/hsSzv6EcdfSXhkdZuX5D+
UAtN2pRNlj2djE2vlQBJmmIqRAxpHNuVkCWx7jt518OHledrsjwELI1LxIHijCK2+5+YYr60K4nK
E8nS+iEww+2jJhvQl2Vr2u2iPgD9PlDvzWNZlZnyOIcn7MxXCZzKK3RrXIVTeWHwejJ2PXPbew0y
MW9F0388g0CPcajulzDn58hmmc/WXOp4fy6/AtZ9TWpYpZLodKPiS51z/FYTOjjlQc2AAT9HfypT
HYvbDkATyXsVX30sYjfwAWdo2AWBsCOJbxw8+wMA2phbqRAGqAY4lNpFfjMv9VoYobjVp1qGzO1M
opbIq0jrj74vAPF5gjCCeqh3d7VNh9wwH43FHe1OkyqJhXw2NFtyx6DGAcbYbnh8+jTYVcVWYS72
onH4HhginQWUVR6VXxr1nSu5td5K+wz1VEiZbq8DcRnuljB24kCOgCnPOsjjQgx7xwqhBtcoRE7K
8gWmETLD50V3kyoDyKJ2r7P6fvlz/4OjiSuP8+G8OvGNd8MR1FxQNYR/RKOCCxX8ItbrngHHQx0R
35I8utRjF/hFl3Tf0ULuV6QZ1uRyoV+Dy1Ownan+xBkcrREGq5YZoDOxdDNapBz+g5UVXXIHCQbZ
anOQF2k0plSrzaYit+ONlK6zzBJUg+bIO2EBVVDfBEarXG4CaEB1w+sAuPutJS+5ADrHlN5qYH5W
59bvoNu0KHQcydknKXqRSAy2xGhERpQuDJ9rcJsr4KNjAB9GU/Bhyj4nqzmDrt/QOArv9OCXhRKg
BnkCbxMV8mHy9CmsmbDc9aVojge+2YsTLI2oxSn4zbDgR+HIXFikoNCok5WJBJjd6cf+D7uzKnpI
LuhvmE+gSVmcP1rtGdhWkXAI2RFEYC2uR3rqpDA7Nvrv+LaHomuZkE0K4hH+fKgprBtbVYoMf6QX
XTMbWs499CjKV0cCcid+n7O0RbrIvtIZIejlWNsfZZ+yzjxu5oektxXAaycPCutzjJ1eYEKcDGm5
BU4MMzS9WT5H1VtkYHutto6824qcDK503s4dPllf3Y/3O1lUVi8e7R5bxKmEnoraJF3D86jj7xZx
Z997BmfVLNRjRFHCYGrLvkBS82uD0yOYGOcXYxLCWUaPrk3nK6dWb4WqBa15TqdfyhvKqtzeDs4u
ytx13DF1VW6qOnRb3QZQwq221kntJE8fg+q6g0ZgfWzaX2N9JymYE2L27b12+bBpeBR8AkyQRRpn
+pPCmrtCDFeuk/5eLbaRVjVgN73xkSVbnvH36w2m7PWjyHcrekXdTf7eLlrBYgXdPn4gyP3WsmNG
JdL2gq7KuksAoaRUlwuATt8+Fd1ain7YC2g+Votlwg812gyJwlkrWCaTNVjS9diDhGt9QDtFhiGG
ExHhLJYr0hlLmn8Djzt15KypHfkRaXhDv8GewqdH1kaHPLp7rB46FUi3JRpwgeSRAPam68NO0Xbm
/m4FrPpmmOPG2OE/1VLzUWvhffWFqqsunm6uxPUwss12bPUO/ixoC99avRagUVqRLYSOYOQYssFH
qxGqy2c6318OPKozL6jQ2xiV/zPe7TJUJC0AVeAEM4xXD6IH91eiQ75EjJ5Zt5jrIdSkJtn0IxdZ
rUNl+nSBwmqE98aQepTIfVaQ65Czirc6YB34poG4cyfPFS8m2Rjbms9MWhTy78w9KARevnNv+qif
D7Qi7if6DpWCgVihskaPrklGyWX/wZiYpeuy4y0jfYphUlM0Cr8v761dKH4ij4HDVcHuXPqR01cv
6QudctiAybxznHDemmS6YX+x9BFESYiCARSX6HIul/jwxZHTD7RAU8D005+TTnon6ZqL93IBpdvl
YXveeOLndEnwjX/yVyhr65A1bNB7Mp5Ei7kJ09DQRFNWmO8BTsEisxn3FNhejC3KICPEx3YhKza3
WwTTI00Nz37mFdiK/NEVLRWx8eDVVoXKrtJ3KEDipCn7YymKrBk31xue2d2HBFbA2dQoxwtRDbtv
RA4x4L7WGkSoLRcRjgLDU8u019euqmgdOSgK4Njk8Ubpug+P/8DgrRg7/5NPBKCx26unnpP9gTE6
202LDbds3P2GZCuD4haFgsIqTErFAjFEqiq8gu25TCcGtlTYibsxBiwpTuL0RQVPKXZqaxb2yqi8
fq4pgdxGpqmmgyhkypoSyYPUhSqoxqgZHre7y/imDu96tkTffUCHStdaMheX9z8wwfnUYm8vlk4d
8zzDvsq45R1p3CxAauhmyOrH1mA/x2HbOE3NavMiwODWfxllRHtYxGTXNShpMuKqZPA2j00grP/G
2lHqHEZ5y3u2mIzmiyEktRPrt+wI+kBQglz5mjHNPrIX+Zn1gw9CUglkgREEtcpJ4Z0qGV2kGUqL
vqPIUh+qTFKTJe5/sFVm72tffpHkFyJ94xpgiByYISqeKO+rEqxbc5fO2wk1lAwwf9EF7ABbk+Ed
RPGPgu4sHeIuB+hFUQw5optGyfnmzP7DDFRXKRcKWxbVxTn3VncCrbv9mbfdX3KxVauyH31TLJZW
2gLKiwnaEK+e6cPClHFiTGIAgwLxtYbUpmZXSjn2fBidhBpVkshJl111Ek0gjRuMLaNLGAsRCUjL
5/+MVvuoFnJxmCMmAn9LJ/f2h3aiKbVHlWidCzGEaZdEIJJb3y2U4MlfaxXSYaqAq+cOXcPJKxkP
SwSjC4/6tN9+iORnB3dkFrHiO5qlJF88jmqCF3J0AZAPZYuesZtGRKOn2JXi8wGKCfTD/C9DmaFk
Vr0MF1dFt11C3I1zFDyAnIt+Nuf5C5a/ICRs2xm7L9gln0TfRLINihZnL+qqh4CG5si0vXvhEg/4
OJ0EN82BB9B/tvqCBcHVQZqheguHwfIaypTq6ccFawmeoWX0NeWG08ZDtTQaxAR/XuRylStINoZc
WrYmcswRH67BJAiqNHxCkmNIuY2uLP3QjVG7CJOSy/LO8F/fxQunrS/ISkz5lQOHZMlggbmSMuMl
kkDE0DOC90NHiAOg2uM/KkOg+7cxmp5mdS/oy5KNbc4QcaxBdT6w9phe56Ql1Fw4iosxdUB85xKp
AaqiRpa2vFiChWP4QPOKVoZXMzS4r5s3O7EByBYzd1cSiz1kxbElXM5DS0f2qgiCE/vRzaNr+cUg
UWk2Dml3s5hJIHl7UwGl+RlIdoKdyoWEYBo8DEBBgMBsRdpWBWTdCVobTcqofjIGOKu0p73/i3LU
0Q5UXnSFO36+fy4bsaq8uzouUOplzlnSMnt6KjLjJju9fdOURRc2RalTOOSgydNWVReF74TSJY7+
LISQDgViFF9gNbTxex6sGsu54Xj2unj5uJYp8DShyMtoRZsYJvl2WWMHN2jBrIrQKnx/EJYqieUK
y6i0euM8qnoRpjdY7nei2MlAGEW/PaF1KPUGckKyMuuK2tS7KfVEun+n0KG7ZVV6uzbWdihfIfCv
m7Ep9revy/1FyEhu5VIK/WxWtlxtHdl1AUuOa24ux8mHvTYlFVuzPXoVB5ozC1Cr50rX8qlJQwKY
apuMPcRab7XhotVwFwFK+dqsOBrNksHLo5VdpYXZ4aTwdSeatHnZoknSWzxa0HpPFZkOslKYJAbx
syRkMeoFX0saf7zn4X4hapmv5QfwYPht76APtBGldgKXbJG5V7sfwpx9gg0fr1gGw36VxOvfz6xB
uLU8sV59MTBETCfKaAqf9c1ui0MEo4KuphUwPIbFeZ0TqYthZ13mtUxEjg9iqD7MvYC7oVW67aqK
K/pxzd+BpoLwlmAHpiRxZymddaid+q+keZaY7+gphynhj/NUnGdfWQSwlz3rsB7yCKu+PT3ukntC
zkQ2mpz03gUDsHwQAIpz89WUTTTyRb1ha5LBRXwrsZ4xRAbO3MM1XsasHvvP69dCxZF/Ypx/T5X5
7skiH/llhLgqgBFswr+g5uX4KKe3UstZMHVIFbAdli6Ui8bJSUr2jz7eeb/6KxrFjjA6jGi3om4k
rDQreiOTvC3jTk4sNKosXiWXRxdU5khKOGLOPPicnXr3d/JSa7tsm9zcStmfaORVJL1vtd+1iw9X
3Mo+fCIX07mAFaF92HMf7ZsT7iNzMLXBt6hrU8KVVKcQ6e8fuSggH+d1qKME/BcEZE70RomU69Zq
pFEShsFCRn5oglBWwOnP+R7Dcg2crTPN6z645QW55zsRobUDjngojUJaIGG7IO1vlLlsu/DAwKSJ
2HpH6gDU3xiZDcoHyZQnJhu4qfWK3BA4fo6bB3jGjvVRM7XY6oPFW17k6wJz2a4vlQ30BcPpkVXk
57g8wpjtwHFwezLJawzq9NEZWiVJF6opS7JZqxV+06UnQzKEnXk/xk+fXI4aDwLjg1THAfwZyyCI
dCI9/OyNoUVvy3u5sV5ItMvuBzov7RjO4QKlnAncDV6EFVvJaYAQH0kq4NfCpvxS4H+l0eE2+gF9
JzmsdLzS1cvUPuUZniEcW3VNojKu9vu7CjwTmPX6+b0E6dgDBYzs1H7Gg8TJFgn0M2A6TuSo+Po6
dxQfadptVoQ0VPlsQSX/fN9opOcunlMrKMW6/ukejdEnMCMKrPQZwmBsMU+S8ZDX2dtowWIB9SYG
YRhEFpSpbCtE5VNZwHt6FnZyOJRgISzU0aFSSZTDqyXHS0Ok3Zu6TaP9UqyWU4o6EUOM8xhqVRS4
0eI0zAMHfh0TKEXu1sLkRm2I4nxEx90ItnmqmfVFspEJu1Ee5YAGRXrH/AwuRlv+zZRtw/X+ZnQz
Lcg/DD5wXamfrlr+AsU6EkRgjbdoGxgWUW7wfGTQHQqaToXlYD9R2yIS1dYXdKvAP44t/gGloBXv
HHxN3XKaH5SCG+mFHLxBdgZpdbSFzYwnit68Pws6DBMjh4kFhSjhJFxsXjvUulpBW4VPH7xyuv0f
qE2j2R9E+t98rcStPu5wetqke1/ScUn3Rg/w1YapGxj/J7PeDwejEe6hyfrFreR0mdWSYuNp1/WP
tV8Km5qCsY1C7O2WIGydhfyolNkNiifwRkvQ5DgxOc+1fK4AR5rYhaxu1SGF5Zqfkw/tDCdlFGWI
sKMAkmFVosSZSkUbHXGq+ooFSO14qaKQrRI5rjyHV/OP0++GKNCLLaQ5RWaTjAAgXyBvntOtDhF2
SDAMj+XieaH7hnWU+OwARMbccO9hEkTnKEsIRl6nnif+wMmsJXLq+W6rfQ+kpERha8T4hu+USn55
n37ANguW51vNX6Ma9EJj/tVtEtfUixc1UgsbxlkO6o44zOfA5cXRwB6NA+vz/JLcW9qQj6EwzJqc
J3Mj/KJGKgZ8D40kwl+YMBltXTO2AhYk38qYZf5MBH9vytQ8lF4W68klXeiqSCcKijKawJHlhfLV
0JzAT9EcYdmf63xXPLpCc5AInwq1cjcKII6iBbbRS1DVz9AisnoFi1U6o2GQj59+1MYzBu2GuYUf
gQdkgFguSq7wScTP7Mk9vreGUAO3HSi2t7wKCwq883dSbaARD+FiqqF9LTe36x18IKWoNFTp0Gbd
brJEwzOtM3nYoLm3/HhNynC5sOxTSeazvSFkqv/Ncyr/WE8v3QJ1BfzeyinqJaaQL4SgMvO5oGe0
+nIWLoleyM+ets2AKwQBiCC89sAfGMEDceSwF46vgpD3sykH/cT2si5k9gimpMueIu0JoqY5zPHE
zqBmqmKPR25DLKCepm7cIYO9gaA1yr9W7xEFG3cc9k+fcQfkyqE5UOBoLVVVl7CWwNQLG7tdFfSJ
x2cV8SegO3luk2XTRA+OoBfmyRfYuu+vU7yB6iTWMO7wJtTgMC0soVhLvM6A+NlgAJzr9CbHKAwm
h1MFMsQVsACVtcR6feyHVe2G6sOory3EH/KcH8Xeoeb7gdtWTvLGtgcv+jB/5jxrsdMftqaFz9CD
xmRqeM4mOl7qRWv1dbCFj70RHQ9KRAB64bItDUp3/s9CWJWJzyDEXC7C7ErttBfayqsn5jfkzI6h
ydRu3V3r5nUclTNZ99CBgNKIFKKzUVxlvy6H6oRtyXrZCbZ8miZ8MOo9H06E0bLk8ZwTqkmt8GBY
UJEXzqSoiBtq1gKBn5X8C+2PvWGSVDfJyISsekSFNbWhHjpbk0vf+XLks4mzxVHWoUa7o9lvQLfu
I+6tpNwoyBBCBqZvLQknZmX7fmzUXuqbr4MBmEGy4uoW66KBRlu9Q+4XFm5ImeFlyD1gL2FCmFqz
e44zzEjFUMnqFLN27lPvaPSvcJVFEGgASpelpOanBDPPypmeHQ1QLqU/9Z+f1tgYhonZ5aewRfIQ
oTXHD92mRSgIV1nfoE3p5b8JLL4nzx28szWDRbk1CbGx4+VMVgzXIlkK56ZXJ+/TJsYRGv5fzirI
9zIF3/iq7qSt6CNd2tONMGlg33ZYBzPm4Iwy9A57hLb460MuwyodhIEdn90u397k21MO8UyMd3Mk
RmDXZrDJuwOsE6i3DIkVVaUMmHIPygPPS9hE4sb+9nwgxAxhdmo1iBW6FKgYMFvupO3ah5K2xoiT
ijZfhbUsDMpHdHVRtw6ih60KSY+EepRVzUVjJZUqsUb5QvpD/zKFFaBco8IuYMqLveC1vvEufdf9
iqWVH1G8MhD8rpB6rUW+AUkKY/hpTu1t4Qc90oGs55tTdSbYMHGbt5XVkg4dPQ++YK8uS1K8qzMf
eb2JpV2LKk0yLzDUblgcBAlSEB3ftQfwoSyvBn11/+jMeMYoJPCukhFJVWEQCvLmmJYDmW2ivRAE
yp45puJHhAjnG20VoWyTPaHkzkC94xqiUqjnq9Gm0r8qOLsue0A1EyPReuzeKGSw5fc2CW5nKEMK
7xS/qVv+hMTDl4kzWHsThMBOhdc7ZXeJRrdmnHgPc8jY9Fg1+KsrZ1ILi0QJt5ahdznF07yfrrmB
YLazYBw6Thx2KsnAOzPoYq+tnWWvsXh+YpqUd+c+uYy4txl3xUAokTi85UrXIjQrPH0EAi48dvNv
hrecGfnJTasU9TdJIRp+3joCaaEQUXc3TJUnlCL+U9H7W3IaqFMPaqYxPG3gEWSjN0WVJEifqx6U
aE5cDaKC2fKDFxV5x+pMCXfIQ7b5c2QjHBf5/IrRVTXCgyIaeCpvtHvQp2UEBpyKkzw95yUbp3QK
3Rrw6M8wDFnLp1PrV+JcyRpQ5Bt8GkyexlyHtDwlqeEZZ/OCo0iSbWEC/SCg1m5+7h6kQKXHWRC8
oZ5YDOogSRgN4lZVZcRwedZMAyd6+zhHVXRqAuwRj+HHbOOl/O/zRUuDLsyhJDHN8rATMbTtg6wz
ZDi/ZvmiRUKNu/K638t9XsI6YN5TjO0CXuNUJX81Jp6zcduAWW5ifQ9uvwRvexr9fqyxdDwZfn5I
v/fIY7/RdVNjXbW2lbYCPjfeDWyqPXWd43Z3zmSYlOSkVfP0BF0JfDSppg9FeykWft1jWBvH6Cw8
qgVAWr6ZWD9bL4TK63QLQJGQ+C2qGe4yELezxxpsO2+qJKdPeYTKL7B+Vb/zN+M+P4JPkm/0XTLU
N0tn8JqmT7069R9q52sq7KcpNVTd15Nkpfn69oIdKTpUhRovUCe/vx78eg3bXOmwGhTyAppDLxSJ
XhnXuaSqxDsDsRnFEdh5ZNvzi56+/k0MUoEVKt3cfFkEOKuWc8sRxTjbNx8usAOcJ4HOhR61YeqH
juTwq8WtiHIQaor+WYLKd837gyLrdXEVoBO0XQGBZ5YiFl6h7FRmC1SJDf6KZXbe60Sc3sRLfxER
Y+ROg2p2dF1lq8w21O3sDB8ivo4jOBLWdzZCzWRpnXTUmI7tnxXU9WptzpKnkOCXjaOZ3sdzqJG1
nmF6yHLpc0djMpAc534dNdJ0Y4Z6gslYhmpncr6Quc9q0i7t+7q0wesyzPhaiQzBF/cAi0CZVU5W
3kc1NONoT1OxgQxvzhgd1y14PDnPqCOi65ggUHpmuy8edV6wgyG5MSn4Fii+4RWrcxo3CDByw++n
YwQMWics9AmHQfP5D594SjhpZIWhsbs/gEUtpf/NuwjHmjxfXlIjZkyPjFUfzzD0UT6YZiG3Upcc
LACe9LIaPWBt1iYSpdTlBKZQQKHJKt7+b022or8aHOEnC9zdvms11NodPExdw4c9XLLDh0BOjgbL
uIFK6ZLjwtUxr5z0c/OR3YUHjMb5uLN3BuHfio5eMG//QmMLjYlb3WoNl8szYC7uAGMvjt7XjW7d
LCUHvFw6OCyyDg36Usty0bwaYkv2+MzMXOyvmFF+XdfMyZoFkoOm1915jTCSGhTBOh1rrdvoEu8M
qkMaJ31vPKqCtTd9+OuhyL0XoHds4zUwVPi5GAYXqvO0XXGb0q3BO0HHIL9m2vMtsDo7oqxNyDk/
8hBXd8RjNkSyrMavwtOkGN5eOdBOco/K0IUF2C+dU4t8Xw6yEtDxNtomEu15YDzhYkoPbpp0B8Vo
8qoxDQhD4fHum3cJtLiq219vhxHCCKpDvWQU/WjASDKgti4YCXYfDCasxpjKU4xadB49Jd4EONyj
Tbq6EPaO23sRZonrlNfcvvG6fU7MrQJqwPYABjvnl+9YI4VLql01NcV3L0v7QtDfnwkhJiNxJU+1
ZRB5K2EZuZaw/TdiNKA/OmJvnd86pgFJLGYqKU9sfCCRvO+9A5KyCAGml3toR2qqpXiIPymG1RZs
nIGopvtRG+7o8RLKzYVh5Oj+fxXRCWIfv4vbcU25PKstEp6oHHWh4OdLWECKoxVGfNgfbncJqoTS
HqVxIk3udTCwdh/B+vGxUOPBjhf/g1xXE0VqllqVlowchn7iPY0drmGfi+FqcDxxiP3oOykgiODP
ukZRx2ywJTjtjvSob+bOoQ4O3yFmdnWFD/at0olByd9zGgbxYjrU3Md2R3Jyk2Qa3Gu1NqgvLN9e
tuzRbPKhLd6KReGfGre82LTVkznQ4NLqN0gr9Xicn1/sn9iBDvdjsutJIuOY56aPDWgxLCfrq7tX
7UnwZrT5Mp4FeTwWYBP5e47DjtFsm45gnjD1Ig3R8PAf8lEC3pRYWOb4C/dqE0EufTkITH/dhhtX
EvSF9OPj6NeJTOF+Tcp2HTHrkkB6j68P4VaZhVbZHdhzSYU2qVbukyZfU8XbaqEgEmVkB1IB1pwg
IWypsWEMPxXB9tffVK5W8jK6nAwJN+0qcO6FPVmcv3+14zNhvkhd52Vz1LOPyvNPWKA3R0FgIi1e
0m4zZc0pSXI/jdjPXrnAaPCv1q3Us7J5F37l5BKnpDl8hfRkMpT8IYZkGQt1GExjaZAQlwj/Al1M
roYhARTnbdMqbYz0eF55eqQbm/QlfF/S+Vly5QXreC1NWH8P0hMCA0skd/CJDKJigcn1ShUzSPLx
TtkS15NAy+ymTu8PvQd3REVvJjmNyL2r7qdM6R/gKjhD0dJVUAABgJ2buLso0ZdgPBo7jxeQbcsY
bkO98oyFQrtffVD20cxTjYMy15Dk2yoiWexUi/Bwa5itL+B1ifLcS8A9j1Kr8tDi1gCBnRVrYgIK
Vqre/exAFOxh8lRKulDRyKipAK6Eye5+1ifiFk3YlXDTCAukZGlVXdkxiBlec5M84HKCKS8JkYS/
Rt2XobkObrZm4xDnp7UmJeDj1r3+uY5CYobcE0Yc7J4J2e0hzIixJX1wkAcOfc49ZZjWXSjVcsy+
I4eZETncql9wrfYk1wb35kcMD6sOcdvq8GTAF30BMQ1lKqa5Xwo7x0G0pMjh/ivI8gO2XcvK6wX1
z0iamo9Ly2tdRxhsQI88O5iC/FDWKWZlj/MokTjxC+PdOz/RV85qE1FnxS7gaVs7y1eqqg2HyJ49
tkjfPIzlHMnu+5k5hZ4Clzmyvz9JmD2dpqBR9hRcgAnAx07sSJyMvn3sYHVshZJyMTAH6SfUjeB6
lVmWFByxsawAxthz8PaSBZN2BdfZRYAePpgmiOwTtYvM8N4MnuPzANStd7ZVX0p7G5vzlzTEcmmm
Q1ThuEXGx2RhE4EfswEEsTAIIKF5+jkWYb3al76juQbYeBGek5HvrB2uRdprM1wlDiOt4pIg+syu
JlvxI+Y9EY2zWJz45mSYCMZaGU1auFWj88Dp4YLhQsf1m3JEKKKkE9dkRF114yTKuygKWhScya7W
N6UFyXlIWsJuRlydVGaVnkPKN9PSFr0LwtV124SpvNlii26SJxucb8VWqNkXIwp7lgQnM748kscF
0qIu7IJep7kNTyvD5dWDL/xCvQKJ8HmrzFagk4WR24iUroTx5PIr5eC0k+Df21Bsosb4G7Ol4mem
jKd3yCScFVLwCLpG4egcze4w1TnFEHNhjpdHyVuYOOqogM124+A8YrL/11aXJ9EUTBSDtftTBO0A
5CPv3EokhMaP/Lb+QAH1sg1nmCZA3VsunsE2uKp7e1yansoecHhiIr5oTLzh8jYn6ocoQiwLju+y
YuUSitSEAojfm19oq96kbs4pWPN7DqackEmRN7u3mU86kb8jS623mk6SIy6x+huk7jgk7HecIFx3
kdapbL4df3Eh0Psyt9CCCZULMhR31R0Y93yWT9nzmnewXFPcNjtMBdvOyWDZm+0QOr50QwniFnKW
mgGnM+pzmNM0DLu2VsY4tZP7/11fLs2j2rdZFFWpp0aPIx/vnwoPAfCq0ZCYpWLzYoLFAnfFLfm9
nhzzosJKyAG4dHsw+gGowqc3buw0HdklCMXWHj/zRc6gKmoxhzQS7p9l49iAPV43vHyJPf26gPKT
pvDZ+PDMme1l6l5Ji6LNyKp2KlQO8+9vJTsMCGe9ygyTNdnmPxwmjRRiVBuHOwvi2k5gkJPme1FH
93209hqr4o+vtMV2e1Q1vQeZ6inrd/ubqBS460cXT3ixcEsVXMzn/YCXn2+LEPM44eBfOzsqdj0S
EGor3ouT9nj6GN2RLWzOuJ2yoJW5HQ9eShb/AyihBj+58li5eM2zlhLjXRlTWQ37xtSRigqZJDue
Lt3QH4P1e1134NQubZy9laSCzYyKayLO/XIO0G8HWhwrIHkNzKSq0r51nZtbLGW2hW/dR2O48Z0+
LXIziKzieuIgCUexzzVlQ0KgXq1uHH5U4wfN/5HzdEmjwaTlAc94AKkQFoTpuGPYO7N6ObBceK16
hYckcY2W2SB6CedGknK5eXx+8i2au59lbKToLN8ecCOuFPU7WLacOZqRUu1cl9HqiAMxXnDEAYFn
ZE49s3t8EqBhCxDl4ai8vXJwoKAa2eXWLy/0egE/MCFay+4PJlz4oOz2OtYqGVVGqUa5ynuj6G2W
fgxJKSIAsGjba82yK0t+NWiw9Td0qmn5xIBg90b7uz5GamFS7i387XcXRwC2I3koPKFj0Oy6yeHG
rYLNLJWYiVB5nilovtaffB7goVgV8FWgfCgJpVs4dFjg2DTgmLc5UK//SB2SwREsdyyF52xj7vnS
zi6gRcEyOzN6Nk5CRTfdaxNvyNjnEjcdrMjI+c1xavro+WjWpasHjoQr1Uk4j6FFe6MQd/Lb4yn7
twRm6H8hAmhF2bSb3lGfOHvY5cFXvaxKupRUsayBCpAoWeTFEUgco/2nDvibBbiWNnaSxF0ckvpM
Bu/zsNVBM8GCGBIkhaDCoKZxyQd1daULJD0M626rFoYIT4Qr1sYotUfHtI06XOgDonAmLOV1OBHp
DcUWZuLGGQSW8hl4nIkfFcUioyHJU2PIiQfKriQqPrJ0pTfnsrZwFkaIPFUbgZGkoDTWk5xB5YoM
bipyU0pDcgco6AJvO5dplHCpQbthOkMmWHXAOEV03DmAssBfDZ3RY6uy0yfU15TcEgSRrioXbFFZ
bXEF2iF9iqYIQ91FOuMFQ1QAU+U8NSxiABKYL/TsjYGE/1GrNVocNH5Ec+Jjvqk7FtiQXqJYhFhy
k6fixb5Vk4k2W/UPmzk1levFVLfZ1dxnalSlLzkiiD57J9x65mke/WLM4wBRnaKEImzKrgbWllpK
9pxp0GOe8q6ObDUg4x6kDSD6Dad7s4mr+4yNlNowxf1zSMB1FBiAoVAq1mIlhmHttNc87o21uLgl
FCFpkub83p9VgBx7fR0xc22I/CihbHd3ms3az1I74oMaverH34f80w66Mf8g1LAiCjxuQ0fKCm0P
9/njD9iuciSf/uudTEQWSM75IoSpFoxKJY9x1QtrmsM5ZQAln2U+7e1JeqDrjtOV21tIdMpvO02G
HRzKW/hbFtVWNnddcc7+JmMUXyy4WqyQpU4kETv3C0SrVa3LkJnIxkKhi68XbkK5w4DnN8cQxonz
efSQlp+qiv4FNXYvN/a2NtrQaddcFzLV9kFOa0i5evN66T10kNaTA7ntX7n1tNGCCTWL++ZY7hvd
RcBPW+rdSzMLEDEbyI0+hHntQ1eXbmQrZjgBfpreihCuvKMihZ/cLZAx2943irOIJTRIb8kbrlp4
E+3ALvsfpvGTNEZLAUyb9FP6IqJCrzzu1k7JSHMObMN4hGRG8KheDlLbEWojvD22OCRVS9qxfNyb
GNK7oByAIQineXliwFHrFp2gApCohYZMwwTdPoAperpqpDpSBpQKhnguPbfrOjUCzbEZjsorlv/C
NVb5vEoJFAjR3WKJtuRh9An8BELphRlGh7j6+CTzWzh/qH1gZSyPA8eujSuBIkt95yG2i+SfRzCC
s3qTIbCUmxnbQYcPZsCDdhSWAqD+uIgHLn3EMhxJTIiVbSJk/430lN6J3cpuv8akWUsk0K8TWHbA
m6vDnkzuD/4K+6VAID3qtQa6iId0Ew8C/WtJ2jiXVrqeUpmPejlwZcU4YZHwAwhf5iQyZFKc29XU
0CgrUbautBIXTDwWYpFVxg/+uKMQlX3GwRjCrSBoT2gCEwGkIEj9Uagei8uL4YCIifu2jvPOHQr4
b/JNo+SXaKtcmM3VdszqTGuLHiDZc21Y5LVaYILS/1gb6E4tYdJCeOEJh6FmE+FzKF+Wewy7K2Tv
rimnSIafKx6Ir5qx7FKWVrFCHZL5Cg/g+0g4arGVzQEY1DKvm8WFVSO4vq/Qfcp2Xf6CViRt4y7H
ifXFBg6bgSYnBpljnFfob3/P4SDmihpyMWYERByHFvP8KvbKmFH0xV8IbCwMQLCtXjycvzAAmJzK
AN6wlj+QQPNkTy/iJ64TOHi6vUq6XkLMR1nRAT5/hy6G5ZrJePaVpVXoP3AmLS2RKgY9ut0k0EJK
Xg5zwbRm8zJdsrMUfUpC9CSEkuC/1HkBTf44BPP72WGVx2sOcFtxbcJDqL3GQfuJsPsrwdJiFQsc
g85RB8Qig9mynnn1ozhqm+SBk6qxt+QAcBLWbnFv32SR5mWpn3BG2gCDHdtJm1KLMBDeciGLzd6X
MzBWj6YBWsXOxks7APx+snqXJI4bqOV63TJcu9JHaHXSLpmBeOJ9S+mLhdKieCZxapdqXftWGllU
7kOLSQJdxtAjwlXI8JPTqAI/2c7mm1xRb7/+thRjT+C5DiS8baBEzXMxWXDYcrV6vtuYUDZ/EPMD
1P9ZUGVQ5hbQQIZBLtRrpCzcviKxF2ngXQ+Z3hdONPVr2mMVevdG0VNCKeEd/ONKgT+eJ9Fy0y29
NMPck9NpN2qZ5LCQHDwmlTzelSfflSiKumBOQZ3qEUbUZESNlGwVgFPUHGDlZwWMuzxIj7uYO0UW
Wa/uyOgZlEcOOeIYKoTt3E5nPWWPgqA6/CZW0Pk2J7GQXjR1DwreN9D2ch5ckpEHfJTquTlxOwpy
vlXI7oqcA4QM1B/F67IL8vxt/GqztTNoRgjPpb0wiiAPB7oykKw4VemyMO5SVCnsmrkN8Hbj5IO5
orXg8NAiq9UjpPgIEDpvX2i6h08DCqcqFlhHCxF9+2V17fLVvWNvH/rLPs0pB4askbh4U0Mfx9X6
BAhTZZvh5pt9WMnbYlNHo4jySzU6KAYpv2qEEHF3r/oUPGklW02XKe4TdRLxEl2Rsd9wTnDjxjON
DmoyphpkZ/9cuIabsF67i7bi6Lr6CNd6lCCPKCQOZORwJAzpp6/J2XMmfsvUMT4qUoZ67lHHTTi3
TNu6lMjmYIgWNCqfGXNrxEWYdPnpK/SiZmdTSvQqp9v4690yXNv93BbtBiLKcB8KCSYmaS7huCP4
SeOZ1I+Vab/ICQ8emDMXBak6D6xe6/vc75Z8xP/EcJJz1FrtRYAoi+0zytWVCd+FX+FDftSTnuCD
zBLBCtBsgREj9+/Y6i6pNtQukHxwFq96Y2fES+d0pEzVhElEGh/U97r8RpQXb+Vl6LuulomncekJ
l07Xsr2STQ6dmlm8UmHVoA9gCpbPrRcdJSAgtM7XuzPrVGo3nbMG54z9WeEJDJnycUW9lbCf+2x/
DwAJjdTNJ+wlJYaOo5YO2eMDpjolCM5j/Lk5JWVer14bVQYsvNEssdEupABA3adBe5wu+C9e04fJ
mgD21ZgG8jYvCLI8CLeCEk4Iqk9aUqGh5H7MtJ1Ko8ipzrEOPe9j1p9r1rKyn8LHO6fJVZz0ltty
143VVWVX6HEvlnEZ8Kt2nhj/T4QcR0sEXD5n8EtIf/4c27WSO+8QTyWxo1WulPgmVzGr/aIIQsJ/
sDVwwNvAJHmmghMSbNpIpTHDm4AeCaYNcOJ/TN027A3ySTcT6pr1h/mr2J/a0fRGUh3ljRGvD2zO
K2HXk6HRuDA192tmA+i0gKgEwrEafLhmp/pl/TjxrK59cmcQlga/BaT5d8j233DsJ1kCB+pzBOdW
3glGRFBYj1rKhQOq9w73RB2WAbV80xGsoAEFHkPj/pEH1v/Izmgk+DN+TOGXs1y+XB2n/lgcAH8Q
sPUpNzuac7TRBa6n9hugZgz7sM4e6mXB3x3fSZ3YlxjswvdauG4+r0IP2dXVudC/hTFnDgPYW1HB
wONZyZzYuYPnlN4QXGrG4pKXL/65IX+cAXdv4/7F60+24IP4IkUmyQTiWfXTWxi35XZnlr6B+AMB
Vpmk0VG4Eq8fDko2XgLWFtPSLcn0knML+yOoV1kTgOzFVMiodJ7YmK2iIqv+bZeTdFWS1sFVRx8M
RZKw2IzkFZP/Px5twRTZMCOQReoKfCxhDGxPogTbaChPsUExCBix/DNfoOkHNZ87vVmGNKDnsVIb
tN74tycWnymg+ig0iyhR7P+4FUYqll151E5EOqvMegW9bdpQk+1LY9MJSvVVXuG9+O7jelkBPVdY
vsBx24zOzORcTuh4bbptn9jgWVhxhazh6/fKTnFtR6mv+0ODJjmkHAg758bcw5dh+vi49K5BkT1g
tobgNmmPelklKP6RztESsNpHHLpmw1MlKFt0yDdP1zQ75fug3NKTKqRG4gOc50xSQnryoKMDU6w7
C+Kwf1SveF4O0YPAPPOMltCWamoVX+ABX4eZcKO1lImd9qH2UErgsd15i1BEcrqS+ZjW+3FFDKQM
Ad7j0dU/H0CzcYemG/IiH1AWBVZX9YeSPiaUAd+pomHwSIK/RiI/Pz7q796vbNfzG2xe4EyIA+Xf
uQJeS/7q1BdbxVM7wkbuphnTdFhMxJ6bfjao9vFqEIOTa1avZb2RWlABw8auA9KbzgbsMnWGBPOW
fEdaYfC35Km5hEHCzmvaFgaZc0752QOUyauIixZXO4w8foxnAEycw2pzlyB1y6Vr9KTxyd9rLLde
b2GD7Hs5Mrlso+bCLNb85UKIVVnVBQZBgQhzQHR59cBkqXXXrdw/ekgLJZJ9ODuXce2ZSCelE24d
xIbPJzsXQsoGv9boD/+o2G4mYbvgSOh9ZG3APYfUMYiXPa2XRUl1IJvuEJ4hpexRAXw+7PkINoN2
GFsp59BghGvliYi1lJWrUaNOIF5194TZty3u/LsMZYHDBMuZEjM82w6E7iV4Ob8pQNhVnQkZtGV1
XMFRL29zo3gjhgm8wtlX4jXGgzBNM5vnn/t3upRV5dUNK/X56WgTZ5lr0UEK5PiBE4gwrVgd16+5
u5xVGLyOEXj3IB5wkuaeJc8TprNfYrrbMREv7Z3tv3v08eet+vL5kDBpFvXiRb9vtzK1GUsw7q+o
4XpIhjWcORlSwrU8oNgwyyk3ByQhyK+q/UbsR42usuFEXHcfezK2r1mFRGWtxDsKq4aHV49ZX7YZ
ZXokkq1Z5Ump+VljxUozZgTRQOUFVh3Y5DO8O3+UvUYRY82AJlXgk4NSWyujgzm1TDlIn95n0wBA
N+5cFF/D6LW1t1uPLtEIk7mJJnAAOgsj5NCfr6Ju848myr6sU2eh2gc7K+3/DeJl5ykJoDJABbpX
7OuZnKaBwiy8eyIPSDqo84Moz5y7pgNa2rcbYVVMkDSkCH9y0KeMwqNnTVOPQGcqluwzxWnwd7QM
BSMxfjr+UowjM0q5n1KUWUG2BrQl2Smp7NRd4uWB2etOQUE51fUAALFyiBYXtTkPEWJQza7BaXwP
OD2o7IJjYm+NUsC5N7cMbhJ5flaymYCKPyJf1lvRbQ2FLOjIY4u/Cp/VU+EUqJ6qY1fU0MQfd7Iv
OVfllUKHmKl2+OrVCqvQG2kfO5lkz3ZzzDHO7ZpRKWtGUK2VFoWsj24MohOFbr7rRrwOUScW7OcG
B5pjO/DXLIaGO/yuiyXtYU+7zcSF95xABXkx6NWo3q1UOesuiCgYvGJUvqai14MK1dMz9/NIIw7y
DBcBgUwUIh7taEkd2yPznYCRzWdEPQHmMSvNp2/lwEyqrHiUhKrpsJg8yvG9m2PGRJLkg47ZFhMP
qL5okLsx/laVWHVQroG1sVXrs4Ut3rgqUWelf8smMRl8bGh0QFoKXIEUOOobaS+Zzac8m1judIWp
2BG3yVDSEsRfO2UaHu/55Rir+TDjlJPmSmtNjp3r8xLC72RZ7WGekawMzfbBK5ZY+h1+6fa7zP8H
634fC4asZJPxWSjbMM3LviRogw98J/tDhZl3EW1pCR6UePezZnDI40gDC82ikjkUfh2xmGFXN5Lq
lKtaIsIB4lXg41VfWEH+7x+HTdu2a9uhryJRI1TeqeUmL8sfTw7VkeM9DnuUKqByicERQxXHUfOE
EsLqbi4P5naxFAkRUEIRUZ4n4lTCO5y0rzJSN4dGfPl42rs7V2XA8gF/7J4YnGs04vzkOTY6jF0D
Gqc7g39hcuuqVRKfU34FrgtotZTIGCAxKVC+aX4jLlnMRNwYDAQagEDQWq5dvfT1I4EAmjJ3yZcQ
vnQBFZ0YhdU47is35R3HAz0MRj79X4LGz7De2qNdTjve7fYz76oQayPK4TclviAhvD8nD2Iux8RI
NaY0cdgMa5gwMllvzI3XKpecrBVmHxArzlP68YLUfO1+3QPxDSAKr9bq3nN+pKIR+xMM2ZP8ltbD
EVct/0kuonFLa2mNqjtAV2uFcNLtH3eo9prwbK2C54cKHN25tBH+pJFJc7+cRv2pfMtpjJ+97CU7
BVg3hPYTV9Z9YVH0oLY5h3ha0Uofnye4K0bcYQLiTgyvy1ZSiuDyMgaYdh+VLaWNRzWk+dLuA9yl
UyTDFJbgRLQbwrp1p6KvJ5WlH+CW0YT+lEDECWzV8PFCi/E5nxfGOs7w5OeaxAChCvUQPwjIRK1t
3H45xuO1KAJKFvZJvcdaS27h9LQxEPdVNe7AQL7MatMUyTl2k2t4BuNOIpw1b7FWd5j2EKGvwLO1
Ng6Ae13hhv5gaZJ0pMHz8tK9bGMK1STSPkcZwSF+0L3gc01IdBfp3z/kO5M79r39pGnKYfR9tNnH
T+h3oF6GEhTvDsQuahSE55bLtk8mlagNomeujHjUCuJFCABL1VCB+f9Ecc2I8N+FZ+P3psnnLQOz
wOhaXflBIppIVbnXFsUjw39XGWbuVzkHV9lGxV+LsBo4FCkcfjK5MIU403Tlr5DjsZKSz/JTvVZY
MvVIzA05GhLZhwkpsTXuIyJ36UOWxj+4PB9/DnYnSDNy1kA31sKkPARp8TxHzsgP/QaBHVl1BLxt
3g8hhyUFxpzG9ormuGdkUo6236BFZRxTv7sRzFf4mPZShx73IYPnHLTSl4KKU9F0IDC6YDuBwSVM
DXMHJ6c5l0lN+K67Yq5Smff84tP4YqJQe6SfDjHrek/BAAjGuXgEO/zIixqLPg+wpj7SBi6ACwbT
PTnsSZ+vd9B2/LNTgFPB3ATmH9ihfzJ4Zki4DwM9u/HCuOC3o8zxJ182i05xleAH3LniPGJz6jVr
LtXxLtH15LJs7kldCCHUVhvsHzfb7lOJswL74YxPxSQrRqW2wQUDB5S/h90lktkR0zd4rj4Bi045
+ablTiMWtoJPDKwmnyXSNuuI2T+pcpDwsQ1loCAcddy2tU4VqcLGpc9I8mu0sO+pdINbj4GaMqdg
t50LJdb/VqnYGmYwAVgEJxRvAPxmh/lpfLwrXBqd7HYGzUZ486qaUGu3FhfYGYelZA5D8k1Y38up
s/4e/QG8LkRnBlVnuuW2m1Z+r5t4+iHTJ1LEpPzeLRPxQcQlXnzULqd4XmESzbfMlxtaV2qCO5wb
bbxHeQHeD7Nt0MAuB5cozs034KXz+xBu54xN4Ma3S9tjD6zU0IT488l5RjxPkCv23LtMlQekkuPK
jR7cHnMmKrZhJNngXBWH1fP3FgTOPGpkVVcMjfas5X+ETwxL56daCzTyH4Ugald5NXcBcfXo2jdG
7q1/tweH58z8ThFCTt/LR3QLGe0n6stlGx6xAKnudnZ+F4U8iHfQtuP2SIzfj9cP0mWycD/kG/I/
vhxqiKeVihnVBzI1jDI2daAwQ+jYOqLeGdBWpbhlBSbBcvuhOoBmEnFatQQsVZ9CXUkIqJ38F04F
DyEDpFWLWnyZZh/7DD475tHknR6ZmmDOHpMZA5yRoCM/rnNmya4NkwiafUa9vzqVsIoe1eVuB4VX
Nm1iQRoy7r7fhM8ISa7xQB0U0KkCWudsboGMwpum+8bS7HrDHmCQVsx/kxCqHZV3VJdE/d+7BE73
G26l/lEdJRSWn7+j3PC9CTI4lmaV1+9OkTe8EgV500YYRTsz3hbb3pyjhWdP0Rgwyp8t6EAgs5Fd
pA5qK7IDaINMKqO0xz8gKnky1jpav/9PwVNv97xl/zRt4ipYz0Is8c784OcANLPMRcCPgrrXWV9m
7nB4MU3dLi6N/bNlff0vAd60F+FuogMm5Ibn8PPb0w8TiFset+CNMVZ4A29RSJ0+HhlOMlZz1bd6
iZ/elnmnu3ZC+DtIscuSbCAfPkwlFxzQ+bzIf0A+APNsaTgwfie5EJnViziDYxvYMNk4on0QsPIz
E4KKnTgW/k0bMsYvP3PXa8IKu4nT/cN1BJlMOw1xK3ek3tecYLfGrDSAozU502/HC66a4Jsm7J+h
zhb+yE6++v0FR+5VAnPIrUnbTgS1eSq54A+NRZU/73Tp0w7u4ikhitcqyUtJc4Qa5u2bzBQeX63Z
s/DAxjSIbcsZLoXrnxWyBCwJ4lACfk+XAGqmESiahS10ZY3Tv/o/W/FLxfzRyvkujZ1mxI/U5OfI
RLdOkA0Utwdotd61ueYE7w7ltT0QaY+9r7nHcNEyKcizcjRxRWGlmmyCSrcuJfnKnOn1YUttrBz/
KFY2pHqjqDbx1sefACfbiLylWPK342VQxeLHtvjJBpiigOggjO6PyZeJDekOJv7mG+9cWdovtO7C
ujxruVnLzgxfZRwhcFza630N9/dZYFE348dsLZfwYA3okSiQzRWQy4G0lP/MNQ+ygVfwfIe6WF0A
fiwAWIRBGK+iaZlN1oSuB8ufq717btu6cBsFhmfWXiVofEw5iECnXeVDr5jQ8iNBe4QqpmIyM9ax
POO75gPHjQ62gZffIcfYLcDyANfm3VD5HpcCdrS2gPLt98iA/nT6X1Dpwp8drKDzllSannjl+dUu
AC9p0YsvEYNxcvqK6gSYzbEVhG5RzXmk1/GPyF4+Noc0kpRlurgMsK/nJ+FacdWVrZ5jmaTGwdtV
gK7yecSs80QwJg+GcFs3WPvJ+n7J4xF2BF1jGUg6ixttXR4M7IPyONDblv+FAb2xeJfjmrqhKghM
nqWRyf482VLraxn/lCc7EGyrvRjinV/kYGaSqdb3Zr3Qt7p2mThUnsNnyik6C2OkDP1jvFwC73DU
3HR8zF1zFPeyH0No5wRe5rTnG9UshaqJNVOozMkWBpBbxqFkybGolLe92xBI541KDNJL5dKz9Tn6
X5Zwp5LfD2bEpTX5CR/3swlcaBfeJ/dOWsc4ro6tM0ANwAIkihx7V4vv+gzOjtsCrxTnEKRsGaNe
V8tDCOM7nSGe8hbGDc5Be7xIjwun3qAa8e2dJ8h06sjJk4mWC8TCsV6f3ChuDmg2tbimRQXGV2nE
JISaTQjAjxwnvk/QuiTQhilwuatM28/HjC4yE5wpTPNuqKSNSssffek99STMYZyLGVZfpqo0s8RZ
jSXboJTjCJlgaNdXOv675EPAt0JE8kSJavY5KjsdPR0u9+7x3o0sqfVZR+bFKKZk5hOu9rKwsAcM
YguNniFMigRwCJMP4oQobxXSEf1Bknuw7aSi4VrHwmht4lh2DhLXyd13M4Ha5BrT5UW//ZHk4K9j
oIvjFrA8zLO7Xy7eh7e1VVZaNIPwBL+ldY+EMtHqijAg3hMnBtxNblOPkA47xJsmGdvUjzQG3ro1
OsCbVdPfNbfMOhSrmjX4d0DeqObLd+pGNd6bJL9TJmuduv5kC88oLvHUobEZqW97JqZ3t3/gEQy+
222/hfs5lKvEoKCRS8f9jHlbuSuSMTl+112RH8J7rZI0GsNlomxfjwvoEcje+2Suv/5Zc7AjDsDq
21gDxkOakwPYcDV8Uknbp0i5PK49zuEXStefoUs07kR/4x9udzuBPUfGKlWUJq5Vbal35iA/hka1
aGLd+Y1XQVdRmIdGsxeoGZIVoXidrCLtPgJHD+esMGURipcJv0hfQ5XmQZiZBFS58PZjjAfAs3TU
YnRdrUPFlRIbQHGlawz2q/Z4/vXWlQ7u/ppD3wtcRx768Ip6vjhaks6AW6bJlS3yoMDWqV6jm8X5
6p1vWWkGG0cC85h33Gf7bAlkULa+MP8bhPDHZhmhvuHS8PWMHwtUbEhLAURFF5l4S77XdYe+77vE
2gokKr6YJh3Z8v6NXAjt7rDHxapBPX02Njl3qODQh57ofh90Pkp5FL5FvFE1x+l2mbIFD2xhmXl0
6ZIzFulx4SqQ9NztUbSt7SZ3nUBN8BK7c4o+maakALbmWCnmWoX7NvEwVxY38Ex1AH0dgSJSoM5h
9OCBtk2PcbZq3DUQ3T85G2DR9OGnPt+XAKCaM2w4kImGNlqPuRZrmpX/5j6swuPxiGB47xQiJLbv
r7W7WTd31SPQFWig+sXgZXPtoyMjsrz/qNaz+iWYoOvWAdOup0X3GcPpisSJ/BszWBfkSdKq3prh
pm+pl5AEeaQrXPbHUYr2cH/qN3enVzdykzT17OmFV1OscXMkWgMBRwIB31M5aAKzgUZbkuuvoSg5
7fjdwR/CTv1xKkO8wpH6lj1wAv+myc2yNS5mzrEGZVLg/FLQx6+S7Zfd5BK79z8mIcAZj5PFxYc7
hPayh2ciDzXFeyO8ENbkvdY2lhwU/h8sCl1vbYe29wm5SCr1QJswuZJyE5YrUrhDiTS/FNrhS1tJ
5/4fLMFOtk8KyBgj0o80d+t9wry3NRCGGm6aTSCp0iPjFGORy36m9YwpFLba/XXHXPUrGrmqNPTQ
zqcXnBohY3WoNU05wdSr/i/wsJzxa+02VUxLd/fjHfM5BCIqkER9UxcsWavSYT5nhY3Gz4CSrUaM
d8r7s+TVy7V8egu7KyAJOty8L2Xa28EzmPBrzsjfNMBnJGgPcqi4Xs6lulfxrb8O6GYqxxvK4Gba
1M23z3x5v67z+eyuuZVgG2S8LFofEz4M9EBIwNRMzDOW73G4N6TFfQAi4v26GycbRdUHOyjR3lyi
gODPJbG5fgFFam0kXGPDe4W6W5QqwFs+x2qnPy7t8OEikWJeCMVe7C0oXhRhITz4+eFY34b7Opjl
yrs8cv972hrkpIW0yWPR1mJ//uBJX2IJDq0t3w2XIGbM83ZtuO9ZSdRkG6sJAcM+gVmPmdYWh1u6
SLYu9xgxYYvHtcq6vnCFHmgk1sEZKSr+VyuqYwgz6A/j84LIqkY46wn99dSpqv0zcYHWcLV6YllO
A0bDgqEARu3575jn3FoSPqMnP9qj2mYbyM4cMvnwP8C5G+hsY2gGYrjI4Wl4+dCULE8/6kYh1IQv
PYLz7HMYx0x/edd1Cq3oPtD7jlOYfj/VTyXg7BkciLGFcg0rXrUuwWrXIAYVCbaPyvNIl7hL3RLj
lc2sy66gxXDY6AuRmcMdOvaODLy4mmOvIW/lrOXhOIxQ35R7c8w/WmSKlMbSvEIRlIVHPCf0BpUR
8/ftfMAI0AfgqTMWYkfEVB796dlLwECuiY++ZkEy/hmRJptzoGX0r9N6rJ+9UlFIzPXV7bH71YKW
/6xcmJcIOweejTjYLuCy7Zf+GHwD9EP3ZDIPzuXY8/OzTnFHVbQEcYYqqW5gSklDAEX2JQohWXnC
97Xsd3khE4ojpXiWwUPJ2AuOxwDf0HjEGNzLH/CxQYw1n2Sf3eYePEMohXwrR5EzxRjIjRwDU/v8
w8hL0JrvH6M6LtqDKJ0ewoPq2JeS8hkfG5YhrxITbXaNVqHyuvZaVmwm81zHmUD+g/2moexhPhN9
Lq+29NTpD2HbvBoWIASw6P+nuL4ltVCFTj5jvuEngxfAmOL7Ol9XbzJd+IBjzMfWUiyv/kAjmsr4
9CFjMZmcFbYgYMHbGfyn8fyqL+HX9EciD8vlRMxhhKFoqIA0OPlIrfSTyVCgWlPhcyAXougfHOSM
x8kxoZKZr6JQQs1TBeuz1CFnUb1UC0VQOLOt6NrEfVJKEXPeb4XquDd8GUgzgpwkTyHRYQuH4gkH
ljo29ox3lE4x2DKeyg8oGUjNEqH89C/gcKfsBathMW0ke3uJAjUmEUmlkwUG3Zx0HNigm7KebvYE
Z+BBPahoZmlwfBkPgmpeQs1EHTu5EGh2zTw5B9ToJA+93rKHg0uCaPNKga42Vfg1TP9s2G/ejgXQ
ZJi8PfFlGSRqF6FAB/6cuKhFDldkbYfmSFRXSIv5AYQvdHhE3+z/nbwV6l/QM0v939O9t2+ucSjF
TzFIE+HbiXDi77TzlFCBXhShWYTuyz5vbhSPDKCxI2sn2yhUfFd2Cr7CYCHDBaXVndKW0zxtAhNI
gLdhXkvndYF6/Ugh0Zz6OUzC+Cq6f4+Rho+hO9NssRcOnzp17gHVFG4Bl5FSd/nvQo8i0CvUV6Zl
P02eTwc0nlwZ6uUSHU3sCN9B/PwRkDhSclInQx+57mA49OjKNtExgDp7h2GStC6biEu+8+VZH0cB
mqAvrcQseMfWtmaSkTXLCh0V6Fuho/Bk5KVfn6qN8VHi7Ts7ckf0FSgoYiOjgfMSSLNDF2G0jnT5
BmwSIZ0nQKx37y1BTHzo1TkP5AFDPPSuq+8q5ur4O0+7TLCcpBHjGnQJZhvNbl2h/V5uwd3CX/j1
LtVPThRiM6AHg5FEn4tDSrf9VU3ggPRkqFuFLgE7BAnsceRbjOsa/Oki1N/on2M6LM7ht/GYpySE
ITcmgYcLTVN6qYjAx/LWD3qpj5PW7R9LIfpB9pYOJaIGfsesmzZTRZHFDM4NTkBo9i7I9kkqwAfc
FNLulNc7tzE9kceJ0opOMV5zSTNDyd0Cdok04IPYTW8LYoPjLpYX6jQuruiJLsWk/+CEmTwlk3g4
Rx6linchd/7wocAmlR8OpCbCJaXwQ7ewyO9fLSEE4tsX77FqOMn85NcWcJ350WynlT5LKGNsOKxt
YK8u20K82G/nGrlm/9MB4uHCIRighM6uCmWx6Q7u8OdUJNuH5TiyGko41k3oEiRBYIs0lqB1jmda
6Bjt1+xltEkzt+lkGW/hueqkilenHeXesS7Nq5wRD9yPYgH1iCda0ObX9DTFyLsLExAaP6XnVLX9
1iLt1qTXC6nmY7YwnwGUgMmYTqi3bNr2vu2RSe88GDrqOeFiPCG4X/wY1F3z4Cgz2b8q72+MHX7M
xr4fl4oVevxEXyARXDT/YTgu07jcBCUmpOkV2HegEtmhBbReWwVi5yV5C8p7v2D8ydA0WeXFtVU7
0bnomtRJ13cYbgcblC9FvGDQltal7q7XGlxefW+0LO4z66Zecd4ImkcvR7M3x31yB0h6ldmPPEMS
P7Ar2HaTiafbARnzl1QsDWC1p2CNrXrwYSgZPsjo7j5aA8Ng3uJLJRqjYuVCu2gMdPENwW7KvihN
h6wx9OU9vrVK1tgGgSKUWT8SfNTa83t+7SDIVaTT42Gen3rNKV/mOMWVFSDSrIry47hqzN/NC/wm
1VDlzDpCci8FYhU0ByF2vMlqbyh0g95Ne1La+bRTPHUt7EOlXKOPEd+iTGXKxZiJWpCzUtoRGnas
oFqBGMPTJR2Cs9jrTvsx3FKtzxVU7X9MT0VGuco9CV/77rXQPi16zK1rx69xrDdUlKvkbGMizNfU
xvBS4Ozk3S3tApJRdR6PrHqv5ePMxHXcg29fsOH8F9ysLl3jkW4CDyA5RNGya53F88aUS4Xgljkq
tmx6SHUmGRKaD6y3QTZYxS5KZ4qjjTJa3x/ytDZXcZn8EL6Slu/KjOJERj7JKyIGNCG+LVkkUE+C
ZxPCuuWFup/BLDKQc8En7l44Gyoru3ZPRfdVHm0o8gmXuqj5iDBDyeTs+0glSlmye8WbpkpVOmm/
XXXSOFmIi5zhRXaX9UNo4FfZxtFBKZPRoJT8xZ1YVFyNvO6SOqw1/MjpESU6CyQDcyyzXvZLeLnz
muV1dI/EW7xrx3iMQJubcvyOPcDoNvNY7+IT28ITVrUrO6oIyauYi/w6pLeH/J7Im46CFaGpdd9s
ilOlgBi4cX7kuTn3tzJzoS6VDIDeZP9LkgyL222O2St6+KCalMsSmSiAR79IsEKp+B+/BYbFnTxp
Xy5rrHWMpLGm+XlHHRaSgTdG3S4YHAyZ52HYeb9CvPgLm+lle6QNXjA9neVO2cQr6Yd66hMSnA92
u4msoJv6te5kOEKXIHQns2GnRmK868Hyb99JmKqMmOL7wa2j8VwnO+tZgMJ6pg8AMpkidW3Fo22t
ZhE2ksr/VPzuQqlvitBMyYXKZLdrOpz9h6TUYyb9CNNfBxanTTijJnvW31GCHD9w9FNYa3xWhVQ+
0k13RD23zDHW3XisZZwjULjlKcvVlspDwNNe0H06immkKDvP3Yy22cgi1RjW5pZXz1e8AiWraD8q
7xcc5VrjGU4DrypS4IVLepAvufNSvCoDfmvoUCLutu2rzbrcIACRkTPVHVvcCHfHB7GnuwisLQ6E
UdKx0VV/lMu3/lQZwSfq4X8hgQyRyMzmPoOVCLskNsZ4MMNPZ+se2K1X+6kpjHEuoiseGwstjdpm
aPJSiG62JUkEbpGgBrsYVcxvYxrvB4eu8lTCKuTWrxG2aEdM9MjFZD5P8E50c3E2FjH7IQbhZBgS
bvvs5leSjgYM2rR+MkYMzCG8fzWwQGH/lN5rQLJY1Tvi5VQQfs8kLfodu23tH4MfwMcvpETbOjEv
MjZ+OIHJ1VSh0JJdPO55dBboMLiP7MmqA/PUWGi0xD1BUvPJlvDeqzwT2vTERsE3Xyh1M4V264vb
RRTkmWMgCpDCpbAkqQ6Dgspn+UW3rtQPKMVqETKfgq0TohjDpuHK4JRampwlzseMLS6s1VTkwvc8
I5fcJDoxR5wXFrp3zsu7y3n8H32dKOUKRpq2+LXJH1uxrPuI9Lsk2SfoGxOJFXDTHHD9qy/x8dmQ
mpEggzuTLby0AUgTMLvTaTHca+uH7zmW0jVuLKnXoGl1DWJx1iCvSvO+zHkQdwN3fSJoHsPiGcpc
eF9bJA6sct0b1uRA42SidNGKZkpqARh0l8qhankX7gNl5qWkunrVD9lztS9VdzsPyGhTZ6UyJz+m
Mhkxgcy4A+uttE3kR2l65otKm2WB98CccJiGd31nvFy5O5hDVRMgCmCP4FW3U6wOioh3sEsIvtDl
vmdEy74xisLxLdRHVTAZxHWfzumNPMxTAv3OCl6wg2AKPCygEL/brEN0tpml8ivKoYym8PCWevtb
/Tucnk+RSZk+90RnnONECumQGBvhmCQf+lCOXYiQGcLceJydYEdJvCvQ2HgJRbo1pzAatjs8NJUW
pR+Vc/SKQxHGTnYTt5DLxD7h6E6IGVbw93bHkfHR5PHzWV5M9SrIZOqTCCa6G4LhpGQ8d91vb2MA
AqOkcrFg28ByoXZGRRTA3FNz+z5yYFMTgmagiLOUSp/4pwhQvGfAYj96bmVrwtWFFRy7bRjSCfKP
8kVr/YxJRVA6fsYseP/wP5Ub1/7InUg1nocUKY7KyA8B2mtUDpYfO8Vw/PKjwyQTfF+rMBdNeX0s
N9BpksvsFddJRKO4AGJM3KTGp0slaBaEgWYz+gOxQWvSVfCo+JIgoBqSQqOlg8H6a2yIMiXxsn/R
/E8EJhgAsS3Jn6k0QUtC7gcOEqxS/0mths0wqFFQCZqffO8sj8At27sIPgLrrcmii9JYADSoX0Cq
2reqpdAdbjby7/wXjz8oduxbwmHPtwLO88FTPh+1dm7wzQF8Yna4JuTH/rZ2tLFVwJmYIYn8cX7v
gbK3kqAQsE5m5k8/H3Xz8YgWbMGy0PFBbZ5ffLZPtZlizJ2+z8Jy2yZQwdFfY3LeJazQUxEZxgyO
nIwXOEni6i14X6yDy1bB8cJ4JA433SVd/gDZsYn20jYgoEXiPMRTCOwQYKOuNTcG730Dd8i/qCLM
j7gVWdLIpF29mecL6xy2S3xk8aaIKUzJhWxxoC8ymEY3qa408LjITLwP18re4f+Ay/1qyLGPb2vM
GEwG3q6XDUFc7B+xduUXR9UkgRT8gR2quKBWJeeW1v3elJL/BtRxZslEWjavj9YSpyuRRajOetdo
DbQb/6prV8CxKOgjVc57Mt110lSTq6bjhFR4in3tpsdJIbrAUC5PKEYr+Z/9j5alNVnVpgB1CI1L
bD2nkmH2egQdBXUg0MfEye+QD8YLMsOGp7UUyn8gqHZuLxogDHCoy0pfmrMzSeVAj1uxtVfl3tHK
51z/13MUUPHYmnVFhPBWMGLeFkDOD9+QkMe6kPaGSJV8zXYM3FHcFsLRCqjEOwIsdI1edrSJRgjs
zvu5LqNpkl9ARIpBbAbngTtYLUIoVQtf3Pke2FEEyMwYuPWTTupcKVMUBhWi+lZTDKMMLmRV5894
/ih9fuWq02SqlCg0P/zcyk+IdpFroxZo4CHp5ON9guHxTwhW9kTn/JjrmAaYBo49hioD+PAhtM0G
4i1rj86WkCghLvf5nyek51NGaGScIkgUEVtTkkEJ2ESFCSPOxzgV5w6YNyqDdN/S6xhZuFH2z3Vr
q4K9MLtKmh9fKqCZbbZWjXeUNhrbepz6yzAWjTDo+1qvO74Ij7J8/JkgmDvf6Y2+acZtnTRRiFuX
D2h70+Mpi3spbZ0u5uBKZCIUNTsPajfVB974n2o9UQuiP7OEWRjZiieoQ4ft3R4suMtpWLaEpEhM
rml4Sw3n3/rNJF7cDWdW7ZmeJN7eC/wxUgzWd9qL4GivyRXwdIH3QxLq74QpIVhA7i+TN0mnCJCG
6NfHCi7sfYwNMqZiiD3NpgsBOza9oc+EFztr7iuru/y/gI4A6ZjzRi+M6h1WWpUw3aQi0qYv52+/
jYppysMbROhdT++efetVXWYdNlh+rqO+9i9niQijHqYiD7M2DmBVzgTPn9ptu0Zv0cZ+XzEgs6RO
C/zLv/PpK3jZUejTt2Niqf+An44N52B+YYUwzTMgWf+YQnjHvZQiciWT48lBaPTwmNaRuuVqtiZG
GCsCo4kPnYH0jY16TnrpRDOUXSNHAkudEr3X8ZIgFkLQ9jCSK2E6o6eV03fBWO7kWkMU9BMXXKYA
bQMqOLk0JBcJP+Zk51y4kWWe3AFQfK410+EbW6/xDJVd2XpBteG+XJdOoyccmLj95ZUuWLuqUyV7
NstXhBdTQKfRXCY+iGrSpS6FSkSej7DGdzU/MoSVbN6/ZBYUL/NTChToVjXSoP0gm4oSDaYuSVCE
b3LHgiBdw5zlrnkwPetn0Qs9t+CXlK5CMOPnEqEmfVU1jPe0QL4ovpHR11XPUPDWRKD7q9APyy77
osVUyYH9kNJQfMN1dBEXtffETeqo46PMWN1iZPTmHCYyCnuzl4VAQENIQoLzSLHKiBKqJJds213G
/Aqt6OFEja5ExD+fZ4raSU6syXpS3hUpuRuBv/LjNEu4iXbf3WuqdDoq0cyDawWO7Z0MbDQ4C7Tl
91Q67nOGMZcY2z2dHxa4QMC3h9Ou6vu9XAE38SXa6WND9nt0qPTb9vZH6J8G4vyp9WKaAU8IqbnM
CSPnU7RbhNK/JRANg8CmuMML82Ucyvt/c5ZRcK8hfKu2+HM+LCeyBQei0SewhQEHiRP1S1j4qm9U
E6EHXfExHRmNSNkjcc8Qu09jXWvGLk9djjUgxhLXwNJjWL5pwxSRWbTt0BgTuvHA8wmi3rs2gM1w
4HYAbi+bKUHNb3ehWFGEMyKYrVrVAy3kMX8vHu578v4pBPVQUwftFhDYvHIYQJekIWUyxpxPgJGF
7KYOLL5eHs53VdSM5fMuBb0WwcVw2K2ejCNlKEHBQCP7ndproAgZEVoefHSRSYlJOi/eAy0/LTs7
Zek8Wb5KFWzIWuNuX01Ms1f2VWym0dRjqE13IhM3Ia78ACxFUrt3COdTsHvKV8jmVb1DAJGNh8rB
Og6JX1BxjwmdRKeaGQrFjTXxKUdowKuoJYkwkE/SABHfNRQQgwDzdPnDf5giwzGgmc6PTZvjBEsj
JtI7KNOu6S+HibqRm5tCSG63efdTNYUNbHrEWtBDjwehKzzl51AscFdI5h5hukJGexXhcU/cbRWe
Q3rnryfW9PDN0E4qCkGmjAzzXvzOszexAjNmlUNxorOcrPKfAfEoVn0YaS8bJ8WukPoUMkZC3h+k
mUzwWZSEntGA0OpUNK0MGJSWpgQc6ZTczTs3zBSfKtgfNeS3nM8D2/SqARMeYQeIwr8+MIMp9tbT
Iz+1QO8PjnZgLo+N3b/EWUJfyMXQx1vhTyvoeDtgPmzio2FaVQzyhGIv+kQw3LjMSGah7+4L9bbn
dCA6/IHNmBPKdqwyuUXr3+aGX/EzjQiuG8M/eIFqsMkD7NlNqnrfNuDEXL6ssieZZMYNSwHDEbyD
efht93C6oYYu84SbxT6YNIMMVpmmxLf6czpz8sThAlWYANGk5Pi4LTXI3D1CoqKLYXe3TDWE5asY
FdCnLWwoq8hjAZwT27ojuYGblbteB510lsejpbSTIaHt454XqI6oqvShySxMtz6WJGMDmmBPYnPl
B2uTbFqKxncpSl9DbgpjE6W3ClkIwEa5OrzNvtAZK+k5b/ZzCdwWbYv5fw3TJFBXyrq3LCaapNyg
ZUjLI+GOvoevqcDtzivaDT9s3LhMOLkop/CLajZp8so0+Gm4ss3CgDse9ioZYHl9svnpvuxu1LtB
aS2lLtDJMkJI3bJqRUCZxFYNrOrP7N4h6gDz2EgMVg3gUdq5kR0XybBxlSlGs3qeHBGwfQ/fAikT
mVo0QyJikKpWemohGYndIkqnWbiaWC8aNyIbrY9T8gU7bgc2Zj6a6ZPsDF0sFgsDchYVDC8ak7AD
uLq51wHQlDUVZpXBW8o3Y+p4gvV5DdbV/sp/RXsfanvADo/jCo6SMPFYFfaAxRnGh8YeUNN0DLEj
VBHxCyDgphltCkeAE/HZeWuc+lrV5zR0FHyhB8zJDGASa2tQE1rqbPwmH6a6mT0UuFi18CU5Qrs3
wjJ3KAm2O6zQaLnsoFtIZL/t0wTxqTvLHEcKUTs+EJni4vroc1WmNiym31usVGkZGwaXRdLmdpkx
d3qbGACi3ML7xiythsgArBjfGXQbFJ0ukoMN2BSRchfoXUkGGG66wR3ICmiA7ThZ6UXc+K5yub+c
qtQEGBWsoTnu7ryl/qntlgAmDqsawcgA2Q5LlIPt04MBRjWDKaJjhTZ2Pn64YwVX+d7vBOfqYcJP
J4wwY3ezNSfkZaf331NzkglI/ryHZSq/i2wrCd33OEaPiU7WirVRqMXTGRd91fmX2fZdVeZ6q5oz
dYf6+qKUWFhRGMkihHgevLjpX11oiix0v6Rb6lJMBIufO+z6s8COUMcOnX3nkWSkJWQI3lJdH8fe
+693s0r9TKeIlY8XFr4SBFqFDmeOv26DPD4CW6CMaO6sO7N09HT/4SligsQ1tFe+L822jgwnaRVY
j03+h+vl4dUqpeDZizC8YSDpAA7pQwoXBPH/4Posix2w0slUHb7T5VGMwwFZRQOqmLtGNV9hW0nt
aOfLHoY2r9D1yam/E8Zva+tlss9aAzw7uxyyPlhfsYiIL5bLPAlXHinYQGTwzhz7b7qlbf4alfLr
d7O3GHsRGL/3C3vcwxR7mDhMgkYqbsV/eEMvZNSKBYxkLyTtZTcG+9auWZVdYBkd2nYYe7kR7Is+
rZKSlOGI7evXRp9N4UuHIs58QYU5KXQVHzJ1Q/pZHkGGfi0BjTwYw8hXZgDsGNLG0BGsqprQopBI
hHitMNvWb6aDIJCZp55FxfaAEGoZiST9cZMehrvqucIzb7CQID1ClpGgLdXRfnt41D/M9m+UJJoZ
i7DiAblLtffAQycuowZAID4ziu9TQSe9g/ef/2k4EAOIYarL5atpqcHvW+tAfRkMUrSPWne3ZOzn
fCce1a3oEblZwFlVN/JE+PYfYvkZR+afBQtcZqBudQzHpHnjIizmrhvepO8Us8uXN3a8qp3BQTPL
8ZMJ67PMSaRFPZHvNYuqIYPj+2bPb/UiOgz1L9JK/VnKuXuqvIDMCPb1MmGDwBdmRX0dPJXt4pD2
He6lfaHVdOEDnIeqmfS21Hgvbs49VJfmo+1MT6tpkIyRSML6O2FeLKGQPUb+7PGkB8hmpkJQwJ8i
II8x4fcJzkiE/v6x8iGIQ5fIvQJYyS8dn0++EQ8Op6Qqf5xG2G8KD04uUZTXK9YvkowwCnjgBNo2
o/Aadio1rLtDrMHlaG52ucLJ7RKkLXJvHZWNWXpiu9fAy9KusJfCDmhHYZmnepINbLIL/lwKJ27u
namCR4GCREp2Z5MvQ+z1wL1K7XWVXLJERhltv+1SaCVRnzlx84Bvkv3yPOQRBtbRBU3oMPutDA6E
vqAgbcBbCqnG46o2Bd5ASjCJWZz4mZabRH3F9AdH+uv7+4XZTD2tysP1TtijZ0Nud2i0nT30RWOn
AEOouYnKrhhgQx/jhG1p6AfyNg+a/1J7m3/NDJI//v9/lYNh3NExy/M4j5sCJ7RIKRES/evVk/lY
6zs0ynZQ1MbjrcgnCbM8SqalDGMw3z72mP3+xlezo4yDmubVPEijKS6otd3w4edu116Vi0qrydwo
hPmejnvVn5fjGGtt56RzNkHmPY7dwj6r1k8hULb1pAUNH4ikYLMdGUqi6XYNd+9dyW4nGC+PmRBK
IR5rmiqFgwX/SRvlJihjHWDjSHbdcYctJCscjXePcaWnWeSEMn1WUSY5+ebcdy2uggtXdE++zF3n
lh9bfb4e6K+pLcT0nBXYDB44bQbsXdUlrgga2MQQzYUskXt9jSMzmXRmHKmfcKap5tPYQ72i7q/0
CyCxHhX3l5TZ6MGPBmyZO5+j4b2IZm4KVV9uht3R3Ak7Adv/rV5tdhvKxogqn7Q7bu7O7WtLiuh1
LbHwz5VK/D+R9IB/OJZKHrBFV1cg6wdiat2+me3lf1BjzTZao1FxIcTxMVytrlCzj9jQRBsKQchd
cbZbmVdHZRJqsIiQp3k4hh51yqTL0Me8t8yF5CbGQZfU1/nooXNT2o2/fKBvFHyPcfcBPduPowTP
zrBjwfPBBsjgfTZvKnYLU9lgwB1laeidCpZ/ueFn5fG1U+d/6iw5+tlWSKXR4WIHdeSofT2OLxBx
+Et91Gi2BZtRxko7vtS/alfB3KCJDlRsyAtFNR0SDfyNB546UOHaIaMLt5GkHb2fhwFXN54xqo/o
ELKqKLbqgaZcGpOemIhh3+4jd3uHwA/UpmMrWw86VxOXztA6BLVRUl2mITCFIQVVN2+HEaBWYVxs
H6taIGi+5DaL+ZxbrYr9dqLwQePJ04aylU//IHYUwq0sanmku14YpRd3XYeaHH4gE/sQEuqVTFVM
Vw27cw/p/xeoJGJ881kQbS5R3OlIUqnax89uq3mNLPEwIBySW8322sbjzpJvfTvEh6Y8a5vWPPHT
+adDxIWOnPyZpE5s5EL5bKe4zm1OEyvscOMWONxsvJnlE6Fn/q5DDhrewdqKh0QNb2FqlXh18Gpt
bggDLMglV59bepROfWGY1ksqrPDvhoIGdGhhMEmGKLp9wf2Xg5w0mZd3gGxOG/2+96izgeopNjeh
1sXXloszH/V21nbyEgYOA18yj3LxOKa0GDmbtt7P9QwcUiPm+N8PxQByli46rJdQsEcDXYmT/MzO
CF7VcfqFwZvaQgp1IKckZ2ATu4rR+KGj9GEkfGnvTY1NMruUklckGekT0JgCJXS79IbMmDNXwd87
vnZoBZPiuX4esh5BJlrgT/ZrWNTzaakp/PZZzdlCbjOH3TYBO3SUdqUYtfFH6oPUsw6pk978mDxL
9gQcdJfNvUqzwR+AIV7XS5AF2WXYzoJRQXcFtjLsCdH/HYMbPgzF/qvKehQrTasefycQf8nA/Qq4
p1Qj3GpxNS9ztJBrS9is1Drh+Wbh+fpnSIggRyooI7R5v6V/C8SAVAPaLp5qQe2v325kAuzqBKfg
5yLHdwfvEPyu2WQ9Y/daWed61VXZeNfQpG3oLe14ft2e99DsMljHG6bjEuTr38WAkSLFke2ieA9s
o4W4jHBS6cn/dya0TY2HyPpr+77YxsGjXR+Ge6ixqcgj0pwlK9SnsUxAlVy0Mo92Kam1HWQWR+pf
Aivpv3ma/GVIFVR0jsuRjuk4M+Kf/MxUo1ypIQ9b13sttBMiv4i5HhFLRLzabqskkniRaAV/zmKC
UJs94sl1njwEcWN1W5haI9n1/sdQBcPATjXkEegRsaLE9asmJpmHKsFrgxwPBznEHe/ESc4YswdW
YFS/DWxhDmRIMrxtDtUm4nJxkgbAuGLN2RdKY5hMrmIDhOOgxblPhWe9SMLy3a8de2wPeCM4Agc2
k4N92oYsmY0WJDx89SX38kWqBlHQ8TOs1jC07KUv2DsHDNsZiak/Nn4/3MeN+37mstkkbSolRUFA
Sp1qz1OxVbS5ejLlnffZmWY6Znh9rH2sEWGr3n8Q9hC3jE5dtMJ32o3ZMcy1nGk3Z/Errqmd/fAk
D4WFFcYc/9x7UpkmzSzrwLUiD/mh1xG2Lst1JMvAXGJOtvItejKSwhpPIx60+cPbTfQPdxFt2iM/
8cvVtT0ED3icdSflnteyFYBiJ4K7W4SDiMVoCCsaX72FBniKWKXllPN7wK9y0ZXGvsM6hibTQAf5
pFv9jDxIGZkyPrsTtTC9lJ4d1FdizV0cS8sr1464kr3CyPyWkR2eXZDnjvUyjvibR6Bzd26XEDlm
tw74iQy77g9AilB4vS0Txsw2GDzeRVtI2i9mOatHKfg+bnrGPhxCi7xZepLAJB4laNF1OaqMCPx4
577jx9A7VfA/m7lytZ4OMbVax8TJreAWYLSSuNjBuqolFGNrXRzkkvQxRoZXBT1Bvv0GDDq3wH+Y
4YzE3bz+g022NwFOSF13yS79E7I1O4ejrxv+J83Mk7TDuZ//mHEUfW/tTu5buo9646om4xR/oS45
ELPWY0lyRUW9dskzfHdSI2vZ1yky8oKVs+Hce3QtvPi+y8iNw+dZrBrjwMSjF0ICGy9F5r6Z3zyW
ze84kubUwk3Fki6uhKkruTBN0N7FiyQkuMTQwep4Dg5vlCMbWegYd4LYDjZ2VqmlkAfb5qfmaQGL
6xU6Nd6WUTusl2kMlrp62Ko50eDEx6Ii4MHRZAiqCJOCyXvyTm4I7uENAUnKn5OBsrXrvwsDLa8F
UZ886KudNYqCWEdr/vCYYoGOyMxfsg/HCrdpBvkmQGol1zrsgCMQQqVl6RvcZusqVXXCpqaN2L44
23eiDTpSMfZWYmB/Y6LMGvzHMOXZOwB2jmgKV0cZp2RunYmjH1MOKVkWDvAsJ9Behm/o5jnvIaQT
yWv8hirVkMxhIBAXN6tUhNCQsUskWs0NLBX0Zaa4KKf6pIQog1kyp5KfbGofRSex9IpjJlwdNemX
0DSgzBtTGmnHYxqfOKka7xAaTvJSG5ZvQelD+cuNjDFksQWRrqaqDn4SJo7ABVg3fCIFctfbV7ks
08BWUmGvAi0KuVe26J8ewsf8sCKEChgK2MsxfBLxT7DjhRU8+1/6BTZs2Re5CD1DwKB/GboqGgKI
R6+HIA154NwgkVi4XGcI3XAJuDMIdRH23e6xNtK5AW8n7HigYiweIly0Q/Hz3fXPZggW4pWXN1St
nQRG1T5YUIV9tRhm9qN5gxx0K3Uj20iOmx1U1tCrac0WeuFnCnE26a4DgW2oOjl2ylQhPvH5EYwB
808tnQKIkHYXX4hjn4eE7Q6hNKy8AMGSp/XyG5DcmlyDIFeNz5r/fvzpzP/qr8UvImQ27FkC3frI
vkaa2Qt+LCnuUf0fDSvsl+I+A33kC86gfMv8c02Cfy1ZE0k1j3qc0ndv8KdVau10YsB0TFv7Z4Ea
hW7iSQJD57/mYxNfQ9hTnawUJJgTPRnMKmZvHAs14s01/zRnMfwp/ipY9utIYuDqhMZPelnOyMcI
KycgvnhU+ORYlqvIDmIotfsD77J/MgaMPRnvad6Iex12oEkOwZHYBsWJ+PQaqDj9Bli30zDkjb0h
XnXNzjwA6woDneSEaZI0MkefyzHfxM3u/v8LOJdynMiOlXAdSv8kT9JvSWbCQUCyyu4AYExnis+q
pt0QC8z5vKeosNwcvZWn8hfCOoFpqe4QwdRe7EsBNrcAd/Rovi1YUElBOkkR06fsnlPmUf8D5TiI
dzgjg+9xHP0kH/xcb70PPk5YauHbCfcBEQQ1zhLQUKavAaWgZcg6vSNWwlkMY4M2ck83XUqXtbeq
5wAwHNGU1nL/t5XO5iq3DC++01GlFKxFR96bm7uy/rfEHTSeWLlBUxUq3+M9ziFYVUDxUAIM/TK/
Hb3QKnjPDOwMM/0ph4UHKqZ53Bax7AuilbstQCEyr9IVU95dpVJ2sfSGcqitLD7FtBFJnWsjeXwT
XWe420aMSgKmyX9Cey9E6fpt6eORQ1w/lo5qXf9H0kUZZ4cYzpsLOkHpQ9iiUBMAMn2HzY9x4vmz
6P6K8AEFXRqlPhOr3Wtz5Ywc7Nl+jN5x2lHKxiS801AvxLBoOVTrcQ9M7JuoWa4X1aNDSw3TPsNW
+aAHlnJ6GlefQCw+Bsr/HmIByU2nXukXfP7Ap3zignnC7LawsGQ8xr7VeozN28RDuftl+efsGmEV
m3cG2uoUmonsfv0Az4W5qleAsXb5BUaaix35A+aZlLRuiKfh6O1NZNWk0M7n6Zh8yrWIN0eSucoW
Gw3egz4mOuoGiBS1qNJDaNM3zuYe7d/f7oLS0iOuBOqs98z6XD94UrleYU57sXpjNuH4aXDlatW0
++nkLqGvykS5QPh59H1svDYbt0aA9as7jSKxyOshn5j/22YGQnrMRce7Q8FrdfyoI5pzmCgd0TkY
pqZZalqELAoD2wgUh40Rbk/gEV1YOQi0/r/au6vIFcshEw/kVQTpOBwPmmeEQ/akxP7e6+IrKWDx
OLVGEeL5B+feXDzhJGHcklkckoLrZAtlwkMD4MH0rEcUvOrN75/zyZgzj7a9AfHthnF/NpIxPQx6
VfloZJqXP3PXyhSjaxZV0KVeQ1hwpXLzoIT/rmUEYcCHiRYwf87Fwn8ISdYPMKFEGlhV8AiPOhm3
wBdBEeOx428Oq3fQ+8ggGPnFbUba2Zb+zpI7N60ZFjuht7RVVh4BoGKdQKAahqOMwKaM+/T8AMR9
yuCX55mimBGKHVlNEubF6OYQ/xjeRcA0MMLz9hzkJmYfJ7GVw8pgVSdItoRR+cd5hpk3+T4hWaqr
JOT9wgNnXMifY9pLwdfky50Ftaw9yKNOpmPN4cCHDN/jlWDmqBt0s671pPBtqLreKZNzJnQha7B8
VlsmhvG+/RP6eM4G6RK9MX+oMtph7Yw7BJ8o1IuKShDwW+CruNmxgKu67JFoVcAqBuYUr361iXbl
cD+FJwPqLpY4lyLhclSivOFQKOd5AhcLDN/VUTo0lmwKvAaErMjo6AlpjAHGTBl5rOMFQ3umOyrm
mr9EcDGslMrF4XVpCjDgtJaDnem9CnBmRauMPjsN3aAqsaciqRiWlfKy9zBPbf444LUrgur5mxHt
Jdgb/akpCxEDNYgXP0edMPZTZHpx2GxVbctfYsjqItDp6Il/YG3x2Z1gtD04LVadnd2AzS8LMl+L
aUUYi0up1Mgzj0x9nPISxwwNnmesdwboW9Guamln+SmodV7CkQVv29UvIEvUB7a2C3iVSKpVsntJ
b1pFits+hxXYI/vgV9JVxXIKFQX6DVBiXLS4yxYuNrfiDZtcvNkbrVC0Ip+N1z7giVpoaKOIRyEc
1aLxBR5/lTrQ9NLoA1lai/2Z2RJMltzOVvGxBnUdpqiFWm2IiF8iZLeEPSwUjX33DpzB3e9XvsIG
lRA9Wx7aDZCF4agaSvyvtcf5mq1s9t/B1ygrfd1UJ/ZLnYjq+Sm5YKH5G4tAkoOnKEpr0HXYi3TO
RJIleweD4+yjXT8tFPrwkOrdBOyd1TNDsoSN8OqyXFTPLqNqZbS+Ac6IT/k8vbv8J9YWkGxs1D1M
BskBgJf7CfMFpAvZsVTAxUUSaoVVF6ZQF/0H/sFUJLS5YKRTCd6pavN/TQ/4yhiKJ2fokMRK1agW
jpF4X91572O4shnQNbmrWnh/Zt8b9sSlC9EwU09c23MmBthwjnesuyyoGigd5GBr49FIjTqoNhxZ
8YfHmhETpOqGNu6GP/zJu8RF7c2vv9N1RY7wqcLDdwZ0JYILP+u1jalFi4I6Mz1/3PRGcHjPGZYg
ojlO08Xez2j2laf2wW5lrWys53OU0+qNUJbz/uGHpRYMYSBCb7S/qKIuQUt9tX2cBJXsrpGg8EWP
eYjFRDf2CL2a4f3ZWuud+T/S9CeurunvFEvoo+NpvBMkLNGQAryW0obtGjH5ZfOde3glEmkrSuiA
krEOofmfl91skGeeY0xqgRBRXUB/ot3JBBVChwTEpIzhmJqm3+PrUNT4lTNsIzsAOfMzPPFjVNmU
vJyah4XOxrHv9RIxqky9k4+/l7HRcWOoMBzw8LZWnsbO7xoIIefF6uGktH/gGEBFXW2t6DIqUkT4
5h7cYEj8BWZE1Wrh5klLqVIN6S0hks/nq1dlR0oYfQTD+ycOgKexdAKX9ED0YBbPqkwawqJvieag
4hKhCr+y57ZuKg2aVsmZlBE6+KA0LRB8l4tGtap2XNv6Ra1K2PSYQfiFJpW0iSedd9FFXGUWjDxF
cxPM/CZFmkD0lhN+eQf3ercuYZ1dLwOtP08O/tpvcuL6QNsK+mgNmlwWn/8l4lYsgEYFY3QDXoGA
KQM2xvOgaXsGgeAmqqmwndEm/YMRnIGAThbTjRL8ttf99ZtJ/tJxOSOlmhBsvyfH6c+roIly6EAr
eXh4eYz0U/lp8ERCd1zBMejvvTBvXwr+JthMrafsxkU44B9TSNgloiquE3QL8UqleJPZoNfS5g/h
Hak23Plv083owttSUbThfSUupmir+CGNjS66FgnZaI67CCSIah6swmWWaAjiCY1Y0o1zJYec9q24
kOLCZTTtjxok0riwK/ijdXJ63eYvsIjDuDuY8AycXClf9ML3eu0zsuTk9HubNcJ6TFsCfcY5Ojza
aBLtuHablWpYVFupZJhorJz1Izr8OPO1INfpmDbPDD6Fc7aD42pG4WfZX4/poIgMTtlZn8kBCZB+
BjmkpOyxTn6UrH/iEHw+xaiPNLvcFU703XMA7FHTN8Lk76wvolWdCc72Y+xI6y/hiFefwRt6jWHy
8GoTKgT3TXNH+1Uk3O2NGsITAbrCRCMdBSZN8VEOZYutnHQZ8jJH8Xg7Hn0bWLi4Seh5DWoDWYWu
znT1TQihI2qYUGRZNs/44ONsWcUZ/HabF3z6KbmnJi89srxwahJ7A4inIQY5rRLztmcDbv3DHr47
o1pYjUQm9dqezSizSiJ7WEmQMjxaogMbOmG9AdmSMTK/mWSFUrFyvgEMQajgvzaTbMMpKvNW48WE
FlvITwrfiX8/bzFaNZXLxOnwKaynX/V82pdlYdz/wb4FAxc24Hm/acA8IA4KaQovjTBc7058qByd
qlXeqVxP/yKNUAWf1NfwiLPIlmmzDjKEFeHDeYtIyHGezC5ApztAj5bfQmdKY2FBKNy/GJDPOcEx
VnkRo49mxRVsU08baPBt5tYu2e6J+86k/wuX40DiQIy6fRmTreVD++KLa8Fi9SmCFicvXraeuDum
Ov5EaL/LSIBwIMF3bu0/dIj/uFt/VdFmvrI6n9Q2HthPW7EaBFV5PN43XQDcpZeP4YH+wrxOi2Mw
mf41MefyGSM8a/C7RAosbG+xCGeIiM0EorPrl1aakgQN4U15zodxaX+B5iE2DeDW3UE74YmaNp/3
JFT22OKN4wOWs+PHvLVy7MQtkKsFrUmqLgl0DYAhj5zF0PdbmcHP02EkWhEiaOeHiop2drNinJDL
WAu1G4pYkUYf1ATB6EAjTSDUcdknpGFe2LiaEIBLGa3evWwRuFjq3E0Pjn2xWPqofercicOx7Us9
xsSHg5A4phKWYFEjVCdF3Kmb+GGDE0Ghe0aDLpukeZ8RN0HgaU5THTyXDg8y/0QWsSWowTnHvouo
pgMgqWnrT9PxZQyd6kbo2GjbNF3B1XUk3U8TjtN13IP+98OzQUeAP9+G7ONpo6dQ9rKjm3nLeSaD
7nzAxefDEs4JQ3HoAccQ6KDySjRomgLCqCUcExR+p1cSH4R+CZJ+luAhZthidvCCDFxiGKPXiprK
ELssPwg54ZoLsBhRjkwjF2qGKXXyae7Db6EvyGvIL9fgDY1FwV6Q7/mzNfkvVI8M6X3HK/bp0phB
TE732m8Y+dTlpNvxi7vTig4D/epnmI2eJN6fekhKX8gyYXHCsmfJ05RGOr2G5fMmgULE/5pywryt
OZpTYQIf2C212574QYj9HU5suxZWN3UaPT15zuEWD/KDMul0fq7xbUdsyceT7QRq7OghKqtYNVV3
Zqb6FvYbOZU8LJ3mHQLMhOgyvQmyrAdZv2weGrCV9br6lWDCLQfFZ3XG0TpN6MXcyI9lnn6x/6fo
FjPhW+DwtVVEovBM4bs9r+hTdS85e6Qh96Oe73fz+fjjo/v9Qm5MLb9yqghebJmH3moAfMvNb/JY
/SPovQE6CsXmQRdyA51+E6/FcJZSEy4W6A7ZeIcQBNBxK94EMpaYBAsdnM6RDRlBFAMKWgCCgA2M
XSY+44yWAmymwPm5peX4e7EtM3xF4dfymvw2DZuPMQRcoXW/V/inNYjyqGJQCq7sNxbd+yP9HNp4
TJlId6RSYredTYj+HVDqCJA8STMTx6x7p33vn3wg0xS8UMjyDqasegMxfKlFRHs/fT2g5JTO4kRm
lG9XHiI4mcqXx2HhIc7ZyeuAaXteDlkfBe+c6hN9jugmJdZi1GA/QhCXYpPd1CTEDQ+Bh7joidIb
SA5scNzmxSC5gbIAgBxsgmOgAd77l6LpwHZv+7prhmd2OZGHUECRYLCtPaXykFefRdf3Gs5pJTT8
qiXylyy2gpwFiz2egs0UKLhFCEuV6xWY02Sh27DsTeiEvPr/j4cpKTViWdTTJ+aeDCutoIi8lDTt
7vowfPZLoBbLPm6o1pKYZnWp3rDDODUJKHS65OogbB6E0uxheypb5+o57A96ham5iJkVOj9Hsm0F
b2ALjOT4m9JDUppaVQ5fOw06yirkRPH0iPYD1U/2nJ3b/98u+iLLW/fx2cdImAt8nO+jbqkhM83G
S6Y7rX8EyFO+JOwqDJ+WDFOXftRpBDlGrCg/crgNiYG/qN5HLskTldoPwm2uaCM7Tae3LwQyHFeX
aY/xOcVHjsVoTXZk2BPM5HwNUz869uoWSXmsNdtFd0qnd4R7lsf5oZ4l6+y2n9Y0VUuf4awcxLAz
wEhG/DtNH+JRHWQaLvyYUN60yOTOcBgGbg+/2joFRF74CmAdEkwY8YvLKpcsRA9+VVX54Mg7Tq6K
FGuQghRc7r0xHoLzjKU7vwy91kY4TB4sYdK8Zm8EZjivROADQ7hfhxjCTR3ZWY3itcT1QfmOAMhA
BlNkCwJ1xcKCsylovQe7kfPL1LQjEGkTAQ1UzNgs2g4nJnX0OZsyUclPNXX75eEOx8M1sSSkRGbk
K5ymyvTEl2tQXTGZn1+rsqHQhvHvcvrPn88IIxGS0Pj0NMbGVeZrsz4TGYgVBdI7TM8aPtMF6lgJ
cwgL7YC0zY+7aiC1qVeJ+lZzvlfSTa3KBzgsDGUaloYhdmrgPeCxoMPPs9gTbi2VQUDtwHwZBeXS
LoG58GaqN7QsZ8Vnxq86I6QIuAnxFA8niMU7Jo9QwwNO3jDNolz/nsOb+gazjQJVSjBVBHuGVqgD
ZFvD5BizrzQ1x7ltkMZQeOgbmC339QcRiumm8Zt8yzN3PT+Xaw1ZM9NlaUfb2us3jCwsyBp+paX7
zYLFjXrzcvlz7KXbvI+FQc9mjdJ9U0MyNRzIb0r7JgbSbTKqzSCPT8LUBzyn/5d4zFKokthh95AQ
Go1asDn63SF7IflOpFQyxuans6glmMjWteMs6Y4y8bZ6WEDdlFKFbTURTLNwblnZA22K4Y730lAS
V0hIlVPr9plJrl6cv2azUpy75RDRuKM6zdwffAUMl7Zco8vmci405qS1fDEgbFC+MHfepidbPQD5
B2kiTBpuYeJk0QVwSiVzED24WRIXtcawmVpVIH3Q0X82K3dtjr54ceiRwQEvTRa+TDkpc6euWxqK
mypscEgxVALlvOjm0uOo9GHzLgS7B3c1GZhyxrarHuOjCfrIahp1zYPQH/pP//NwNG5kA4GkTeoq
lTo/SEnEK14x21oEovtJXMtpZNHU3fl54zzyNA0a0sLx/SPLhSVaxjXMBiJnf81YBhxjIqIFvwq8
mB/JekjJ6pida1ZkgfUcX/cMefJhaOv5GBBx6472KGgF1foxegQKnxZxlMiE98PQPUI3ui/rKXdH
XypeedwoDDuhZK5QT/69uGxM2ZbuZyniMOVT5/MUMRq9On9NzR7k9OCDEUw4hLFIXuBIk9kxsJ4x
068pFm9CN/t18T+rXQuYDDtAvbbsG1cXhM7M9YjKmgcRgXrctcG7nXSjGihlHN5NVRfCd9ttkJu7
jmVIppzQk9i1JyDA6BmQYyjOQCg+b8zIysoVguhKHOsycsrXrr5+0oeq8ZQggbW2pKZJHCk8A79t
O4wq1tLG1Cksjh7TFPxud3lTD77ow2bh/N0OacYacC8L8Aajo7axldqwCZMl8/TFZQqAebXAPTzJ
q5K69JJ02GGQk32Qeo5TMzeOwP7EX5pFQ7Sg6LusjedsfQv1bUZTRuHfeRSpaNaAf8M/e3flQ5PI
g6oUuNBRKzIt/oHaSQRkCtgCWqJEuP7b0YV9TMFeQaQUOnJIyO+UU7AuTkKZyfr7/6cSLMSW2eUE
RlKjFX5V9q7KXkP2r7ve3r1AVGoBVrbFH2b8j4qufBX1OWNB9gb0331frOp2QbS3Zp2uzcsbxVXP
ehB96pXWNv6/yWaxxsbxc771Y88hLvlhNU1sB32TJ7PMnWmxhJ8Kf6FKUmgDDIx9CO4ch3A0YW66
RlLcCeuBFWKbGhHVaKfHmqQCRWXRlrM6wbL0oLcjT/Q3QTHspThV0kNNNPcdqE4pV5mPUZZIToG2
qela0q5AkBqMGVoOY8sUaJta8MVaIClXGrOqLonyI+kK1zcdfZlIFYJSTBKA2iyEfkhSLHmd5iwK
Q9TlohJHTCfOsx4a1LNO1grfl6VOC1GNgHZO9o8D9v6RWx3IAvzs6rXPW1RLkptu0jhJ5Tb7I7fW
XCB1EdGqcQrco55rtskFHhGhULzFJlyC/iqMF4oWV8JnLT1nh/HE1sf0JO+ZVjyaauJTMRIBU4Ic
gsWy1ELy6B753e62eq8FuFr0tIIpOAgiDQeESo6nXHGvKs5oZeekwxuWWEnDszifgqTUcYiSbdcb
HN9iW49EnMzMN5YHwi9oP0O7SYi4muuKbi2NsZPlH9E9cMfxKzR8E/iG7md7cj2mbLmM7oBpOqqf
EmRcYAl3TFKCFMuBf/mYh9C8gQzZO0CxJCf9or1m0002/rLShxSIMl/dBbch2IJNE6CX96OcSNLG
jyfn+HNsjt/n9TB3oiPpdb3RBKMhTeKPLRhqZd0rtviJvwa/MHxpIeyMEoHEs1H+Z7SPzAWbrn4l
TztgXjTA1L+NVCKfBNLW2OFzJRFd1Y7/m0OdSHMUocRi8+R5EgZp4jFrMHsgLFamYxwvcWp6JdI+
86PkP/20LOc/ty9w0jBSs9M+T7R6wX6rDyT3wSctODyK9WpwRM6yNZ/YiWzuFsepZilVLS6bI+MN
1S1i/hMvURvB4UAWvEqXO3+LrQu7X9tEva02yczzMHd9PAhzFeYrvPevvHXtRV/uuxjDO5S1E5Wi
YNSAb/Qd7qTfhWoINnptCeU/cUtmgorEQdDMHz26duOgPnyjOfV4Kd4OzOHqq8jXplfgMb7Oh4Ee
btqgbETpm0S7TGsTIYPEGDAYlv6xRvpTAigPKSmlgRRsN7fpkjSBeY4OpRNuJ0/F07uVtX2JfJ80
1T4w2Ixx0iSV9pDDEBPJbxg+9vJNyyjIaR8/TgAHpVCunTSxaavW4MKdL60SObJSAj85Lv2SDXKX
32ySogfvdBxAyUqcGghjdf9U94otPAmMeSumvgR07maJW0Xz3SUCiFmTj2xQpg8AU2xlDOD2LTvK
gp9ZjDtrczRHnrtMTcwbJqi5Bghqx0usSLzp130VJPTCo+9J3hbBiPyZhU65hN6soT8R2Ed6rvcI
Lpr9BJkCrIn/LtG87LdqTD/8II0DgEdBDHVVWwJlW+lUx7+YH8q2yiLAXtVrPy3Pd4aZ0zfkfU9q
mzh+CasWaxwSY/ZShmasVUJzUwGFMKRWH96X8Rckjb3Bb3oYE+UKZ+mCzAOclitNcQunRQi//rny
LrcEPN8n8IZm1QihJKcENum8yYRnQGtdCnMEkTYLY0M5kGpyI8QwfXvCZFb3a9XwXiYCjeV4Tbix
2WptarjX1KnhWAIuc3X/oc+PrFxgOtiWlKICvJFPsZhMEMevcRb/Gq1cy8y6+wWeGxbKC2NniZVB
Tnf4SVCvpq/f1fL49xJaOrAh5noLACvG/ZeQegYWFQ7/0zmrYPpkTN/IdkwrZWXrwt/j78TN5YlR
Gw+KGcf19qbFQ2ZdJnOv7gBR2ox3pwhUghpEOhUHWeNvr25jq8RM7kR/klEuRXzA63ZTqKT5mBGK
UiJxLUUtqVJeDGgP+Qiog8ErAqi4NIkM0C83repkxCgo1YCIpV4AcbQNUoayTHnEcBWZHCQnyz3N
UhJx9xHZEEXo6rx/Hnpl7LLOEk1HpdyVCWXxlrDHaBlA78A++lERgpa5oxSYZ1qNvpt+AAgbMWyl
FsQgus0TJzZH9mSIAY/t0N2jjq87eEWvubGXr7+CecyPMhUomx5D+2bTWj1tVv+/6f0WvE5eXHVE
x7hg4wqxG+P7O1lEka59dSw+Wwsxo47p1mwLkxOubrfKgz0CRd45CSji3+MGPH7HNJQdGPBU/2dH
nyLajISIrHBpB+5xwaYoNA4Sb73s9GbeFTJ4CjLC5vRR6oXeUP2N07OTuyC3+7965s6F5K4EaSDO
9hZj6nTAjZruAC1a73wHv245zX4SkFJT3QCH0US607pGe9GuOqp5i+gO8+lCsP02nQE7HLU1iIz7
/EjH/nzFFD5XKi6O14BKg7EnGxbAZ+mtN9J+wz4+B4nRfIlDjt2B3CpUrWxbPSJdiyv/OX2cgfae
z1r1TcMa7YpyG62V8xUEgBkmhvxfbH8uI1ITbEe01VGQRVCFZ8Bw4Ep5BKRChnZ6v3QCCYAkymIR
zX1JE5TU+hUgzWg7llOw3GflfD4alnOmeAd6GsHNR/BvE8oj4FjeYND0bb7eRutMSPxPPHj2AT44
K4HSm2ldp+HXnqNt0EaAbRDPdu/uMfd1yParhAw9MTzXLTDwEEPiqXuJkUt6m/MPoTE3uGxdPiz3
nyh2yrrG5fX7/cPR3q4+LwDpPMcWfKtJ+Z1LSEYHoRiBRZh/z/BJvvVVRLH8yk5WTQOQXxMjGLTV
BJsVxh+uHubAvqbh02Hkyu4TlmgV1neRmzj/jCNKIXRuLfyrCrb0DCngLTRej3ghJ5AmyBkf4RWR
OXl5yvEy/XVnzv5heQ5zD1gO5Gou3qI9G1XbEx/R7GEMUNQvDPKci3AHmsd5pVJw5PavR7NQqaZU
g4E672gWOoODMix15Tb7BEzbGlqWzYA6axWw7iiaITm7MkUkuayCtoV/gunF4siMt+kqg2Rcwj8K
bCXsMHRiMZI2TtqOuOJQ9OTFasyVAP0bJl1ta4iI1akckTgyZHmcSsDqXIGYdqJnXRdRItmm0dl8
I0H6TzbhlM4siGhSWQ5oBzS9BV3DED2FBuJKHP2bFcn8lZds6Pf5l0F4/RxWkmctCJI6UGPF5Au9
CqwKRfi3ZJgZZvn3YGPS/hXpxxc4aF2ihx4Xn6XEeRz8CiqanmG+GFJo6exLj/yNLAhttxNPPV9F
hUrlFPQWouCTpsP2yB/vLeARaPQG6QpMSsE9Ml7M+KWjHZD5HkKc6O12pXdPbYlw3fbqxtRkbmI2
p0+Ke1Gv1IsE8GWMCiu4I/CvscubhGIgtT8AS1NCqUCohgsUrNG4q7eVNGIUceNC51KSZA9mMqDw
v2/N8gawtZuaRPrB+VXN+5JrMSpJuolf0PA4skBTeSc+8EpCI+lwi6BA7i4FsBF1WPdtD2JNRSFH
fs8JGy+xKgVHXSGKJ07DQdWcsa3I2AMUYA+vSUkul1fBjX/rQtuQjF+NKkNZGC97tlpT8T86Ijfk
uXXk9N0hD6ubLInCAn6s37cjc6V5bZ+ruo/8iePMZGnMFtmSfcxjsE8v6J66B58Z4EmnvK5iKS0m
RquzIZeSyZFSBHqWbwWFznFFfUZMb1FWnYUju99nFQx88YBep9wiLd8rtO37Yno8brx0ZHF8CVqP
8XvrL94KC4+LFha7eNtoJKYgVQ6LcpGAcLUrJDTTAyYTvxwJfTBda38b/sHALsbSU8uLlyuLCqlM
K7wyNxWhScMXAOLKqO4rsCzAZoKbmf/xK6KJXheUSyXSqUpUCmZSp9famJIoeDHeMAkQtlp7pbxz
Tw2gnh7OZ8hqBQlCYBqrGz/1CpnGsEAjKNYVEnv2k7Baaqvuek2+rFFv2OfZmalS8ys24rIKPnVf
qfV7ek2QG3BocmlIpxXY7CKAqgHYrD99YtiOnUPm1Vl9HZErIBCY4s7S0c5a7JUbQBzBYipJ0cX0
eFzQDocCjqt2bVaV5ViGfA4Z6hsqbbEkYj9kA4Sq+OvQWzr6RiBSAh798BusPqHwg+4qqnrFYJbb
9XgeZ32Kvu3TXTg1IV1ETHLWcWjlntkgWdG7ObbR/mYA3uMIwO2wu6ia8VOamdcNEQhqaeMm5ziS
2Mi0Lf5L1nSR3vreFXwh45TjBpuFOlPBfUV1QpeP6TWVKgckW/EXzdCk9br7/iTH5SfvqHq13EAb
jDmy+pmcULKWJUBxv3kpsPm7EDxECxWEE8MwNT1o7QJ6wjXyDVThi2a4ltvAxSQbH1eXqARoiz/b
NA6k/QLuELHTG2ET5kIHxrx+tEndTZad2CYX4eWPprKwLZqK6/z6onH5sWjhkXIFwuqS6j05N66f
C27kVXgiW4yFDXGBmOERCpoLJ8+/0EZv1H0GTwWV1FgV2Y6j3eiAAeYIjeCfB/u+SwGxw3RipLHc
gRTN6XyFdvtdj+j4zxOYF1JfC4ca0UjrZLVFd57ETXVAXqqHGe6JO2L7EyepFAU3rwp8LGzZ/VA3
GJ2o9Q7HLhC9wL2Tqx6E6oyLg2KbVCfjfGwp1NnhcJDiyuCAzEN6oDDA2r39N1xlmibfOB+d5DtM
nL8wIsn08kO6UQjMtHtnmMPCGQ9InmSk4jWrfp+raiyOddkkNNxtrIMsCpLue3Z3QS8orV8q8HZc
Fubx/0pCFsAXQsfn0ZfpHiDxVVfpTeqIqlqGiekuA1OOIosJMfXB5n6Oa4JO9uQOZLwJjUGy5r0g
/AfUUWA7ulXWWfR3prCbWqLc2/hT3zrTrEXPGuBIBN2ytgiLGCjJb9Z8fuqLDWLKs18Y2rsPiMlE
Am+6GJeREEL/lh5vc5VEy9kOK19ZKRnxeEzNQVApv+wIMJN/bSyhkv/152N+FT/GnQyKfHZTfu1+
ilM5oHmLRE15dBpC7/F3XbzLmLaV86wqlGKZysEdIIpYej1NvuermtDaOET0U/DxRB8mEnYiLsiv
F8nY6CNqHiihwIzWcqn4k3kDLuW20XhJJdNzaOmT0doVJcD1xrfMAHaAkbbh3MpSRKJ/ukVxi9Rh
6EwHEtDyaIs5pGyeUpTNJwcdC7tWc5n2Z8lDZt3x7JAgqWUUk4auMsKWQhF5/ekZttrWBdZfSela
SdYjh9K7pNqL+WwPQyJQZM5z5lE5XwPGh03X1GJlGbOeuFeDtMXRflvW3hYN9yldpbhha4+YEbLq
ucEwPJzM/4LFzwyr3kl0yRSxz2/NmfQCE5DfbqafvLe72Jc0ksUcKYmeAefW5odtqk7mnNW+mqsW
1zjOMjrr9S2o8y6tNOU30He8ueLCg8lMmoAD3x7o3yV1nYVVy00id9+DkJUNXh2GxP+QDl+juSmn
uCFfEJvkfdcItSLtAaITZCZVdaCWrEOl3kPMDQtT6FiYb6atckUsSeWir4IRwnqHiBfi0zaRLbY6
W3JIWOTzG9JvgyuYlOmIEACrbOb7pT5Zs+/sZeJdHLani6F/k5Gf+GcucO048f0ceWKpyI3G4S5k
kCPfZjLq/6BTwjnPiQFQ+xEUerObZKhYSRFej/td+M3bO+mLS7Z8LPZJ+oxI8iIdEOHycFA2Pf0z
tfHS5tWOJ6SCdX1L40/7ptXGnl1zIZid9Xd2dN1uehuMDIHVmdxZOq/ulgGQctkoXJKBKPEkEAYw
zbGkIW/OkYSZfZy9nWPyBo4ePibDc7YPl07MDoUijZq2fHX9Mgmx6k5OvLhM/rRoRDSrKgEyTRT9
Ym83nF7urd9/jcOqe28rfkYg6dxTBGwoeYM4A6u0UR0GsPbYnefJWcAo5AO3TWuO3n5ABcRiqV/5
cuJnCa9gZR8R7IacYCnCHnPo5idaGA2sV2Xfl0QiwR683pFyVMgXDGQPvB1spN/AuDkxJ8CNi03r
lZpSgH+3yX0e++5EdEMaXzbloBqRU1X0qJjSpor409+Maz903XOTxmEzXqGhEu4o5Kxgps3b1yMg
cgBLDDzz6rnr+RqE8MQXcubl3L+gyZZA+oPIYliht/LrFA97wJJMrYblCxMru9O/hj8pdx90IGNK
MH7I+J8FsWGt60rU7rMHqXmNtn9NRZATxPxMAXByMN9MWXWmAV87Xh3FpPSnQrM8Hd2HDP7VRjkH
hz5n6JEWctU3Z+kfDxIIulHONhdwy1Y06JQRDXapbV+lTjMPO1pZ71nQ0nm5eeNsOceU2fU/MGgY
zwz0UtksUmKaqA6wI93LlObmd4EAXrRcJmJXzi627hnolO4rzk0L9FZJ8tBq0v0JrEG8om65FNeV
U60VQ8qYz9NEaOcr2V7QGsNdocGR1f1gpoPy7uFKW1SHBaT4dWFMGOxJpIEsk8wtBZYK+ElTvtIb
VxEoLAcaRnYDgvMY/VC3Rtuu6FAf/ixV8sMhB3Ltn0SMnmdIydWecbUvqCtpm/ImZU503TYvcMa3
fKNN99xiBu/RbHDoUr9c7Q/2xN0XCqg3RXQIOI+KYOLS37KyBKTnTFLCRmcG4FVFDi7PmUmGYWmb
ZjMzWBKqLnrHAFzYlhTCL0TfqXqgwXoRYh/OgAeolIDTe5dsOwATKglre4TY3DVGaRGaDHwn6QMN
ylUnrC0jwHCw07ym2lGdEf6faLlKT+K/QgmUEs5YeXWZz4ULHZML1N/uiHvqRNoan+vPRW9RGN3N
2M9qM4ZOch+iY2HXgBxUZHqT97+YHQNSLVJ17FEZUA1MT6DFixnFxdznbfi+O3fCpqfGRL8SmbZb
G1LHRC9oGEGl7uKwOuwH5yWlk366a6VP5L3KtvjnD89o5eOqjwyXjIKBrV4uu8S0huNEXGCSumyK
uyYqt0DlgXgCn2Mm10GoRsA+/XqCR0yWHnvoNGtcum8cUZywpRlUf4hrTAcmRx1gXX+ViA/oPYPw
DpVEHWfc5B7TEfqNcaGmOnhLAnR7OkAqLlx9pm7hAbEddQoQinrEeXT6QDUa6RRqf2bKP7yFrl6P
fBiexfVJn6sHsE6f4N8QJB6RdDZ8f7Npoqlz0UByILEQy1VWZ4EO+rYvyN0vbNei+y9itzUbfMgb
PCQ4s5mf2I5WkE6mh3wCG2utG9SLOpquto0OEXgtHB0s57VVpsUvv62EeEKlmFzuaV6hEfpcQnOE
Yrp8ZRCarB2GZnqfV/pjKK2IG4nLBrYiL6P24DRltH1LaaUbUGIbJ3qzQvBuq6D3fellYizsZ9G/
KpLCr1A+KO56vWydT1yaWnYnor2qR4RqJIEKxJ+8kGTShHjqKYNlrwt+JBMwVZDxCdqd003UWFwf
FHeN3aplH4BMYAtlNwhyeIDOforfRKEJWWeVXR3wvyH9vNQqXZ8PJ97rLvuVxNTAEumA2P+lX6YI
BR0QAoIK1ksR/KGyGxrrjZ3TFFWmAuDdEjrXyKrnMgt/EbbW7xhqISet5XTIT/vRKc7BzvgyxCaR
9yPWIPPaJ8OG29b07n3a5QcWZPg3DdjU1bcZQC3t1xiFAy6TbGfk7sf2D6DNah8uv7Jici+qqkD9
wzkf2k5XYUPWwsjXIkqkzZJNTsjtblJ5ODtgkXu/VYNbyTxMUcj0V4MQlo2EpDcq9YCIsbr4ZduJ
NT8cyHSb/auyQcY4lS7+DkciFxJeIoLUMD/z20tx9K88qLfmB3qJ2KMbol+Aj4NAL8/wsWcg1zpW
ShtrjtzzZ9e4FbiRQcqdkrdBdIwPmsXqDy5TREYS0DpzS+vZNUxrFXreOjbZlQWhJ5XP2lx7+E3C
xpkEp3pR/+QLxxhuATc8b3VNjWka4lzhT+Y2F9mWHAcSv/U6qK5s3/EfwlIXPH2jEByaqAiXf+kP
EomYWrubwVFcOUWZ5E6lppsSurA3f1ixwiFj3y/jrNo22Tgpw/fGUpY301qmIO4HSjzpRaaHpVLM
AkrPUnGfnPfb+OwYPRKw0OviIC1qHmqcVuwKnBgmobbaLa5nvDFJ8AN/Sl21ubbvFeM7+BfYz41E
EX5tDoWkQ0w4xD+tBViTRXqKP6YwhnW6lqyl3wmP6SyulpZsb4AePk+YzIwZal4h502dOuFCNrEU
timJs5ABmB0HSrsW8U7CH5rS8fWMOJVwrp9Lk1FXDHx99jbVhh5FEwThQ1JGqT1NR2OIio2uLUEB
kmrfD+A2bQI/hlaAkFQCyZaP43lJef+AAqGfP9PSTXc6hRQ/R++0zHyuZaglIR5Q8vh6ZIHhRsns
UU6ylYmXMlysQ8puhJyLxrIxM2k+6AqNosKxHivwvTiWiCs8qgw80dW03SSzuQ8N7lsUb/P2DORU
20HgWWozL2JiXOICsVD4RDrB1pftiX3qC+xI3aI7k/q6Pgm+i92d9OIskkx9OSP5eJCTHethJwnL
Vlp28OybFy5KOPDOLgn8FwjZfrkbvWB4bTwOopADypkJaYbByJdLVCct0JT42922VsUEKo1Xiog4
frkkA8ETtxB2nBOz2gioRfYoZo2qSL/oEa4JOYfUTYyMtP7YfnYsQgRKg92E3qLYyfePa4dT7fK3
u+stc6k/D4kwK5sBVVhNxokn8FZJ1okTmE9SFzUSTIhZoVATHzM/ebKX+V9Y+IOn8Yz17ta1jm2u
kUF3JTWo9YYmou/oB8DZvudG/Bv0B+ME9aXw3mCVKKMnAQ0g2j6o7+O+pCm6ANpxMggPN3ugJB3b
ou4K84itq07/Od+01poXFyP+RlmS2TbwWegKwWhhNqT9KTepHrtUcyMD1H2lwvOcTEluNVArCx+x
NkRR7JAAV2GWGrcWQrlYc0Q8mO2k+JgIMVASN6GookBOnY1of/Odjz2bmw6R+/7tG+M8ZkmBucv2
FA85VkHi/l/vfn1nXqNtwu97Q3w/xMg7pQH0u4JESZQILv8+ktIgaG9Iy7MhjwYPL4zoJ5HHxLaV
Al3wIJzykXHMnZd8cHEsBTCWX40cQjdHrR9UVJREalR+vuihuanK/0UK/STbtiHVx97WhRBFCMBE
YY66jM3kOpaoYs7nysBoVf8uoXoEfSC5KZEaWhSFrPdRm8ZeRzgl0akQew0bg3ntje9rd/uFo09a
xk2gGaqWcrerCmdCqaqpbFY1fUA3+++w7e69PyqFRdXUwSwmR+ECibbs97ph10viZ21g94ttVZUJ
C2e+aRbTZ0/iMF9q6/0C2YjZZp04YR/T4Oi2+05kfoLG3sG+t8+9kmGh5VM0J1KQg3rp8bAE55Bm
SKpfpQ+4n3AYjnOAIyEHA4ljfNTFsv/sheHyOXdvLbo66pDyTwufnfs34EBY/OQwp3KmL1LB8gYL
8y+Lf4rctp9YlOfOMjWI4iI80Ny0CCjyOGynsFrKAixwsJ1wEDmTcmEELRkSzL6OJaqR2jXLYcNK
VXLJdKxPqfRe8vF+RaZXGq9yMu6OmwOnjGGOBRgwB/kjo00C6Bv9HxSmlOPbnDwZwOFsVc7OX9hY
w8Q2RmhXrN9Bw5bvAXn8HrKgInFb/3k2PkoDkUEdPBp5cBQE2unLUUXFlvJw4VhWFSNmgmvzTpPW
JnfWBuZhh0hco2WOvbsaa6jSsnSKU0V+jmf1ehKvwGnTHpLOePQp4ZJgcdI19CM2VGkIPlY0R+En
YydZE1rGl3kPipyKktnT3CDd2MGAGQLryrdAT513SPTJpWiFYVnTx7mgF5guHBPfbXOgitv+1AEG
nCplmZIYSnMB9S25Mq1w2AnQvXSgdCRkqxRnLGNfr/51ZpGiehUFSeSnjnmHCSF4YFa6H3zigCoF
wFBUSHARU2NCTPC0AMflJM9YxkJhO+ttR/KbecuMVS4s/3NcDxMON5xs9V3UTDXm0EhyFxq7vd6/
0lP7izGXpV3BslXi2ZhRrFOcbjDNH6xj4YvxgIKIVSxZoSwQrn/t2nFF0M+VfpbM3tMnaw91LuXD
MmcG7mJUCTO5kSLszE7T9vhP6veoklvaSyjO8nfCZqPr9Ml1iWg92jgT/RFBNouU0gcnO0Zba0U1
i+b+CJr0ffVkkpRxUDANngWffxFPvhrNL8w0xjx/wcoeLiR1ITu+4NQ1VtMDrfXkCsnvYjcPDVx4
jWHNisSP6LcWfHBMdLK0iC9SUq4moyzDAOF8XYj8hUu36AeWc044g7Ag93lZhb2AokN6vF+dXULO
ocj56pPxDFBb+ijqsI/L6UROx6Ed+5a+qrjSon6PQHc+9Zz29/NnQbsWeHoieCTwuB5Mr31AB71K
zaela9BaHTWVTIvRdLTMAzudcCqL7Irydk/+ecGzjz8LBNH957kWr+opvthEjRS/4xYQ3Bzdc3Qk
oydvpwoiv1l9UYJVDrqJcTmETdWlEdMW85G/rbHHeu4rCtnMKtPEPypamyLjMymRSb3ejwkWATiK
vQlL5AUf6IXpU7Zle/NM1t/Wlq81jtWN80L//3j3Sk2hTsZK9GcaTFMWECuxikHXsOn2fp4jDuBb
p9PTtg2UUZyilJo9gvinOS7TigsysW+KMwp1WDlEXkZe5X0JMP5PKP7yAuH7ZSMu8O4km7T9RGMg
NNTDCeBYXST7rDB4XeVjoS1dDkZPO2qE96XFPj6RklXumHLJhcYVjvEXczpKIi3iZ4Yiq+jQLDxb
BmNjQhf36RZAY6uf4l7Jqd6QzDTCQb0XBm6cI4r0YMzbOlbte7xEU6zE4E79HZYffEczoP6PqCF0
pU7fQ3ukkiVN2RY+kr0eBd14aEryzmrdDcdFs1A1DordK6xUaELBUNOhbVgZIq/LQl0RPBWkrQL+
vPptQclALcTR2C/USI1mA2kFaL8BI9fDNFg9ZQb15Dais0nNpuNFjwJNslV+7fII3B1bwbW/K9VZ
Iod6yc2WM7OWkJgjH4VOg2gGebUWUpJbeNEzl0z2DZW25S0SKMsXeylxqLQ7m8r2NtFfMrGUoVga
5BcmnEMrPdHRDCf+32IZhuxjvv+iRshgrTms31IgD2leWBqEX3C8+MxqWnnZvwLoXtbS2JqTHsUd
nZkAJXZCZIP5XkNXtMROdoVXVyLIAeNaHhJ05wj1IhyFMEgQ+5eFMaPkj4K+3c12ndVlhR/CXj19
lC8Ybi6Bhs/NJbKRKIsqJX0eLZ+eJRth8S9eE8HKMfrDeFvLK4+3r3OjggGJcs7rzDNC85DeHMR9
gEBns7SDIcFXW7WepVLP+ge5Z/ZyBccXjEg26xqLSejDLyxy91n8wpTo9Xfk6s4Zr63mVa5K3yOD
x3ps9ppne24C2XT1q9vi/SOM5c9Qh+dhk9u/41luQn0RZ1cUYuR6V3PvmMyxoStFGZgfoRQZyaIa
iGdBFSV0dnZuZQIATUTgDNWb5JUavFuAdFy8DVkOjOrNFG15XAmQSfZPtbqhtRfLL7LT/+YVGouP
0ako7+622YwuDGLSCv/fNnDAWgSenjrF3xyeg5GS6dDG5kX+kPWC09tGZiBJbRqY4RRs29cIxSuC
2Omb1Dz4k82qIa7S+N9l8s+5YKdedIdL8qPXiPTIwJj6vIODP36+ga9ZyobK+IGPqUchv1HPKvK2
YUshGCWQMTQGuDtER8JL+kuFQf2fL62PA7892hPDc1diuyw/EUcpQqkJjzComYNN4PfoG4zZnaug
ZGovNLMi3eNj69gemD5516YYKz9NK36TRiXSPGDI/PKthday79wUN8sp0lshNZyT0vr0/a38A/nt
vBRJlOoH57ZCW/z/Iud3ZIPqk4ge8owjnEYcVNkcnrkTAF9dDLgQdw/hWkObOrpFFk8E3EVhdJBn
YihsEXufqqN3xXbjPm3ptmIUV+4SF6kqGjBHV+2PZjJw3K/R9iUsya+Y+yi+f22cFEvk7SXjMzsv
qyBWxeFWGCyIdZnWW9D5V07fVlyH7l1NSAASISNIAteXIsd4o+kj7iLPjEQeUYMsnItIeXDRajj0
aiqyXLymi1xYWeuZSixFho59ZZBBoTo/be9rdafCY2yZlMTn0eCZGr/LRgDy2rFiXrHEUd2xIHdt
ZaUNFGM1d2ybLIjPjqrPMBxzkM9jd7ZiU9isGD/e3RN/m7z7+VyLEy7BwHJ9bITGCnWX0VvZALX/
6y6iRrfn9naoYZWt7CiCp6VG6D4EKQ26UJvuCCL7+9LrRvxbYJgk2NDgdjMh1URx7FlxD3y8XLH6
kMv4Iif0fC11SC123mLCFjNav1CPkZYeuwFmmDOew+T3hnkin8+xP1l/NYt7Rgc385O5V2lncQyI
moC2fPjYeUfIDKzNGY6dLOYCKjZlQp0A3m2Gi9AV5Hj0W3YHU8PZPn8iY31xpdod4qHuGYpLvRwb
1WnEz1xlRF7sD3nZHDKOKNTGWshatBPLtWN9+er47HPfCuw98q9Sonp6C1m25PxA7wq6bxYc4+hK
n//CET0GJiIL/DLdFbc7NSQ5q50AKGRZ6fbXBOpv24y2Grc4gIz2X+TQ2ANaEfufQeKeD6HwEra8
gpjE5HpFt07f7Xi3iDDrzorCNe2mx3syvZC+ZWs3NrgYbTSJbnvw2aAximFQKGP4BVmUvKQP6SVQ
Ydfa6afw/JGjddhmBbIKENHK5ryzq5VSK/b1pMTLFbaNKnS/w+ULQ6JXXYHxArkeSFpOqi7vFo+S
p87ZP5AUz+cp8hRosMdXXmcU0ZEtP+ydjjgURjWufOq60GUiH8Zz1rA1k0VSE+Q/IBQ6Q6Shx475
hZLl5Os+4+5Vl5v1MrWZ+vZH7ZSkPZNaiv1z6MMQPrw0ZnEWrqgeCyxVqHwLfXoI9XJAR2szMn7P
FL+/3GZbeWzypnY7GkpUbieP0sLPy7V9zsN5dBIqHl5efomrIubZL6lfPxb+w0g6tNjq7G8JgXaX
v9U5GL+PmlyyjxTi7bQtirDbvxd2pHsxpr4JPwn4Pk3BzH083LiDcL1jMkC6Hc2pPxrU4Hp5Afc6
cdfYcH1fbTyq1heFEX/iGC36Ul7cz7Won+l7UF3t29pyfBpont/d9DMabcrCkpsvNg6hNZL7loZv
BW0rwABOh3pu2QtdkNzOQpndNnovcTQKaLrPpsQEgIL4C7hu9iNeKjqf51NAzwRBuSxshlQaSHsA
5jX5Qg1DQBiT/cAmcv8eMLw7RKzJNVlIxX3ykQjDZLxlAZVM3i5Aot32MfoRVQ0LL9d1bdHdSh72
bTpohnx3Pjb5GzADtuNAhk/kpBBjdE0hgluLmbBCFQZFiyWYb5PW15kR19KqDV2GrxTKUe3a+0/R
7nXv+aZIaSmJUjMq82pAMhDZiNhNMm21t7VkXiLad9yTE3k+V7i3Mpy7tsaM2ZPcTa7Ua3GQeonB
xY2OTWGRfo58+47e0fUAmMj+kQvB9X/Nr886FOGHOBbBFtZ4AO+dTfVP9VxtPXiEugZbnsX6IuEH
LNrh31XJ3Hx/CyxRFvhTwSJ1gFg14anuz289sFRqLNXfuLtSdSWCoxebKVBi4GgSBJLOxPUzcf6e
FzK5k8f/H2aQ10WVwAFb0N1d1relvlQq5vpSgoEDU0vEd50UjqIU1PfSVMdrrMz+6RGRyNIt3xuO
sE1AzE3EOsYjm5a0XlOj+QaRyLCGoeH6vpKbelVliNJSm2xBXu6vaWH/Yi++BVTJ/FvPoMCVAhyZ
T5oBb9TXClXld9Sn20aV7Svj5Eh5XyKjG3dtreqQ3/udGVvrRfJ80m9DIdrdqSBwxrpPG7B45FJ9
XydVG+WCfVVsuuWHz8Vfa9yEr5QKxVWGcUffFnscGPtI22dbWbSY90mz7SN+NF3fKFU57mb2sYLs
F9dy8ONj6kdPcBb1bxy0ylc54zGzSm1Se/Udu5hU9Yj8AfvLzxTIZtCRChF6beZusodwD7/KHeOs
XnFhdVG84ZQk9oKRL5+2RHWnCGbfw5yaxO05QQwvw0L4p0iARklUfLTzof3x/vldOEjUxHmD1zZN
LNzRPojZ+Agh5fXBYDLM0xiejjxmFlvgCKVFn8CuLFAj5XBwQwDRiK6B623qGB8jxIhKd9svPZsk
Cgh3iflYJacwKMfwGjXNmpqNXLSMsWlRYgDE0MR8kU6A+7X/NMgDtN1JPzNwJcv7ElVXB/TBupjW
fQ9WP5K3edVryaQorJKre70S9aSwMAPPQJizPjLUpngS+azXsP8CEODn2p7XDo5sjc5y3Qcxmg4o
YgUP9qTze/UySwYs6qTx0UJTZRB+SB2n1hJftrWUaThzmiVMoSLWc9dMWybChpqQWSNpJSxDqmx+
5Bb5Va5HwbUYvP/q+X2pFvzu1UFBEwHIhW5q19SEkM5gHKC0zDdtIJ/lvhn/2vKyFp7aHG2pV1yF
Y6UuCUWq0hWOtI4+Fxvrc4j3WO4GRqbD3cFIoErxVs09csg0Rx2ezvxMbz19AG5Y+xRohZ92oq8V
S1Y+WbHPMFTu1wuRTFDbKfSk3zd3ZQdLZfVSfyuSTxz8JyXdtCxl0ahezdzkrO2qrTwWr1OGgXqe
YOWb4vKI5d0lDN29B0TrjW0Gy09hRsVkoloNNKE3WhqYqWQnIOVe/KBwJeSbTJRZN+NqGkcrir9B
zh6rIEdT8M4JKJI1LRUqsM8LdaSaRco9zqVBj/sFUY6w/t51g2hmtnVPRfNE0+F1Ymm6AtOO1tlV
6onbK7jI6n6A+l40hM9B7ihjO7blQ8Q43CrDnqA0EVH7Fv+SgkEtSZBfuVL8WqYvy8T4of/x6ZeV
hxHGpQ3eOVrqm0572NDBLOmBkdveavt0ZmnaY8PWd102PUwUuIkdTjry21Yj3U4pao+QZpyqw3lc
ss9WYbHYfIx/YMAJ2BBZrAVXPhZgk8aWxPe65iyCf7N8zAT2aK8piDzQG8loc2Mh2TT0eh2C4IQ1
0xtNgDSZEzwArqrM/jh45V029gdkxBH+Zh9m9nOayCi+bMZ+rdNmCu6zvmfiaF242OPVtV3usctH
ULVbtZyClZAEivR0bLIkGaC+S7lpb3/Szpm6sswFAhFg3YEjIBiNzpnlIyUNU+wAes34J8NymGUQ
oHGaxSanFOMCWrAzemKW1/ScL7gRRCElWCsqWNuIadEn3/iew6OxUjmfbyFL+QVuT+z9iNFXi3Q5
tejvpTVd0P7V2rywWqXkJLpUVx2Pf+5arPAy2g2svw/k7V4VUhG5NqoKvRdXPBR0OOgvikpy2W43
nOR9qX1Hy/Pp8NoAOJp/2WO9ZYAR0dsbnMgFDo+yP/CI71ruuOKuXUx1yNJOypLLwbgOOZ0AAIvW
9g0kzVJEiooTHuqjprkBYcAR7GAcEcgcLX8S4frxNnop+wqvVAocEeRN7Kl/KQibTdz0NaSpfnqq
xxYdHu6l2mX8qSlDDxlmwclUmWQuE1+zlWt61/6dhUA8wf4N21nVAeCvYUDysvpY9t2f0n5x+fFB
X6Zf3F2eamuKJ4iFgqf3ibfvmd7wT5fBxOanssiqzIuYOJkVPyz9t1ZT5zm60ldj+SuLJTiz43NY
EDHVuLiMKv3OH6yuI2EKHSWpAkGcQUU5hAmEc+qJOY/jWoMS/V9xb86gJVnsNzjcC7IWVdaBmJ+l
TjfEyTW/yzFg55raOi5NQ7lBkcTTpJR+S6wP7+DfmaIhna82OCN7B7lvNeDJNgprureKbjAZBiCs
tCDfRtvOd0ZYTWq7bNeNsfCKJDkJ9nftKMCsLo+uunTDcUEa9KhCEuLV4xPRvkPsSxQnolhza7CW
+0ZY9cdHAVqswJl0roPVIUMr5Lm4bzHBS6uOCeeMxIebiKzHwyAOCelepQqxjaNy6lbT+OninxRo
EYbbBLIAYghd1vltfyarIHHHVsdwZVqyppyCc059CVhV/+9YJ6j4HdRCTUnaZ0JxFkGDCLOcDZ3K
g3BsfJ71FcqML1MhIx7bS2leOOoICDZq5xjtXCPFytHAB0/2lXVTRVd8WWV5PnKzfEtUCdGZFz89
CxzbG4MLt3qP4pn2zfahCNqnU6CLMxNRo/MQGUsJv0LGDSS3bVCY/eTfh8WtfVsR+jLqCJ20e30l
b69nQbcq91KCQp8UkDG/YlCYpEWF2P+9Qv2q1/baVXSSJPvFdwbKHLiUX3/TjcQSZVSA940JBjeB
K4ASmfhJCPJUDRxzpmv3mvYNu4GF5aC+llblQ+4EzSirkaJamIi2JFOGif4n2TyQsDuAMG9QbcSe
ud5FFcaE3nhNtOCSQetco0dACwVi7caXH4B5C9DiD1Zswvoaaduj5YzdRKulw7q+Bk/PhCyFMphW
ZfnCrAZkkuC6o/6cEQ+RAL9ExbWKl0yous/PhPwh/KnXJZVEKXCN+A5dOJMpS9xxXdAMAJ/N5kWr
jiWuWFH6WIK1ssKm77uWRLmVOeRZtrohstXsEwfoZrODzsWvyuDBArqWUVVNnpXzSeSpthcCzkXG
L6e0fLanPNWqtMG8ejgHCk9BfCAn+BrjZjh4aHx6CiNlXsvtb/nz2dC1a2YgFx0jNRFyBp+8yPl6
KXdb022Z9aPPsYDuI8pz+fIYPk5fG+80paKFiB7NBksSRi79yLXNloXUMMH/Fx2CspeczZ+Ml5Wi
5xTI7aiV6b7nqZ5ebsNhS8oiRa2I5i3/xImcWhA8K8M7ISkgojdk9KqmTxzenV9Bghq/j2cDF+iZ
hfYLLU4TvxA6e/aMgnfCWcXPo6YWleZLEEIoJHY7kz0pw3Fin2k1BFNOlQefHzrRKwnqJamgRTtO
AMsCYzmJp+SWpTDiFv8X8GrAfw0DpZmA7f0dNpDvqQITWnT5x/q/FC9TW7fWPilKr7eL0TXHgT9j
AY8XbojgjF7cXMeiUli/CrpjEGIWuHlK/syzT4/NDw1REErvL2yBdrY8aSTfTEZvIoPLOkBAhk5O
hkp2sd7gIZeOwrKGWoroW5sYWYwzPLJ4AVgnO9HZx3RjArpcE1x1SA6P3go6T0GL0yUEroqBu0tP
yVq72PcDTbtJSvrLpbHr9zPQfcYFymX2qzr5I9HDD3ZPJlCwNTPrthDpjEJ9TIlZ3/iH2/+FgQm1
tYahF3uBcoD7ENUp8sp1ZzXkhGOB/F0NNDCrtekcg5QANhGNYubu1nJ7sEUN58IbsZlCQmX8ss/n
+k/bEeomjnk6KrVkAG8LS+CGvCYsHq1QqDAUVJlM10FINjmkkznqLX+eAkkEQvoeHr8jBcecc7J7
S8zBXkb12N6YWzWa+PAXzAF76u5odtvNfDlGCWzD/9JxMD4iWWhxt1UDu7Hs7ZUNjCUYrRRCEfJb
fOi9MABwVugxUl8QvZXIzJRkb8TBPI0Ui4lDk4mmcPolfXLl0mQ3guHFy4SzCc26rmfssYPKoU6v
LXwZ7O/IAW+B3Oh8PZRwmvqNGrH8O5xjJ5HYhNm/NywvJoZl+p1Q8CsYy84OnHMwk63CyeCCELBk
UIj58YfpxNJRGMMehQW3b0ZYanxKnUwnA8eMsRxT3deAREznruSsPFqJ9KjDKIo2pRGfzoZ0o4Cy
Jw4IP/IkrlWtd9HhFuBDZtu46DjpKIdtiKeXyr5/I/WCgRavFZcQ2et9TQgKs9TQzntDrLUfziWJ
Lxre9QH84Kz3BXU1QmHFdpvbTFsEZze4K/oECcK60o6Ty5Bx9BIBkuJ7owx4cTrg+iwG84jXMkja
in3Vyrdy8gDDRSSO7P6T4YLWRML4t10laomLnHhKb6w0TfVRzrD5KzvnoNoRpIktM+geBDUEq8OT
yG73YLKqBK8eadguydJHb/oy2/7t2nbsOTk5LiqtR3dGosQczLsvjnRu2+tLYVS7TSQn3DApM89d
uziqowRYM9XHiCmlOlenRwKajq1YTMqLirYuPkoTJXIGOQlVPZHqW0Px1dzUDIzKgTCc6MBhGH7S
jE4XrOc4lOOZ/ygf//B97qwQoHb7yUd/s2W2bd3/uGJ5QelK/SykaPQbH9XZvlZY7xBTGUQis3f8
oB/5p9qLQwxXJ1YmjexB7dwTE263XWXjDVE2CKxcqqoVhs0tjPKGdOuuwpNqSwEcqNAuKxVaBid5
gJqxRpVpiNC+DnObxdVqyX1xyQ4P7CQ9/rvWfj7MFS6RNh1aZ8JDsgdyBPd0+SM/d7AFmD5eEcW3
jv6uEzfYgDreAHkNEio9Q7HHL1hc9DsU4PBLtUCC2zT5hJoZF/o7n/QzMNdcZ2hpZd8zFFafg4aB
yZufdYEE0w3ZfevRnc1jctFu6LWY6w5RW8qDleuskGaL7Nn78UpGUG34cJYFED47D4eARcEwaAWu
Rn28MX6d5MeyaQcFEvU4KJAZ5k22N3s+zEo7ymanI3ZA66xqV+FMbaICPyfgnv2Rmt2DNSjVFLj6
bphdJQcXT76XNYB/6DF83nOWQJReQVKQJLKOUyDh17s/OpMTwAb1gOGwngUxAfCN8MFYZ0vJnYno
ACm4GkVnI8UDsIgczFz80b0pMdGLRBRhNixBtXEZX2doIwsINm09npYEf8Zt3E+gniXez+G3/CGB
5186PUOGPcOjvvXdOs8lvFlZ6mlHGXGL7+0nIHWlkPUN3MAS/DZeZowEV5bwXONP6Cly+vVp4sNQ
8ikA+yTzz5BFwFC7V2fsgYlFBNrnB7pQzH2Z+1sbfrymG+PsSz/NwuN6d2cPsTB9Gx0CoagWfM+K
9p1qIvcsP/AoCvtQOgqb3ircJSJ2UggZQ5KVDt6DD7049s3GBfK1TPtE/BczxWY3XF/E8RYRfsxs
fpwB3w3phzXgPTpumQ1BhY4I6kCSGS6enANu/N6Q4TS8cUnHoFDSQVneIWC6BzIN0p0jZ9ruobag
X3jgoINWFAg3SDJiz6mgRd821ejTQvWVoD6LV7HzaH4H/bumsroVjcBa8bufH4EGSLvny2sv8pmP
1x/2AvdXI0/qnSCQD6RSHWOJCPnMSCuKflER7Chy7WMMagvEiYLW6fW5o6KGGN1tZ3hKiXVDdaIM
KGFFWYtnLPNKWWJtZ7xxERxRQHOkZdcu8WvTzHxZM89g3kVoCxrk1+mooidkWNVC1F3feTN5eJs2
XnrOmfyNJxea6LOtWhATPRFYPIE2S8QO/KKfUvr+/vQZL/BUSSRZuSDJdnuZJZI6sFW1jKIp7MEU
uiG9S222D10qHBRUkd77GgWPdowbWZef3W5GjE06nFRLcKJvXrJ2z1aljfATqLgXofkBQIE7SUar
slb4oHV0ZMqu2UMlpGwp9w0syuBBNrvvnL6aDK9FKJkcplDicWY14uN2mK+q76nyJoWgC45w4VIJ
bBPsvBa+5BybBLSDu/gefURYEpGF+/eNYcxwkjApAccHYt6y8wfKQO9idqdJnOaPmeqMJ8rm3fiD
TiaKaeSiMvkcoEPRATGjnBOm0SKgqH+cVW6LPsUtfRy6w2JX9mLXQJczf5XMl2seksqu5xlOxgcT
9ZoFJfb3xfgnZmF2cySh5bCpcVV7It5lnzKXrKoWEWNzvv9PB8T/eF7eDNFfVM2i1zLqCQmckixv
geMBkXIZ9GKMn5JCeeWtoVvkjDoOAFgTi9FVz2xsSRAKJjb/OiRW1cWukh/Flj37HN1y7qYKG1eZ
IRQhVd8YSt+80d+B0QqKA1QUy6jSFM4npa1aTgilMoYrNQzSMUFPRI1TrWXotxLDiJI44qmaYMDy
Qq5BCSgAF4cx2xlcCcSmjQ1WSbrbj7Mjx1RlG1tzX9N3v0/DcvZgYcCovJyw0d9IWdUqIpQ+59lE
qccHbU5523UF21q6rcyhQJzdWJtff5K8wFm4sMQSJUYRNDOwiWYr/CHVBLu4h7CQoFeRYRWIxwPc
z7H7Q1j43YFfozYjwP8RkDmUVnAdnRaaUWBG6nmiRtQDfk8q5ecRh0AmCWN2zOurhJ6aXizJmE/F
mp2NHOP95iHHiVVBJBEuhQlKhKHpoyAFAr1eVphbus2LoMcFeuWzY0TOU4chCH+EynkT1rHPIye8
3b19hA0a5LiauM4cFMftuRftMUHCktuUtpbZEFjh41VFRdMoaef28+GpIBA1K7ouZOYhfvY2kXmo
sk/yM8yns5f1ZdxkHrGaTNjDmt2SUlfyfuCKBN8VcUTOr8vSTztIhap39kYTRCQW8kVMIHVrJXl0
vxdo2bhnSpfZxItEY3YP2HOBbbF9lOqicJeNFLAE94PIlEXxRaXoi9zOssZcXAnLuG8XrnPNmVhq
MGh9mq7choEyGqV9PiXpYL7jhSWcT8Oec0Cm/jcluGM+MeLntrDyLDTVA/IJSEBaDwkkVsDUB3XW
VHb5i2sb/4BGLpPWCVnL68Mg0xZ1P2gGpt4AgPQbtOytmZEd6B+onj6iY2IiLFUA67kPmAtV+HdS
oZGKmiwyCot7fOUWQfdPK7NMSV8u9p12zSDksTZ+z3eLj+t9HASyo3OdYkf5yzAjCZy6uhnyIP5U
5L8GrkFZNSvf8BSLFU/g1SXzGTjkFbx9FTWc6YdWNvP8A1yQ1T5uNP5vAHyMaz7rzKpXHuabJOTv
Uv5fZutxmx0zDgAUFsQp1tkQz3z6Bli3/Ag9fsjo1cpABJ9DhqIT2gviM5XGxaNQQDe4AAjlzwz+
q5qnrTNVX6gRcFwiOyTJVSVB+w18bK1Ki2KVXPheayNccywECNCx5kPYvhX0Pj227+EDzZuDs33c
xsCj2qsEoAOb4O8zubKc9x2bNuPdYmCU4iN26na5KGac/C3E7OHimFLRqTZuKDMB8WxjCxaJ3v2i
s1OA2YktcAMB4rb2XJgVhyv5Ds+3vBaNl7XI/0XxeUL+aAiIYD8MRJDRsl3qG470KOq9IuLVHYZI
xQn+T7hvcIszFBCg93zsSmUBQjvCR54hSZdaSLVZLy+nhKaCECGSLOAC9LtX6+0poqzTg7lCLSu2
rDxRXzomT1pgwZdfhmZMLP4u+vOGklzs/4KtdRD5FkshvfnHioH15dw7NM6mmfwPXi7f0SfbZ5rk
4Qu9l2waZY67qOJKVyV12Xq3vi+zvKJj0w3cdcpBvBvFPbzjbT5q2/yKZYAGH/a2rcR3NWC1/wCN
KPwyeYPw6FtJdIqt5uP0u/56im96jQl/7ctd+ZYf9l9HRlIm83oAlvgVBg8lR2iZmengkEsIg4jk
d/4CTESM6Y6KWK3lu2xLb0dSBGgZe414DMdSRgUwymm017XcKDKYNcPnj8hiPQxKajI38D2Rsv9r
0KCfS7WfnsrF3h+T0Rkc2fOiWVpt2G93PlyI6YQ2MLiPuJELqMsD7udnqZ7zMTeyrfhQqLW3v+q1
gV87jYNPJ7Q7Fnf71t/X21GIwI4D46+NM+I1VVeIYXIrqxEyatLs21hFKDoo3pVdUCUOBEgjrf2I
2sinAPCCy9NXBmjMnnuSmMOYrCk1GYAnlAsCkBqL09c8lV4qTDTNdNvTxqHzef7mPxOn7HBE3RUh
3PnwUrJwFQ4WeUqqqrZHxR7o9GfcAbKOJrE1OIASdNm414l0TgYcBSdZGBGeMVMphy/M/bVponb9
C5WEpmuvppcD283O/4G94E1Xsw1ClWVtXoWAJBeXEdFRWdEj/E9lGUlYt+1usG2tYODq0pN1U/vp
l8A2VErrmZ9/ev6Y7zfrlhcFzprgPv6tRJmZxYuv41nTt3gnmlt/pXxI83CoxYJ5mMNmxK+OSR7k
0C3WD5HfAgTEdB1hBVA8lnp9h03SdxeWSCYgok4kjpTFid+3i8aBCMAXRI45ZO0usRr/MwlfrtMK
c4tEaSN7DDFE3EqsF7UJtUCa1SZic29MY0RPf7B95KRD66K9ORJR0pqVW4OalphzWaV8A8AeBYm1
L8RxzuDIH42+Rblce2T349AtuT9AZWJ3cgxveXz2Dg7sbF43F0ITykWAqHius7qTCzK5/O7112hl
h3PQA2WDdtrRX4Ywg5Vdv18xOh9DKI4Azaa/70Rz8cp955zLgq7WxbdMbu5fIme5eZ9ZInqMrRFZ
jrDO/tdj9Dwj3lKyaG+0++/q8Qn52veDgPSfskbbZBa5xwxv0CrJNE5UUyRMbaBOuKIXy11DZC2j
d5yBzT1Vxcl8Wyfw/VAH7l1VSas/rjneSq6TtsKMbHCqcSEPpN50xdKSE7BoAeWNlOz7ERsRSBQx
5L18sKaVQ3ZriEvNLJExQbM0oUp5qYe3IcoJg6vWYhcW9redfjYIJ7pkXXQxb/XEB2RQBbZ+cc5i
1iznLN1jMWIlsa9DVMzHrKQLv99isd0KqcMTBjRPT8eQ/wq7HpT8U55phAVm8JQoqNUWnAxe1Dh4
PqquSOxRb5o6zzFd0ivsIODkb7ru3N7U6qfc+tBWh9Fi93sHr45QUmFBgkEGGurXAEwHgURo1iMZ
+8A+P4QNg83yxAEqXibFqlF6fodN4lxNAP5SZVEv1yMX/Wnwu6Mel99i28dpOrJXrrZQn70uE3gp
5Bd2YlFnphFbGOVmUNgA4I6MzuqZHFEmabiB4ccwBo126PKhZwLB9CKbNNzgRljuarRQ1epip1xm
OGbc/ZydsikAxYEj0nsWbAUXAAp2ZE38RCRSI29u7ACphqAaodQmxb8zvsJdSSRkIIJRFGOIsCLN
ryhRcP+RB8ITOJRJk8GVg24RSdNfihS9dR3H8O6K96AjwuV6Vhe2yyZH/drB/PnWqTP1CdAB5Slt
HjbrJussmMvsF45lvvXLaexC+hTSf8IIdMCSM1fTEbQlvHh6As5RZDWNz6ftLFGOIOq0PsOU+SG/
ZKZ4Al0hWzo6nAfJs7aFBFifL/r4ycVU2vg+u1qUBGjncVsoPDoDTSQ3jayHgRFzF+xk244eQ1Xy
OPwIQfOuFq7bppJAANZI4sPFnvereF+GtdRcspB70QzpPVf2JmarnfHllsamIcl/IY6wxgH7cKl7
QEeKn0nDz2RvMZS/ZzAEN3TKEm1ffblnmL2IUezaP9UCPYsESe+h2zh8W2yX/iPOa/M0U495FGwK
JoLoLN6KwrBl1RRzMCyOQBKmuGeXXV5Jyaf6EuewxNJji4xtCW+lya0HJ+N8gUCouBirXfn/jywS
3CTsbDhZFfeUPIux7lYyUZWiBQeI6vp3aj6lWN9+l4j7Fm2GZ46HSmNZDaRyr+vqYnwGxEIvNajJ
oyo2IrYlGcrIoDA36jxy5T3mR+GM4iJvPyY2gRTtvJIJGL0OYl1CvMdSoQNDStncMvGG/eLtnX2/
2uZ+CqZm+nYDJUv5EQsQ2wRWmq+5F7sSDyH5AU3uEtWcUlPbHQBCT0MA8825NM3qF369qR3uBBTH
WfqbfSL5FRf7urZXDkzgK7JtlKl9O+MolnXNaCT6rlcgEtw3t5R7dbUHsM8OA/6AJlPO7zt6GEpY
lgdoFKeabxuuHv0lQRDM73xLGVuK710hmjXKzhfbP2nGLXI62th50J5vQ8Pmd+BqEnhlv3Y99gcv
sZFyixOypCxnt92tx8GrvCpK8hB+ZCfpNA7IhpcOKf9sd+GNbMM8vosIMkQJWZs44JRMeNAmH6++
1BhAE9AWqRchKHVvtHg2Qhuy9hmEitPLiO2CDSalB1lb4DPKcXwKSpeKAGN4GasQgum3KpxUOwOQ
4LSVs18E1La17Bf3uIIMlg61SM122cNyTjZx5G94y0wGa2jc8VHZ4qZTVuQAbd7Czz6erPqpw3j9
GHscbUm18GaGYZrVsnnPdX50WTGYeuwoDpy7/ENhodknqLu/RvOX3eHhGauPTwNc0Ci1ll5tzaYx
u4wfnY0JZBrqAifZjFATFGOAqRIgQjtiskoZ9BSF5hNHKiKlcj1o7G72oA8j9UNJBW+TkgaroIlV
iR50gmztzCb3jNc5WzQzWJHrT7hxjUhzFavI0SbrVDGWaDk4KrdWKsS2W/q7GEA1vPZHGlKPv7uj
TG4qbWOdvZ+vfdlwiOIbFfxcgzFejaWPqQGjRdV2cv060w7WCy8IMCusvX5Qg5LB/Hfq5b5CjDXZ
gF+nEJeJmNwVcgKEggWMicK2pQ0GdAGEVGNbC4o6y5k9x+xe0GSxICQhPNlyRGnWtdn6kDw4DW1E
D0ThcdQ/bM4W7IS4RaBZpslMpcVfzt/yFbgyfoiVcw5DTaPHOmq8hIpUgXiT1czxcFg3AQOREmeH
ZEjzyWONBmQxUN52og4hhPTJMbvzqEXEcoxh3xwoqie/VLwfoPTtljaSO7aXDoNtg+d6D7ovjqWk
jWUP/FBYtr9fYLj3G/VspePkAGHFKSczotYYZCI/pGxHZKMU4voNcT7VsihQyqQNBZKcY4X0bYDU
t302ox2V5heZMot96pxHzvO1hEzkK4ZM2OhMYwd8JK8qMgsBAaTyp1CSKDqALP+tlxuO0iMhn1fD
p5tj0uyeJZpj098fEp+YaXwk/stVoSIWLn6Te5zKHACUYGb9p2e0EDkiMSWuzscFhbDSHbZHuqeO
tS6FygU2GYIrLCU4xv4J+6vKme4RtfOzgAcbKo/rvdEY0L8A608V7ZVHyacZZSQwnQY+roCwXsnx
WJqjrP626quY5DFD3VdCQ4F21BK1TmWoZ5HDockEU7Vy9CQSXc2UlRcLx1cMj2AkVWm33sds+Mg4
4AeR7BgOUHyf/uB2XapU0c1VIozOAoy9Uo4NdoMu2zBomwjyrwNDV+PWcy4YvepWK2ZXFzWea279
ddl75nCCyc3fJBkphR6rHMjz8kDBJEMd1IJ2dt3fkrj0TybS+YRQizrKVELQB192eM2InGAOuJ0F
hsFLBSd8Mlz7DkAjRNWHrNzx0e8AAewKd6sZnBeugqfAgBpe/aWvcjMuaOTByJD53b9KlSaUPryg
tLP4bWC25ce7gx+VicQtTSkzc7EGqI/B1aYFEDiQ80LKEkHZsMmTvXrtF7qk5/vVNWUlHGzu9d43
Q/DknYr01+z5BJGdUXWH1fKNt/xUPze4PECUEvryHorfZTuQlUEQUd7M48rKpun4bIbF42Rd8J45
pVMnNnIOfHHHmidIUyB/N54yVkTmWWRAP8XVP2VRCGFstc/aoBqrPmgXMLel73RkFQTK3VOLP8W1
lnDN3/Rtz+rleIrQETpLuC0pXdQEzdM9b+Pg+mN4K6INZsN2bA5cedcGfF+nxgFz06t+0tiGh2+j
Uga7J/Rsm97VMVrap53a257H0osxFK7Zksy1HhdlwFn5oLzQ9ZuQMqf5nTXz0LwXfI4O0WlYW9u4
sY6enBX2A4rVV5WWfsFEOjRrNsB9L7bvhuwxRp275rMzY7ibTzbNe01Ijr2AW9NIBeNcXlojYqp5
Z8a5UJo1JfilpqKoHStHZ9RQFUyRcqs60sXHg1HeODCJBJUGFnUEBbZFfZc5lPD5ICJt0h17ojvz
EdtyAn0lYdn+3psne3ZyQuia+fI+rCFOAj7YKWAcUF7dEq8XXJaYxu+TpD4k6alT5SNSZTBlpT1E
2JuPiUSDVjo7zN04SsMGGUP119S4Ra2VYbPQZ3KLU0VjhOdT7d3GKaJX+8QRJxfwkvEkVXd8hNIA
15uyupVfpI49cIrL4cgYVPdutUhAzx+E8dAnGaBjjp2T/xvr0Xy12eDYKs7zGL6ioZp6ZeCFEnIG
klOLhMwS3rVpcpCaluJa5zeLy+HVZx0E+H6OMdoL6vSiKAnErU8D1tL3tDCK1KhKE/UM1ktSUXKg
W34WPrujW8YCl++se3uRRbU1mMARIl7vZfWjylVy8ixabwVUpWnUPKl/nLl+g0zC4qz/gMAUN6NW
K1Up/LGAUe8FGcJjD1z6erMEcOAogC6MB2t+HBC6YCsOoYHxQH7nDSXlkZaGY6aD3xSNvHXZl3Lc
z4cZlTMTwQDH5ZYpB2aVxtuWA5HU4+33TzFkO2NPeiqlhuo0srJDom0EiNwvfsk2TUoGaLwZcwoS
evDlNCv7GY3r2PD5t3DGxkooa2mwQfGPQlc1RAvUu/jPJyS8oeO0Mnd/6Xytne0nhgXgtCgO9D25
dZ6qWeE1zM5+0/jo42erA4P3w6749RFGiPpqZJJPtwFVgD5VBjBizzMfGYrlSsrIvnuJPwyLPAHd
noZ0IJ4V+M31xpiVyT9ZaRaeahXz3fuZAvQudoPKOJF+f3rkUEv2oPKMxTia7qziPPjND+yYBeCF
gYYsEbhDgJXmVxEjvoiPAIaly/qpUU8xtInsucObn07pIglMdqTnGb2WZ56AI9XKgfg1YQ94JMmD
Qy4LBwtUj6en+v+jAecJBOn5zNReJjrUtUuSZt9+I95VFclekm4+J/vtwHRf3cHPCyfxwfVp6rOk
zZigskYeAKrroOnJWUG03wpkW9IBhBlHSwvHbSjOS5dCYNdN6Cp7iW/oyFanvPP1j1YNq7jGxRYl
xiw8xKQqnrzJdQxiPr/BU7cP2oPyv+k8s9KyzLN+qh9GOlczTuRUMuaoKCz8Mro0lZdoIl4lUoqC
3zrQXiEjoC9ngrxeS9WMsWyizALOb7MHOu26Tck+gx1naSqgeJRUw9YiIskOKEU31u/eO1CTirzd
kvjKxrdhWMThSrFQ3QQBJTwJjzQNu32AXLB6f1x/BDso5k88SJpW6CsFW65A1G3NepbiY24Vv7vz
RGtZnTLXnyJWm/PldDFAtxnpZ1u3uAn+e22JviXCGM98W+31ZgC7BdQJiFhqXZOXAMET2mOUbrr5
FWPAGw8A+kKjlZVtTmfROiWJGA0YQC4zRdE+IN5T44biL8UfWgM7aaTDwUHIls9jrgR3WxS3g7qz
lspSUv70t+xVODlDNUtFs8ru8XMt6PNLJhEdjOgZBgy48tF/FyExS0zPkFkFP/NTP/24GvHIW6yA
hHHHG6rHWm5UhCvh1tuW5tnBOVA9vZAlO1B4JlmyHJUjR0UdPL4B+HScC7LsmB7adTrlssQRUTcy
kIsMx5XB3lzN0dwwj6ECEqc/U3vJYK3FyqdwfNaHRyJjBzMZrYA3Z9MY5CQSZjrBGcESo+/gJuK1
YfeEi1/+8THpC5Ubvb4OXhOigSbNdTryXCbloxNy3l4vleaZlRI5ecHxkS95qTEMp7orG8sTIU1V
CJYBzWpc4YInTzzpFiVHOWmkxB6eWVzF/OWYDsV9ZvuY4lfFehVJBGlQrhSYkCTsz2/vKYj7YX2K
q9xZbLzGDBfnCNVwCK6Ri9U9uiHyJmYxJRjDhaRgSUhUzakDnvMPDJU5nhAOrVWbYpesjJCuhzqf
5yn3mrncCY/DwV+p2i8F/e4CIxFr08D/skmYDhAWpFxdoIpQf1oSbTiQJMWKc8bsirXv7CqNgIH+
bDsvouxfWxtdL0xxzgXAxLrbFxmaIgEwd/4jGworf6vLJ6hYIB1ztblSnl8coxkdVwe+qzjppzOq
lko1bZFlyDZHvmEYUs7Sdj6PNYm6/+T0wLELcVl51IXqGpHfz85BmUquGyv1HP5AZKQwru30mo9I
FUkGpj0pKvWhhriARsxHi69BAn4zxQdltIfdnI28ayBTM/DgNKPOkEon6v+om2ySq/xtExtMBy6P
W/DYAxlL733o5XIcJ5UsDS8ciMzX2sQWlpv3hTonb1UzrhbvCu5EBCIVtzEwJURYdpI2NNvcvatO
PrhL5ZRKfK6Ka/41cRZmU4lw8awRDii9Nf6d5kXTB3JUy42stuca1ta2WFAiudJpXbtMO/YJFqsC
nKd5O/qcGqY/BcLNLverWAsoI5kBrCoo4KU6qP49ChG453qpTiCQfGabEUiu3fDECqdkYynHD234
Ta3IDfES9FgVUxAAwKkhtf0lJzILn8fRdqUeB5IVOOq8M5ME6x3zFlqkws/CmVhlOzKrP5/k/btN
31A1MVSAz45Hd3hI4NvLwIJHUC2Y0d4AKfaFd5uQa8bi9oKh6+iEJ+9vdIpexdHRkA6Em0knc6Jq
7g65NJADDXtmKX8ZMcEB+AwdEI1GFINwiHlDJKQSsgIW0/4KTYTLW2vjSfkwwS47Q7KwFkSNAbx/
PNKqXIyof+6/UZK+QH2E2eqeZoC0NwzV86eOEu6EyuUVqPn0364NKmQrvslhedi0Rlb0hFcIAroC
WAXd6zaezj0AYe33GRovlAaN3157fa9hUfaTzJAvDzxOYYdXy3MKrsEsJgPLnG74FXMTSMwFEukY
5/xwqx+Bt2EKJDpC3tQ2m3zN30G6HAII1k9OvAx6DpKL4S6QPzXZRfxs/ZPcYxosX+wjORyVaZqs
Fu3kb3q1zAxjCufuoldcRBAfB8OW2HlURxntH+XEVy8bGPXhZGCMM8bnAnpEcguEYNnIyMH/NkVQ
QObeGh1MoIOyfVy7jDhNbCWwGuMDoe5Y1zfDLNOpBTzxa4TgAk2rL5jt3fD3Mwk5ERAxCuKZdsE3
Mhqx7dcDnikCiN3TyqUlQ/jWnCyYqWXXWj8Y8exmTq3RzfHPq/P0jsynJ7iRflALPAGB5vQLaWlb
AmY0KRzOnRBO9Man71MmxS2rheUtbOQUlDxIKhBX0U1gNBEV7YD/b6bVesJxDag0Q5+VqdXZq1Q8
Y1TUTc0P9en3M9wEwHOohHthqbZOQa2reuF/kNv83BWJhcCtPIUCfaKUEcoGfLVJn82HoxdWihnc
GmMEdLZPC1XkyGNrhcy5rEoabMcs7YT8V99z2Pz8jBs2EcHwBiA5+sJ5ShTevOUlATASOETWTWlP
hj+s14EJcwEiXT2wYn2wM8B+/X2d10eHsWTGBCVFSfmVyEDWVmvnupegQ4ERG7sdJRgNhGnuBBgW
GziIuBkESoHXST3pIGgb/fVMroruqwG4jfCIdHpIOwPlNi6v3E5GbKs3uuUQkU8hsMWU7tAwbY9i
nUXcikJG7jKywP7Dls0J8BkVYlqauWzXN+zMQXJTJXcjg1QczDmQQzWlrnWI/WxY9+FvssHjvZri
ZXmHTxHN/bbG7hiErNpn/WvMvBqRgBAilIZWgj/Sm69UpwVfUlQ2WCKXREU7mmDqt3IEMOgovzxj
r7FCnqU5Libg0SX5mhQU4I3cxj+O6coPS1bLt29nYCTILH8bfOSOEorH0VbC+JwyvYuA4UbSzyNM
3cksyMwkLHfFQIOnh680l99OUohhkyayYMNyci3cugm0FMSdiEgZQBQD0Pa3E+2k9VNCfwWk0Rus
suexsL1JizGruQVd0IWocXMtkc6p3Px76it7twNjVwP1S80buo6q8PaafaOR7FQtZWVKag/rkv7O
CXwakA2tgYxYLDVtlXujZalAVZcePA+sgxAZwu1J4pcvE6A97evr33gVbRcS39czrblJ3j5kbvUr
qTrINGC5bwZlpd57Ne4Z8PD0HrE4JKB+ZbENqlLn4fk9BPM3hj+xUmP8hUq218hbTBtGCaazmx5a
7Gz2bB2c9on2y4JAQEWTY1PCNJX7UyxTDDB8SGJewBFIe1tktgINuVX4a3/eFwOvn+Ir3zm6nFTc
GQxfUgx2tkSj/UERRbU1hWfVujGLQD3A57S0wr6bPGyX+Peth3Ww3cVI8q749OEBEPLVa2jlbBYa
Rb+JyxKxfMsF9wuLTuCo3g3NOxEhSBZ5AMTgtJdnVNpf0aOA2xQ03CPeEXy89GbVla3yYHgR3A3y
fkxzSD+zFBADFfT7u+/CaE6+Bu0vlkPLcJAUcxSIDCQOe/ty9np1NFh/2CCUJgsIy1Osg6viMEhz
7nwVBbVhpqYV81T2P9S8RbKkNEg2sitjbcTENDNqBPW1Px4X571y2kJrAryur/5bOYF+I5OOicU2
PAMBmpErJ3OPCZyraOwbp07jKmHPJWTiXXpeRferzF4Bz4MSgdBWpRhjRd/jEaxCHGgJztAZz1/h
z9h+UTGJvCPhOvSUqkLGzBHhbGYm7qxSYdC0AMMkGMNrsDN8EZAWJ639m1qUkAbugN2rV8TiAPyX
9viMSPOoY/LfyXF3QaG5HTKOuzB7OXdhjsMRZ+/6Fj683btwlkj04Dunz/+QAtnz0e2QgUSwOw/J
0OU8BBmdES9+iqUfUYmuVdc856FgcZdxrJRiGUYIjeDOyNnkRCKXUfaMbacw/mZ3vB4VC81ZwiyT
WWP4IJR1zryM7Ll1XKL+5oKl5jH3KMXJoQV5xtiSzoFUbu9GSHPRUQtax6nDEVbfFpv85mcrMypz
e/tbzpEzgY07boSLmrd+hJ3OW0qru5XOEM7jsnYM8uMHMI4qBEI2VcJ3AzJ0diKXQgog/Qb3e8aE
kWV8tHNG+tsqAxxadk2C9iJTOMno+oU/LzAUurdoAvzO2cU3rjeSyaQ6+ZPl5Wu1rCehy3itnIWK
RFlwW/irdowOqZEM0ZBK6Hv7Mz6oDM1cHKoUUZVgYjvfbQ0wd7oI0zSjz20lc0EPWb4Hqr4ju/WB
ojC1XZPUh+sthDUkP+z/t2QlhcDctB4K0RQEy66M24e9wYFvek3+dsqTuLSWm0jaLJGmbRX+FAZi
fyuXmapPsE6PbglH5jSE4MRJKdtTnaAAlxHgVMcYX7WONXzunVmid9y2Co9t4HNo3R4tY5P8Og5O
nuXyxbrCAsVAj0lZNamj7BiJwq9gOEeNOBPnOAO55z3t8kEuU4gYvfdSoJ3VCLB0IxG5LdyMTGNc
t7rhoWmKtY6llACGIqdqkalT9MIKX0PRIYuYPaFBYpcTgdxcUN0KaL+UEZuIJ1F6N5RLh+KBNUIH
bnYSHo6pX5tc524IYkcmQYYBy0qOJ2SxXmyrtBhj+GvdF/nX6KpiKbTy0wZr3YtgtgfYKrV2Yrqr
zoKbmjFg03LmusQHBJbud1yPq9Hr85tPCLVWebyMn6BGfEAOeISkjue8sRb9jvKtwZO/FWd+nMzr
FTcLrxYRConLRrbjkmquWtVA67psMx+Ox3hzMpcjVJWZqYQVw+Fwrcka7TtcXCoaS98u4JEx73GV
FRrnyoanUAXgYI418/zqDsr/AO0a5vljwwq1dkBTi6jBNhNRYcd5l371BpIC/OlkxM6JIbF5g3s7
dnVBAUoLQL/mqvPk60/2lxTD6y0ITKLTyB+LT5WUIiRcoGosCDY0l0WNNLGUx4racSulZzXzyi2Z
30RivOT+4iU48e4GBJkkiBRXYbadY5hQUhdxATiWDHnGcFeajfo1WQooN+WnE8mD3oDyhY1AT8mZ
Ssb7A8SveruHgAPjwJPGWAPC6n+Mm/lguJBJ4h3Ya+tNkhCaTHKCT30dSvTH9KUBDLbY8rVwSENl
PqV4Ly8Mq2zS37JQ3csCTCLA01NaZuQDGkf8b1vTap3dV6EvkbzeJ1ruBrPqUPXdi3rL26JSY+dv
deqK0WF13cY6f6qQK22DsIq8Jwx0XK8Y4NT9KbrfiVcR3waZyMXzkc7tUgJy+vz4QpAd0sSu4ulK
7hQ26CVoOY44W++t2fo75CHTXOVxub+lxIBn3nG7eEfXv3pqLh4Hz71QF/uCS1XKbDPVW8RstEo1
ZT6YpkXM3LDue1zA9hF9AGIQRh6e0GraOOK971SwfGehRmTrE2/EXwFfcYlQ79b6JWpnKhDmxqAd
D9fRMdjhUQJObLQHkcAscFPCcflAoWYVskV3YNUWFC64yiyJW33T9pibGQnSl81Mx9U5IuMssU0v
fkXsQOBSDgYkkXE3BItzv+m3SWAJC9yzsbBiEsYZvC/rllJHqp9pByEnUjkgI+dXWAVrUzIMfv69
T/Ep6GFToDptrueAt12azkrcjEmfs+9LlbmWIA1HVFh9DNmlivyRxN4DJBLgyA5l2Xw48lzBVcp3
18f96cYS5hlLMd6KXudj1SOi3w9zTMUAtww9T4/J92cE0MI0Fz2tS+K7IAiC/m9kX97Ta7NcwcZF
fySIYOEIkrAASXnwoF9l1I8AQdAEcbo7DvN5Ghgbb6Qcmuq65O8e6eg3rUdS9+XMfEtXBUVAOYv6
NQ/43h+j8rUalK+R9IvlT564e/li618Ih2RNMgC+85038YpjzcLueyo3IjsWO9UFMzLk0CAcnuDL
MsFjCOQABhd/4slZsipWjTX8fGCIpTxrwW0ESqRdPVtx7N3JhC1pVkSvcpwxr1itOUIjVHN9mNUU
rPT1z6kwIiDKk8EyHFsFAJZrBdz8QNZbB8iu8GRwq7nkLdu5IRpW1orrP89pGnICFOJhoUmRpgjh
D3GPuKjBknLs2fhsBmZLHboE4KJXdISY4GXuCftf6+pmSbiUfF+EOOpPP3zMIpCJhNlree27iF5Z
Znr8U20za/y42c6OoOhWH2zA8RoIzBjtCFOtEfsXcS3il2cGsMDS3tJxMXpfpkmCeeXygMs+neoQ
yBvt+ZHtxFZLL2/p1RRkcu0wIn/jnSS9612ku2pv2jbPXeSETKnPtZtXPDuA8DqeGVKEaaPndfjC
NEMoOXYmDaJt6qc0LXqv5EJpPS5poZ3fId6w2drJ7G6tDMNNHsghM88CITacERwesv0loiTnHOFn
jvMruNNBwh273wCbFLi+GjxgNbwIG+p2S2jn0qTq4vKm9EFJsYEbef+W35wDeBOPMwE58JHbc0/Z
w6AMLarqf1AqoAnql+DGYNeAlefdXpbgSp9sXWnN1EoCyE6LOfRmp9xLLztGvlmU80h6HC2HQE63
QqmOsA9cl3y8rUPRtUtzZzoa8x0fVLL4iP8b171tWbsX/R5QIlvljtVL/UjU8xee7MOQB18gYhkI
HRJnVHjezH0cb7eJAiXPwdpbf/p/DLTblKSzEvLjedwpMeZ/Bb6e1FN4H1bY1Ngire969BvWsuGo
oBG9uzjkt9voTpYrM7xqbsfV8OFgvsdgcFLyf0mRu80Hk+QZm+Aieu9NoNxpWhOOCEzK2g1qegD1
QPsCriKIxxsldxJpMSAn7XelFgKc12brdNhJp0w86gAuHsvgdArNfb6k8tsfIZmnEO7kYuwWXggN
dZAgo14C0uOxQEvy+6nbfoaHg2piY7RO3yas2oStG7+HtKiHeaM/W+RxBU7+3ib6kC56ukN2KyXg
it0buKT3WxkcnDw3DpFlGPn+Avhk6KTx2sttpyj+DWa6qKlLj4KbBT0hcA0lSyIkLM4jj2fFoM3s
Mo6BfjSxyluzBQNc1+VFWCTBPAEKYugJXdz9h0LxF36m2Q1k7tDps3296AM/EqAPl4u57PA2PNNH
upa9wrRZn+ZgTnnQt3n8e1ej6E33i4aY50IW/JHNzvhG+K0D0v6UAAvSQfiqFaVrro790sOPbCBW
ONVfY2mVi4qHrtO/g0xI3u8IRafpd9egBakABjLHO5mwyWXqDCsu87bI9I30go9YDnqFvL5wh70H
HS7GIT02yRmHGGveDgwV6zz0kRWDMYRMusqTKqmeB0xk6Kv6Aw2cncIEaN1leUTqrJvdQVJxZYta
LaRWBb144EIW++FhKpUYE6K6rhQaYhkWZtgQ6PARCERS3vwd3e0PFouKtS168tfvR4/abqmtO0tK
yWFBYFiIqfp241KVBNLqC2qsDwe+f1wZBWpwqFU56iDdmnW8T8u9sxpg0VdF8ZCH26DubaNTx50n
IEkG/cWAlTsPHnivwXg4BOMwpzeq1oFR8Urp29FrokQD8uSM6YvWwEHcX0Nwf0ofFOxYtQvnPu+T
8P8NLJpdWHU5b3UQm4aNzOzQYjHQ9jbEAQxpHq/LsaTPLgfV0y6WS6X9BBbY3oi4xgVR1gKqZ1g0
mD8W1dWXoIlLbydzByLNZfMCf57DwnhRNSU48adCq46MdPzNSe1wSEHRrYcBzfbtQjTbfJyKirwe
Ws3dwgnCW4hCatBIGyypPW8CJrqh1jpcCFanZjeRe7nKnj0vBvd7Oc2vCMOAEwY7iWbc3oWSXdwG
pG5zduMzuVjjys1c6ELMMyj0/q5EwDaclqU4zYxcpJDriT8UCJbtD8Ij83SoslTRXqtpSMMwC+XH
YgeDquXtlhqaUwRTkGaOSktCjSQ5Jy8sa7vEkI61ue0zRss96orGDud3occ5/i0j9zlbluVsq89p
zPTRCNwMzmjeeg4WLHAD/Un4IPGbYujJwhva09TEVpMpRx5lLIKP4Pl8rf5m4LmTnTOSVvepYqW2
tS+TushPQW4z6SR+HuzxvHfabBJ3CJWQXCsQzDEcd5ZzVxdVUK646P9eIbm91UV+8ETmzJZkCQmL
BAVM+QDZh+v8aNR/nPbs72gZzhSgJ/gNQJ3O/Y4HVkFjcs+lDkjWG6j2EveegKqBWa73evQYUG85
EZD8EGWOVx+fVZHvUuyoLiLlgF6UTiwm/qgF0H1+sQZufqhfsaB1lUn0YgwDjbNBCEypxXs2f1xj
KpQC+Rab1wZIL9VGSLc5X/Ybic0yDV4TwvoqfFwsAp/6TyipiWofyMRliRlpYjhqyiWNit5iJLA7
eQ6XGKT2gK8W4r+0HbiESPYvZTHBJrqjHVWTG2I/mCPMq/dLKbv+xqP9uvpwLdJKUhvjSXd7m+mB
fBX25L+PfPXehvhBZa9R9tTfojWWz7KwI1+qg5zOtJThY2Ah4AnLtVDqt6JMf9Gm6JaiyoEYFjTF
+XXeZaPFoKp+hCQADUNZHWE/Ytd1bo3uyXfmI+8asErfZ2ksmEdg0OC/TGSp2WGzE/hMV+D/PZ7B
bJNzCWCbnagelyr3zBXQ0xIUy/Ufq5qlKdStA/YXRkQYNZO/5oQLgNYaGLIGusXS/s9U5B+R+21f
WFTxGt7gnLU11U7IbY1wn3IFtg9VGFMxMzic0dvDgW+71nAytxT63SqnTEGmAb7LsrudpETEPwmE
m9m7LUdwtWBt+KLCVj/n5I+kiczgsoxFVSVnzyJA1dm+/mTV4+CrkaBPoP1QyPYf52SF23Aj4rs9
wi1flh/Hkf0eS8kGgl6vaxBLCioGvRMZnN9uye/U/69apVSbZ4HGDb9HjChOZ5D67wLuGYR37dLd
uWvgyUkQV0Z7fPeIb8c+DyydUuMMoCc5/Hz/FdHqfxDhRNY/eV5vWQBE+LUDUQ/DlKeNeJLLwIYQ
QxCPBqZ6HqIWzwd/vCN3pdQB+Utmxl/L9YfybCfh4L+2TfQkHUkgpKOu7F0Dj5kHjeYcxxspS/Bt
VVf6Eo/MrSn6qZlff8Ja5okb31Z+Uk6Q6cnimP0XpHMokGcLzjke0vEeT7cM6aKp6q0oyJbpBqH2
RCyW/YVIlQaAJD4fHHkB4qMdfkjX69k3+f6MgiN6mPnDcJQNuq7KN0/wv3O/x2ZW4xodXhzJfVRN
q3cXUR/r8wguzMn7XVqUudjZl/1L8WbcQN1qCrnjVK7FVs1boVsCLtyxz3cDZijr1cdZaP243UKz
d3PQ6rTL3bL6VyWKKPN6LC3LBYYgLI3nnly2ALf3tLtv81G5tAiGErpjJLaG2XY7ndxL+lwEpvDy
+dDUzgbwUd3estLi1pFaNKdaAwCz6My7j8z517V3L2Cx0TNksEZJIKh3pNObdKEPUsM/Xg7BeFGJ
vLMfJOuJRo5UX5J1u+J4Q/qK1D4VabyJDkC7qU9VNTM85NSY7YByl9nFn0P63vG6g/W1cuBGyv1l
lmcPYOvxMulh5WZMidcoFnvexkgkpwEj5eI7Q+kp3xZaKj6ksjjyYpFWeW0tF0RF/A/u9sRSB0JF
IyXnA3r+jGF+wDcyyCOu8EKb29QA4mfiWHBg2sLEB/xNVz49VXS6vPp8V1ZFTMKi0A2wvxVErfTs
C6F0RgReiJFoen6J/MHjOCEAo7MB0SWcFuddhkC9A0NUQBSjdB1g7+xbeQEe4d4ryroGZxqfpibD
0UKoJpx9KxDoLO9NukplYW2ToGzAU5ypKVvyC1S/BsmLFiVlLbw0wyWXFncu+891JZlt8xY0Y8K0
gLhpU5L4tbXbXoihs73Ozt8ePGFxTfJBm9V78AVOkOWwvfRsF1+KMFJPMek8xIRt7YcaC2jhkQKw
XYpHLC/H+TKaIVYmzn+FUFmhjCk50eWm1yTAf5nx1DzEoZhIL4ECX0omfT3Y3B7x3P+XWijPN1UG
OB13RCTFT1y7/ferKPV5xUi56ULz3N1wPjgIXuPRD8oMpw499Z9ikhONfq2U23vOjt7rm3vXGc+W
3v95qn4/QX+r6bjC8ub8uvV1YuImCaUZOYNkqlw7PkBZOKfgHWVEXhdaHP/boyNi1XZDNUHc17sk
Bt3fb36QZ6N60cYdB9z+dGYetZbCwmqL53KDpGz81zHBiW86AuxwUlEmkPrYaGVFNVjaPlKvF8ti
P/iWRLf4Tk5P4zVJ9a1tCakmh7OD1/bQj0TGalBigY8tu0g0G/p9MXH5Cbj5qWIhbhGArvwxFeUn
9nvM3NnSZz5BY5iWF+nqMbOd5sk34k1jkUO7zMbymZ8SjjwEPs+DHUSWZY83i4zsyAdf3hd4YMrP
CHb5idA72HqfMAnNSEATh9jVx2r7oiBImVBSaavz/uyc16hkU+tSm/t9pWa5Wyf6dZIkO1vZ+xBz
JtK8idPeevl4NAPFLmdZM9BPXtDJaA6TY0At4AySZyYhW1TK3Ox8BDsWJ4NaYClgpAr8xTiv+FK1
bntUO8vTenN/WXMjnu5jyriq5zkBeripkK6ZRnP/vjvApJDbmguAvlWkNTFQR4USOHzSOYgWNq2J
zA568oiywGxE5NMl88Kba4kfuipyf3NyuuvBQ3/WTV8IkzaoLZrzvjLupuCqYZFd0R4WiQ8rxDYI
14YaSD/cSG1R4Ok19qEwmvdkqsuYkst4EFC54pdoyiwfN3d4wtg5LGbEnr7prVcA0E/J/U92qyMl
oNWtEv3Gyn5ojnH+ROdlIndaA2AG0L3tOoWCHv/NwqedotxFLolkJw3C5mnSrdwYw641wZAGjKIM
iLfOZbqOLdwp++O61x8YaF0pMOIvTF5oIBz9Qi6xUcNOmgWTzQH8NoVTPbSTiBUYr9M/NUvNGyx4
TjZtbRztvO1W6NQXSlL1IDpg5cbeOpctkrQ/wq0UpVrKHfVqrTZXbXdTbuz8VyECUzgRvWdkA/yO
pUwICr9lglIgAul/ApqLCaPUB56nPJH/hBlmPY3LrlrXEVFWzqYUdTLBPsvCHUp69GIgD1/X7gh/
ih6Rgbme3vNbYZ4uWNygeNXtnWOOXgNFXZGlZE/S3WmofOf9uCUspW+f1ZU33eP0mzSswjcsZav+
aO4v8Q3M7mhgVnlPSPcQT4vmV8eIqOIfuLezSdDHfeyTrSzogKMnrlgSKaa6+f3FwLVtdI5DnhPE
dMlwTJ//RcWJYB58r4zuU4Oc9AOjcm6lzY0Rl2rKSwtEENtOBWsrNtRadmJrrc7Tbj507OTfkZlj
1FUTHPJWVANg7T3LawhgKepG6lWOqRJbf6a66lnK/OioYVJWUAg+JrDtDM2W/kDIdl03Z0E2Jk/2
g8T1W7FcYcEHLjKOV/x+MoF5UDn44/8iLsbDDeJYUWvMu3lFYTLjz/s1CdB4FN8pp2Q9MBv322VA
IUdkWMEw+fgd6s1z/prjyAKhOEeENa6q2DIYMcv7xFQbxJndaooXjpQeuB+vGLZzgJ91tKnoAVl0
XnsGYlUsU92D9BBOGI0mNX5we9P8BSctbDoZEtwuP45DfHnfWCiJ3xZqnXVDm0bad3hZGW+tgRFg
fB5ZjoCnwGZD+7QAoYRDWzIXQJ3IRJhsZgLt5NHTNNK4GG5T2oQHmztryWDVLdZLTKrAEZ7e20rU
/VJDcE6CQ1teEM7avDobGCVOiZ4H2GVMETXHciT3GiZBMaQ5rddPvwvDcm3XiIRXT+n9cxw21iBr
4xkuukVLsxmE35VaDSchpvUy0AwFZT+ZfaAGjTnNVXkuWIohqPXC+H/tLRZ9PW54dpMqbI3T/GVp
IjkvwsgLiIzmUUmqlm1FhvkYwaJ4aA1AOO/vsjxWcpsw4zRJ5fOZ/wg1NVbG7/TIQuUt8J9BP/F7
KRmwvTvrYrHaaw8w85LVBtdYG/kSKtZ47WpT4VU5GkMxdsSeoqAk9THZKrzD1Es34qpw1D8SibWg
J0wOxCFWvPFSh2aZkAX645fTR2roar/MNPJuCjlwSnjxHUirs70zRgpgewhPYGol8KWqceE4XqZ1
Ua0CHqWNBNyYCGmKUdGqKVmI0iTnLzt1JTOOJX20xNQ0f7Oqf7Utq6DPp/7Sfp2Uc4RpsmrznP4L
SOxu6gMFEbqrnXnOAQkjDUchZ01OSjkC2AoVspNTkXBOZITW966clhmFiWoIvaGhwefr8UN2ByeH
BzNneNXhGRxKgmZdy28qaJUEhyu4XBW+ISMx0IjVS/nm3gFhC41bqkGKc1xjjLJNKMwKtnBQW+17
jHZ4za4XdhxzAJ2DHTbPsqJAIe0xqdMQ47yZ0EcQ3S3OeRt8C2wr0zKhbIaY5P7S3udm/OjP1WQQ
LcdNdhQaZlkpvQXGXEUGCQ67FzxLpzSDRQK1xAmOGnxetSolZhm6BJ4cdflt9JdGlqnbx1mqjL/D
kX1oiqW0aoKFjrxGqf4noSG4/PfL/WoQRZe6zZ7baRw+jenBbljNHdBmfadsx0jcp/fR1W74f+pD
zf1V94NEQ5CQRiVqEHmF8Y+7qpBvc0F/sfA/HgLP3/zAh2aawJsJhWUjEpZxOJBimV529zAN1V7m
6IS/7idcihOzIXMrxCKEq9Jm9YCH11vQc2AnTOGzTeNAlE8GLh1JpkXeklApilHQz+coLpJJYvXE
JZllWOhuBFZGHiwVOY38PdCSCG4Y/xlWG917A9hrHo7HPWoWPM34fEafKjJoUfrd26OkFsJVW0KM
ZQ9EvRXC+f7n6KJkbKfDNc4mG4oFD43MReU272dtPpq5UJCcDzXQxoO1yOCVwwlp7nDS1pK2+zOX
DeoCNPK+tJAk+M7uFpyX6iNZjBwS5I4ItcCvS23SFjlmgEH154ckeozF46FDnc+/awik9oaBKjEY
b+8SbLn3gGYuZ93NXDATboi3ZXnrPx/EYFdYF9xnJFdlIHfovpvFXy9S+pLxBwwJPucjvPoyFW1q
JAqJZEZlTs1h3q+wNiOS7m+7u8FY4LaNn54L0PFw4bLxp+BN9t5wugOnag/eAVtpE3axA08QorDD
wwjUokCOwGu8lW0HPvZIfkl/QeD6e+2rM30wcmiZr3kjyrm7V4NR2Nzbkwsg3VmwXL8fNH7Udqg3
end29XSoxT3Rfnyidfb01cxQ66Gh1Hq1KZdqLIrABPcc5Wd3EYYOqWmmgqof+XHb/m4gNkASvyVY
/QqH5kS6MZ2dRb+u/nWdOarAzPkA7nGfWsXtpdaXAQVsGVd4KHzGKE45AuwTEDAeWQ4309Yem9RG
YKFpA65S5HK7kDCjpOLolJg77PuARB5mMrzrQCEU0t8khr+wbooAEzshlsTy+/4M8MggZsTwA0UH
zRfCEC+JRvezeUhE3BwXhAjGQzTzxDdxXb1ceh5sIhF5LjwBBWNUbkKnzcSBlYilUSM61bxFg/zj
RO5hCsHSdaQwdMhaL9GB9ZfrUhEPSXN3gstxEozuptH5Eqr8AqNeyTcfgX/GgzctQ2KwP+rJkY3T
AU9dibdAStoSzGK59MUvB0LrRDTNV/F6vFwed81vpu8+KvNwDGjzuSqIjdyikotQHcEvtEE8McQc
US8M7fxgP9DbGopZ+3vOgtcCV1XJpSLwjcuv7JCwLmiAdhL1Y4G2K6qp+8UAXGFb4AOXQHvFm1GZ
9RYU1VbiKyrVNKzuHURh9q0YoWTn4VP7cngKw2T8e7K0H3Q5irWQ1CmYY8Ex8NGFkBION5pn7nSl
cVgKkkclSZGlzoJuEgWRpc2I/JA7Q7zBUK5yYMUGWJOwaL/cN02STJ2JFIQh0pBQvIUZNVflEsVT
9VVy+VsoZNXXT8hPnVm5uH9znO6hezlUCu2oKGQBfyoos3DhjcDr5ibYq9jmE0bvLLq0UurwxJP0
h9Z5G+EJ8gV7g/0W5+VbWl4z6rfXC+ESyCRq1xwU7m419LdMp4UlG7yhbfd/G8vYSNeXsJJdLYge
9j29pvEJzkvs5TWGwYEKF+4tl6CCLfBw+w6q0XzJLGwGToAhlz/2G6Em81HrLLx+foYKiPbW5U90
8ACBl8l6hSKN5sXWBQkoQTqMXJLrlm6Ypp5oJoymHhD/g6Ncq0nYcG3uSX7kHu2JRtsHLO5m6Zvd
BLyRznoA06usx+Bg5cC9F0iYeuHrSJqf8pC+4JvH/qbifAbyMoifwkFgCaaO1fXmsnptFEPkkQx2
IQlzYgI6OcZxIz/mPu5xPE2EoP50r1d1pVQtQGDhLdqCleYix18/t/sC1XhV9vVgKCE1zFQLGex/
fDRLxXfGmG9Fm6Rs4uIjUBzmoMp6jMFG+1RiozyCB14WjkVRdpfrPjM60Mp+oX3MCcNw6bNdwFjB
kSNk1v7oQv2bW0zVew4wpjSFiySfkz/gSRw1/ncqfrjGpPnO9jMnmX5FRafPafIMaPqhVKzQLpbX
9t+GxZW2FzrPRwqqNtHACMdlYK0FZC3PUvc0d6bxlqnHcXwSYiajwU0Fc6TzEEOdFqJdBITj+WmS
B746D9QtesRZifl60+GEhNs2WbAMpQerl6/FiUoVJfUeF/hv33hBLdr0poPSGo3GNaQqJVM0Htj/
skJiFPVWCm39jO+EudTHo5+sLajDZziRo0IVsDIL0K6aTDIq1ak8vmcJrqMO04HYoXDWC8XSAkQr
USQ06Y5U66ytAiQJ5Han0dU7fp/UXaeDBLIDuPDuHTuqzHgqJfzFADvNKrKmFQnRMr5KbLdfRr2e
s8K84m90dAYpLfoKsDvM0DZ8X2tZsVs5EH7UXG/5Mmt3vwatEX3JG6jzoTH4XDZ9k3A+dKOc4GCO
mkN3ahXqL2RjgTcwSJhk5y80fbEUWGUApsMnUc9rAlYrp1jFCGIl58TvOA7Zq8zsMRCE/scdOd++
whinG7XJzEGnto6OcWa337nxDQ80wXOO006fK9l2ho3oDPFpkCw3T8P7+hLIlsRlKNieP/chFEcd
krKvWWN0oOgSnOVyGpJfEZPhr4qyLaQh8Vr08TuF5AqdLx9l/7LIzqtymgMPFjUht52kIzoYOgYo
MbDN5i4AVO5dQaZ+BKcdROHtD5W4ykw3VivVN3e8gZQcSJVyLv5Mm55bPGUK1W2cNOUy4CSmvLKo
L9bCbj96+l1CzkJyjrD14wjfQe8SdNo9S/CLkuEOsDrxM7MwsP4HLuTkm08ovwYlmndCXJv9yce/
T04otM1QClod4g7YD8g/jvYIaLhC0muNakOCGkkXDSR2HtyHvFLTqSBwxcavZI1Ve7o8LP5K8NOn
m6oYZGKtDvOyB31jCBsNDcPjYwVCweRXg/JfsOIRPamLhLqOzCr1oNYp2XYL/cT/61HuW5d8+iLu
dcRrY0roVSEs2VT5xr4vI7ux45PE4fjd85xcLJYfAeZrRIlO4X8TpndbGLU0C9YKxf98Oq1B/nBD
LmT53AxXCibKS1OBMQcEaiS4gEUUla0bQqjk8yqD7QFvmcekNk+l+NUpedAjnbkah1w3dYH6PjUN
oanK0aemE2XHKk5zLjgKc36sKF3I533LuIpyxxsJ0rv/f+cIUVAf1yLmcwmgfbAQKy6ikj3nRMeM
XL670a1RF0gkUoOw58zHLvwdr3oaFtWS982x/rdwjoadtTNWRR9eRNawD/uIXD72pEpxAqqq471O
IKaAP7l0NkeuUfS27HW7tbra2P0YBst9lAT90uaG45OaFI58I0q7jtRtthITfRawctbbYnpJ/iYf
lejKXLTNgdoiKLf4NFBSuvs4PMLeUKr1tEgxhAcsZqRjYlPBkpZ7jzHPPaylrnAV6ZQkh3J4DukT
P2rA0TT93L3m9rp+22Q7wD7sr26NhAPQu0QSkZwWnwEOOizUQvEM0v3Z38km7+RGgatPrYvMrwGv
yMtLN9syR02F+AfAdH37HniaTpuaHilgceT8VMAZkT6NNwWntL58EfCWUKuaNJFG2+r5gCTeZwKo
0sr8sp+UGqGL3Du6032JEIVlk1mWA/NHz3YXAyZaimDRMIa5wTtH8+hFR9ndmrXzOsy0seImprl2
Nr4dYfSCNilV3B7aIY2/6kT2RYdbIBOjbBjDyI6LXM/e0qYo/H9H1zzelXheh2fhWc6RGVrr33S+
kEODGoOFen5+LVC6sW+zf2yrUKvxyTd3Ef/LIsUaYsu1Vy2xnpGBYOvKLIoyDI4uNRP8Nmg/GBFj
pmpMPwv/6/N52LtG5rV0OSeYX+Ghkqx7PK3yp8HenNAOiPaquTU57Tt+1FjDC9YGWzgEiDFlWNsl
5TuwYbSqu7PKP73K4S12wXu0hFHpNdM5r19jsVAMdlpoJbOM/4Q0f9Io4htI1q2Lz1OiMqXRV7S4
aRECT04d0cqDiX38casrirCraMb8ODmunn7MH6FIWC++prVts9JHrzJ8Wt0xv+Nvv/bITHMjXJnH
fjF6LnV1GxLocpQ8OIQUNHXd63COSsVL8/gIl6CoCMwcB/MbK4gbwAH1C2oiLdf/gOfUmEmj7Rsj
TVkHkcsZ82wJ77faSIo3V0rMjNPMCswEXiCaZnQft3aYU9kE2VkCsN3dEdCq7ugAOl1gKQ4NFJyP
K5M/kkFur8B/iN5mEfaIcbDzdEfaF3jTUUFV7V2OC216AOxusdOTv9F64RHTtIk+oD+wRvC6jN31
vniB/cBHvctPrZEHxdXzQUFhqaxnBT0/NWclhXmWL82UHZITK2g0vIaGKoqF+0SfOBGrd0IgE/us
kXUW+59guuMWz0LnZun/Z4m1rrjQj6c9WxAIHN+bqZxwaWl8EmoT/kkATK40/9SVW6C0+OB65PRk
lo0UWa3Lnoa8eeY4rVPO7BNnGT1wHN6O0QLesArMmnW6PzPKAWkysOhrilp/MrM0Ta3iX6EqqUTf
iulJ86g+pkR/T7PGyXR98O8CkGHlGFHrvAms0Y9sIf+YtJ/1sBJ/Cn4QM+LFzDnZc3Z1dcQQOtNj
6KNsTO1LXTsUylAGilAdqbHePH1m919JbCWTsH3V72eOrWejY71t1k+INFhWYI+h/uutjZ2/opCs
EOEoGfxoWBXAv02lEeiqQ13ImwNGxVMDiApCtv5FMBpKGYPn7fKwngaJx0IslSAoJRiFI1d+0scU
3YRalNNKAa89tWdzXVc9xV8FFposCCie5LlZMLtpPaVbuZ/ybkqnM+7mMbPMAZSUex3iP44NdB64
0tQpJeS3RW3DWg9l836abvqvUPTWyLF2RN0levYkRHW1o8aP+I541xQqDEGa9+zxlIS36OuzMuDZ
y5NhKdOIObTHBmT6slrTdYI15LD98vE7ASYbBtYm7VAP8fXkXNVUrW9j6VtIyOiCQkdnAUIW4YT7
zYgIE5cmHW4ZY5sjCCUJ8cHJDRcwaBvDLbzbWqo5kk9Z3lLpae0fxCSBQaggeUTyrN6mg9xJKrHt
hJgebQzP7NXDF8ygg/fBL6Be2yRYZD8qr+xwFCGvAEMMMgGGzy26XJ0I/x4aFRHXQGAZNWC+gH2B
0qOKsWc0HDRSNg2cfzpgkAa1VRfAa8GJKy656A9twIX6dHCi/EAHpCz5Zuc/ckStee+VPS3MkbJz
Ima51Sab3E3MOut0yz86iTyHbWxJuYJO0YifqRC7LW109Qmye9/SX8L5eusX2Ol/A3YPX1CBZ/RT
h8PkDLXVLbX0fg8UILvLbnZySDyrfg52Gn19Bz9Afbj42Sstx6Tk/KcwzY4/n/BM2O7fEBUMT2mn
/ah/g3FXBqVf6ZWv0EeJ160Bm56MXty/liSxhBhSGn/uEyc0fcBbkhAsb9tPaJQDSwFZhVSQ2l07
BGKUTvm04ukKcjeWXKqwMH3qw4rguob4422eAkYK8pxAk1xmUohLvY/Xn6oLpzFIOZsaF3gM+F4M
Aq+x6nVecBlleCT824h6F+khPvRDwlEs46LEV5Ebd0irC/Yj1FAG5H4r3l8tLcr2dmrgw3uue61w
u8yOoZfDmqCMglkLdZ0NL/oeCjGNvaOF3xVNV0IYgAlOepjgqpHZWWBAQj3u8AUOWNfmyzj8p7yH
ar5f9aCDNCRq3IH8hpmrtjEmZIKF8EmU6gHbkLtCWI4dBukM/MnAnLbO4LZCgNsy3OsXv8tk9PQI
BbdK3kV3totnVe3/SWfsn6XpCitUnmEb0Ot305CSBwsCrmDsDSjbriM1CCFfqvmGyohYS15EZZRK
QmqBxg+8fYi5b7swEA1a4u2mNLrGX1kBvwOMnLKO4GIzTy6XVJF2l2esCmJOHZtkeGWiC6k+n0P7
PazmR8F+Pc55HQOFbI/n3bzIBwQttGZ1nRtErmUOOskIGTjdaK226S7+1dISGIChJ/4+NqSWQcJD
y7vhXGZ8X4m7+rdlDVUOrAynHn4Z+PD5PGaXW7+t07ckZIqTbjSbEzs6Ss+u2pfw7vLwz8dDy61C
h7tGhwhC8+hvgy7uv/hxqx4YhI/NnVjkmZUNHHtUr8zbWkHC76YCsHQDbOy3YJnxEb7I4JrUnbQY
gAtP7JC4bC0wRNM69f1wXy0VS0xosl6C9xJoEOqC2QpSsEcmSs527EjPTJE9dYy+mhFhWWZ2QgCJ
+6MQRx8rJBvJIT3M9/7PAmnf0OALMxGT9PBaHlS7hM2X2V/aPmq0tWqsfcYYbXuAskux0nkG0SYC
B4qCL+IYBvsOUbnth4wgpIzRsBnMU3yUTytI/QTEqpzDYI3ked0icEINWlkZV9PyB6VBiXywhZAW
KHAMHfgtNqlka1UKnDJpahyVBSfvW9bwJMcPJ2WkM4E66u2U5BKBBvpe7j1FnLQAawCiGZargCMf
4+xMaOp3uLm35Z+Ko4+TkTGYY2HVAHvRBKTQESQRwZDubp0JcceP7ROiKyiKb0quW9+uwIChbjsb
NdjxcfSsGDGxJnClDy1QfEAA2+wdV3FpBvjMYi71KRVCAOUg2IWaI6GGpwuCRC8eW8lnHLK0eFvl
26MUzEtseQWoA6SYA67PZ/xVejI8+fRq+L3KFkIDYsc8IT+BaNTFntihH1I2yt7m+GWulYEdnw1C
n+yntc/7p6DTlQjloD/BYMlTBMlmKVvgm1VubPu5tUuWDZfRGmgtd0nimYRkXIBJkVt+fqMCrcl/
g4t9YQANGQKOrSXNLTIsq6OyFVuR1/WE8ESfCYT5v1Jy/zoIgg+OzIUSy0QPajHBkk9QQ2Hdaox5
mir2fEvHx+lklMYNYIeBAsw//G7yyl/8hy8WIq8/FeTJWa6llHVSnD8DAW6xER1U1y3mN8VDsdQm
3fpYctrXLjTpx9CeA6Z4W/3rWinsB/micGJ3JZ8s8zPbzTUv5Hj9Lbp7/9cJiHKk0k6wuS9untf6
k7HDFbwW0EQYhGfiywMAz2m7D2XVtmPHFHJiAkcyQhUdhMa6ZDIPDwGfxXROZhSRPOEWlDsTWWOB
6u0bjptjSoMEQTqsqImh7MFJNq4St2HY3uYtZz4UYDsxKfXwYy23Gp5GLWGsBCTAmmXRxAk+AegT
p5c8TFgB6QbjXZNJ2mQ3sWS3CaVu50cxvL/abZ6b2WpiNW96+lU37jS5xytAjg6BGJGAzMsMw/0u
aSo3uJeU+fx5T9xWaFygi4k7ng24uwsXmxWLrO5RLNrSOdlUPhpQi3xwaR+zPyeAqYMTovfOOiB5
5U2y8c/OB5UmGl1Bu12G1+9T02wxVTBp1wEl5ZsZ7OY9C8BLfX7cudOZVJ8n0HXACGXx0z5UORTM
0JE3moso2jUmJxyZaxDdlk4f/U/edoB1JKq5cc4UgcDMpo4vJ5wmR9HotkH+VZGXwJaW6tCirwmJ
OnKFC5kY6mFW7CI4kkthP4V1GvYfRXqa/Jl7YKSxH6f8UZQWzEaDenvocODAwqtQ+Awbvc1rvQ9P
5mTlGL1HzuDuDy11MIM/Al67vh3J6Fw+uIpB0sP7bJjW25kxWIvAjPFnFaA58aAOYDkr30kEuZs0
q/CyW1mZrD8abNZnsQaIPTgih290TO7T+5PQc7giUv31DP6IFHSI+xCGpFQnS7vktnifRRTvFFyL
TNWaoo4SCiaLtMXtkysFKn1JuxK/3H4ngixALhdACepjssKlREcuhiP1nNF479EvRTGEYRcI5R9J
gaWirMtJR9K9MS8RJWviImrj9NoJANw789Bnp/wXqwqC+ld/UQPqQXJu/rkXSrjnSUrL8KEo0LHm
fVjFfMDc3FYHT6nmKDumsfSxss4KhnB/e1LexFyZ0bFIMFWwuPKzQ6CVN6L6b4XwAxnuFbUNlN3q
qk4D2HnmDAJQzv5Bvbj3wAZYX+GtB43CFrlmNmRHP71N2RPR9ucEy5/kdQLxuxJuw9XLEnR3J8oq
cZurBN2TS/m/zh/DU1kLTFAx3o3EQBkQoEmkBBUy+YEx6OFbf1ZeO6JehLlczBKNUaPgYstWt2OD
mib14LkD1tUe7vRdP/6nOHMP/tXUpwV8YAeyzwToIRCKvB94owRRLMFP0z/cWIOJPtcZ+IBhzor/
GPxx+IxZaluONSuZmbv9Ot4EVS5CxXqveLIQrxRryefRvxPE9eepO5oLgp2rTkwpSdFhR0g6r7Bv
9JfamWome/F/aeWJGBcCupeDFmu+ogp4+5I+fh9XutVhmM2NBFcOl/DSGi4+kXw/TatoRtnT3T9L
1W8G3Nlt0XfSKklZjRb+BQ/CvD24kDPguor1gKU/dlw67htDZjDM2ZcQvEvWJaq5vk0BqdheKzUc
rkG3cU97q3WcjqEXbos081P/dz0uJkREabt0DZ6/a31xPX4+B1PSo29lFDE8k8oE91V3B7/APHwz
lShWSE0lyKGzFZcQmBcA78mV5So3tdO2xClS1rtrZ4KBA3QpvBmVf73sf62zuR7YdgIpLklYOZOQ
yiIrCPuk3pclGlFXMorjDM5uvu5PO9ruU5rEQa/nbFFAlT1OS2AQrqDDeQr7P0GQdhZaGEiH8hox
Ibyu0vNZfYSdStkP+YOQi1u0UZM9/lbBOfKtPNNER8uV9EskQDqdCjKO6UNHPBA3jaHl8MEpc74Q
fHzExSArrJsJ+E9dpUb3xU4U40tjxa+2F63JRMnWniqwECsAshYvPoxqB7KtWNFzLXWey9ktwROx
KQQqTwnD538a5JVb+n05g1MxmludeRduaImuR3CBl/d26QQ47SflnP5jkt2HPEMneMJ9ONAMk+iT
O/Q4n/zkjpBKTdkoqv3t/LET+OoziPlgxPLL1pgDa5wOCBWViz9pzRaMyc9RAd82hN9hpKE+LU23
bh3jU5f8qt33N6nUwm9C3GKUGBXbqoegPCHEgry/ZQyQrLcEcZL52ltL1Y+Jht5pElFE1Bq59N0l
Ld/BAR7mlhFlACa0Qb0Az4EZBHiFLGC/RBPkVbXcOZWqtl4RfBpZZswf3Jt2wRTN6iFQ7+hnQ2VA
Vieh/hjFBh3g6LlwdWPmwgbMh+l9JOmUIMf9ma3ep99S8PGOA23f4Nj2J9hMolf53DWgaOOkz7wT
PVnAuXp2HhGojTnpLdvod9Kezvex8Pl9mRnpikTN+3cXirTYwzQ4tbxCTfoXtsuXBJEJQSFpMl66
8yTiM7z+jylwLOniov9bEF1oBRNHzt1Ep/5zDQ1hooCi1LCCbTzbC/HK077YhZ2nOsop24xzB7HL
sLvcCC1zPEErhQ5OP3ujN5BDOlS4zBmpjK6ypQnlz0Ql8Axrt6jZks8LPswumaRwWylz1BQ4Rpcs
zYpD8S8DJY/53YVhmlDUow+tboF451f/NH4UQ2ZqaIJ2j0j2c//CeQowVx/nPy5Ir/p5iAbW3ID6
xJZjxYyhK3+pwhn9gdBT1wokfNyQUTFCfF8kW9+7I4HFzMid7qRh1yfdaiOet5In/qhnfi0CSqJm
JIh1vdV3MWZu3EZoAPfSIqBtAmTP6Fuglhzub1sbDFG1e0T+dPw3S/M4lyBpDxki8VTuI8mhYMAN
rzoRZfVTmDTvQmsCM92Sr4i4KJDhMc6yNqC+KplDa+7OQDfGHdGeW6eQ+34tqzwCsqaV5Lztn5qb
IZEkN+amedgEtZF+0sFKuURf5DUi8O5fDwI8KElHHYZjMlI2kEBvpWEMrv96/nAzU0Rh/cXuHzQs
q26uMd88RcfyJZQWgsC4pUF+COou2I/qFhEZElAN2iNOT4zvquh5nj5xfEaIEX8ESTn0t87MIObq
Xn7ZxIM4OlSt67hg6kWi/DRdd2ZgvimOUUHwwQ6W6hNXFoT1G1lJU93oT27acezlB1WePcpvBepC
ETArAEk0iINkkgC0TjdHRoWv2N8BfQc7dZXwbv/wGLzgDyuy7KPTvvyjKLaWVKGkpojg5N4ZLzI4
5xSQY3+JwtDhle/ytoYPXfjcVBfRtcG/ywddyYyUx/+SvTC88w4VVEVIBsBAxoY0fxuOFEIVh1O2
44+uKJ3BHA8VdZ3fOimv2XxwSM/Z504ZK6Tp6aJUx/NzSrfGWx+qRv1Ffxc27i8Z0Et8C953hJfE
gPltuGjNVgvDn+k1WlxF53R8WRXrA00j9iHHVhE9iHL66lV8ajsNtNnhTt+9nGlSS1Dqg/y/umUP
VZ+zmg2wlnV1xWh5xbbpE20A3WL5+B9kzACl62wNMSUQhtet5aMoOxA5vdpMUNrE6ooNGR5AmYSA
khim3MMy6ChGrIYQqkfpNVYrrQ0N2UoTrjWgcl55BiAUSfaKJpG8CXGntWPc5h9lGc2+zSM0agt2
q5uBLu6idJg5Zps4UJWIL7LSF3mwKfMNq5LJyVyDOydrPeZPPFxGN+cS6Nd06Wl7OEaGizr49mNh
z+2SO50IGiV2KXsEW5QSvgYEUrCSjwj0/MCZwcXyl3UWWkBL0UFd7XRaxejHiN9l4kQtWuSOyCEK
CtrxxwnUcX4SEx3mdloCQBUWr8p0qj3mRpnc6wCSkJz8LTf+MYNRZ++UhEi4yKJ9GSxbxbYSNxew
0QC8nkt08ToC7aufGHDZdNYb4Try9y0hse65mVHR8LVkT5ql1/NT1JR/cIqrj1vh2InRaVOGyYsz
I6cKmkRCjIp6GuOrLI1Q6EtdHLiEUmbYyO/f/KVLGBjPWi/2PeuNWy2nn74klQ+swMXn/1bOc78B
SjDvsVOoR8kc3tT1EjTYG4R9371Yre/PKQlx09wXmgQ2sZT4DtKNZkDVOofhpWHD33FciDODCy2W
irOTv8VZI+L9qo3JCmmmIsK0nIi3v4vR2Awb1snYEeetado82Pfe0+eYAu8L5rOmuG4By1QEDd8K
AfmQjpzJDeiJUF4qssCUPpbI1W6P+r+a8BWIBwFQJssWGuisQQnCNnNHo3UjFVILv92MgxEJ+hXC
9b9biL/dL/RKJRtL25aEuyslrwHUHv6uDuq5iVKip6U7obAhf0Ium2BAfrmPa8zqe8TajqSp/b0d
/QcxFYUSkAmiVlNaBUjAiPcBlC7fvDRpKX26WKezJ8GrDF93oWe5MvppVSN8RwhtAILJegFy2hVW
lMXnZKM2cQk7pCNC1xghMVqO2RCfVKv7YpZtnfsNk9GKvhxrbkB3VI2loCIMEz+fe0UXkykz+dcz
EdOtAvqOILGp7Lga3JGz8/NXf5+PKm4wEDp2mtxxXMlGYMFaH+VuFyPWWkgAABPGG6TE5x7HuR7S
GtWsCocxVeQYwFgvXfVTi39hTQn8c1W6TS2TgG2EU8g1RyiUZ7sn9YKAxR8CE70NydaeLHjfkMsk
7112TcoIJZLJVQSc/ai1PeGAxGS36W5iSUHVv2jU/dXYaZDO2/Sw2kkYSIcp/D3Z9jAqsC6CNtKo
cr5jsxEt8JqzbYdQ6grTh0FNpTC9/0uwXS2svERM5qhAP9Xq7gEtxE3cOu8xUsDAWgHXfQSOnWhc
Kcb2Tnh6iNQZt+dpoKZ4efrwZGzUUbXlEHd3u5flRgFcOv1L8k4e4UqADnScz/GY1QvJd+TZpgKp
fBUqw4sOM7boq/T94QZWZ2Ox9Ub6anBuo+cWk2IVI+4dB8TUikkPcPrO/qm923lQZrv49KBJ+v7m
v8nsYdhscCU6xcxTnRX3CylijpOFkfevy/WZ/eovWI5RrXgD+skx8uslOc6ae5ArzztDliwGN9J4
Zoo2sROz5zV/0KUYUvWCRz+YED9M3Hz595nyTWbv/9ArlqJlRJVmhM37PS4+r/kEPEPBSEE0b4RK
7m3a0VKAHF2kMkpG/Xd7jxe+4oSo3pqKJhJGRyxqgzAIWqilFFpcC4fnZTphjuTkDic/B0MOBbwZ
onT3Zg6eVQnQisPrG4lJBQFVOJHxGDO07B8bBn9ci0QRF0xHpWBoskqySEgl6Bl34mDZec9Jngf9
bTVlTmwWAqw/E8LtK69968DWGfkgXjeAaGJhIB4Ww5sQAKJzbDtNxi7Qyd13uc689uDvULrD7VF6
S8X8tczRnJrvBrkXaQYYzZlcerUguqJjTeuHc+eBtvp3oVvynIz95065UUbhkOMZdeVVc9XztZbz
RP4/VqyUckXcHhqB6r7d+8RIP51YlSDukpYoUTWdYIN6Yhh1NIvS0h06haNQIZLK8kVgXOHyN/oA
kXOf7ue78pxV34nwNayIhObozK3tHnOyiDXW4Vqml8WMJWGIn5wVgxFx9NO3CqkShWCjvyh8QjcK
7iXv/EwSp7K8jvTZncX925HXLiZ7u7P8zZ2C01M1ff/Y1dpE8tQb4MfWtytc1RtjZkGKQ9MIGJyL
XmjKniDm9fJRldr+rxB/gC9THE4Pcniq8Jnh5atE0m6W94HC3bWbM/EMXVJdeFytrMDhL0mpsv7A
fT93mZ5Rf3YbM5cDO2YTnBZUoHwOH1atxwi7ncsgifl6dFjGPTQ6QVRijC5Pl6sXgah6TRiyc7Ta
5Xs9gTVlQy8A5DES1wOH0tBqOuLkbZtcxCtT9lmqSdxAwk3ydYIm3WsDKLN2vQ+uuEJH1eV4Vt57
sGzSYxrUhovl53anSZdrO4dSOuRfTeVzXKbz8eBtJp2D9ujuALzkHnIHeRXyQoyFRAvJBYcDqWLc
ktfb7F3DiLXVoiNzxaKdTS+6Kf0rlLGTGeBQTfPqkH9VSV+hvNjIZl6ve59b9lP5MCM7CgWdhpx0
qP+nLKFJ8BeyfTRg/NuwGp9hflDromOYhnPve5GN3pXeGwgbaTpX494C15YGG9+FDyb3ELoIokuN
b7watsShBSHFaHMsLpNxopVCff06xX2GD+QMABjPDXHYdPK0F/ryuBtST5VrdNhDgYNNOg8knv7F
ry/Sjri9sjVmzKhwbnsu+Gocd3wUeKUGD9EymaZoK6wleJuwM5PqDjAOR5hoqk2zehPPi0BrVijS
uFXKPGwN5wXr+ugdo8ibFIlu5pLw6NOsqSMRixCAerZvMXzO0CsBNw5TKxYBD3ymQr4wN784HPzR
Vk7Dgm2v941+8kDcjTXq1GeQXmVSad3jGKkJBO/RzZGHg0ILUYDDFs3Bq4YkiueI8EHcCOAkgkA9
jn5QTcmNkAIe0MA4G+TA7QIlmNjY75P4kGpo0loy1T50tWjNHtvHROlRVdbPOPokB972luoyVupl
fhx9uog+K+SU7S9TZFUeJHUrYxR7IVAYo8joJ+820Dh5wZTcIKVSKsXuqMBxL3eXFPLMA3Berr6M
HEpL7hptxsaPNWR5/5rF8UC4ctj8x5Tu37WLu26byiLHPEjmhVyXeEQykR26z/A9UhF2PWbnQtC9
oLsVEJypihtS4LVcMd/OYpbvHEEvOBSbM1O5HVfzLhPcdpsh3uJ31CfztJwNs/7y01tPuQE0sp6d
yqSSL2bV5ZLTJi8XUbyiQNNhsjn3cs0L8Da7BohCCnK8GPpVkI1jiCgYX5OdhXWL+8zDb2k2nhLo
jl/babXrEpk57sKNunKupMBJxMObepRq0pIG1205L5OcWun6UiHrz4j7P2SEW8hCQE1Fem25ZG+F
N7QaqkBFl04aqlW/kpqVnykePFNfGy/7rBPRMDVNhf6H9BzcITlfzeSBvBq9OyZDidD1yTU7EKup
RkDYEFfs0ae9p1rsEqKHSpDoO028hcZDypYxuOv8FcvFfaP9e/TDrQ8gwPZ+XpthuhWozaS/rqsy
fMRRms6uSIGjAN104BkATazu2qeYxzukeQFcBgv0eCb+7//9BP8pJt0zTa3iY2t1iT/2HoA9jGoN
BgSAdW2/gfWFUjZU4nQARNfFSSGIZAbfo8wgAGinGofZ4mYQXDum+1YH1h6TWY/u/gbtdEQ/Q2k4
e9/senCOPh05WDgxpcdSup/H291Yef376o4xSYjlGzSK/pE+gsiO9Sa0WA1M29JlQYehQ9pUjpxt
gkwFF6nh3zm8N4/lnjaV5Zgy58oxQnj6DHa40ylXxNzGJpoedOTR1hXdgsVmp3yT2iObKrQBLz8l
ZsZvbRot7gZC9A6Mo9F2eWMjkNQnET81SgDz8J95WS60rmXmokjsnWfHNJhIerB9zctjpPuBngjw
U/qS4OgMGgaqJ9CirmWy47dpNYbVAV5bSnoLUou0MNNKy734HbAOD8jU+cZwboIRlPfDThstidF+
pv5zsXkdKu7tgAY8SYU7OnfHP/j7JDhR8nZdwvECuf6V0baWktANa+5uxHMQYqgMRoK9EX9gcKIU
uWfxzRoTFnDJ8zzdG7762fbgJeYGgN/Pgv+b72QgDqN7X0AJvbi87niX7uUbdP9bcNYqkgrOFRjA
D4KiSe9YVJHctuqmv+ZaAv0OBPF7r+gVqWUvTWQylmNzylx2RunT15vU6wbFHA3WaUui6GqicuSJ
qa+vIw0KAdIj93UqHEMjHXAxCud1CqnohnWWJUauV+wMmbCRzGftTNhZ4MD15jGyW/e+qFGuWcGi
5o71UtEgkqIN61jGOoW+1y0p3FVC+Ox+9audSFyqNSUayh3/Zc2Rsyzk2UeZnN6l48kD84nvpY91
WYitp/5SKJWpiofP6mY0GFDhZsFlyZHWNYQrSAgS5EBTHyIwXJNHjZtLuJ3XixBnv0AuZ3MzIA/u
ZQW/MK2QalGYdqBvbLRQe57738vlwdGBaxLhFF6laxUvGNMkEr4W2Q4gu8IIsg3yAzwWQBOlf0Mc
p/vfW6Ir0Iyej+4XnqvBT1EoQOQN0H+kGS/8rl1Sut+AopYtHHzQwoHcWbWsdrLE99p/VEltSkgI
PLD1wmM9hP7H8Ld2f8+4pefmITiyNp7/QVkjsHNkNpMW9QcCvDfgL8ze3H/sMaTKvsqkTG46tzp/
fuIvQ74asW61BTvefhgVfQUL7SxSOKvO5wWNiXEIeys8cKMV1+6wcmZa+0GZRJ4CvKr9BBDHBPln
iayDikwphKDOva9Cfv3ZYAzt/qSRMISPR7uhbiUhm4sH8rqzn3cPKSWQfrKXOF5zPX92rEsk6+QP
W3QM9AN4eX5DEFW2/hfAZ6eUpn/XDfdSelIHxpwjwixc4PUd8QiJ7yQ9KjSWg8OfydXK6ERcrXGq
YWpn7bDX0pVayJZX7idiBABj+XZcjiqDg1mdhq+VY0NUgAhuoT9QaJjIdJRTad/U8xDO4uqIVNYe
O5J1oN1z+om6O9HvZwHEgvpnJWU248dekg6KJiyvvAYHeHxit6AUqJsY1u/3X4NiWxuNrwLNHAEg
t1qfX3dgDSX1a0I1QOmej+FdUj9Sa4afebybKAY284HKsROl9x/8NtapmFK3IKV5AeRIsSYscb90
500DgvF19rsPOw7sUkIbvS017ElpLONHfQo9Cxo6uNwJAq2eUd3+i1GaHfBDP0/AzDs5wvO4YW15
MLzgOBLjifEdtFbNppt8ekF5EK17zt0BbqeGw8WNPSPFL2Y1trjHnenqgRGLJhzATANWtOHVRBKm
7A5W01IlOEtqjrMee4S7vbn2df4EDHslY14Q3A/lNByq4/TT3s1J4ryV4fuRSzugNG7KJ/wTU1Y8
/VO/UsqbDbfRFJL4I7fzgVk6zN0RRwicjP9KMACJfOxNfcL7g3yTGkDb3Kjjw8dLyOa92A8c9aNe
4QGCgnQNoh7mSgdPPYSUbg31VSAeaDSRVmXSBwsi8/8f+wzWYbzazLsbAml4+gUVzLrm+0f2qixx
RSUTktPY8E7YU2nK0N52Q8Iys+SoAV72HqBPrIV3rXiGiGcdeej0LFTU/PW3KurvwTayFfYqnwPA
tGcGZzFvwxxkHf89SY3gIN10mf7Ue6CYegqdAzwtHnRZehx6IwSwVP/wc6FoHR9mBNaCwUwTmO8H
L4ebsONdPyoMUWRNQfGGc7qcXHOaiH2UXJiYZMfiXupm46xwWh5SsCDH5UoipIT536LSeisy9vCw
p7cXDJiqYVza8mX5W681emHcd/GoV/uOZ5L67r4u1nInNrMbHSfaA8/U4zFqHnlEunPmb3gaYcTm
B46e03uS9108O9Ra8NxqzgKENDmhlB2HsPKbiCemRhINEzTQZl6adQ15U+mgMAoFY6OE7NtV1z3r
kVW9fLTmXuZHYCL9NHd6ge3lKSSowNXTD8CExUfFlSXlg6zFS55LxIrwd41OwoP+HVwnx7SjdqoV
Aw8ESkS7qjDJI7IO011qytCm2xqcda70NBv46HHS5el6fzMwnQvWwvzH03n7I2YhfRkB0q/g9eqn
jg2SBH08MODMSXzfCAiNNegArbt1PtuY43gzsRGZNqWX6f1xoCichdpIbCC4TlqGfMxOKggtCnnr
eGL8MysdhZsvPl3dF6EmgUdmQCLky1AWOgVR2iuyONUQrfvC5cn/O2cpvtoIvMq0ccfP4MMggzsh
tTcpsAKZtmyEaVMpYBLmM1ObFe/sd8Ab5pL8UIpCK9m+GNw52VuboOLhlpC1tLVGkzK9/CJ8CUEV
9TVbgs3hP441EEsKdcVzFzhV/WJxR6xqQ4UsWLD4K1GYy9hGH5VlwNGV2rMpLBgrfX+vvZ6/4l5D
yTdwPGkZMtGX8B2f6rofGBFKx1w0VrX4XbKKHgsDlru/miWA6/dJ4HPYVV3HoxgxoE4vkACzZ4Rz
loXg62KO9og6SEhdvnFjlvrdq+TMkVV1SBX0+jxyHmanTDlgPRqqYg3QWGcc3+fFymTicuiu3Rut
Tg6Ht3RCzB9o+9BmMi0UeffelN7yHb3A1hE9b0Gd215hNBH70uUhQLc8Y9mBESLBoPX3O+trjK7F
fKFw0/+NaRcGsztNZrbG1kfWLkhSs2YZowRRGiQmzCJIB52h5FCloFN6+tAcOyOpSDRAF7k2rQEV
uBm9DyXOVZV6pSt0li+K+Yt4P2N90aqWv1wDiDIdY55xV4/UdIRl4cxG5jpuBjv4ltKnpK5QpkSb
Ni4QI0NJR4qet8sFumGt940emygDstYDegldxD5spCmCse9UoEHS4jf4N9P+fr+w+MYcMXyGOdOM
9mmE1a7kgmIWwn1MPrhB3e7vJfYHAiLFy9jwAe5KACKcQLHZV4QZCZgeOBUz3jAB2nRMrYDx3nzR
kcssukUbsXRxTkJ/cef7SUfc1aI9vsQo4gew3RaAIsynxMhHxgPikDFZIiS6e9sGBhQk/qYtENag
wMw6NV7zYizU70ss3ng8GVetKrFctxXsYbRAOcWPZrPCVArwxxmDqGws5tZDSL8BqF1/R3lzjLFv
6N/BI+BVMXVO0+1JLD1ORMTJnsx32v2t5wRV6sZE2usmkBFs/XljaxPoxxMqeT7czTREGr2B5yq2
n8nrA5VZz0ioMQVSR+6JLNleDVwt8DowGn9fnKv/fXwS8yfBh1LC+RpCYoscMrFnPx9Ptnhy0O56
IA5oII09jSv7bzVCgnYbKT8kqyANLTQcy0KxMALP+IeIIgk7rb7k3CcSPnZhQGOPY564uYPoTw8h
qh7pLaXuYOVQfivIK7Hx9u/GQ/UaylLj/UfksYFVcC+7PvQn7nugqCPp4DeZLbJWj/uTT66jVKc/
gOIHY+kLx3CfMKXfcSRaAsKRaz5M1uLMbaR4mYUgv2WgeRGzvMf1hAFuhBdU780uFaHGmANdw0M9
9gCBPPJ5XMA/NIhDKxb5KLdBty9mJ7ZVByi8x8mvBQQCHBW9aBbbvHGEXFOhwFmUDoBYrychP6EG
Zj3h9Ic/us/I82gveZH0SpFTgzr7CYGSGSbSWiKXGgRNymWot43Ac1ns+eFylGn3Dbf/q28819dB
vpy9Cr6CF1Ex0PMgbZCeeaOrdkTnNARcx+H2Hlb1jZoeaPm4lWWyGFbX4feT/06EkuELD4/ZOOr8
MkbnBIELilZ78pxubxiANHADwmqpojP3ckvLrcNsviMDdKjPlxUMElSL3AELu9J/RXgDhsFg5JsD
VTxaqPmgZJxBObjNYLVWMXikdCjZfF5H2+f4h/qmoVBQvYHT0xsot580giDKsfjTS/3kKcd080Hh
A+g3ppsfnTeG/HMIEysl1z4C0QHuzOKyiap11GTjTkz3AMKUE9/Ykc6pOeT0kEifUJN/S6napJb9
squn2kVFlOWkUkB1gCpAS0BeKS+9V2YoD7ccF8u4cMiF8Wh2RJ+IScMcQhjANszYQPy3n94lwoWg
QCLH4i1VrYSzy8w+JKPdeP1wBOI2Uc5+Av68Wn1L8maJdUcrOWKfuuz14g9JOBahuDKf6a/vG7z2
hE7y7sza1dw7C7prgGFRVo0921ox89IY08zteKFaJjGCASiOr8szx0qskppknqtrdkNzgA4Nuv8I
RXItpQ5SX9dT9nmyvyR9ayAQ8ZGhRzJeuKyvAM0CDKwLtUbgAPZLfAIUUrTNfy6aUEHf8IcExE9l
sox+ekCtSRKbb4fArAOhDA7FTasa+t7MiIQ/QTrFl1T9LOEL5XmpiUwLe5H8p34OrnnYS0a3AHSo
K7f65EKa8zJnjWiJNOolVYFBJ+YgxxxkaHLigaBaKnMoqIfStg487IEAp17CD51eYEEOKvpGJGEn
IzXaX5PRTL58YESkvoCk1jJAUfxGP0C0oRIlQQW9X6cNt94Z9UJIi8xCg7iJq+UhpKXHuj3AxNPs
IWJE5VbzZZ1auNUo5RmzBaUn/NpK+NgPysM5oKHVaF7sKlhRhnulsWAPG4ZM0MYtfyz9uiqEiQ8g
MCryeNuuoHcFjxwdq0kevKgsgLrua7prxajQvgvS9gw+iN6CbGpNfbDC1WalzXviJAz115UEkrqU
AFyn3a2/7mEEOHNnzXlDQNF8dR+qA1ub6Vp75Sp7dsK52RedxevxmdMD1qH6UvUa43jplwrDuneS
ETv7TZ2mDikg2t3h4e/7frZaVRZjaWVObEHUwe8tPKYWtA3vxLhqNAKEoN9GVViTtIwLPj2v5pge
+rFXj3trli1PQ2gMUOXN7vSJbNV1JWO0a4In/Jc9qC3enRCWn1ys9ebTcBQjiD0ftUNm70YbxKMq
J+IAFYOBsPFRhX/xmBdO+NiImQ/wl0NUUciV2ULad329M0OVYC7UlkyScbOaM6tTcbPKiQiCvlF8
T9U8mvCtwyrjz1SeM1ooS7yXjEwpFbVr9asouaNGxMbzj+pj0XBKP3HvjdiOPSA1Ylj145x3PoiU
esorNUEWHAc1eRobD3XfOGCXWQzTlnD0vCqo5CGOWlv/zc191udWPoawDBAFCyUKZEjlrwUsxC07
muPxgrSNaiWjgEd/krwgdl2J0GsuG4f9V5enrxwZ+Cxj/XuZ7sO1VaQGfX3WhaNC2oGnVZtVnPOg
wumrJu/gkZ21Tg3UgiSqg+4lIIMts09E4AHdxUT6++/zJQSyS/m5AhTTT+KfOeb9X6xojdzXDv8I
wq/KCUjLb78VPqPYuXNFlky0GmE7Wk92bXIoMIh81oM0mPg8Cv0fyy6wFO1fLntufSgFfsrwSL/V
z5Bqx27GE7pUVOcSz/rR+gSyeC3eLKP57evldpzP6xS/XfFgmjny/PbhncdeRxNfqvERW1gIT8cO
H7k+G+TSUf4O/Yb+UTH2ak9aVeAEkIlpv/AOIA5Sk4oBlxc8Z1CXCym+v/b+2NGZazqlZ0nCKs8u
PFn/7SeHQdKSfh6ZgVcOJiDRvSwF2xLIakpjHJWvVNGmfeDwET3V7zonbUyseZRKZzPe2xukEGME
0FxAkuHOMAH5xdByieO3dHhPTHIraRJGBX076IBCfFWaLMLSrNJq8HFjN7nN2YU3PDix08JRYCoN
XO2vAvri8w5EOfY1tk24tnlW82DOG+M6XafHetz/SBtUq8iaEcivUhA3v8G4mX+7N7RCraFz6gsi
ZhqjP/lGyVqVpiyzAlcXfQN4QO7MwINXEexTNAZ9+9rDNqgAlwI5JomlwJqkReJnEPLZLFyaADII
XoiFnbWH1BboKwLXslHaHieQCmSsfqGOpr0kXoflBzQVfRJRzTxttvDLrs6rR0+Ix+dY4HLOwwGt
PFoNlVKwMHOjUT8F5cgDW3je0QQdIzYN5ye218C/0YJRZSNtR/ax9n6Wxsy+LkOVk7d32mgBJkta
NmjRURwN5p1Um7E+V/DnTLproOVVHawJwnGgxOXXuAw5GE1lykqwPKCHZpFyQqY9Me91Uoaa8CSU
Qk1uBe6lkO5K6ssaoc8SacU/BNpLKpyz8Y0EtgCzllzuPTraa5E57xR38BEZmN3QAorm/ksYtnbS
uJ2s1cJrt1J8Aj8LzQOXQTSk5CRkNn4xUklesEn4gWHnuUNHFuIC/VwG8Fv5INdHG8Zl5A6QTqAK
UHDgAtP4LW0Hj6ZxgLRX0tXo6F3zsqiE5myoUovBhGhfjrgUc29JcFQLDJS5VqbXMCp9Ma0xOvFH
TEGicqx4uGCt+uLu85UI3Q58oyIaN06RUZ0cK4gxpPSygPTCMEEAGUlkc9+MUfpQH2BijmyEn90S
uyZYZqxPilxVYuRsh538Z+nebqo6MgiqeFPcRWlSMYUWjhqNfZPcqyYs8JqBrm3nSESsmFGBcHOy
EV91MriBG6OLESk1u89YnP877ovHzgm4vg0ReGavt26n2uHDaFAlAWxnPl6EBRe31F835Nx64mFE
noQrANacvfy12nd9eH+nowCkV64UbEDAlFqNRR84SnQZM/pbw6vkptZlwc34+wQdSU284hTUNnA2
rAMfeUpwQRHstqRO5nUjQI7U+1aiErtnGkFGdDQhyFY5rN64etVzcsalI/v0Pn4VjQnzfJ0SVxV3
3zHl5unwIcuKCVIHeBz9vWkZFVnqFYtmz90EsYmxGFPz1W4PI0nMCjXsIAMxzhX5DA+8q+lsU9KI
6Q7h0XHhAtwkTvZ8nQnVgS0kRaSPeqnJV5i6D5+Gp6YYIs7w9si+jiIu+PcLpIFb9sIfW/duMaKJ
EpEGEas8XqiESMEALd1MWXmMP2W/qIq70bE1AGrHC0xu+lTALMeORDTeDQd9vo6XA/SLfvKy5R0v
euUmNfOVog58kYxVPxgkyhmVrwMVYnpKl81b+ExX2Txcd//uYTtWjIM4+KUvOfSRrb+LAWL1gAa7
VCvrmmd1g4fTKPtROjefISDGgwaQEL2eau6E+L9PzNReNlJi2TCYTBluK4XOysgnS2zfpXLpjH/j
W2PIxhXq6igRWUWwzSA2Qd3+gLN5B5gIh8nDgOl9poIoSC92DYHTgmul1L8EbOqJAE2gyl+UL9X0
cGAH73zOcAHVKjyRcQqnZ9f2xOO/TYx0qfE1govK7Ov4GHoTfWfjkiVrxG2Levd2dPEJuqQgbBYX
pcF+Qnh1v5/KPxRII97n/Jyw9CmOIrRdRXsP7CDaLrCuBlRQmVLDqir/NnMrWzKN6trfxj9YOS9E
q86m8oTeT3CnjCA6rsm+gpB8ecntpAF4ZUpWAZqZi3BeFuj/ywHZZIigpbp/sxnRRh8Fj9kvdF9C
k4IZVfW2OuDaJFSvLFj3JM6/adWVpefBuWkTgxCBJnjwrdjpFnzYIok8iSS5iG8JgLrfYusCiaVo
AsU2xT/hX0ek+yv32HLl6ui/y/8FA97u6xW8iDCZV7jUXRjsDjIgUrDnNJFZ7CHDiD0g/tyDTcpr
B92HrDnIldWPWja4pruJkwVfK8Abf92SBLd/U3jMQiwqOPemi1RYV6hq4mmnJjOrr9xn2zNVQopI
zGGH5v0GbOjkWn0vHVSddx0cMmYbXygDYjDEMsmGGD8jSb78vXMie4oS3iB4vB07LpOpn/uehwdx
zUfe26dOfEvjqqvw60saq/pQnaauHXuco42d6nRImds1oByDc3sR8xtoIqcSGC4/EWLYK0xhPIfz
KoKvKoSArTcCcxFZLLRTJW5ACbC6xCEje8EQQs0eDNq9AQENFVl/r3bAtVsAfDE4jQPEBTp5JBu2
Oh0WLIJ7YSso9qov4bWc67JcHdf8Fo+1Kn0PJDth1gHuuQjBXGVKaBZrsREW6DreY7ypEaLBSM3F
kms5yTLHLSAxeXnKEvHofDWQ8MbRTGuIRo+6uqr2lMOdeirhfDYdn6I4WBlOrlN5AjhXbhQAjZlq
bgq6ZjAuPiF46M5haTHFa92wz8uKs+ZvmkPcOUj68fRvSKoY3kIZvXo4kYklHgJCZ4A1XiyzdP2l
e2/UYun+Efii5hMbWdT65xbHQG5TFMVujeXMU9srqjzXxkSDGNq7fIQgVhTdrZlvqicXMUocIlWo
hb1tM5HR4EBlwcjl2gBbxsMkiOZq2jvGmapePO5WWbQ6uTKXnwOgSGqN1wHDERI0apqb0iXzj/LV
tCBM3+Ev0hcOIemJzMB6g4oJTOccfk1DSzP5OkRGXfzMit8uZY8aunQ1gsb30xxkx/5uOtFCcpOJ
MvYiECXmQ2L16AxeGAYluN6BBM5w4EkrgQlgOPsXNX6LEgAv/rHmrWmYjrgz8qt69znPZotmmdk4
Kg7Mz4nlqCl8zJXilP3PN4b4JdpqrrgcqS5DaNxkRC8KpCvH9L8NhavvX72mRTO882vDzmhjqGWS
Bc/RDf8mMLt+xr9L/Ib8Xyoh7d95NGRPhlh6KgjD5Nu/4gBSsAoUyrHfIbcN5wO5799Hs9pLHxfR
VyG1Qxly6fR1MHtTL2Xz5FS6DNAhfROQS8R9L6OuLSV+mViYoyxjCAy4o8gkndlPYgZ5buaiaW1g
Lj9x/lQ9vX4Q08hGAv6vFO0gO92t9BpwStofu8TxMl2fibUzlCYNqLms3J7sOL3AYXd0ZhpwLjCc
hTCh41vJh+btLg0Na8n6UoZwN9Vv3pqtsV8QwcHDsZoOsSbI32WzlyE7TB8HRy4UP5uqE59EH6wG
pYRY6u4VearvV48gmBu/TImSMWVE71VfqgmVDe1kNaH7moD9xAGLiOohaSPY1QqGnmvDiKldC1mx
s42Fg8TXrgkZOP8cfAO6YD56e/JjpSneFeGu+ewgTL+cIrOUj3Vd2dgO3UXdkbXPD7ltfLXCMOKa
vJugfEWWqj3M4IzTlNJTm5uz3ZqFInKVrDEPt8hTZpwVT8CTdbWGczZ8xqscypN9xM9MVTVPg/0g
BxtZ4zoWFxuYzvutrX7QLWgB0L6HWqkn04kIWp5iWiiVstu6ZbMT0RRyUsRPfZRgJEdTHix4szLn
hgF7zw5mQ4qdANGJxCydd0LEQwDlMFaFU+HxVkXNY6EsEbKK0n7opMT2thTxqMaysEY4PC+aB85M
0oVHIcsSB2yaLX5S96D0fjv0qeJCwNrYFOUfA6hLglizdYeU6STUBDRa1nj3AmRtgiVMeeAjik+6
h8JdkXNwmq5ecvnQBOpZxF7j//LmNMHrdVVGr8ZfQTT1wrjb0ZaIuxXnDAh9v20lW2ojztj7popJ
WE4wJtBlW+W5bxozxM/2JacxXfiiU0Js4qt0EFzdchO3ZUcjRd9xEZhTj+NrGlp7uXvsKVUQCPEi
8rsSjfwjAGOkYK7pwCzfareRs0npgzL5+Bvz8d8OW4KvZEAIauoG2/8+EBr6mHRoBVdjrFZza7wG
Aqz26q9efTcm6qBzPifXAQZt9x7zK8jKjWsq6DW71YVC6NjNLk6QgduZyHl0mcyzxY+uPNkdvy9e
DBjGT9kU8w7hKlMVHKbKfHISnyMLWWlBWdT2WAM33ropmEFguBsBPLkvicf80562XVA79C2X/yDh
Qu+BS27mabkp59z8dYYjoYhKFAK6dWEPWVA3todGm6jNhey1oz/1sUKM/TX81mRWhHlYcuVkQhDW
/QU7bRRVQaXp7iYMhKjGP3MWHvV1/Io0k15S7CwQaqo3KrcWqFWFN0DCN5kzUXaCrKvd8fbU8mwI
cko64Hj/Om8i1+8gS0pbbhm+bGhB6K7RcFIkkJ9TP3q1r4es/5Cps07PWYYZx/yTL6+JCvRQFcBB
CRFBk5gsJ9imWfLNYS/PNwRZ6aFPf/PGEyjIf8Jvr6NDuIyOODk5Mf6Cbg+EWI7t4M+4UOS8s7n/
ix+qWimUGNe2RAAwXTMjIUjEDigpRzsCjm04Bx7TCbB/IxQ7CXUZb5Q8KI5qarvapGGJEha9elhy
YeZ6YGeUXMUxPjRoCtJ8nf6YSl7QO7YVQHXIW9om2eEitgEaLkwnpGHJEPzVHkjEns+It6VJXLXL
run0A80q0UIkT0sKIZNXe6IPS+IwXJ2J/l3XQ1EFVcGw074vWWfDDqJET1atZr6yKtfIF2qCloHS
+BIIc0yKD2EZcIMKF4DCpg0hhMN/uM9XZ4YbOEfa1rnEkXfxTUgBXYx5X5luheDx1acFa/tj8kxt
o28B0AKyXWLpyjfOiKH7r8/osO6KeC4QDCn/eNN0LSR0BKARVt7Tj75rEeyJofpE2PY4LV57A80e
BEhSzvrHCP0Br++Jy6NdPnzjflsrL1C/j/HyWA+ndyI8xZBztfqBhcylCs11MLxkNilRS0AOPmww
nSNOMLaFsR99dbYlVtjjb0PMUBEf5VDJ106QtM5noil2yPiSBCLAdRv/djr7n7Vda1G0C5UJw5YH
aiSU9jf+kPNO/n9zTtu6bk4CP5+E05SVqcY39kA8L0SAwrL1A2sIh8mN1lL69bfnjtpKnEY3WdiP
+SQ00FdAvMQbwFj8WrpHNDbHKh/+rkGLcXHnVQ33sahmAav0++Q6UPZy5Jk4jGxPC9bHGSayKi0e
lzamyXVfxpLi0JCOMFMeseYDz5W1o7APO4ly/MHlcfdSGjNGNxe/kIUA+3gFx/KipvQ0A5DHmeRL
UEnfRcg9G1ZuzUtieAVMCkwSm96Wt93kOv58T5W03+WebwOyRDSzqPdIHp7P9nXSy2Y2rVnLf0tI
xj4fd5Bl5A1aatYeBi3vbo6Y5hsbLkGybe2gYYcn+Hh0N0Vu5FyfDB+lj578a5rHMEVQ7LAbhHYF
MKS7IsG4rP5nSuL1q6YmmrfZ9d46cTKxT+r6vL7tFa9D3smrY/Br2gzl66kUH+ipgBZWXVw9Mvd0
7Mwa/HlNlZ+CRdgn7hHyxcYfBuObIgM+ckpxZVU16G01aZws8V1YxKBzzF7/kvH46Ba9FcPMVm1N
elAaCgP88NjE0hyMSPVYj5rx48MUfBEDxjJcM1NtpNBDa1TcNGimJxlwwKvyDqrBrc8f4xL3T3GO
eT7qo/Wd5Doym2R6hdEdCb2RdR7n8tcZYLzyvoOZHWKlk7RGWIJ6PA+mojnS6u0fPKEfL347TArn
KDtkzqLjZO5lQ+2dtrmyYYqvIBar8moeFd15C1mdca27A0mMCrH4FwfDSzrSsAQXIKFigYSf/yTJ
BG4eQ+yipZpJKaNnyKAyF0z/CxcsTdF8XviXoctLcu9eMjTeP1iMqqK0j9fC3RYSJ71ZhUdVQs5P
NPuzs77ClEHz+PBD3OlG4QERThtTzK8Q/kAAVTPKIBFKhctKdv1chcVSF/+jCLRe09kkSIlZUbwx
FRw4nduHuib3FO04VwKtsJjq/3It0Qx0AC9OBysxrjchC5i2yk+OcMUj9C3oyRwTcToAx2ZoY2G3
sh+IBPAFOK8pnnFpEhVaJr3AdU3hMFRhJ4htB93rwy4IPBRog2AQ11iosbkvWjJI58YwgRyvv9lj
YLOGQMoXuiKXXwkN4x2A6jTSNip5aBsnKI5IKk2AhNXdPedkq5cFdT9GEZdqAv2AW+QeezTYOE/i
d7KuT3t2O2X6pcMnRshPIdCx0bKUqO5x+qG94dPrF08WfSVyzBDmiohbwVZAwM0h6a/GMgt0ZMTE
sF0MGePTkZRbUa4IlguEN0xiAkrVek0q6+3Kver6H/2ap0ChCxed4PN+10k4bQVI26LoGjHxuQ2M
eee+Mn6nVn6eyQEwl+FXjk9AFuG0jbzqNgM0OgzgRm4yr7k/mejvUtpJ/I3iK4eE7SU+FQ51vhSc
+Iw6/SCD5W7+nTZHk5gIMZfXHJhHrmhNimUYKGTsrPbCeuLPqrpB/FeF80anGxJ7OWE35GyFij17
yrQ9SP1ioj+rlpiG0MjaG870hjMRLTlOjBIk3TuvnyxNZu0VK8r+ivtzPfrBEerFL+MIV9dHHs+k
1FIjE4pVKMVgUUR+APzsd5sqn4hcuqbkVFmKlVJ6J9G7NR0uHtjh6OKnm9sIqfLvd55iwC11DXpP
Pb+ZN34d0TMn4mWABr9W7+fDqu3Tgnb17xJ461IHXUlOzqGnbjpbjJt3cC8ieVjwOm6b24mVJFlo
dzs8UMwjEH8MIvdjFwmZttVCsnBKmlUZrpT+V9P8F8hs2XZn+Tvl69x/C9njiEbdRgGihERLScUt
FFWgqOzelTwyccthZptUCH3AfxKB7Kaq5H5NqVFCLK+qPdEFWD7cF73FbkZSbE9RKn78ua950BBO
4cweQCiapBCC7ovlCQIaxzm/PoDlqfqbpHsb0EIuIXsYxqqT7V4QdtntfxpkfSaAEUIJjB0CoMZH
mwKrJSPe4Plu7gJ5Rdza40liXjiGnPc1lGfJULSCPn33x3gYkh5vW1nOZRHBN3NsHZaowRdiJqkH
38+gSQmaxEQPI8B6RO435a60z9TwiMQpr7DnQyofcu1PpJ+2hlkU14UNj1IXjc07Ym7A/s8W4QJG
wQ5A0Ev00cCPTZK1U7YIzWZVDJ9/mDRBlEvdR9Mqe8s5VKuXOWq1Alv205+o9JZ62Q6Ni6rvokaK
5ZdaQZJ3tHzXzjSKh8+mWFQepvNxRyB5/HD/yk42heZeAOFUv8RwH3xFEuxF1ndckjXWCYV9mRsW
+kVf1g5fBwY1wS+yKjvO4eS7S0C4u/3RUGb2YeYe4BVp64Fx2t6gf6h7ipMzvfcXHVTM2tG/sb6P
QujzoPbnsTb3mpFftaJo5KobQnbK4p7TExzsgUA0705v9LX72O7AXvY7pjpuyliKmdVyeU7bShke
33rPa6D3nenBYPu4xt0QRUPXGRuWOzzM8NgvGfRNwlrZf251ra/PEKaN7EvV0fvPLgE2CdflR3gA
rWnwUHtgg7eTeOuZPoqVjTULBHnyTbeYj65ZEGGYImvF017TeztJnULItTRMcK9fiP7QdqR+R2N6
29lpqxtGtwzgeJ2LT+hzbSeo01vkOpkwUu/+wt40JrDD3AKvSq2JU4fz3OtgoycaUbqRelY+AWCR
LkTI2tvtmFbo3he/eWNQJ9UNKrmx7Dm7rOxjIMqB8D/i/cjWZs7hJv0KD0xsD2cWoQbZVeVYXhSI
drajh+5W3tIRg9W8Hs2P2gl8tKAH+fbcVvrmamjwG5nVE8yw4MNimoaLchA1QEKBLUlCLIYEuoGc
jMGOvj+h/iDmVJ4Yz5ByekiqBkP2VcjbKItpF8kHVbqeqO27/jt79EqkpHDjWXG8phBjH85e5TGy
+ZjERJwtoPzLqu12RfgR8g42PVcX/SorLZv66YX+Lx0APe28aS5I3MkhZ7vxNHavioA8i0in/C/X
hy07xL5BA+g3JqZcB1gyTcegns83r8NkiL+muEjoPO8FaXFnEH0CYFn2SXEgCE4CNAHSAlkEwASZ
rMF2T+5yV2uLh0uNv9KItNHo2S0GRiCW0LkwxhygZCF4LD3JhtNTtAzeYBqfXjWbElGXfHE/2nKL
SHZOSKoTu1T6M5HFUUe98dL6CP3fRPPfHpWyX0u18isFdUiGosh2GDaYMSOMpWtwser1761EODvq
H/rkZgbccAqqYRryJKG9UOqpOtFAvNtQrTWGBiZipVfcNVS+fME/8B6Z4KUobBR8eoum+WhQmTMn
hTO3ujTbwZFXj1MTwRQ6q4dj+4Ja/Ieg5tPG5ft3syvVylAASvbtdBsh61Rbqay3Iye9KK3exWIA
Dj9wmSEArwp5NPrXvABR6co14q9ndJU7tA8ZEn17gKysQvKj2dUSCQCeC4QOQmPlYsqzdMS+Z0dr
vmU7H2GRJdGKsWF74jREov71IHVk4K6oYLTPKsIauN3cgQqEO67bBb7nLCU6qft7/i1MuMAjnzq/
P55/lXGOfvHtnF3REvlsVmooLdEt0RHRdSYBN9ZezA5KXoYEcF8Sr0cDgh22YcmR1gCVvSekGBGU
6+BZc83FCbSrpAL5VAC2G56IV3qOVPYlIW5QrDu2xa0B1ZujfyZAWZIdbJo1RlmBOaxrr7F5FeJH
9kNGKMAuNb/vUSUN1h7Jk7/XZ0lIR1WvcIIu3/979oAyd6Jkwf71A1VHeQmGQtz7Jq0jUrfoYOsS
tAM8VfDmxO8pjdkptZbutU+Ym6ZhltlTztcKWy9OHKsWyJlEvNNgujGg4QY2KtQ7ALZRTzJnz1T9
+va7vpYKD03LW33umAgij5aSJ2MiL7jm3grvmRWHlioA/xNbyelZzh02VKpvwvvpnwa5IWVRzUXo
LORyC5iM/Z7uSrhrOSiDXRcyEovzQrJXl+OwTaezKgFZPi2xs73DJrxafU76vAxtgMToFl5BYokp
zdr2mIVfXjoYFq9oaGF7/puSPUo+h/6OfjCxACh+SNpcPsE0XNnhAGSlw7RxNi8w9L7LqTywe6e7
w/vCBwy6TtuIGRHd0ok8mOL7eGc3P8SpYazdxoBh4tqSFl1XAYR1QDLhHdzO7KHPnuPOpCHLRkhO
JAKxKTcljHMohvQ9/HXCCtdycvfYXstAVDx3rk+0xxU0hUy7GP/iOjRARLD7XtkZjnw/noBJw7Gg
oiNq6GQGSUdoemS1Ol7tds0A29nnQDlfug24uekjLBoDlGOHkoNDVcOhkKEKoSrb7MrDDj7t6rxH
gVh2k4FfcmGYuVelNKUEqm+GO0h7SasJgsynWc1AO/hZJ4ZHNaREXhtp+u/1HBVuM4g8Tpv2UDtR
n2DBG275jp0FhZB2IgkihxaaDD7xYvRYFthwiddRqgjNKAso1efgk/GBpndUfT5+1sXSk5aObzu0
0DE42HxOsoQHFVfZIR1bfA3Yc6bCYrL8o/FA4Yym/CzshfU/xI4v5rXNqEZaPnGEXNolRaepxHt9
d6dsnuRhx8UXuC3g1Su203hsFjn2n9otGneZknsVP+CSHvziAYaDGNfPRwEgqUDtDXI0Zwtz2HZ/
7vu6+zErjVEit1/m5GvXVl/Yu9U4Zco7/zAeZ/b4wrRStPILIhb1CxFTu6rfF7fZjyTFXiSSsx36
NwWAnJY1yHiuJrTcVzvha+GLZNyCKf32LY5Wm3jiLAly1IKepcddStrgReIXoG7FId+CuUbDh0/n
fP8nzCKqzWgUa5EatMXwQvVddCRO8qgpysucO/ztLI3mHt65EB8TWNLVRJqxTOAhzM9g5pB9qd5S
kxdCiZ6JrTOkcZbP5MuUHI3qlfntPvhJzNyXAcFYJclylUPG3GMJa6lAxwNrRJCuWHMnP5VhjN9S
vzt2tTDgykq2h4v+Tl8gSif3yyEA4TvaCJoFXMp+v8TDzPmAR9LFGAJGaa8Vu7JjYLviXghmExKZ
9vG0THF8+3b+9WQmUW4QNIZ/1plg7SFzTQRhzVtySoKvUL6uSNBT1oRKptRtIsBRfXICznWNUGF+
uIbeV0tj8MwnsCtWBuAFh5kCs8FpfW/6ySV1wD+jn2Rt4OVYN+7bRDEuhdzz83DKBye+Pe2JUoL+
9AZmHk5/8MAx45jSQ4c5BkmzWKSuRKGoFFO69I407GEbz4a1kGGk+c04R1CpwCz/ZwLY28J9gzsm
T9WYxhuyu065Kk76ldOwJngzUvazKM85+VQBTRbnvA7lCrPwXqUw/b4CFWevRPc1DuFnHMlcZMDk
vfLjADzPqTcz1PwKLCfcmlTXuqlDtIesiIPw29UI1YOhZa8TyccXqSA5W8fFd16HtKFVgzq/eGjo
PAkUIlLVhN9eHIZjePIsWsnNAJz2cUliHREg1EhWl5e7tTlaiqEz+hhSU0CeYkf5tekJ72KGAU4D
lKrVDAb48l3i8W4zBmeWrVbsautQYX8iy3t5gmHxBfb62bE4Xu4BMB1tIGJ5KqBXqhrLsFaB34CX
bl1kGyq9F+2zTmRTprk//3pr4tLrIRj/SfkNOeKr7DxYdy4c7lKDe7pCdnomnhQvKiBiLxVGCjVL
JqMHhhiNmiQmdURLS3pnWkCcYXn6cVV+OYyM3ObYuHxvXx41hRL83HqKO63TYNDnpKDXlPrSVQjf
e7cFe7sGzzB9c4iBWsbLOxjVxv0r1PUDQ50Faw1Gqyeg0ON6+877NDvRCWJSVg20qjgEYrP4BrJ2
CwI5O1t0jxRd1w5KAsPdj+g3NGBzqKVPo6yGKznZAXiCs3BhKEMexJFLhChO9zwN6hXkmmQosXMd
I+bWG94a2no/Vgi4C6oILzwXwfKqAd4Fzu8z0Ynkx36r6nK4nXa0Yc7YNcfkZ+yYte2HFpqV9GRk
byOShDwSZdtLah3iMXqXVpzpEipkk6PdzbQnLzLBj+KaAZj4dmGMOltcgp3qH80SSx082zJxyHvj
VIFjnZlfuzNANR90kAstZmOJMZlP4I6FCTo9bxB56amXvjdXRpJqCaXPEketY7Kw+7iPy6aBWn9S
DzaN8WqnNeO+LRVuPaYjzpIEQBWVaMFhXAwpnpWX4uGp8Xv6nNiQtRggtw+iotUP1ysWGHI1/orL
uqQ9F0kXnKhdNd9JuEICJGbO4E0B2jyD+GQ15OLGrf2F/KFDZYTNA3sof7JsoUqzmOL8Z8j/8pYT
L+mm6+4UyMtp/AOmfGcELt89DUBqKLscY33OGG72qpK7VKgsi/9iQiJpCazbEy+gBOReSEypP1q9
m+sV7shpPr3yPtsqXvdM6smILiZp7OhQPfzF1CQaYD8Q+vlol4fnwSI+AR7IiE3zqsJ9wVKDU+mS
VeZFY44oTPqht6kOC3lJz3m2qEis1zrqLflJdwzDNTM8fOQS2g+DHEi+tukr4gK0cKXWL8WV+7p6
uxNlUvRiGC97JHWn1Gn9sahFWvpAehsDGxZSRuTKGZfA/sGzkvX9RTBWwDkhcwUjBEQ5FLscebRO
n1oIdXykhxsKS8CwE/3cgY9Ld1T2ULWSBaceWFNwQqyQlmG+xfU8bGY1CP7hd6k+7CfuYwz/PiUl
DYMeUuIZWVnP9NuDo4nyrMbtBXv08zaC081Xab/Q4KnCkgaffl9QS/ZBXH9/RMQs9PJKnrQl9FyP
Ut0XV5Buwfll5fjbsGAZGaXjwz9H/c4NqqPOjpytugEbn0hoAXUTF09YzlrRMNtWB+XHeL7hQ3MV
79eo1fSyV3yp9EzA+f9Av9LXJzXWAsfqXXvuDQatiuoPSRzPfmnM8HAX6DFiCVWcUYPhRfoNx+ft
9BTAsLtiq7DWKKtxcpJ4EEdwSqjho8BKkU0z2H0k6bOldqlioBE4kCKPFIKNBy6MGUAdQ5cAYKzr
VyrIUYf20hqQUxjuobj0AbW0ISXoNAOL9qIO1wn4OBespdIY1mY6et3qwcwi5A5Syg1u25dhyfDb
2iekMCBkGvjlHLJ1tE5p9Udi9Zz/eUkyirGlUN2dfc1KUuKZYyqtdgotbZfoyyzwshpSXFtHehD0
GpY8BoCjppIGbwFnv9prdjfRNs8WHCmQswc2psG+bQI3JJ5e7lReet09Eop1WJzZNsQZgS6G4b5h
nW8XL1snG9xQ7a2R/NWaNSdNBur3zvVUKxLSK//3KU38EG7/yrLqa1duNTytA9Q7Y6OlZDARaIy4
VD6ljvW80mr1XSbBSQ6pNfi2YNsvGM0Kycsa8mzysbNW1HYnWw3NkE13Rjvt7erEqY7cwCuWvHw3
INuYFiTEND4PoPB1PcAVjChmIWmqfcWj1AjdZk5xQE+8e0iYY6kwR912mNptcVTGS7QAwGx2LbSh
oXaB+kv6a8tDU6WqiPRCrpRipslSSsvwQcCSxKC75pit9Xf7Bjge9WdeApRlKSFNNpjx3OZpMW5I
oo2ZupYYHUH6KoLN8unXAptTYHeE9n1Mfg+t1Fn6yiQzRkl8EoOz5lws+P1TVtWGp5kq9Y7DOTkm
HdxvNnV/VoedBMeE9tZPe9nm700PRlkKZnjuHVrZ/0/by1137kFcauUyinaZngUbdBoUPuFlHRTT
BPSOv16gM1pc5wBZnBKfN5QhOIDTAsgEPnkcwA9nxiWXfatqO2mRZE2/CaP9iRfBgnxuYlKfT2MM
yfRh8tltHeTRwMULwexbz/F5i1u/7e8F+P5nGcoC3TcD/DBkfcVh1zVGHwqbJMyU+l7GVVkFvsAZ
8GKYAPbObtccOqlbjApq8VYXDbxAyYK93K/7lR0XqtGx4NKqQA/XJgzYVa2YTmGoRW4dLhKOrDSb
6v4qk8IwldmSpYkr11fIl3O4++Lm7GKqubcsixcbgKiK6aYaJbTOQ8PBiQ9O/W29SmuWkvEcGIwQ
MEoGi8DkeY+knKwmpdN3M1DO3Ml8Fwy3UXtpebw4r+VJym5fGgEbgCpb6f7FHDb7zVPCgYED4XnS
7hsW/BlTHk05RiILwLL1TGI8VzeYeIP7S6EkvDoCQg/wpF7PztLdUeG9y1J5o5yrYc3CRVUOhAXE
1LJP/7LKSg0BfAFX9m0+Zbfh2MO6dT1IYfqTxM7EhYLRNejSSCUAVebH88iK0Ds4pPXGJ8Spi4Ma
aSgq57BfbzfyUnYyT9t0h59wl+aXbdKND6KHvD5QFsr71qhVASvO0U4D72YIYj8LnpE8lCol3Jem
MNTYGQGy4FQjpkj+AqtWbD9VETT3pSVOupBQ/FpkLgYTzovKyTtSFy6yHH5PnXLvV4jqT0tr6Xlt
OCGTL7TAyYUFyCWLZpmOq+IBZg6O9oyBzLdJ8gTPGVcyhpWhfoCpbjAt6LFmWrOxEd+VtlA7m0Y7
QBwHQVNBftZyGY+gRya0IysPvIe3PhEnyqfhMrNL3aN+DyaRppCV0ZHtadsMp1ScHO8VIlYZfU5w
QxoVa5xyF3Xs/fe2HdvcybUsFj4zrMLiZs0yiaI3UAmDO2VOAFzj8B15n4HbN3J28THhBiNvh1Ok
MrDO02fbSbFmPZ/Mf31TMVEP5/+JGNRdbuA5eGFhSccbsZwTgeoDDmVHnCnYCzgvrP1bd6gBTj/M
32woZqnm2geFciXWr4Ft0t7RqG5Tq8GD6g3dCvUnx1L69QNdHLEHfPonpRleSrZmwixetY+ift36
Igvfepr7xyKdJA5BuVSfPwUP9NtwsQbKcRb6armre111gPdi6wBnaTtMhU1j1P/9rErVbcKKZjgU
/EA2cfgWxKf1SgHabmvfgZ0lkZIT7c6hd6xJfVWbTyuvYkAi8+t8rfCYV3aDOSJ2DSS6uEtatRDl
B6Of0u97JhML0JmPlX+ohnrKE5lQyYcl8dloyoeX2/AApjy9i7s/AUIOx0lCzCPhp0AhubwR2eoP
T4ZtFso4nuIWqN0Yj6fulcKXs+PV70hJ71klIyGn6F3Hpa/d66FPpdrmyzZVmgGsWAC0hJ+f8WuN
RgAyUZ2OFFGLAs/+U1aEwRBl3nXjXf260ANYF3yeAdtosQxwSjfSGg+05Kztilge0YrkowiwMhgj
6bk2xS0e6DpLbk1BFlwLZ4YCcv5hnF++Sd0wyhPEC9XF+2aKprleyF9vQe/0WHOE2dYQUze9nRlH
MRNM2siI5OP7yn7YlzbhnZrr2WajhuEyTdLFScrxgngSfqzMee7TLmXxPtuVe5cM6FKFJAx46ZRv
Ww2YzzGZNs2mAE3ahhHsyN1SzdAQTBHY2hGyaLGyPmPqgzTvkuyPcEC02XU2F5dCjfqxfOmW7EAF
K+5akVI7o2Wj8n5w4ydKhIHodI/Qg6nyFbgDKZEJBsi043KWnUykvj+4Al7/3PJJRG3/zJ7Achp6
qbuwypAyigC2BlmC6qfJPMNH5gMuE8S2M3PvRA+t1MTS33PS1TzLxKigJrvI5Y9OABd0kbHjjEr0
OaTPrXHZlycE9VGCPDQRO6jU+lLiggjTJMbOMb1ZmX3AuRxVFuof8BvCUPeF7+JITFKlJdOe3q0x
wg36Duh32prksKuT0xSynR6fC3PypkrGPPDy+7ORgHAEaqfaWW8sfFysEooCOI8l9xAw0YKHqFNK
KCsTkkuRnZkBfE88dkfXQLhnn1eRIfSvVE+bRYboqEJoyKmTHjplkWUqei0wlM3gguJ4BxLAGczG
2HEtQ9q9CN5zMI35t9ZVc0xxktaCyKd1xnpB28BEwxJTAe4USERHm77ZN9Cfe0jLNU4eS91osDb1
4I/PCFy6bAsilszkgFtiLDofJ8cDeMZ/OKKRXoCt8TD5ZdjqEnrBLnVGBxqcRm5gv1TJ3gsOFQtz
y9SWRwX9aPzGRiOumt4/2XGNAXhde7H3Lh0KmNUfNB+XYJ1JeLtU5Jr+JlaxadG3Ty3Sx3OhzcTz
YYDKmZcA+AiO/xAmZAxo3jXKwdaZqwFuofs1DrEaIEyxrKhbwN2a8jkzuwLQgM9zX/dDalk7br4B
0kMLqEz3Xp97IpJRTh3JqATwI+ZXLocAxpR7YXsIwO0rfuuzgs012cmJKYVigDWC7Jl4faq4c+0L
7Z0dAl2Z2S9p6SUGWo2OEnhwz3B38FdghH12b8BMHpkzjj255azEl2NURPv7wnUlnFytQhDNOrHL
JunlhDYM08nPE7VhGAwPuQEV3CXEYTidAWehqQfMT2bVVhJQr7YOAFGnOSDOqKAM0zAXSudnMjud
LVR6i330Al0Rl63u6BfdNFFr9d+bscMHrPr7FtitqWkEy1fh8KQob+Sb09cuFF+OZs2aJFXXDchn
1Iygbw4FB5LLBqXXVcaTEtsH92J8Nv83t+SGwRv7dN0tF6vvhzbu9dkgEH2h+q2OPqtUiB49Lvtq
kzSHjBaBF5n8w1ITD+XBCw77kFesBUavutsHkqCqEN7p+yKeHNgzd9XeQANWQPlrDZ/tg3Z+Rd4z
IcqFJq6Ny/mdnaCqUq5cd8JAZRatJe9DA5R23Ld4WBSwyvxwMXBlpH4eou7mEA+hylBEB7/x4lQf
UCXa7bNPFAeQDIKBujO7xlFv8qERwbKzQeI37giE+bKPXVUbO1sbofj/hcj/kqdS6VBP3xm/vJo6
t0V1tu9PU3P7XMPJ6+4vmRyTX5/yZ82amAZMPY0fJJXr1giiRGvmNJxesrGNjlF0cauL6WSzHvOv
dGDwMeCl9vQWfq+48gmVq9+v1LmmZfpTa9ufKshIg1/9mf6XSJzLSujNUVMOU51Cjj6UHG3YWGkv
I8u91ORxSnase7sy8fGnMhUo7i6Nzlkyjy8XZPQ9OD/Mj2W/eiwBBjHQxFnIiNY5XpHaaE4JWhLY
hjo3MiaBv60s8I8MrE7WZjULJ1DzWkQ5YUsueJ3i4zxBdzcBU2NtlvplyUPwSMunnkKVJprVKQ/d
m7E5lyUtnV0zJZ0mP5hKGRVV1h6wTaR4+f38k5mpv+42DzUJSU6/kR/Q7iJ7QJZWOPjNBuURbMdG
7xyQjj4jfb3z4dSelMcJOvy/E61KuDSdI8zA0F5o4y/J1py9DSYgLxeg/g2qm25uxw6Cyn5AM4J+
mnMz4cr26NzZTN+Jb3SxTYNnQfSQIqtxHbo66XxOA0wP8fzhudQMZTuhAYtT3Vr2g7MVeQFgWXm5
vHVEfNLr9+E2JmRjOwL/czB3vsoBDdVw0YhZ9tRTrr4DZ6AfsUbUvUd6/tbv+hOY9Cv5mApVHlpI
++XWUyAuPvUeoN3kquzTU8GTneqjn/8Taz2rgZS8RTE57Cl5RW90YUTG5mNQn8TpZSJe+A2llKQ5
wUfNPcWgj8Fw78iuuZa1eaj9wlgFDsTtB0KOzVQF6s9DNeKSufe7bOA1PQjgXO+Oy2qLyLRSaFiE
9mq0ywr2aQHuRJX/3lhcKWQh2fsyjOaLQywxeYsB1bd9hgNg7n8SdC4ndp4F0BBm5Qbsd3NSHL2f
u4+/ndgkKFN8hmdCalZ3T51Fk/vhWUweo27OO1/gRfj7xqdRY8+o3eDJIEM5x3Q+Ya3wXfS1Yrez
GBE0OEGup4MJekynWvSaTykhgA9MnFC7mhHOzbrVBzv5ZUiuD7cFHr2gByLAfMeWI68JZ4lvc5wi
bGEXwqA/iWPu1edp+0HhWqtshaAASWbLxA4yIEDfom/37OGPiaQrujfEFuIP0dUwMDQF3IMFZ3SN
kkF9R4BAdwnScfgCDW6xtmWOZ5XM/i1DTJaN4ryoAreYV8nH00kfvpwp4eR+pJeLhnApXYoMqYOi
hZOxu0jx8adPR5ycT+qF3LBQhqDziMhup/c0C8OojtdcLM2EcsI+nOUIjf2Lcw9WHXzu/3FL4xiv
qHrhw9+Ms4LVOfNhOfTYq/K2EPpkKUpMpRm2/zuq3JjjO8G6UFyCKDwm2LT6ylGrYVanzXIev+7J
/XWImnNTcNpQ1AgPYM+cKwiBK8/PuEGDaFFm0m/d4h3hVfmwj8zhGA2O071AWED+86S+tT/J1r55
HNXhYnfJTwbBouJ/OGtPeIgkJOanCA9nxRffIl3x67M+58i3sN1t54pENAy+xQpAHtDOLDVlYHFg
q7l8YlknprSFQ8GF5kU4i3WdMihsv76kYj7TxRQe2bdIIh5XgXR9SqKSJOmaXGbcrBX8a2/W/23E
ZJsEhiCtJA54fniLdWGu1vHOGMoL/aGZgglD2fzxGwDiwKeqf9AdjvalGTzpXqGZKvXl4hBhB7Gs
L2RYEjUvJL+NqAW9QNcqdGGpsfXiONSe8WORvcqzpk52OBAzLQ+57yZxQ0RR1S9Nm7OdmXSYOCk0
2IniZnhJHVWxrbqWMh6LL+9UKD6xda7aEBra2/aERJkJenhrKrqpNPdUE2jBdWFgmNd8KEhDzIEH
cs2+tc8ROkk985DLMdfcUErD2KFKsmFAc7IyljzbrZl7UoBud+NwZN/ZH0rr1rO4XPjGfjPV7vMv
7Kl0Rk9VSPO5OdquUozMI4ND8O06J9xDiMTCRYto8GrPw49eoH0o0X5qFq4phJaweuyLA8cmkaGQ
n02fIkoZjnkCZazt9YCFpcK9XBGXC1t1N6SnIs6GHciWPHtMv5OPgsEkS2j+MAzIgKpxDQvdKmNs
wIQngGZSal7u9STtSaXfPpOBfZl6tLmUjCC7F+VpUsEmxGJ0DbJTvn1dyrr7nQkwuspNCwG220Gf
UOIPI4wbsMTO96f0mvTiKGR5QK7sSLXTUkCh8XWCn3CVLGd8QguWp2tswbdNAgiYiO7ynSe5aRLm
+xXsbGOa780Ai0Jp4KcaaEXiH/8bU4ee9EepLuBYkKoLsJd1N9XVHfgE+eDeWwrzgJvaPlv4mQv7
vj8BQcbL23daNx1p2+6fxcMBvo1uD87d6K2sV60Hz2K5aNxOwDoEbkIdaEWnVAKr7ZWpKMq/sUxS
5t8gFoAPuHt9PanCG6YyDwmjDH/WHozH/OsS75KlwX+A+cwOsPML3wBZs3m+5lkqIk22EDjEqrSb
IiJJXDJHp3iEzY5nyQi3UX6L1EuWVzhAHvAKsSSM9KogyCy+lFJ7T9idaPcH2MGs1u4mCC8tOZ0b
clTXcjtVKO0alKTCstw5QaUKjBp2BbQKkN6G0bkgQH9odrGWElAQI4ghBoEi57yfsHvJOToDhKD8
ML+haTojyl6fJBttDHbjX+ODyieMEpEGpTX9dVl/8v/G50ubgkAQ7KK0Ym6k+e+TaRdehMQlNA9E
pqUHaiFHxAd57SyBRFJJhxwmZ/xV3tOrv/YaedgqfXgsbwjiFeHko4trh3ktBEDIzyIbkhQXqs7b
KWxiv++gWeio8Niu0/HKnNxe3RKBI8ZYjd6T4EVEYtlbE7BFC6iScB3tAV+wbTWkEIP4uYbD0pLD
haGGsGeurNNkri1VXZUJvHIli8SUtyh7suEntwUZe+RwSiRoB0yMqnyl/VF2NKUbSgX8VzWZrBR9
7Wfad5F+pKFgK5SM3Afj6atQXAFcGExGBU6qqgu+4GhxhUepj3uOoRu0Q8DjiQ2SLzCKOsDCyYpJ
H/JNUOWsRnpU/7ScBF60Jv98x5URKoTQfvoiq1oVGsDH6F+FUS9QjpRug8UKEHG1ROiaJWWx23ch
2M/7TAY8QC/ee2xWRLfU6rxPgl+Uqglm35ZRTyY+AbSjwmmY/F7R2l1gijZrxTyJsNkrDSRr548/
HXIVrti632v9s7xMV/9OL8jaZAGEY+LB/+bVKawPc9A/Rm7ogqOJ2/1oCBlH5cU9MAtC4F2xFjSC
nDxBSKe7e7lIz6cV/hvXzU/F3dLTyDPzbtbDaqmWwZJRJtEMaiJnEOphMoycbdHWgmAlPa5QYJIC
RFvJWFvJoIpDHx2VaPqZIy5zE8EpsUCA1IU8NF4uRXGB8McofeEmP4YwLoByqyBiUP8eqnLLC33E
OWRGM3oe344Gxo5WccUs1ZaN3HCP5+LIog2IxTx6XKqvpA9w2uT6ZUlAGdMk+lUMFTmT0IgbPwze
rx5L0kZmxlPBLu+6PuucwpMt+R4/LSvscYSh5E40N5nEBphcaLeyJfKXhborqvwlacLXbh9R1Gjd
W6HThKvsP3mp2Cw3ErA++vHlv9NqtHayOF4d/R8L5xZ3C7Oj3efjjnkgyaLpJuGyKds3+O8vsAqy
nvfy9kgUPJSjOFZ6jIzuVE1dGShO4RupVEXEErmxyPuWAzgtVpKacqPqfel5p4MV6mFIgS4t6Lsd
lzpxGYMUVO6TWEnr/0mQt9jCkbGJ+mJzIopQvCBk06nqQOeebFW/XzCCe1TECHNMXNVA448eMfuv
crjQf2sPyfsh9hR8bR1WKXleQn0ixBQwKwZUJwBDbWKprMKlWTHQ7Bh8ghRvmon5gn7sAYQ6zsf6
SmKWjWXoAYyZRMnlPlRxSdTDNvJKjj7lNll8PwdaiAkrrsciJq4Fc2TUQyPaTM4fe6F1yFRyKdWS
VgKLYIFujmTofUdPrBn4AIAHk1fkrxRbpMfEOQSpNgelJaC4vDhL7v+mIVdP8HTLVCoYpy9pebnR
2xM2f/X0bBAzjTc70XNxMS0iyjHH3TC3a8ryiHyGOX5YKlAsa9Ljs3CGc98arr01MVYTmywj+y5J
COjcy+WWCIclEhBOY0nZvGKOdVzge37ycNLX2e+9/IvK3Y8JYB05tEaT/amlOOT0PKu+B1kYp/do
Xq6/RPQwj6FbtJcP85ReU2iknnAezKdYb7cvJdJhZOblpcklm1CATU7MGU+ea0ooMWhuiYurTOzF
hxsxg+bkQQyet2Z9owkSVIyYYX6eEt8wfuEUSFM0SQDGuw7Upi2q9gSng8/6gs/EG8eHZS9PMNRW
zDICbUfyyO0LM5JAK06YWCozKFtDeA1alE3Wwdse8FpYssstApmT3A5yGTwuzxAOybwTLgHq67HK
TMXByGdf6VNHBbGKumX6QyYvEq2zJ+yo65cYLsgAKHr4qo6brB1uphJZ2ORLrBz94KE4NddWc+dU
/pPqgda9QIijAQMANTT6ZDhpziRW/8xB955gcFNGMKuSTBWCqTKA6CV9XFpsgX2EtVMXHYXAU0J4
Q8Zs8/lDM0oodziEk8kUnd+wCQg64YQeiYLukaM0XtbKunFqfDPqi9JVZlINHpnjWj7Q1rwUUoa7
Jnb7AwfvzqxsDVnsXoWxFh2V5uQUZ4r3q5o/46Dz6N+s503JE9cCU2SSb66cS9z+VvgDFAZizlKI
zjfEEHITY6Z6FAl8Wcuy0WboYnC5u0Kkbgh1hSEExtvJASeXrLRlPAVXv2KPvvnVWypclEeypqko
2cku3DEJa3mjYffXvWwmOgC3XSChz93BQCYdu9EN8+10plBm7rhCxBoimL4BH9bxRu477PWppzdt
yeI5Kqtl4/eWyI18EMA+818+IEMW6yGSoPnDcP3xCAnjtDjGVOwDMnPfDSAdiiDR6Q8H7/2iMOZo
mttm/HzwgPFbHsQcAZpbX1jqsk5xrdz62a2+LKxErtgIM1VAklwpGPeAOAKsnVmnqlrsMvDWn7Ih
2f5Cax75RZxZok5jdLCDYjUq4ix4xv2v+PolZdwNHKvXlG5s8/ytOrf+rQ7Evp8ub74aSJEb5h3Q
uuT9opugElxZlbpm47giEPQ+Uxs2X+F482doJJ7QGTJG5+NsnO2O/OW17cV6cN3zlXTI9N3Aez3t
+V/OWMKmmxcYZEeTvOspCURvUhQXsLRbRZ/LSP48j2qNaFvjwDyEa0Hyk3Guae3jmlr5BYcu4AU4
JIpZyMFXaCZvJg13N5pmSMOtKas1/tANpKKGfxwOmkEOxxO7eCybRg2wfhoQUb4aXwFmNUxqmCZ1
eFf2nyzv8rrQMD822wvcQDNuEGKAab3th0FFHInDnwC/Nk9QihmFA581XBT8irwVQzm4+XiA4wjI
tRt95LSoFUuDJrDGvHma0D0caqXr4V4FqXaFYM+zU8gxAJKMpFn+OdzukWZEO8lUhekrkMyiHwa1
Tx3bDRaON6vfWwXiKh4T1/VlD6And0X7S+nMFPeOPXwZm+0zyjisFZ8664+ojlMZ0qBrtFpa4w01
2BMHaDhR7uYF0lIdnpUqQkRTSXBV6+d+MGnd/2IbcfyHCwuwd+cRNFvWkIzvfIkyezgj12FjpK8S
+8hhsm57fsN+xdXQjPD6pib6KuWn9RM0bkaMqoMwhucd4abAEIL5V1VQCKv2ldow8BA7hh0B1k88
KZc46inzpfo/FfFmZ5lkekJ5nCmPhM6ZmVWplDoYHTje21tAyzu2jxrXF+f+zcDeULQMAQGt9JaS
O49ADdtxWGYO8trcdha4BDKObc17vK3zMy/RU15n5DVTfdS4L+Duo7sOtP75w6Hmvr9Vn/YTyS17
JINl5xrZj9OXhkf9U6eh8ZMeWBNM1exU2VQNeWHniQD5oQcznjXlIeIg6ixpZz6bKsWTiKSu3lX6
cShQpOWw7UbVg7C29NPtj2OLOz7R74VAQJxXuvXdZtP1j/hAZT7RucFJLAs3G1mmBE/eDoQA247/
aeYnviH1GGeKEvs0Zb6m6ZzAtK56hO/2H6OzDFSAw2ejf1sliKVRsCAsRWy7qKTJiWqPwpf7882v
xqAUZKKGVMFpPSuaLh2ggkAW5DrG4UdH3j5KDo6C4YiR9HHFPJ5iSrtw6g9wQPOz/BzqKFTBhGpN
U8yySGcCTUudths0GCB5mg1G4uSr0f625FraPja4Bfp6QyiYpHTgZ2UsA0aHOFig+GbhcjLOgo53
2gS7bTL2gTa6QxUWbZd4Ds2Z4w9+B7yHSHkJKF0YduCIdYBfeVSiZoGs+FRoH4lHurTdUeGxiowv
9L6iGkMx7LbkkotBnnZA+oUY0KW0q/Dv0VOpZaC+Z9/dtZRAR3sQNa4JQnuy59nj3wAgIjwVu3de
Bi8Y9yQlGlabUKcvqHt3PYwTyqo605j6HhfGJnRA1zSYUhcsPeEu+UBlIAyKyvMJ+3pf1bChNvmt
LdCrpW6X78iKh4lPt9utWselpgO/1DnGb3xrKFIPoJ4DM+jBNBN2CSpeK/e4O+jq2AUhaUN6X0zK
ahsifqSjvpjFASXyyX2E73D0st6bAIdpwpFPsb9PZ8xHdNu27QkpsBY22wzYeQKiKwa4f+jz0lQM
ap7zFfv4kyiLfWA4szaQoHQjm6DbUZhCgr5xR7Foy5ywLDDGIIXpKSneIxmsazsyUwp+zVA8NVrq
+sASUNNiFDK5De5Sjf93tUqd7a4gMGRgXvBuBaDzqcMGYyPQgosrqnYELstuWuSa0LnxTujrPOm7
m94YWtzvQBGYFaQjuG/abyIg2KTezfy1XBeEIyfoe639Bq2YcGwxvvzZTu2DCOD89H279jM9Z/Ps
B72WIC/1q6ECgOGm/uBsXKarYIh5OcpezNQvs3Gh5mAvTfhG7zEW0icpf9tdVzuoiHkkwV4Cv3TY
C+Bzkg5ZhVbIalQtHULtuhGqnM7ctp514hxn+YQmoSEXOxFk+GvIzR4phhia0cD4wegnHm+hW4d4
xDwQmiGBU3shBh5N6EsUD5P55K1QMqjvWhyoAdqDzP5WVecHSvM0tfg4xzlB6Rs2/F+KSdRa6wOq
gpslMunC9e4E5lMbR2DV0Gj2MHdhc+tmE57ABPI5jumbYsm6WpaPtATNv0ouQcHLy21z9vc1MO4h
QbG4GWSILR0n4yk7wtEU+4DmVCISVc3Wq9Rp9khSkR1Xg1ot9+X7UJ9PcWyebvk+5c6xGYZuALAA
CzpBHXcUzJ1QnaiDRXLLYkZbqpGTUXitI7o3mSwTJ6oIs54d/Dm6ElzczGsejrr/ePAQ8KeTo3E0
nuvBB8BYy/2krH6R3nU3mWymjwzGpCwKOhsN6UiBg5fBdXkI7RGSG8RCGi09uy1ou6cdzV9CC60o
V1zOuTrD6eSELFkQb03BId9PzC7wq8DlWUxJpyuNDLzkPSH01yOEM1WxjVhIKJSFeruPr1BcTdQF
x5akP4ZeHLOjywm6su+VCrofJQxjaYiTjdI8SajORLFVIWsOW2hNLJPX2HEwOqYRqgwo+aVovHgp
+6Jyi7y3+6PbWZnYWmh7/+3Zabh0IdGBk/TWEYj0Ln0nc8OQjuvYaB9sgDcJuUgrLlVFyx19dDdc
bE+KDUqPh5ppgaNvfhUO+0bRJav4XCDQTR7KrDcGLhl1OEcpsX5UaSWxd3ofb0Zyn4AojGaWjc61
njQ/pYr1OX+1vMaof/3LIPIQMShhmfWhudVUCEheS3uAz3IVCX1ZpEQclZ1PjyYGU+nF9bcBhOJS
jEi0Y+x5jyGh15xWEAHcbpSae6OMEMgHmcSV+n0DK0ObWlSUV/wwvPAHhQkyVpmN+AoBTNxw+0j3
fK/YZzdo4fND7yvOasXWMrBfea1nExnmkDbcEcLzr7A7GwnV9KiRrymBg8pWaqQVWuTPfRlXtWPS
0f+gH+PZMRmh6OWFH6K8u+/B3lqU00fsDIY01YZeQ7YSUxXkU3FcqRQ83J/XppWBAqKJTNXOVoaU
IJJtyzE8I78NvbO8nOr8gCQ52hvVN8TayFvjSJvSIOwpE3jFJnfPFU1Ww/zftohHWzDZXYwHwcG9
2YBxJFZVgRhlhA9HMRiyTddpR2DYMHV9gZ2BzXJFpva1/dwIa+Q0lMmvbfBFE77wdNE97B6csks4
LFMnosCZyt3TVmT3/E4fdLWreYqPKuHuXZEWxJWVZDjg3X1T6pJM17bOTjK5riIw1jIj4TnHVO8+
iNn/YXNpZ2J/zhdsAgWioHgU5QTWf0BxHwWv4dV9OlYwlPKOE/fBsGSDsC4Cb14owXgqBbLcY+sb
p2JaJ+H9tWEv2r6Ft7SJlEeuOh72phU48LancI/ViOHpN/hFv3UR70u9ancUVkW9luIqtR9TxCEe
AS6uOwg0VqVh6d2so/Q6YOOHZ5pROrX0YTcUOaI5G1ZVaGicgZR2Q6G5CeFohQHG1zFC4W36MO8C
VY3PcZdj0Ng9E2e8XumiBz1xpC17ItsQim6f0Cg6hrHBVz/lOkG63CODJ8FTaDBn319wBntnuMwR
XqvQhOndXOGj+l81xW3kaCJcL5eRS7T5fc4RptnFVl1DUmEr1jxODcfFHtk+Nr5w7EcpJFK3hSJg
C2PCbOr3jpHLFi+QHHayTYYcANhxUVKifO5gTo/w6fzuFY840EURsiELEd1bF7Xl2MMUzHhO8zwh
CCKeV60GjLmZKIoJt/2xe5btT/wtAGv1rsc4MlyoZ0l1EMKTVBMPUp37IITpZymzYuagFGk2SEJC
wMAbsDo7aGFJyfZsiKkcBJJJIsPECFdoH0vZlp1qmeY1PmsE9SZ6ujoS7dGONo/bPGqN6NH8lmsO
WR5m2/RdvHkv9DB3Jl02evQkXrwfW7ggV2joBpveFBgE8J1StD8cbnl+gw5zmo7ZhVtN7KbUoqlK
Jew+lDTzGHvzXUxEoZtEcQb18t2ftFPQvyoTXZzaFaKpJKb5RTARL/BEYWL+Bd9kFZgwmkPD92ax
ir7ZxMLlyZ8gwQoEeyrbetL2GWQx1LkpvDUKkkHJXFWqaEh+de5dSMs4zI3XGj4aV93Paq6kEJMK
ouWBEChpuxsJwcZ40HpPxlfGGy7eSryFsHLg3XWNA/2RXeYqKw/zX40i/v51arv9uJ52uEKcaaKW
0arweR6veNgx5DdlCaQoLdqjs7gHZsiG40SrVdsK8/MaTouo4FclqaWUohiAWej+MxI9H1Dle7yc
gXS8/X9lYvaz/dovDBthopMB+RMr6znA4rd0wsX2wZChRb6Sybu577tqyQ6LEekdlNcoswB0F4JP
OpymeUF+Z54lEPQwbxzoKXHc4yLEtLmIFYkXf76xLMxfuIiGgJEMoHaH1JxNC0SWhIt7TjYZnV2d
aAN4xEu3x2zYwZtxmt2ceNRlgV6CEV4qstNJrtShLiq3IJRxFdSIw3PZMQdgL6jwILbPeiGoaawP
tUt8D1NXP0soDNoUu0JzP+PGU4B7QQ2bldxjNfvzGKlAkF2r2flwfcwYYydVjPTV3oETPmBaOuSh
g2E0Xe9CkcOqHZzBfP/CEDGBbTPIJGW8wLdXkODPk6IMUin+T6quD7I5BbotI+6x8BRnYPpI0nwl
9f9L5LGpzDu7PmQORBcIk8701WfbZmVUzhT6sqCdKfXwe5L8lvnSkvvzqd4ZLWkjoOtrP0rToJ2U
LRUU4TVn73LzbzLXpglKpRW6azfolMU2EitNZoR59Sdyo/kAXNGhkQ+1NMRRnkl3j8ay0ShCjUgI
/bO0/ScLX1itQTRdM9bM0iEtUW4DDErYNgMsx1ZahDpgiKVEjOa/5mG2EOlnd1v7uU5ZLtM5fch5
fgoX+fR6OE6cxS3WD5RzPMY7d3fIQQtnKtnozgeFhg3loraccGlqSwweL/4MIUW2XNoLGkUbaN9H
405EmV1hfmKzvR1eYMV9DSKkyIkinFnetuLsdkiU20OTWT+/tBl7I7X0cGd2kD6G5r4sVPfoz8Ip
YhxoHGi6lBUCTVfEEywwwraRD/PrDsmMhldrYQPIeW3CsF0el9FGuudAFiXYYF8NOLs61giUVdTw
Rq3Im65IeQsfL7/iK+ecl4TstzqySJAfns/HVUBlwMJZmaC3RLFsX9P3fwDMXwqzOZ+fL42kTty2
MOeIasvnDIpkB4KOG/bGTEDfbngYCh1Fy6c1Sq963FwWHfj4aWvVYH4HJc2DPpPpR6q6cTx9mMs0
bnaEVqjlnMELWjvwoaBo3s6ICersihpoVE7u0oLIcQOiiUydZQPtRWdjmkTRXXZyXr0+/iuiVE1E
zvuYsbBb4AqHog/GMD+VWBHh8InPGtxx6OJGq2gjHvN8FhkTLriCPCYxF4dFpu+BNinaaMYNKoM+
uUlMbSLSQlGkfG+5ShB+6mbSyG87F3I1mrG1fltUy1KbZgJSN9dFMPQVTyMmffYLvqn/CLDJK6GP
EAo4n2j0zFrsgo2IP0XcWJ/K1pnOq1bjUJo9ZSANfIPuvuGcs+BZyFbSo7p7ZhxOzBhroe4dRqId
I4saYbb5/eDjxFfvrA05uJqpdioiio5echo8i20afiuwGF/q8GtRBLZi+jaxRJznAb9x0iVwkI6q
H3lKpR6tCwapaDwMwvGwVnntkVGd7Z1bHdaPVLj4bAB5Gb831v0U+KJeHByb7VJf+KKb3MQesq7y
Ms8rw1pZlgQ40PQve4wMukjxLTTF8o9AN4dsN1t2iwxnhCrhk7clKK5UppU7OWQ+FwbMETsoxRAU
k+8fT0HDEjzUdWxFD1lvBgSMAQ1Os8ByyKDLiidPkmP1LmhDPzB7hYg6BSEQwb+ovZRmfuyiPQ27
eYAmpaXHUN+mI7LkKpg+DkqVxayjmqIujzrkqDRqBJ777gKi883PVJk5AghW+aGKpkNzZHxnSEGt
RSHcGgL7S5xbnJ3DfvuBNz+mTEuuzp0QF4+T2Dz5oWnB2o6Q614Su23damxIhnn5H3Ovf4UOVGwF
7yaXBlnTx8AAmsF5qebNHqgXN275qLIrptVutwkv/WkLak8bz/7hWJLZ82pLH8u/YpOe6q6Yl8kP
TBO+g4hBU75GOyCDZ9qYw2xlwOdbayV0HmNlnrbAKQ/R/TT3hZZ5OiZvNTjzql/YKHbz9YdNRbE2
QsH3k/+QbbdQrzCDUhR8d8OODnWNmAy8i7tGkC1aJUThukd1w822Tqs3CFSbzrYLuWSZP5GqI8x+
YUXgkUIwalTYdxSNIF5KpkMwGbVa5bdrRCu/fJQinkXO5mDs35R/Inv96ZxKIxGvp8Chy3XYx5yt
JrE7YdZHOeGxStjzuBb9H1PjyJB4Ro1++F8IcMAa5WA2aOg2ZIC43ej1rvwwaho8XtbLuczLrdaB
yEUkCUY7EGuXZ3wOToR2FGc/dPbF6rNw4NkEc8yf3QGlS/lVBd0nBchAwkHu3kE/yOCTFxwyjOKu
jMzNpwrUOgWamWAt+2gjex0U5TaJdDyDnVerRGeYGJNI6KZTgyA8kK4KqUvkMg2t6jCslOibBU5p
/5LPkdZHOXhQYeUuthryCQfXZ4H+KNqA5nxtxpvES87uaY3Ce/Y0p+zIJpwx4n4BiRqlPHbsKyuR
RudMZdPMSRz3nrhuw1nvAQq+Mxs7kLgHogZke5FysbBXu4loN3uXlvEyxK6BzvZDHiLzDetKK0vL
oo3KEyyCkbBFwWrrZDrTHqzgunlfnVJSN6ZBP/oioqF9B13k5J7n7TUQ/JF+PFHvH7GkV4XlS5ND
+n1dZgny410cLmVBjrISSGB6m2ToPwRozuDdXkWePIsaH/JArGN/BjsmDnof2nTJCY109h/5s/my
pMIToRJBeKPj1f437cQ0b/ratGMCGkpWjQFmRk2dKCuAVJjZgpcIrajSch8ZyTb72mtmyJ4A+nif
/DjuskUzP1r/NwBEmV6uCtAO+8bQy+eAq/LIGPapxD9FfE3ueb9F1OVJ3WxUomlA71G/J3B/5HRT
CC5kMJ0ew6JhbHAf5QpHtw9yzA2g1YVnv1BOzX32vIJBeRH5FVfWoJrqqqBCRpxwwp5BDzGwhBX0
f79rJWnAnDvjN/nxg9guR0hAtqhYCoRNaiq4+5vIRmSngYfJ0yDL0p4LLU1XPnYPz54OgH5Sr0wl
slmA5TRHdNPOH2f86i92IEHb1CkgFyLuKOH917kzoikdmezzMHDaki8wDqjJAdW3Jipd82hPluoO
nVs43mXt7apPudhBHKSSUoon/J7kLH86EZrLuNc5QBPKSFWJa9FrjhHw7BKFFzPa2PUr/+o+Uwgw
HX5oTsgF3m2fqkB4AGtFvGvVJp77pxSJsGdVQR1F0RmQabm6PmlGuTLvywknr+VMGH0Cscp3+F/d
EoCwlHhqGGNh13oMN45frr8im4lrkX5DUXqQnx+e3J4ljHBk+jE09Y8yEa2foD1zXD7i89oktdVz
HE8EKr7B9HfX+aY6kwut8o9xXOj5j3nGggRXpeyLHBSVjTjtMwC5hUn6g8zrsaWIDsByBWgqExf7
NWvbayIaWH4qR8Gqnlv9en8KYysLnRvESGbOJrGjAxewIcnPsL7YGAa1khi8IlL76XKqasl8s9D5
ms67CBzzDAhNF3mh9j9ehL2wRKsgBfX5isLV0tCojOaR0FlEVpIENvKOXawTeaW0uoX49CYcW14n
NplnErcq6oEvK5Ywybrq0Z3op3E51hbN24ZwVqq6YkhaOOMUAzKOR1rwszd4qYH8avTHQSeBuUY4
E+BNZDMvw3x0JLtTY17jGtd1X8vInMn5VnP53sc1EiAbZlavSW4v7A6YOxnAHUmVBct2HkLDU967
HiL3HIL0g3YuJ82x7BPiTln5PQnzKGs2k85NmSC2Z52pdN7KlvkHVd6me7tk/J6cCuty9HP84AGW
gYxhobO1P63teVsHQp6cN2EbIYvdko+4OP7g1JqAEZyqen6RNtV1CDnXkX7mvnkpxInBNNnMjgNB
JnJYzcUiMJiEyYMWYYlpCAmqpRubLkBrHiUUCyxCOuNxu6QV9kvMSflfCidH51hMBnU6yOTJteFU
hMPiUdAzjrsma3sLHAzV8PXHibn7L9rg4OW+XTwicjPXIkgG3r3walKdNEsuEUp3mzlp9NTg8PzG
kroNu5Fq3cXVBAFftaY9KeRcuris94Z1mfYy1Qbd33QgGSqRtx8kiUFKPFOIMWB/HTcow8kOQCBf
bmGBmvf/lhhYfQ7ZMM55fZ58F6tvISrfOuXWkP9YXgPhd16LnUpOWBofUjN/i6kh7D+b/hkkccid
yK9MuPbbjDoYDKlr9mRrS6XjvGcpZJtU6e2ZeD0RRO1MGDNTuL3SxaWchF6QwV7f0IdgHHj/Nxlo
N4VbGMdUBu8E2Kt85GPykYT9klAMZwtC3a9KMvuY/y0Gg324Dgs+hqgxOqErBcij/8BQetk9PTEK
xcg4qWyxZWVhjeXeIjvO08EXUJ20wAohqprRn1cHEIkFIxAFKzRplBMx3uImx+N/pwaai72v6VhP
4mFUGkR1wZUX4FyzhSD0QTDo9yU9ehEu3+WJwXEJWpWTehd3l2rHwM8h/QaoRSKIvCRGVXKKHFlr
lhLE/ckZwsP5IaN6SIJFM6y/U9w0msObLnzq61Yn9tm6Fve60xEg2M/RNhvyzimR2+pg83IqTdbp
TRM0TjJKoT/5bGkeHj1Q6rajX5MBJT1J1iKiY42+QO1L9VleP3Z1EwRgCYzsXtmLlV3ujlqDtpqo
hf7tDZMRwKVVyE9200kwym7aRmySuCyqpgbkTegnVdQLV8l3L/pBguyeN00WDVzsS1wSmTyMYgp2
HWPyY2AjxowTTOfRDZNdBVjOt4UG1p1Hy2ulMetwsgi1qbVX+y60PPwlXK40x5uznsNIO2qN421n
PKR8Ic4xMIzZi83DLOYR8Io1T06JT21zL2kLbMGmHKDcuW43CsAnP2+8Ra8SQjcaBy3mVhr5b3yr
rIHhimAo7D6q2VOMpqyPHWaELWCH2M/+nLAuVN3b+WSmGrgy/dghUiX8c1QTauCbZR84v9ew5Vrt
7nR4xu+AfSpuHB18Inz+R/Ej2+7CpVjBGUw7Q1Zl4DWbvMRawjeBSHQt1OvY/pRyem4sm6joLZ1d
slXvYs6LornXR9QnAmqmQh14gQDUHJ4JHm3VY3W75rzbVwa0skJYlTiGdkoy/aop61p+6dgyF16Q
Vwgr3XrX44N0IDvWcCEYmxW8HT9WcHB7zUrA7Xn/DJVgOaVNXlTUtvCUacHEvWjHJF9cJSWkd5UL
BbZDbnUxbhtBnhk+m/qEkf11GvEpsHs7gKA1bJIrI7qYr32Q5akuP+d8L84P4OHINV75TW67/j3q
2bxIyOT1fvhufLV8REnnvXr9BvrtG77w22dWpWc9940HhaqK13E1UWe2UDK7rp1wo40tJLWs4J0W
IvNV7RJ4v1akqQV2gUG5QwcKWjtdZn7/F0k6zV9GViH/xppDfNgnStjZq/JhvrNfmaP3VAcRx1HU
m+ghrW4ymMLJ/LKxDobya8M0Uj8LjJRE6goPURW9sFrsEpNjYHOeH9mVhklGzsOssvucBVlTY2xQ
uucBCfLyEc80Ekd/FItYdPDRX6BP4lkSQogn/o4FNBk862HBWyT9o/EO69+/chZ7/SXSnAsLwZ71
X/bBr3sH7oYxvXdmXX62eeHSiBDrniZHn09CPEqn/A4zq0snV+YvPgNmtUJ4wImyKRtLx9tVw7mn
HX12iCY7fj1c4bfht6Ms8DXtqlDBwO5YOwuONoO0keqLDZKejUL9OpMsHSKaMx9jWJ4ScQzu2X8A
abNccw875HJhT1uWjksu20rbcxeLGwBSosyDEBiws5+MyRe150PYRpQMYyb9vLKH+H0pgxUM/Tpi
26D7A8pNs5lCg6xiZH5B2Veei0/buwN3Yu1bYIXTg65yjS3m4Z+oHtg1uog3uON2d34tqeZd+7CC
MBE3pTky6X4DkdyOqsukGi1KnfBVOBcxg1aSt2giLL2k1tzJGnSpFRwJcGxCbDuWjeSzONt0gU5u
hESR1m+zQoW9V56clR9k+AdSFSI+tUQtjj/98xIhPCHUvewwxE3FXWlEbjIBNnBEryGapiF6fUAq
xV8D8NgKxxdZqlMngCs+G9QUNs2cmuJ52c/0YavdmFuVgO7KjqZ7wJyZ8SSPqv2g9KMwz5VEn5cb
blP0sUqza+fe3tYFN9DOsiK+0mjq2CbKcS258ewHkB9nKpVPyBd0+hgzvW2aMdOnh3mCi6nZp1sa
xkBsaWdyJnQ7LTuktYNJq9pPQHmdULdQYhV0kcWqlE7nCBfeJgQNyESCZimqbnY369qKGVtf+Q46
LnMNGf6mY0qJ4CWA5hgJeFrjM+mmg8WYl/8iugfcL8i4Cxy8Bz2tb35dmVwrHGCK7ko0oEhDjfuh
QeVtoIfdIxaU9fyJ492pMs8ykbGBwXv484xmfdS6p0491IsVhHbFQAusNJklrf2+Elg56Yr+GRBr
YTP8sJ6yzX2GfN53T4NHtSmhPfbsrzGDPXq/bpMvyInBXODTlO9V+M8E+rpfJ/oaiQBYXOUHTxEC
TLTFJvlFNdoE1K7u0mKSZwjpl+dbJdhI8ajMi+np1ElCSrD5iLD8VkImoNXKAJkeX7bEOk396yGV
gUUIwAl9dWa/rwRb/paCJlK7QgfYWSPU2NH8sAwwRlA8qs+ej1NPzcv3Fn0r27oVkwPp8uM+WEqt
p4rUj10bP9ZayjFwpFok6ZCKFMXuB71wjRkNhy4Cb2vn/fkjV7BMXw/xDSnXcUbk3hr63u6iY+pF
FpNLddZy45WzkJdUPnQBxJl/GWsEGUC2xpT7/9w20XbQC/fmjabOU2poFxJL+5yjq7SmPbF4t4kv
s2LLgqR/yH7W2B15iaL7MWeNXBewb+lDBDnfy3BMHPKr2QNRgqeg7tntjAxERVeP+FlDfEJ++wl9
4ysPY1+jYztv26ZbdPNWkL/hlLYd8TC9rPKy9lq/YEs/8VhOAmOjGAyCRbRs6LWPyQwkVcl1+QWB
FvYO+82fRjsdY9v08Gy5y9qM/1ObvuzF4atozSFLJxUZNolMNBj79+MyQ9WjAv5F6lzIcJ0mDiNo
o4GhubkQ5hjt4e87bd8eoAv27Ul5pBLTl3DqWeJh3h6Je/aPc7pzbfKDP+i6yhJLdPa2VZU7Q8FR
nMtFgg6ElBsvAvoUMkH9FCMf9azDPw20pn+FXfBvaoyz2WGq25NtoyVyfAy//MvagYWqsaPBZWxw
z+YFIICeUtqgI/GrPAUaw3uwOamivTSPhbDI9ji/51dqTvBao66p0/2c9o13WLbcbxvW/70BglAx
i4+NJ8Sk+hkfLO471BVO0zBaGFTJ+3uNT/JeWKAWSzjPJVeKRIV7vE2rO5dJpjPyFyb1AdVdXrJv
9HzC7k2HPRwwPBnTxg2uWLgZ/84+hi42C6XdsKGAAqrrVzj8HoDzbZTDTWkjm7+b18lbISeJg9jy
y6EEQH7vG+oFwkYHq+Fvxcz2Y/VjYxkXmFnaEzt+LZA7ZKUnDzQYWL/is7r+1gcjxA+6zP9o0+1u
uv/UhuqfmpMsC//MBGs+QFO1JK14RMvoq3vkNljWQ0FRlIiS74ByjmBQ2emtQsRfd92q/u+dgluk
35kZeCdKViG+iZeigDp2zmlBIAQneUQoDrfj4Sh8eNMMievZkukAEEg8bSIdNgRWZBMv+31vaqUr
fy/VUIPlMt7ncqxzJY3xGZzI/56L0aGYkwkidkIJevB6TznubmcKBB7pYaDZFD4HNvd4xCl/ov3f
pf8E+xkcz9hoP0IYHTzXIUmvT7VUNdPfcCT3kPkjrjzqHnAfIlLTnuDZ8nooN6ftqk5QKqqD4+AT
Hgfn3b8uoHPGI2NSl4ASVY/x3/r7Z8Dj5hzb25s67WwxyRnuAfPVSUubTwuxqx0Wrg5xa1M1rOqj
urJ3QywWkxM4SuFcuEbYYVPlE7fgJWPLaDsVkawj3uFW/XBUb8BMxFV7rMcHlDDuOYsn52x0JNxU
NAKQo1Dgip+7/RT5OMq0yWzdIgdE3byHOjDvScqYgMTMOarPdV4yq0bj8RAUmB/JcnkYKfXMdFSt
vq4ydVqZQjvlbYCwm5sptC9qHRBH9qq+YXl2EkZqqvLNkfhrKRaUUHWsfI+A6s26vYtebxhn75Wu
NHf/k32bTridIsGlTkC5ZwmV/oLV3k+I0N6+NCMzVQXVqWZRdyF1ZTWK0wbexBKQ9YTCYH+6Gp1Q
WkwNtvc13EsCdMusNSvQtqOHid82gcfqTxU2YVj4n0ZxK5bQQy+0HDcQvjSWZ/2mAAdYLzeQJCSE
v3cJu8yCOH5ky41T1VtQO4Z3eOgbQovzyueftKfmaxCZrW/lrqWBavFr8pi/UTcNdiovlkyG3/eq
Ko2TBMNwsr+VG52zause/kSe/4tK3n5NTty+gUJi990O0u4E7asVV2WdTcEy92HSzAsWbf8hH4Yi
6acRJqIt0QCx57u1/RDsjyxGJrEVSG7qeoAvYsXSLFAlqjps4DE5c2Fn2HDZvA1u/NRlwdlCJDWw
C7vbRKntrirYPyzUiR/y9vZx+62IOOzkaZOFU9ZP6GEDMYDYovBQgzsroiyFGKREBrXvXvfnoSdS
TEw15eryS8zarKDuQFA6VnuLuwONLsmPyJNo59U8VTZ0+FvnNXLYtnmfFRd8edU9CiviS88nghUW
92BLFOPVdiEvFqEpUSYBAcmIfpMRWs4B2f5J/zLdER+7fldaFyr3wKDXfhgRNU/NU4TUOI/SA6jL
TMFYWIsE7kpkbRO+nH1PzwErwqn8Z/Y9Pq8MQy3W80de9UsaUidBCBHc+a7kBilYoYTyWkdvW3zS
cb4zHOqXNBsC6ivrcNufsAf4Kyfj4nIqbpn3Piu68rYuyHnInmu/8FXbTh3A3w9h7LQDbJ5JQkAj
c8Vdx0IfPr9OwvnaKEOnmTPtz6zcyUWTe6RT9DtcI4zVoBQDLVy16sGS923INtXU/BjVaVwT93qt
wWwFs11YiuIAbG68PaVNA3UxQqER/q1MnLys/zDx4lX9ZAsPcdm8k1utXRp+QsRQ1cwwEKWIGDg4
1MGEZzQI6TZljIT5O1pEIvJEinzHPmg7EsYMWk09X3wGCeMvS8IN8MQG3diz/pFdEB19cwvmFhJB
Bc68Damz4yUHMVQKVKtIUsd+F1FHBkYziWRUtbSR4Whutm+tIgr3gPZ1/p7WP0pUjZmOx0rwnh+c
cXSQoCOCOfPTWy8ILXBDnIZ0uXcw9CTFo9D7Zd3EIFN9BTKaVt4PVgByK1Hf2GXKD9I9Uiw3L91u
ZuQCNQDDHQRuj0EqMvXFiawtgGOz++cIwyPqfx2Sq8RUbGOfdVTGKZpxuyxZhyWNUtPSWz7TWZL7
+TwNAzxQT7FTjd8fke1rPM62SqwkHrhDrg3ojz3sISbVx3pCufEPRhARbs0rDYC/7YABCF83VcJS
mzHo5Whub/ri4ppYfWITONFjXUUIu0cGekzoscryUzERGn8CHoZwFgWP09JJsUK3dALMI5sxqvy+
Xa/2X/pY/sGAGNB/3jh2aTKuGEz0tBfsL9titGe8FMNV5lSZF/I8ToQ8ZomhIxO0J4hBkDeiviYl
zXPkuY81twbiBmdAm1Nf5giiV6bAqtNVX3AirOj0pKGwNXwnwOlky2c8mQDfemOewrgNGSTG5/nR
KQOaQLGG0gGSoYYjcxmVSHrchtpDEUjLt/z/Psvnm75O8WasfunIGGvXlcfbyl2h44BrNByejtPy
4oo7hRUeVyLZf5OVV5fIenBUlXhcJmAgAJEXmogirMRrnlEzPmgk3ByzAfHA0FqxPM0K+UfrDKja
FZfr+4h7eT6Oi2OFkZ5E3Z3jgNqyE0lz6+BdUBnixCrvtsMs0iJmGpXp3LLlKBLpUVCVR6AtTLYt
aEYGrb+M0/mTWyQqdGvw4xZAF0Pt0jv1cZIEpYLYBkp8VSULBt5khPInahxtiZXv86XlvyB4+hX7
BxMLbI/HXNKH2qUWVoyJtG5PpZPJbpyrSJnUIggQmV+BTSlKyOKtByXvIZa6wm8S2UBdXWDfI7jX
Mv72CY44Mws4/NyWznE4DDD8pwH7TGgUUWr19jaErH6YsyC6486cZ/9tnfCDP+H+8HjUKY/ljmrV
cWTLu/2fiUVIeXtdgfqpn2lhpSfPOOtyQah/UEN20Vuoytqqe6nn/FKouobHeIYV8MYL/7n9lmhD
2QZ5nW7A6qknhIFVfMSLBRYsqnjTdV9ikKKa9+Z8FJhlzyo/K1EQYS8u0Xx5xlNunt92DZpSdw03
NvdfzN+e0kme1u7VohtGZXi5WggEP6vKF0gVq5Q03GQ0/XU7p3/alDUQ+zFexhL31jJKgEBmJIwB
rXF4qAtKkDxdbLAQFjY8bwfRfIhs5u/zSG2rJ0jvaUy3e5Eca6slTjaGHEa4foLWZ0mPYbH0s3GY
hxOu14BVlzzpMZFkNvJC6dQ9lFE+BoK52ep/GnSiBf3C53i7oDJ6cJefx2W0C+4nte+anUq+sGWg
VYnhuohL84Tt9DKA4Ap3YzVdn54T3tx40P9Q7tvqQGFYSVv6KTwHhm35RsyliKx/iGk8s+N0Zmoo
oNBLyMxkDcvgvgWDd/Ytc9wylIXI3fe1bSHvIJJM7VWroBTmsk+0nroHrgfkYC2UfGUMG74LOxwx
RTqBl612jvoPQkExT9ryd41T8/tUnxeDmYWkUGAv9IfdacB5AdIZIGV+/6DLi2pneAMVRSvQF73Z
X6DiHy6sNc6u2s9TuTDApqWDfc0qIrohIbN2nUPtnC0+0annIHFswffasTgg6gmbEL1wb5fBxe10
TVbRDOMp1d3qTjoxyf7UC6WOPn5UPSJ/sq4ttNv6miF581U5QSXb9DsNylytZywQn6fK78Nwx7Ew
iYl21yKHJCt4buIikU6Z0kz0tY9B34E1YNhrowklFslq8A0eMrv2m4hf8DQ+900A1C5+3oM9/c2i
Qd0SqCBzNCUJ1fT/yDSc7EYrMYJ0SsUOrx5ypCcvE1oIzuH7pdXCspQAH+peSQFTe8Ztsq4FmkAu
A/JfJXfo471OVwETgDbmnRf0K6jrJEypDEOsc/5jTQtPxL0Gp4ae38ssgdmQ9cdjed2q7SF4/D57
5RryCqknz/qTsGJI4RxC32zbciCI7WWeHZU61eOIae7UvL25reRkmzrlQjX1iXcRtp0VnSh+/V5M
lt3GTkN6Oa25eOB4kl5ifXyqtsnRCSd30717so4VvNe8sK1NNShVWiR0aczSiuonHB2+svlf0PXC
j0ueVkmNrv2+FuhGyxzjaNfcy0+GDNtR+LRid+AWCPOCLAq3+sCJpgCoUiSZQ5ijUJvnoPBiIlI4
3wFW4p0nj38EAChsGYIsna+Vj3aCv5fkJndpJoAiTkSVD0gNgHH+DqQYEMa/RxrxF0uYG5HEElE3
3b4H7B88OTK1tOpad8O6zbCDxL2TYKvWQcbUHdsogDBOIK9gOAWJdfyljhC1dy8cOJapWbpeOMvp
MEzYF34dw5o652vmtYfMSa27oAiH1bKXph9xW6a0K9wTtXKiP+epVbFLeEc3fxsuA0CwY25v+rpl
cf7WDYYTlCNeW24CrvDhMnYhdggz2g+nP7eBuFqZjZEqg4dW0uS6rdCpRSl8qN/zzbZzdl6+VAg9
yHgmR7l0Rx+NGMlL02Q6Eu5DYGwIxwMJZiaQ3QYI0nqNGzN9lF9WCDHiMXVxQDAxK7WNTWPErwpW
Vdrr8BwbGMhs3fCp7i3deIs84n/i83+zOWOy3/xwDOKaiz9KfCydTKsyzMJWBr2fSmGovqzQPwr4
waAQzb4kGm8zV37Ib0iO48C1VN3V0X3Dw/mXpj9tP1TTBVlu0rX4vCtr6Tx6NMTzCkjvMX05PiRH
19I/9VBrFhtjE5QyFIBecl5yoTtVbsXaBDp+p2cCF3SRSdv/Yqzx4BPmGIfiIw90xvx7ENlXzCLE
jYwMMeiVDTJ41SGfhH73aYxWMnJANqBLSd2YH0ZE+ukY2D+lRIgGHpXgQfVEL/XPDDFpQDRWpsUm
yrmquY0sLqAE54Q2OmZ1lZkSKRSNFpTvNF4K99nTCPH4IMCgqQvxqb2h11Um4CCmXBmmV94EI0Vr
yb8Ups1LOigoOnttdeUvhSxPLhI/p0YhEghhqEImEi4VUxqZ9TrNcUungKGT2u8OtuVSGdTqjpmU
oILGqnIovv51wCRMzF72DwDte0I4jAgBAiNAE+N4VS0Kzl2l7PIo6eWvfhOBy69OcFyoAEcu9zas
xV/cocqUQoL7UiKfzzH+DvZY5zRdDECaAkhr2DvdUzrc1wAqoOxDNmSp/IDwQVPtIwqKmRkOZUs3
AG9HaRJDCVdlJyFIXCySMJ331ydEw3AdOQ+Z7an1iUD+k5kBx/DVH/see2tgeJuq7mnUnfLYbMRQ
CKJIKgio4Cvf/p0DvqlW07fDV2HNxcsuGOr78ctvkU+q1L4SRIV/7MlWZA3fTDJ+vT3B98V9Ouv6
ZXA1+DCNrv3Vg5qPR946tkE3gGZE0iBwPXWf9E7pxmy2EkqHp1aPxU+lJPhaLur8hzp/IRPvKYld
lIkbBQoMcJ5IngTsa8l2M64JzRI5F1w7gfoAvpUedJm+tUFjlKmpZxPoDrMmzi5ovAMJu90UtO4j
S9wxEjMj20yNP5wbcnoCHCcnCANaSOZsBySgXxdxalf+H2FTVsjBwo/2kfXWLfNsLTL+YCaowgB9
fbtruu2fQtRi3yNKDRtYj6eOA6Jk0TDeEwazT4PrGRL24mFsV9xzFt4yG47ZSSxgmwtQ8p0CFx80
Po+lWX76HdB5vGOF9FCqFzMpBxjvnFbD4whpy1fzgoNU33P4973xTRnUZ6x6oDTVjpT07H7EnpaD
NrTWEzp4EUQbpsscgd7nzhn/uL7D/4kOEAd3D64dhgKpxoF9aipaJDTVaA4jo3McuUgfY2JmcQuB
/LfeQ4fNLaV1F4iW7Szdw7PxwQYcMeYI3rPTUFZvo4h1Xc0IwLAca6jyeSF/14U2v2/yesQD457J
XYcGLqYf3EoOx1BADx6QQdGTYYdrYrj+JpP6j1xN+u8CCOwTbFTT+RZ6zOIn5TEkKV/oo4XhkUgd
Dft6/xSgg/dda/zJOplgRIxKJE7ATOMd4tdynZirLZVXdPfdEcfK/CI2gbP8cQi5MJWbGk5aMqQ2
ug6GPeb0CdkYbPuMvpkbZAFECuFYN/eJKUTUjpOJhrPR4qD+bKjL4KhtEAvqcLXWywnxVxTf6vYK
IhrX5QkskVRLUyyKWOtUgC7f6M9nR2Z5LnDgdbPaoUsiSQMGooNWQh42K/4k5HBRciv7seXGoi0h
lSBTp3l+QpSRYc0bBkv0M5u82F3YxV6rat+5JU258gU3CaqsFZqKJWr6LF71BfeF+FI3U7Yk4/P4
Kz8o81Y3Fg/wEIZH92tap/rx/jX0h7FnmzIJeIRMYWgh47GKj4tBSmdhsok6j0rIludQCTsOAFmS
YTVzzCHLD9qFhiP6wjtFcrz0Pnj6fihF0CME9MvExJIRUcmyL6QOV5jp5sGKEhulYljmfNmUSRHB
82YRKqPzycoyALG4l+tiBUJglpBUuzYtamVJ24jvwePcRyL/d/dqDMDyeMSZKvUpuNWOnqCfkFlW
A6F3RShGpjTcf7/OV45VPVFAJiK4pPmV5DociA0GnD3uzAbVQnED99B1xhiCxWglw/JnxoD2q6QF
8E3qGba6vguPEIbQuo734l/qB+cr9rZMC0wnv7vOe0EjRbHm0cOD1VBZks/uj4JbiN/V8lJr2fKh
IUbkYztPdxD5c7FtZ0+Jk+P3wE8kAr+xnxiysSf/ha8aW9za6STBZACdfy96RvwLS0zDpwb6fQHY
rYfI37g1iIIJigkZlE/hKVGMoU7/eVmXoa5FOji9yd0PIzDFsOuDWUglFNFyT7D5SEWhfqsX9xN3
mcmX1+ouc+AC7fX8UOjWoxVADIO3k1f3R4C+9N1FPT4c0g3c329GKUvSwgjpEse1FtHYcpDPVJg+
59MbvIZBLosyFyy3tHzcCGmwXE1WFqlVes4XtvC8YrOGCSnlkLzBKVWFtT2f0VpLxR9l9L1Yu+sD
39sWRcwLJg4WR0UlO13vOZMG2tH/fWhiey62YwJCwDQ332XV9CCrlv6qKnxYvWNfU+hR1R61DCrc
skUpe0nWU6j/cmk3ngSwZEzKehUQSEBbc1ejYXF+jjv9ecdfrd0RXZGQRwtlzS+7pUey8v0zDLGA
c03qSlykES9G4ndZ81J667gHBCLFsQ6so+garPqmD1tseox2CnbIMqbgheyzlEQejrPNBEnUx8xr
Rwsd3jpwM9bu2yDibLF+UcyfzYABu73Iz3AusmoXdHT+MTjEMw3EShcBlj+dmM9Ke5LlYkQe7GNf
Ht2K/T2Of4IAheqAbIi1P3/yz763aIFBHeBmcOoyhSZwngEFLyVMNZc1h2GHlgCbdW+3G3hpnN8f
2cDDEWICoocJySy7q0GnaUvwGg0od9uf3I5MsRNwr5/DEoMQnWHmBfHMzWnXgW53jaCE5pGUyNYW
VI/9heBLu//sJClB0xYbHv0XfBEzZzCzsBBap5NTPtZ2MERSk0Oi6ZM2CHoszKwc7Qvf1WX8vekX
179B9ukoJVVG0CpJgR/KQNEmMRyHmr4me/eSBADrxiRQczsn0Grs1mE8hyXwHCd77vUarUYvone0
rPOrDkN8cevtMWm08Uf95iXNYDCfvwBeJI09pRTgQS/ZoILEcab+pEmkKUsLeOQvcFHS735QNeaM
iVdUcqMUWApAfQf9DU4X4Im6CszzmL+2+6UQ0wDQf3OvWiLxvGvBBy8SlQAmCONAKPFJH03gAvNY
IQxDjO3SA26PCYk9eJIFS5zuheAe8IWjgnz+A585sjqO6oy8E50YecYooZilYLo+SC3y5ECi5b5O
/LUqyUrUxG1Spx+BrF2GQSoV7TJFr6J/pvvHaAFEcnssg6s/ZkpP8o613n1cO+iBtEl5IOJFdAez
s65vJrCKPeCFIIawluDYSMzhckdTtTFkoHupzhH3Rr6TCKcSHxZtUZdIAfAILzqvW0kZwEnGSbyT
LheDnUAvucRaLeiL5BHqL7WXiS0FPYDNDmiwnJMVe6vpIcW2owcZR4dXNUkwdHHFeUetLkpN3Rbo
b/ATLnmuYk3Gfp10BDxNyGnKRKppNJMDaaLUuskZaRuF6R9XaomGDPRqT02SxHaQKxVV/kJLQHGV
ZXA9OWlO6V1O1fWGD7fNQzFzTkRC+f+E5AC88xh9R/DHHOw3CIFfcnJ+YEe+3gy3/Koac7/IEkNw
aieNUbZ6Ki7z2aBBUbniN9kQ08d5ejojf3rzBJ8oAbh4mVNpTfEebvJCEeRGq/6IKQhWDduEGrxs
BzFDLpb6M8vZ7El+DHtIYdD19CxcA0D2hYXjf0U0HumTeAQ0/FadKfnGg2EgxLc2iDwSKJZl8fva
2BYIR8pVy257BwNKlV4kUALG270cYHeQM/pL7a3fRLxqErHCF1XFQBDNcNw5e93tgdmEsG6HJ/Rr
wNkr+InnG2pHWB+FRUxw4JKT6/YlVMLBgTmMfPVEkc1m6slpCosSQsr2R6Lvhcoud0WvvQVJ6wzJ
RogSfjHii9XQv+IflSLN+MPPnV41sMX0PLKjh1ANcZ+FQ3dnEHM36RNg5Dvz0XLTmB1mTPzZf5OH
nYTzKHC3nY7pJgD1TCKH52VHp6eewESNqsuqtZf1Ap4Z8031s8yXd5PqK7976Wd53kXKIVanIQK3
YUAOZYho2cH9HfzZ47h+wom81sPwY2O+PRxY5ERwppoW0u+mEROd5Y3wWcLZO3CRm3YRZPYIElQl
EmZM3ubqp76+kkEkv1w1qe2HhoFc9WCq6ZFjGoVYAdgilK9QlxhUGH9YsBhQZRlXd8NyPpnKdyiE
7fnHOYj+FEz/s/qzpNVknJ4L2c9znWW966/4u6TIc03FxKfaVY77lb6NkIYxeLA7XhvaI5kHbwnP
z1Wvi32DIdVDWLXFLMjSQ4iCKoayRExMoBCwUstRhgtO+ZaxLXU33tt5tjKVLRWSMj9sdjoXFkuU
Mcw0b29dOzsBlqdVd7iS1Dmgz0mVPF3LMjGFY0bnOyuunYBfTjiE9FQMqHKMChxzi7CJDHjsfLdo
5MNnCByN1326uBQ4FQvxpkKmoZoAMYn42S++zuNIZmWY+019YiGf+N/QEpoFlnPebi+QEdb1PpTp
3FOK0zC8jYsJ9Q8gcVcXJ0TGC4LoT8E7XFy1w/ZeA6peLl2iECxpTtTv0cQLMxobMyDMT5FPh+L0
Gq4ouraSiZ9gYZk1Cmb3d7MfGho3M+byOQ7G6kpB/mcQXz7CrPxixmAAo/H5DER/SKwYAAp4SvBz
eUehHQy5bj/ccsGxz8awGZdVOuX2W5CR3Zh1BBLDZ+BTAfmrwHSKNMZyk02bZLxWzRrGLdjd36n3
c7r91b3/PvPAPwJ7XxQdfyg7HBqKPuMgSMELP8IWO4APNrN5X5lfwrT1MQ6h3bawHbqFogpl/oVC
vOKxy2vquFKXJ85gBR94lluMK3glr+TgR2t1bKrGM/4Lf1ukQVgJ2HNPjbG/qGkWLZK25R1/lDe3
dLkHJkapWJ42bV1rC49Mbd6K5pTEtGRpZ1iugHXCmp7kKaR0kpcdQExCjPjuCKGpUy99FwAnfIkW
5rnmhBRS1a8+zpckUoHUkt+WgPeK1c9uULXwsH5EzjnpxvPyZhpnPmypHCDgvLDT3uR3u5RncEvr
5eCgbrFIqu001UNqdMLw0vX5i0oymvcDVyh/NdxASPWWQOOhhn4chZLVY8E/uH7dbhthNGWBuCVm
XKSIJNoBt3qv39nrbf3ZINh1A+gDG2GVUrYbS8026FH0FerKRKEcISiZGgGDkeqVzsyWnAwGxeo+
j5wCHfJdqdMvj43sjA9RI65Y/oZPs3rlUOuznvypAKMhJNrI8fNJKy0GRORHVFgS1G4zY5UDCEP6
S/8t3ela+ULr9AJEAFzdXcKYqh4jeNSOrqrwSrifvgcYQZIVvapgVcwhT4BmgKOSd4iYRWJK9TaJ
jpNlgMILaukyyPscStTn8KFEaczZp9FWcwusyi8Be7SouKhHJWEByW5c86UoCAi/hgWijQ/wzRkL
MuNcRWEcelQBsuW218N6gS/sCvOOFCZXzF1jjxjRnYrQzlmqP1Qjmip75AOGCVWqFHYY/DcAeC4F
u4IuL8y/sYKvW8vmNgcUpCFbvQP28kvo8SiB1xBRFqKeDcvpV2ja+RRJ3kVhXEFjNA3ASy4JL8TY
23enNyKI8TX9NfNWbyy3jRS4Vv7RDIho5cKjRvFPmYb3yYcQDEytsGaaVoKcAK6znnNP6cZ7DFXU
0cxOMEMMh5lAWKbMottqxeLa6MttrhXtJXqQ64hmfOKX5vXFxMG6RHcgUofyA00wLLnu8nCsxwvR
xBg/jtnq7dleMJIlqLrVb1mRtb5uvLbm2bC29HXh8T7CVNOzYqzQKOwpqUu8IdXNLpBDuynhDArX
unBaU3tf/6GXc0il3nlEWHMdWPTQOOPKEqpwmOfPs2TRYMFUjVdo/sLfY4NDZlhpw0g3fIY/VncW
lufzXNucDafHr4yf/Ehm6PhNuU4pPfkuzBhHdpo5bYXaJkJKkN5/GDNuz9b46MJlKKoQYyOlshni
qwlH/xHhCKJNyqFLvis6ZlQFDJC+zu/1qRxF2wWtI1ZMFQBBvWSnMpkkMPLfC1RSZyZH2quc8V7o
7IX6yWjs//CV54meSGqw10VktdMU0qw9E138wpF9rdAgMGkHPs12RNcwiSjLyUJU4sOhiTUOpqfo
GAfgwGuZafoDfTmgNQ+8Wc1CzAS24CPuD1qkakbh9+JlpNrNR0mwfNOkxXS7sTwUCZq9rTQ9mJbk
iEpi9yjO8tI71zkQ1BAOVpjNsDmx3qoE64Js0MfARw2XKE1DjsJOEgwulxHlibk6wSxEInj7bj6i
xnAcc9o6+gaxJUzQUFh6MKTah3jGTaSpmSjysvQVUMFE5u/TuqG23nakQRzu941DtezGkTFtZVhT
ICc28mFk4NHxn5Hm7EOjbd05SIuVX6BFFn5jVqctRlIiP1rOIcPfOMQQ2B50RSgP9F3JKvHPn4kI
xbFZ3LuJN+4CdA1hTehtuwIfBxRZv+wtJd7QXcM0dX/n6PcaZz8KoQdKqBU8TSJFI/StpSm83wQM
2A5kWkGFVu+2NHMQ7lxLczf8HZVuQP80kuO9PWTaBLtITUZPbg9pO2uUyxkKqY4sP6Xp3PtQya57
OFcNvJ2Fj/N4/z52HC4GBODwNWRlrSzt5L3bn5/ivowVK8bopqIOStver7n27v0XsR3V9XNKbgj1
kyVAu+T+Zpxk/JKwf7BVegqj3MUdSn3veDbuBf22Z3/uxUSaYCiWYgik0v6OPuzJ3+c4f4eUm6r2
45F7DfcHin8xH/zOX7utGRB00HHa6KPUu5I7KDC2orKBwpVRXEjOIR+Tct8rDAdFNOArZerJ9P+N
JuAWgszGl5/LfLOnDV1EZasUYlyeoPU0e835NeEbOFlYBnyz5GVkoOdtSldrArO5fLcxNKSwiZw9
/5qqj7LJLSuOFZD8dCmmVrNuetsV9aqLj6fTCiFCTyERg9sEk9nOgC/b7x/i/3fJiqgwfW0yTtCk
8CXRLvOInd3ZqCPvf3yy7meJETi7zUeEmBSsl+Te5kkESuJUQv28JvQG4usi5nSQFGkkZycx0j13
CsSd5KhDoFgfjnZiInGexoUwa3RiHarGnqT+kVGjWCGCBT9W8lqpvv5D5+SiH1s3b1Jdnq9s6t4U
V7ms7orDRvNjvNbliWQAsRjQx71mUdeA/26xbQKRdAMvuR2x8kgeeVA/8Hxl5j9GijWPPycOxWAO
cD+psbxoC1IGWFhsZbzgwO1nx96WA11Sp5OB4p6EFA9QSeA09jwApzgawfUXTS+KK8JKS9ObEcrR
v+/FzFrrP7o8dGX9OJQJX9bPofaYv7z3TkMBXED2Qmbwo9mKNJrpfOI9ro7TTl1IR4gyKcyDUfeJ
zBnfv7xOl7/RXCH1475NYR95cuvwPyX8UdpufjvrdRJ5Lk+iFG8yKEvs1LvEO5bOLJN18qnC7AIP
OYFziWQGAv50H6Dz1eOJ3debm6l+9a4Gd2ysyeyLFqYvOOtiL39XL+NHTlc+1S4zgGATzEsmPzjw
casQSggNeaTpQmcY9FeCcjsEQd5x3hLpm28SNUaRVqMxAXweoQcGo2mXt6+FwciEc1Tl9/ydHvEB
nHSWMhfA5SDRvirNcU9WwS0s/soJoEeLfFufMPkDNx7Zney0QUBgvhXK2O/elfbnJFauASwFy23y
XTiIvL1wCx5ycmWF8uFlklRn0Uibto/X4KEUyZK4uHFtmHG2af3gcg6vqHo+P455fIeQlA3a/wmL
D7uACVJZAZMCprNhzUP16dZaaB+6uhb8HcvgZOXnZhaCSbxAfoc3X8M0lcBPKrL3SBW+XC/8ZSmS
4Lbd87Tm1FRaJsZbdnS01DrtrHVtRleaV4ZqND4rOJZberJgWn+dPCJl/V+9GxJIhzwHLNPk1YEa
/iU0EwaY+dYVvIQ9MJvth0PvToFdypkKbkqdBQ+0eMRzGZKOYf0Hzy8O5M+a1ptPYW6FbdzynVF3
F/Nj3jKuj0ZmuJ4dwPIQY1+SmowbJwlf46d+vgkdqkEZrFCVWEyyioo3dCFHV7w/uPQwc5a/es5n
9UWdK7B4Scwp04c784SLmizvrJc7IItBiHtHybIsRrwk7IWFFrczV7ygJHd9BFU17uRexV/htfh9
tjYTABb/ncBa54z181tG3XmPk4clOVQbF9nNlD5Ey01r6Acd9rv9iQTyA6i1bmw42tWEQ5T3qXC4
KcuyoovlzDsGW3m2MPfhJSe+dZDuCotgU35/0bw1xlaU/Zk8zGKlUxuqIkMEg55QO8gQ/fuCD8R3
zJv1vV1AtBV00R+fQi47UUBb0+0GQ8f8vYuTfUauQGe3MYwjGm13lZmQSBMMsMxelDFAntVaPVOJ
RJIALvy6i7648Y77sW51/X6+5AOQ5XnR/2NvlZZj17me8s8xe1IX4tnf2RJ0FwvFxxUAlBmmVqI5
aeQ/OYtQD9RABlmQR2jnpzHaCJfXn3lx58QfjEsSqrZx7cMf6iXcA5UzdMXqOtoTWv3ywyNqLgbe
JVYKrNKOpGTw44w/S/45xbF+5NMw1VzjxdOsLcrnDfQMVRakST360mDzhv4/kQwMx0MkDtuGBmQ0
r70Y/09LxN4rNAzGQgStTbhq1lPGZ9E/mxRiQZQfU8F87wIaO+7nlgyea5LmQw3jcRGRC2qxh1pb
tQMONbB/G2hWIqYnqZaWF+VXAHGf/j+QSUGkgTiqpwUCDwBsBmE4Wyg2v9EOIlr7Bdkqvj9CxMLc
F0mybQi2vyCjwtJsuL3yo2YWeIhMsK+CsqjZ/ZGt++GdJowS1QE+TVpd+URFJA8saQAScAAleT5U
qmbpYBu7et5cNHikn4Yl2DDJkHgo6FJ6zRvng4YmfOWSwdiDXK/tiCqRHwClXcR3o6y+huk5Afr7
0Dh91nlxfbq8m93O5NW70SY2xxXpSjC0xdvQ6EqSQdAm9jR9VOI7TPjdB6zN8yJxvLTJAyAt9u+p
Zq92vlutryFFD79woS0jgBpDCCsxqPEEWaNeFWCPqEQm+4T2/Q696Rly7NVxJjgofILQTxRu+0BL
oaAoMriLKQ276rIysmFbyC/55WWSJ91Ej5fVj06CJXhGaIalcfN210OWqPcB1f81KVD/nY5CKld5
MC/OhaeAsOFIEpyGc0Kztcm8p4RdRGp8OEB7YHrUchX9Gr+fGj/yFEJ1Mi+7GS1RNiL8MjpzV5Px
OuUVUk2nFgZWyrqWYyKnFTnOAajCXABa4Uz55Ax4SuMLREQLkNW8vaFw8hIYjRJjHN/O5eM2vz7d
Y8FrfNCmQQ4qcp0lUtIB+UdgJKOuPN3p4mIq/ZdeLcOg6lO9s5oTicIocMbJV8fUAdrmNXuyRjiZ
B5eXn1j/cV4+T2V0g0mP28f+kQTu5AJKAn4jcPnIK0gvSWc5uL4LyMsN8CMqH/jeKhzU9eRQa8J4
UhOpM8p/hjQHCsFNn/k4GmIWO7O4WH2FXTO5BtqVWYOIL2wPhqdfgiJRxZm0kr67Xj788uYisdMK
HX/Xdd597KcEtFlqHFOAnWin4bDlBpcn14G81DNXHZAqunmAwbKtg14wF5/kqdQzvV6mrTOQgoEY
u3UqPve4JsyE4ZkVVliZ0qIc8ozXYWP8ov4CFvAruzo+SPypIkdn8wh/7DMFLeFlRaQKm29xCwqT
SgMP1UB5Jk6qTxn3kUQ/0ZIfrXP3OZIKrbtPh0kUrVIvQGFI6i/7/O4P0Fbtf6wUJJ1rwu3CD89h
KwPdRkOARpfziwyFhezLCJ5uutwX6So5lTl+wUSDg6VHrZkedE6w0b1jrn0BDrO6NS24ZdiZFQjX
31nzRplUuAFTDE9kJMDcDmyB4VWHLH7QMn904zgpkOxnQhzTf3JWJAPzWXmI7z1Wh6Xu1pP7RIyA
jQBVW3CDr4evAFYKKBrCxM+04rC6NA7zKBfhGy1n6ZziBh5NauXirHpigBB+ZzQy0DqREqHfcI7w
+JjHgBskSy7hq8yWophRj5O6PP7ezVBkA3PtVisvDR6nlVSNAuTC76YY/+ozhf3+Bwzy0B+7NmtR
MSSgpXn7qGagVA83uVcddJA9EIGtb0CH9icHn82hkxB0yPYLOjucC7SprTh04FviQpmCi8Yc+c8E
c16Pij6PEiKoFXjZaEAXtf5+NCW6NJJoInt8Auk2yKYhQMlDI3bS/p7X+qgb/qHCKrYB0FfkwJJ4
pB96zr87luqnCb1uJ47wgReQ03kiIh7W5AgAzkzZcCTo8uZnkYl2TQj9OcYbttS6BNNWfcGOuYRK
WyfZOeEmpKRAhTthUxTczEe5U6oKFdrUWBhb0vXWwxf2pYXAE2SUGrjDGBSmmvkUyl3mZwKqD8Hm
KQrdc2qICo/MjdbfY18Jj7W1/M+IHSDp4NSF90yXBm1PPOrwIN/gO7PnzDpZD7XoZehZy8DA5HpE
Cr/agBkHMtIFXx6hny168WuWqPHD06l2yzQJCOy0gfCeh8Tw0RzzxGudWiU3B1ZKn13faK6K4rSo
4+ccXMNdP6YztjcEuOsOB2aW8Ahs502ZfkkBrFk753s6uCveyZrIZG+sNuLdH7oGbiiNC+RvqiPN
CU15v78zXqC9ah9R41/kBP+1fQhzEcbmwQFp92QgX8xUgS98ZvKGyOuCfoFNWzKb9MLKQNh5TNcK
Ww3Qte4uQ6fWGsEc7HtyypfzBlnZgD1jdhPdvfZ5NmtINoUhJJpYWpmfap9TnFw1pPaXn2HbJ8R/
QwnYsMuqKM8qyc/7u83OIgcA/yiDLEj9ynrj24AqH/aQZJNSAftBck67rkkJcWiw5t8wA32Cipcg
egCsacf1z0EFvlLbKB3mrkdE7AFaaidaRXuL+qggAo+hx230HR3wVvMT4b6Han1JcQxiw9+wiRey
OLZF99UvpORVStjYB7qee557OO/waaiomve9ZYOf4EvAqDbPUFeo522xLOktAJyTN/29qfLm25c3
MxqzCzwuuf1QrBA486/5axkgXReUcaMJybdzbW/DH25QbkMPyBT1Kih1j7/lZdGjOSL+5BoKkR9n
kVP1+Htsnko8pwzm+Bilnl2fAVc1ZXpgqYDEKaaSxcPY1eqo/X3PyNb0WW4+25RGhGZ/bIFl6XBM
N61BSb6n5V4mgqtdVbM7OqUnp8bsDTqhz6AoHm0xdI8sbVZpMHlNyJk95JkSmJx0lwVFtizp9fFa
nzA1F/HvoLbs0+fE9TnUL/D4xxgWiuZnrOy3nIdExQaFXdprt+TpyJnEaahWP1rJYfnYyjKw05Cd
8/WNPwHYa4C5B2evbyLqHXVfdO0kijXZrCWw9IWYexECDLrmCuzCSTqTuwda6VoiLUF5LiUlhguG
6aYIVmGt1R8HDPJlifnO8AEdLyASxNs0f+ahwFUG5JyDEa3Pr9yOiEcfFWLN/R6BDiXGjZaUwf7D
CQVkZPQuVuBuFY8VRqHNxzwDyBGzp1ghVb/ldzSKlgQSAwlvVN0RERFicsptsVCr/r6ukhCnp0iR
03Wd3MUyMt1ZoUktok18lHqxPzsNyvI8kf3WKjzVYOrvAboujc3aE1L9fLZJnGwPhAY82vH3amkg
yaxtNJLCeQQkAW1cZPuzM0DY8hMQbeAKef39Ssm6hO4Pw1qlDMuHOJA26BXJSII9gYPgcTfatdYk
sudP3nyLcaUYSjeY9v4xEqSzTIgnuRv7ZOnzGgyNsCsvc5Atg1koaZnLaPn6JYbOCydSzeVTz7Pl
Ag1fSlfIbFG73qqyqnwF5FplZ5npgRkrJPOxQ3/p7lSMKoG0d16CSEuh7ajApUMozaOUW6EEnQ41
nZSfuqy+mkK/8BgbpFl6CeycNyC2VULOkX5KmWB/vxzlyMykpCUAezQ4kYLmU3ihzBaIh0ZQE7zR
y7xx6LStoUCUtj6WZDlDf9PWbRHDA8RzeQk+7BDP9ZQ0DUg1amyXDjFIc9BILKiTgRbdnV2og6Gk
4qddCxuheZuYgoVNtCkoc+5xL5aVVUTCy/fYPd1M4P8XcP5yZbSGVtNUGqfCS1gwbZ63LA8gsGwt
xIONuCYU4wF09fKm/ZgeoxjS5Vz6qIg2fTl0kjmnbtEy8APAlqQqMrhbxjZlIMc0JVTmE1sQ0ax0
kTOfe0AnnVAQAz8bklSJD4alOXyjOATbvS2aqeeMZavcaYec9xy6sMDfM/3WxsOE8MLWv4bQwvUL
omx9a67yVdV1Q+J6iWj89qKndp3TPhh9QomMJ9fjr4XZsxCtn1RHOP4FNu7a5xMm7GmmiZCYbL9U
N0TnCp3vu9uYJAyR/JphXK28RarXuWL3s2wET87YN/dyBj3aYdEEtUPqxv3ZluwG9e1VXGj78UCP
4Ijd7Wkv5fOTywh0DI/nZyLA86xLazD6wL4AuS/+7Tg2I2/NjFJD4YtxpjdhJBhcUbu6Qe9IuJD9
lSzMiqmdsSqOxfaomNnvdh+4jjQZQn2RXzjG6ZJk2coOLm281/Tgj/CLT3F2j55q4no00i50I97g
oXYGJZij2+7Q+Ka4UH4qO8FlY/eQSE7AT+yukLhy+ZqFGbCLJB0WN6pULUsLKcuQb6/i1xIyc6Li
ynXEz+t4xJEaa+bcXTBKKCAZD/rxxGPTx1lFBt33buchEET8kglIPNrYUYIR19GineO93xlSiMN8
wECd2/2R+/F9f2gSFAr/Wb6TmwXTYkDH2veDrm1MOHEc+Nwn/AUJSQ7MIZLdiJJ/3K7rUnTBmS1J
d2UAbkbE897VUDhK8Gl2is8XhOZW+jglIuY39MA+Dmin5s2jVHV9rkBE4RStxLISTJyAIVRODUtW
4hcCix+xtlgzq5mvBg+eejPBUp0DavXnBZY9b2TOpCt1icFRpBFr7HfixtzAgmEAnnhOkRl2Vx7k
xGhPbP+I4O7MUY0c3ukCIuOr9hTPhO3R2OZxvuAgNVnWf44AxdHnaRJouJvFEdEJ2HyhN6YpvXzH
jazgNufhZQC5FRNDPaP3w3Fn5iljl5ie60u0x+NxL19JCQzuv4D3G4MgQtIlFl7Hr7ALnhNbjKND
jtLDDEm8UtphXhBadpkRIBTbTHU6j4eiMkrhjwkcvtMVZPUcb9XUAFbnEQ11oN/JrJAuLkQqKJbU
KiOymF1dwhJ0aSnZyhdN5s2swXr2W6t3HHwyeIrTTny9tXCC+Y1rAn6RcJPlE4y8KA1/nuPN94XF
dTaQxObflVs+3U0ZD9NZcupUSeNw56YqJNHyGuVF2ZnHgB+5E11XB+XRoq/VF0c7QLEEPBdDeiwr
mjFKg2grAv5kjbBo2cOAb9Dr8k5l1t1a3yhwuDi932fxaAwJ7gpKD5dleUyIDgoJlOufho7XdMtn
goWPtT3C9vYA0A9fIptQ9ta+KFYgaScm4cWZ98kpqzKVxb3D+wSRF+U0gJ0xzmWgKrIP+CGXSGFx
ljFtfk+PiSVD6pN3vQmWHuT8jf+bNZVA7ZFsH/8T7zH0L2fGbPglMpr5lMiEn99Qsn9AKYLFaNf/
+2U4NGdPT9xjj8qTn4NasIfzrvH0JTZxmvcbN1gfwmiruELLQ+xbtln3OzHEdr2QdJ4s46hkAiSI
puH6BHNwNnIIRhQYRkwy4vKLZjmNAY/EzhvcT3qws84fXebeFOZ4+iKyHTooH+u9T+0/IVgRMvQ1
/I+IJ0kvKPXEHN/TXfxMQnwWMMGxgd0Tcju0nfIQ817s/zBjSctcDEusZupy9qPXmO3ExX+QDIii
vY8xRkraP8SaBSIGmQue4svlNEGQS8uQ55qk/zuHU5A5WMPOq4CWbJtIYZhvkhlwOEVPLGc2skHw
wfDQnDSOOKWmPVQD6Hf1Lj3azlpoxTAjzdEscS1Pw555ioVt49D87/t+rUD0ZH9Ix0mFgCDjfmv4
XkVl7e7VXACNkaGI0vN74BLbfU5jlj863RHqk16E0fA/pGnPF1ZWKLJI2Gl1997o5yPVmWhlRapk
xMpGdn8marYLs+dgMbsDS8RbHZkFIajKSpKUU3u05s9WhSrND7sGXQ9BuSw3a7PE93f/yEk7bEmY
r6/Xgne+kISJTYWbedCKvoTOx1L5+aOLhi5qGSIKN1LhtLlFANphwf4ZCK99tU58118iFlZ39xfL
OvhbSY190pt8bKfpnBvkNR5rbf8lg8RWNwyHFstJ/HDBhP2BpJN09+ra6xZUvZ62aihL8oKOYr/f
esHlMzGAIAm63QIIC3NwaSkI3ZCHre9KNDkzwCJxoftE8t/cPluI0+HTPP0iozPy0eYp3JY5RYwO
8YNlkbTkm1HUGYOM+sdDQGHMzk7TqdN0BVILbyvqHBebR1AvWEMZCfuaN5fREz5msgCy8eohjQzT
5hVrbdu39qUZ106B9bJ6eTWsWP5b2kN2jFXjCM4dVZp/Z2fedwDwyeDoVd45rYStOGpDSVB/BGgz
C01AspzD1wgNc/y4pZju7bnDNaZAbP+3vUx7O08TF2CqG9n6POtynDBvZoSf/9SiNxHHsJXRez46
pYOnxnmf/89pXIPGUBLBb/EOVKTmfyXqp1FRKJdU78KjwzomBoX0pddVRh2tWotc+isiWHrYwaE4
q1uWyFHjoD3aVCFyH7hgaYVW0bdBNd0cUIcDUxJLk/quvNAJvbNI93IKYfd/UKGsNJ11g2NAoyyI
3E2feG/wGGU9teE2o6Lbvm4VoYDGBVAnAm6OPbcdsk93n2vtcTXaAdKz6INFl2txOYwYoKE3L7pb
5/GA+KqETVzlAci0589vrAw+6o/TYpB3zBdVJEDRXT6/NxmxxK639sxFuxmWuMkw1XDzidLgoDdj
STTjGLkFkX2EbStxvdlCHLS6AYa9L/LvcCwuoUMAQ3RhjaGgfCC7KzqGMHg4yCjP6IxaqblskrjD
tg2k8VrjWFbEMhV/BmKKHvEGAB5KbHAMvcFrbz5PINLN9dqS2ezzQRSFv/cE63IrhGJum1N62o+9
Do6iR/F8UgegA5sX5kVYn7R+DqZvdBRdH5NrvDHgixN5mOV4yX++2a+cBwERmYoj1PnAsAwK/iCr
M3LzG0d6qUwclbeje9SlNZe6nkEomSNuAvupX3Gs4GCSRnxaboHqkk+Z8P2mtXYLLoPMqZx3EVPs
lu7FzGdRNmppAguCyChJ3vAFVBg+kyNqqpKIpI7jCFtN38v2e9Mkjn7T3S78X2qLBed7eWnDY9A6
dUMbiXMVqVFePmZtYHUGJj+hhO0h+BtD56rlw9sra7AhWES2cNE1DtNQX72JT5O/OKusfipbxHiD
JiedNfFF1ESlSw5p9MuNbo8cmcC7zYlwZXHLqxAbjFwwz8mbUmaLNSv9eOM4ygFS9ssA41JwSIQw
8mQBI4SKB20eBLscV/8Jf6T6H3iGMfhDfB9+WM5VMuKCxdih5TS0av0BTUoNGc/iBhvsDQ0758qt
R1VWYu7Wez14Oz7iWLVf8Kw0MRBzzSzAwmOzDCk2+P8nSExpUpqtidesKf8AdP1xoYL9sm9vKP/r
YN0chpkHVUpJFsyWHcqt+oIYoUOvTJ737VApJOrsJmCvKDDlarPi8Vtr9wzc56+qLeDmVCDYhbb0
SuIihlPwKyrz+kFFHQPybosGgzB3ZoS0gXOmfYpU1Vwj167owvZS6rXrp8J8+lXmJb+WV99sJR5H
dpXyMT9LFTAaJ/IeG5OK1cG6axe4X3ORlPiJp4O9SfU2A/EpJHKtZ5UkyDsuQ96K7aztcUaP1NYN
cL0mFw4D1TxQvGpYnsFi4ORQ51uWgO/ixUDSnkZYbDTI5rcm6RdbZ1/lEz006NlEQsw//hAgeyS7
83wYhT0iSWvwy3/sIudCKaPF610tNr05nm84OrNAnX9Hk1s91/EGDh5s1hj9F1xsyMWc/lMAIK8t
jGZQ0Wm/ucnJrqB55zL3DmEonBpXkU5EC0VkyPB1Rj6wD3xXY0GfMIgB7zq7l/HdcOckptyRsbKi
xMONJHLcuu7UckxN08J3dzf+yRsg+Bo9XEgyDxqGk9QL6kq272wHrskusBTiYFLh64D7SDg9ftdP
ub4KgarYG5hSQ0q+upcjlLKK3o5DZkmT9hOUoN6M1XFRdQidfzIMxLArsdql7WdnCsBy+ouJs5DW
xzHBP0qWk/XDj/+SBRQR5DeF4IurhwbrLP6R5vwnHZM0n9nC7dWUEdDG2HsWy50Nw7oLhncotZuc
1aP8JgLmFnn0Oq46fsSRVrspdHk0zdIHJPu4kNHkAyzJS7vnWM/RS+H5HA8UYBF6r+GToBQYjiOU
JNMjctrdmKLFmJ8Q34gRO3lEzdk/FGTVNXH5Otb+eZv78yMLUozyxMAffGXfrQJ69GQSQrxo7HXZ
zGA3H6uI10GotX99ISKH8B9tqp9jc1gp622C147IHFKQXVFwkiO10jt0WvTaZzS+FD9vsytVlKZT
2CoD9IBnFfBrBMpAph5+Qn0bd3xcJ7a6YvHOp/yPojDRJK3I3Gt3X30A72maVNGbGKhsDKuqaOOS
VZ8dDvysMuP/MQyFhBUX7r0eXh30cstSCv8ccitlaM24dfJJdudvl3Vh9cW8T9iFGxrlaGMH4Pjt
ASGWhnAU+xU3PGx5kefo15BV3gnCF4g+4V74HNRYDqdqKOu3iO3Cq/+qEN3W4LgpPZluAeMLB5Bm
wxKHL0U2F6u8ZL2Jy+0nGj/kFruvvOmBKrruQr8bvPuVzS9KwQu8TDOWIkt0OmhTzaYU0ao+/xGj
De3QagrPwf78VfiSa8imFVEqFH//03JE7FVtAYRJmaucXM08tV073Wyio4DrJEs7MILPbS3c/W/G
KJUdlrJmZp+pc61JaVd9CmkwDmedgP5OIiqZf1Qv25qnln5VEq7c9zYp6w2CjyWIE6xRXkhGosDu
EK/5Hu7Ou749Vbu5Xr6lzaadq1TL4uJMPh+NSV+wg5tsrk5JdGy5KHwoh1EY3OeGFIEju7IVL3/h
0H/Gm4Khyh4YFo38hpPSYW2HUK0JDa4c5w/2NjXqHX5A0DZUtAoD0Wmhn0c8DpsMRFmGoBglHT2n
YHye1sIK+XbLsDE5bnULij0Zn3cXbNmcWRU0qKr29R8V0nS6tgnb3zuG543Rqb93VSufvidzekiG
ENfA/xCNxR9mWII3qhsiRpDtjgw3D+Kmf7VXczs55BebEDgycqfbsMA9u7psTRs3cV6LZOb5zcVB
jfeEZ9pRWe7UTVydzMunZXcMelIbPdwFxY4sKKamVRY0ERVMunqXlRc1+I+IZrKbJHxyQvxe5yyF
871K5S3Os8wuJozFiBvb+zypt2pzoEIP1G9bqt+iCdpMfHdwRVrluM/UDLOTdQNgH7/Sf56JZknn
nBuL6UjydsS0nQO8DvDhBbLJ0Q2EdYFmCJQH9ig1k0MlV87PEmelIDqttCJAVNKorM1NxZzfs5S3
idIgJSf0KtrjeX327dFKw3DGNlXtGi9/W9kx7PlQ5hdrwQwaWx/BWRZx2PtNl/ftQ2FKiii5Wg2o
0CTTAidgH/mysGOpVWRs+FdRdjRLIXpOBOACjhbLT9FYxvcTfZ+uBNGeFeoWREOltQGmzlLAxIOc
FeQTiGo/UwFHGXzCq8KKA9hIQlchf4ymLHpZf1G8p2a9ATjpvraIH4G/pMP38cVynLvhwk4VTasX
y2scBipcI536HrY8B2msU0dkaHP/bulbj73qp4feKMaO3nqFW3Uvqtys67KnMS3iLUIrqn6M53JE
p4zKabCDNP7KTfiw5edKcYODXiea855cE5V67SlPTqSDBOz9oFlfBMXPqU4/a/zUT/gMefN+jl2O
RK3/KLUyuAa4Ytmb5bVMBqnEXkQosd95Jfv6WYfJRMi8b9gRvp9y4SKwdjXowTggvdF9HWeUrbb4
HqUXRx3UVGiJFsaEjMwna7+7ceGa5Ma/Kezzd7tyli8g5BmB0wIWptiw+UoZEDww7M3cm4srwm7R
K1V5w4w9Wng0ycAE82Iy+TctT5JwzYe8gxPkPUpVYGQuTPN3uAwOloMUfy+K76MRkpwC3m0+tn1m
02/0a1lKTOX022lwvk+AN51JWpmrYSaaa5mZR/8EM07FCcsQKkEHn+bjXuPiusErOt+oJNHCqRDK
ThH6s1l73yHQKoJr1xUlhwKjHBzC37PQdsEyQacE++vxktpbedFSOKIhotNgnMuPfvC1A9MKocOb
1k49XXm6zBHhfQClPSd5Z0Pgh4iAMkceL2ripDjQ07DE8OR47VM7Fj/VrYAh7MQ+9MOO8OeLcEDw
0ag5sAZLbVnvlBZf+oCQq4jvE5utt84iJTCKiZVQiAhlsWJW/b+Fv7KuS6jG5a3/z+BZmb39ryRP
139wIivO3ICzdBKvb3PnoamkbyOLC7xXA4uLq8X+FgyRuwLrr8RrLUdWtPKVzvi/3NG8KCefyGJh
ahGr9DWg6dGWQ0ObMuVJxi4MeY30QshN5df52HvlUpSS23QrKMb/ukt7V4fgYxpavTXH/OYCdfYy
AmOkyT4o+RBykyOM0sCKLtk+P2KYrwGfrmpeggr2+sEV5D5FF0RHI+NhAzERmttObxOuxEZFyNOk
iCf8HspQIdxP7NU1sBbY1OUGFwBdbv9TS+maC+msoZucMcmdY5uYD2V3j/IJK+1MZVtFSkivC3r7
5TQc9iswvGe+lN6qZ4xYowah/gKeQAyF+PMm67HnJ8DzaSmaW2OEn25e1W4OpJ2CT3e8WGT/eD+r
xLAaxRMKsCiJSgpsp35P8r7AzPrhXF+c1nbJQPvymgeoih5B8022TgLGTqe5C8WwSqLCNvBxvrwQ
Tl2jho8iwE70ygu3Tvs5ZL7MYrsMqchNb724IdOLPwBJKHxitbVzQMP8idzlrHno8+ocPHkgtlFB
NwsSPA9TaaKbOvGc7AftihQmMtCYzqFCQy2KyZTFfykU5CGDLHe3UE3Be2W7zfxRlPGk2lYgBGP5
77qvUpM+GjeilU3rSifwyCpdw2jgv51D1b17Kh6OMsM2IPEBaD8jEDmA+QMKawGaXr15MYVvpDy/
F+YHQ76TzfmEir8MhSXQc000sBK/Xd2KifPSTSPmSFbjWWgv31ssv1WivSxe+nQWRFa0osVbfPFR
2lhHbSi62cLVwOP6RiFgsRkHvmHwwXIoCxTBBvbABv7BvsHhWigBP4oAfzTx50Cx0JW3Bgwt82h1
nUa0IFD2QlA8lvI0/spb4wGSN8eSLaPMHVoHItuArRA4CpMbQSYqrvgFznopfRAvyiqqpq1cBDav
gbf5gRlA6Mzs7IyXICpYMpk1NM3a6zpfwq//aObOcXEBvGIhhVhQLhK41Pf9CBez+5ibrd8LB6aq
SbZ+dzuT4JnAh31MyczpTbp9UT+9z0ZJDVOXZTU3b0b4jOE5bj7lLD3xYGWW3VUY1QIpSo8Om83T
3jqaNCMswvvoYNmBWJLls6lTQ/ZnmC8RjLT1L5TnH5DEsXzYR19aXHTPUgwW4mARIHezxoTnbMWH
HvLX3SFFwl2tZXsSju65mXqEBHj+9NYAVt8Ld08vh3fphtjDPakq8DlGWXU16PGONzuwSnfT2HC6
fjGTYLcDnY+ZriXzKm21EHNF1uvD+bd49oTzctdMwy7YGRTuf6UrzgROfibqxXdLR9TnAbLL3y7M
cDYLKOP8mUXIjw3tGEPn2Q1jmq/tZwIDUncKuRH/wzTrZcUhDzZhROKipRofc75jK295HlUDop+c
dMuocAAL6XInmVWIzOZo2ee5FPiINCAoZXt1XV932BE6FsuLX0ByxIusq4WlZV+wEyKq7c7kv3cC
tOKTyNLG7HgFTd8KovfaG3FgzWuQ9SIJ4TyxyVMhgOlExUVoygLzTrpICaGFaapD/isrxkLKx5Tc
yi/bGuhJFUxxPAuDUvOWcLFPyc8NG833ih8qmeBdFuQjEeGcGUNhlHyeHQ1Y19SxzyqnOzJS8lmO
bG00GGLaotzuK3suohDKo4WnR4jVqbRKsKaDga4n8MRssM5dZQ3EOXrAq+e1dgQaMYVKRgPkUPHO
Cex0ZfvBHs+FqSzMQy175VAHy5khqFAyr4quEl4F2ViJaB7EU+jMOc5rSi5kRVcn1orvQGZkxhJ7
wZUiKU+CzQfD+JsP6Aj7F5RM8rLDu/6OloEm7MFbWjDLtlKt5yd0mok7jfEqTeV/ShRGtrr1iPbR
euGvGWeGYf6FyFw/Fm7a42QkJUEibazempFdDFUddiNXKMYQsYeojdPPmGB4g0b3O/XQ099HAfAr
QJObLEWmLQ5gJOofJQN/17+4BBfauX+islI89ffDag+25tmwjaiqm7MouUHcASDQym4fQ+Z+s1az
sc/5BIpq8mMsZaxDnEKaC1ZgyYyQN0OjT8OvN/xyzbrEhG3dufNphgNYKm2EEYvxn5AaM5I15lEb
/jTJ4fBbcX+YVWiriHORcue29xGv5Um+AAqomcBGxdq//YwPt41M0F3K3Iv+TJKviEjtt6FcJjbx
TxZ2PSLSGgyCDccnk/fqnB2eFOHEOkjAe5oZafUYTsccAlFaqKqytN5uQGx16aiVMV31FY4MuOxF
LGVymAmdHgoj6T7QOzomWU33x/QYIoQPX+XFjbbC7mGEhSFgkKDOKgT/3gxLtx4LeV8WrUbUdzYT
uzeR82O5Cnp6cPJmp9fMwaFUnNhJHS1e6Tc//MYA57nZEkpJKVOm97piw4J9GCqNGu4/I0nTjxe2
v+F5N8V8mIoJQ225b6l9pSa2xn0mZ3SlOHEL+z1bz9kEw8S2asRztozVyhi+qRdpFR6O2ePKzXpD
ibZzdyEHhpHt35G1854oF1UQxqSqDU6sKgxAlRxWytQWIxB5k4jHhQegVukL+Iak3XUy5jkaETMI
18HwK0zK/ELibch2p+fP4vZKqZkCtAWSkR32dsoOvG+ceC/gKUJBf1By4AfWot5G+X4/pAuhp7fY
CRKM+YDHBLN79Hnnsg+JYmQEFvgCIz0K5OfwmjcUXQ0VCvHrEXkJSKgPODg14jb5aLjmUu61a6VJ
Cfipg5oqQ3M4YeuFIZgbptASk8KeofrSCHAtc+ww+PUriiDBcKQY/HDkcKgohKwjEfWejjCnsOm4
9SLHDFMjdoOSkP/zLyhgw7CjWWyC9yptJX/z/5kbiK2w00vv9wTcuOezGebXw8o+JDntSTFSsonr
RFrei+vCKRkaQ+V2D4YTzeGmI3wc1SYfBOcxLlmxDGNwcKZfBKry49+rbOwvrwQ1Zc8ykgntZS+C
NH+qnAZnwFlbAPPYWX9WmLneiMNTBFADsnU+gvgKFxeTVHIT2dt0dfAOeRHHXjOTCewe9Kj7POX7
u2muj5PxznOnTGE5Zeh9gGlsvHtY9W1FzC4r57r3wKAKOYhrOIwVe/8jFUY6CaYdwLShngDSAWZ8
7nYIyy2gH6asz5jEcJIx2Ie3+hCZTrgdn9FXnMs5NLTBCjmiLaJKSHRUwPNB8YHAZ/vUmcr5QRFw
/6cOkCXG6t7Mdj9LuQtzyNaaJRMxiFMLHzq7QyczdoioIzg93H0ClW7aBQ10u7eVtSf/rANkrHKn
lI5ULZ/Yt74VMXZ9SC0J0sBivTJiehY2c/EibYT8hXHhoPe2OU1bZpNJnmotth4aSYzWh1pYMMAy
aKJ2A/m7FYdsag+okh98vwMsFuv+v0e0OQwagFtAAEG/ISZj4QWpw0AvXyVu5bvZv5bLUMp5ACXd
Tm3KSkc9IZ+OxmUEfGEXNQvaHywpdAwdwBUazJBt0syufXJtj12c9w3ruLbZ8zaPMIAT/JQavP25
qhOh95ltZf3DFy/Hgf5vOqOnqDWftegdFMc+3U3QWKqUeEDK4xd7urXViX2FuPb2rZZLvW/D1q7J
Pkgv5r20F+HS82AokaYuwqA04Ns/i2cmX+5CChpXzx7YH4v978Ie5g9u5ej/WewIgJ0PI2QB3cB2
oVBu7+gQCANAbIghlx3jMZ5YCNt2B0owpWGJHLcrxkLUyg4lhHE58KreYJfIHeGR8NzCkY+IXhSG
KYmj4QHo/kFlYDKuE3j9xe9h8W8ufAvaZ4C1TC5TaeJOA8WO94w0YP2KsCxoi43pW2nKTcoLexH2
p0o2COuf4M1qy7yK91CuMWzSVBRLF9hjvaSy3CYE9iuoQX5lHBiNKuhJUnPkW720Y3DLYJEa/fjK
Pu0TxGVhPhNQSISKOtR59/lSnIAlikqQJDiHRq8HzhV7eAuKXxAmj9vma21BJISKamzdfGwCVb7a
lAYtKvfb4BIWN33PuHGWg0hh6Kd3ReorSGD0GSh6n+14xgd0OVR6WAexQrSoKWiN0zKxhG6ZuLXn
S/9771FZRtjDsR7Qbuxgjxa2CWS1GmuIzo+72cV5f3F3/S8xm1ABVniKs2eDsjuU5Cf3w2Sf/U7G
NBM3sLPWGS3gr9bo0o4e0g8PLN/YmRIShtEDqVX8PfsRYdDj5o1VQylozXbg/HeIDPGbxxDqtMjE
hcVUlXbLNiSeJzXCcXCvIy0EdWRTtvs/Ro6lQ1hb5SV8bNLBS8Un4Xwfrfk1rL7ifhF5iYBlFpKx
I18hWk56Y54K0ZbaSpZhCpjbZUzng5cBh0cKPs4YE2LaG96jGzXvcQ+ebgSYn9yJQ2weuXDqt5tg
Nl197WZYanoaajdjFqD9g690E8Rz8T4Ky/IiEVXO8ETzSQjB5XCpuMZ04QZ2wK6qT6YtCf5duW5O
x9nzmoo/1Tse5PM3RX8m7wTuwIdJtL5hu1okNmh24t+6QwToMYwkzu3oCxfKWoUOVAkA0Kfxiosp
c5Z90tewYIAAfldFkdor/HPgxDihRFjcyQOTeX0BrptMthJaTSGzRZeNGqo6vD5D9GVcHF9eHNQ6
7OTf4lV7JRMRlaBxONgUOOmuns3SrLUWqb0AJ0n+G+j5oZeSGC2q9pzLQyl5upg9/bKkkEr9LBpH
gF80yf0VRsVLGLZM/d7gLXfL5IWgL2uYZ2+KFqpeH3j9rzGQc1ytxQ613PiDib7Ma6WoHTZ19Fzl
660a5cyPdvukmYQaps40D8PRVUHfShEMZ/woVsMQCTp/Oj9WgsS4AVy6kc1p9wFJPOBueXg6/sym
kVHofrxcwRENACWMwxgOV7WfuqyvkRGeylbQC8PRuJi7FMrfUALPUSfIY21PhuJD63XhZqqHnYg1
/V34xKKIaskOSmx5zSk/xUQUvlaeogKoZchcHrINOkP9ZLjy5BJdkf+xrViTgTQ62buRQlzLw3FS
h3KLUfMwMp24ctaXAGyMC0vEJLjsGCATuvyJmF+sLYA/HmR8gH05DimQP0hU8w9wjqteMx5bqV+P
GqzH7JiNHPOvL9zTaoB2uXuxBkPfvx0PFVP+cectATqnYxGEYx3NE0hVpONVezq1HxT7tRtzRMdo
8jRNW2cZbyGI8agPcoTk0qcP920pX0WY97U1jP1tWxQiqhlZ+Z8z5sL19fCezocoxG3M9Tv0LfsQ
kBGAeZr62+/WFF2sqpOIMs/CXix3vCN9mt/G3OAr8vwDWmTpa6j+Nf3qlA5cUP41Yj9o5rYMzrei
7WR2VueiSW+moYt/Je5z5ZrHR4B4UhbYI5fX+eU55OI1Q7EZT/LbtlIfYIj8s5D0qlvTFtqSOoM1
m7uFfIxxFIOq04dgOjLYQl92bV71hGT5/2SxKRQpn68MgAoDtXpxzVb0mv0v3ZuSCy0V6Bf072yZ
Img4a9LhyHSut4g7sgRZzQUHzqi/pipWB3uQYhNAq09cYl9gQBBJWQeBzTk2ThgVPhZ55MprSimf
aGMZGS/xBL5/Kk8rmFAEcaEj3iWu09RMvZGE6QIcW+cQLUnCadxXLXOPhTFsaF1xGp+vl+NR1Fjf
j7u3Z1BaYdMTAXk58KolfnNwsP1qUm2fwLQHTkSy9y433T9iu296Gg+mjlPU0998uRN3WrKEOxDG
6WPWV+5aG5pse/EB01CL3y1/1KqMpeBtuV7PKDGEszLWVr019Aryrb2ZBi2Obi0F9sjdv8V9r3dq
3hPsrqzbdUVqBeE6I+Zsegdu8SOfIuM1+BJ4/KB5eshU5gQCZkix3sF7Vvs2miCP51ZGva6PCpD3
g1vrBeW/KWIlK7auWC5RNsiqFCoTJZ8G/dwm0mViSYeYzmjz89G6WoPCkjlkNcK844a0Wuemwy4k
vJt6u1UVmN/26V0KabTrBalthZQCpC7TnJnZtnlV9j3HLzzfZUJ8Jrst07GElwx09EgGeUUbOx6Z
8gD6buYMMytkxHMFGveQbb8OCbcQWooiyhOr/WmUtb8QHmyZS4Q4zB3pBSvAXZF3LW89UyXz30a7
MLuIVxo3aZo4DSP45btZeJIsmdOb9qB1jxCaYu7lqM/s6/P+AtVDJODZiTekx5+GC+GzhXx9CKVd
cHvo9JLRKRTbdH/7kPobe5jyiNhyY+0T9wydjj5wHsju+Yec/39W6mD2TXOO8ZQ69JChPjColB1S
zKVW5up5mH7w/f3uXm9SNx+cuQpfsqcH3E46ujv3/s6OgB0uaNnQu7yfsXT5slfAui3a8cAWZ4kR
x6If1AoI+/2mlEFKAL4dcUBaAV+ph7U6AlYlKC9hGQq06/5fL7Qbp2aUjZO/RQnLr54sx8CKXyvu
0OleB8qAr0fqi2dtCngVpiW4BpDf9yC6lHDpKPRPErmZsrIko7HpdNV2LVSzzO7W0fFzW8Bzk14f
gzvQvXCSs4bjHA/5nDIc8S4+268lxiH6ZcGPDVi4t04JxNXo/cFCFx3LvOqPQ/RnT1BDZN/FfKSw
XMJ2JUAA47sNcqJzKMs30aRvfNbfeMD/pMbog0Yzv4jqV1HoDgiIMjhixgk7Ssbijy3SfxCnKZGX
wkkhcfwrd5gPqUguOBnEZDKHY0oK+wCfnm/93T5OfOQpFJ/MBCK5tfXUaqTOAN+YqhWMalOXN+vB
Fx0ZJWCQkF67XOZbIhGSImcLjBB7Ku4aePeAZVWF+YSi1noE1udNnhPqg0dbgZ0DjMivaKGVRU+A
DG2ng3dFm2dhzp4m8T15SCg2/27f+cxiymaevpufci/A4DpC80jXb7SPIrURGVjdRrrtUPI1eQOG
skdExezqUyPQgdcm+SWdLAN/UqbDC/+6a/Q1n7u9Nn/zJpb99m/Vnh3k/rP8BzzVNG9wXOA9t1wH
evVTbo8an+pIOY5a+sQuPmZkTkiPwm/Sritknt/aLwTtB0Ytfzgm0qBbcbrEk9XlNyZFmTDq4Unv
wydYGe2bVYhdbqBrg6qnDpKQPDJhVc8EvjlXWJJnH0/j0OJl9hzTKDjN0iPO8jEzNTNHefUmRK4e
Df/9NAYA2hCtXNXNxCqDz8IMYRNmzX99r1FFWHx4XErImIabZfjoNWoLoLzWr0dEymBS5SuGfV3h
YTuJzQymgeiRWDFlZCc9RaqLV2/fehYM79DLFGAq5uzEs3GQHq81WJdMpMDQeKRW8vrOxNjiTktM
6MZNz/p8vkgMg0fiJY4m61vHeqnA3P5j4sfX/b6/9gwt4DxIDytUvIIf5gEM2WNNdBY70qsWs0tl
YCL1qLcLHMTGfiwKdSeH19laCV9YJIlvLtDmoTFof2RiqrueBX1WdwiMBkwk07z0KOUKMuwh9rYY
Tb7P8cgo09Dn4o2a86wircP/0bJ57Bf9wlD2Y/ThbTUtwBU55Ha8wOXDePrdPzgengy6WheGUrLH
MVJRaYayTAX5FPo4AfLsyz+XCXqkwYVbmWjjesv9e4dTn4vYO959bvXZnZy9/YiMru+Rj8zjsqnr
ZoW7wRjt98TuDEGCiq3VBJdX6T3wQKXNteB4BczcFtzYgAz21CdwI/RQgEZyVnJTwpMUg3LyboLG
zX08TrdeqoKuzyp1tglvowq52QLE7Fzd263JrRsQCgvXC98mvhRz1q4OC6T+B5KH1YUSV8fffovg
l9LrzKQmJpEtL7udh55GgSlgnxirWZYG/GHwMcKr0BFvVU2P4hzSDLVhQTzPwK7F3pJRh7COZBD+
nMWuylqOm2FPhnx/6wV7Hdpqov+IcMKN9jQ6N2dyDNiGKT9+iqJZsz1bmad0MIXGDuse6GqPWlAt
ua020GzIIRKGF5bKIJD5UKWMiL8ncOsN6JQAQ6hAVByXo/BNxX2zfvEOpiGckU/zqdxW/y+n6tP/
bh5TZQfPCIgoFRrfdsLZlhG0BssUS10hlAarTDlUni9MEQOPiNycOrCCsXR93v3HPrYiHAxyJF9J
+cuZohrGSx+ihB1TLSPJ0H6Nkm//mnif4ivf4VlXOWt7sF3ZXm7XwVwEKlWpwXKnghZGQE6lh5Th
wsNWc6/tRvtH/ZzUcfIfHQDWrdrBIG5kVDwAC6Ljc3qUKAPoNqtFYj26h0oD2lxM2RrQHGfHMWOJ
F98jLY1z340iYwNv29Lr4S0hgWXYoDM/4KwGIzIhd7vUu3N3C/yKPrq4J8pPUBxLE0iauDw7V26A
b1N3yxh8f93JovLNMZ0z5ek7asQ5Gpl2hV8FzApN0xxDDjIqxxGLdHdM3s08UveTklj52+y/PGel
1ipzU2kJA1E2ypJXQev+76/mOcMgD/7sl2YBAzBAmu0XemqLaOW3m5xEqYjfkIsWXKPd9kpuIXDz
UIHulKBl5/q+iVkWr9T+X8k272QOEPjNy30kxR9kval5nWBm37zEvOnRRZ52xbQ3bFtRXYzm0HoP
nwfUD1E07qBIiOOQjUDfrOeO/FTntfGDj5auLCy6BBW45nq2YbH9NqWd35b/87JSVND2wAhZEHjQ
HFC97YC0JzSmuNAr0PtFc6wU7hGtKVN1gNdTXKmSXio2RjwK/eMrI0XF5U/ymqz/tVgRH+2xPuL0
CoxeAbD8icm3fO+/yMyjcDTLYxPfuyqQ+m3kw1dIbApzfPWGe3o23f6C6u0wPDc5t/syJIHfG9ti
j4ij/hDfCsrNaOsIlVoGhI2jbbRWzD9zM+acUA5CmUmU7ei7WEb/7pmP5lYxYFtxd4JDPuIIilIk
4e5BeYiN1UaMXoG1xfNxdVf3oGLZ4Ik0/qUJKHskZBe+SN+lfmSQOHsHxf9K7o4t1Nw331RH7O47
IXXE9DH9bSM85E2djTV/IMhtZox1ZEdlFtPz8CWPxHdXhT+S9awr1+XZ6yreN1nFXJTlNhUaPKnw
sXYAQxZ/MhNoNbDXRZenUO0Q21WqTF8tEtyJH6/V8k1kJssnFF+rkNh51ap9xCg9J+mct2zBDuP4
J9yXM+y8apRQ/lTQcxypClBRQ1ehP9xpsRGNygSRweYDFJ0iaTio6LGrts9NpKdJaiBEI52qXRN7
GEx2dSVOcO5iwhHKhp8JLsJc06TFZGl/xbBNGApB3FOrWuGdlMJzwwnUPBpMvzZLoJO7u+S9bSrR
ww196MS/ZUW54gCdmr+GCMvLALjDI1TxKxMkmJixV8Vn9fDaQK6z2lXXeKskwP7EFF8V1LrLRb1q
GSb7COhyjjIccoIKlJIxy4EkUukzgmj/syTw8/L/touNQsozI5im0W8s/hx4oXaxxDdDM3M8Psgw
tPcmZxivZOJUO6OkaON2riNmo8OnSrAoT21HsyXV3CAISupmMVWzUlGZ+fMh6IfGvTjKV3OcpPfV
DD9QhRu1HjaaHCKJUX+1x+px8dlHRcPq5jLNPFz+BBSE7d50VjhdQYTCe9JXTRjyYS1BMi1WEgTr
3Cun+lCHVNLQpp0s6hfQrEANOwI1+5JoU7cYrIhIvNKDRHJQV3qClXDfq9pJQNSnf2uN6szm4N4B
JtsndU68NO9J7ESTd8M6uQMNKFcKl5aLYca9TQML1IMg7uTs5FtU/8Lh1vaAxFN79sN8rMYdjZhO
/Lf2u9oWhVvCCkKfi+Z0S1HmDMGxtvERYtu7/crxmsnLhJt7N7xQTKC3MMXW2uVIQ09lFAMQKI3a
Fwazykl+A+6vYlXLDgPoLlPnGQSfitINJYyZb5146Y0wTM1Q/kCdXQ+7mYKfxqlKNsZWsMotJsOQ
y0rwTtygXBRYY/aJVBjlnu8oElyXXcr5EXt1uQmk6Z5KZTSjnkeHwLNIWzaZ5xNvPsYbI0wPxujY
SM4YfQB4kTZPB1E9jLX0u7BX9+jfaoiRcuKeKPWj/acUNmhhKcX8mEHyzDuHDwxexVq0EtdZtNde
2D2pUfH60evpjdB8ol9NfVQuXSlAWzK1unNLqdO5kQEZE4TLoUtJJ9uffv7BZiwU4trJfZsVmElK
ZNSGkJF1CPja5HRzfFGtwL9H3sgddWCni27s6DLgHqDxQb0O0vHgOYgWrmlyWPa276OEPhMCopGw
Gg2Mu8eQ8GaCSqkKeMVlTQsyCy30BcKw6Ys/wEglJEptNy8K/r/9VUfG+OyLQRU6Ez+qbzM1qqZN
Mc30f/diLVlYBuoS8fPSWg46HJK1vNWdp1IPI33E9kGAhl0dm5TF+Q0ch5pt7Aw+F+HU82ArVNGA
XQszEeLCDVtihEXdZBKamSVKKqknlUaLH3e2S8EO69rv0XnNFKg3i2MBq7a15Kx55wOrnTuiVzc3
W8kolddxPjvVWH+OzEw1W1LLakp2vW8rMMKFgi8e+c/PiZVeWRQFDrvWMeTMBkl+IsUN5UrlK/zM
Ajy3c+e909MUwhSx9pnqaSa9/9s4avrRqDUlPc+uI1qo0D3P+K3YcGFL2qFlijzepBRTMbS2E8oP
PKcRG46ryjpWBU5O2uUjjjIezT1Wt1tI8aaAAKC56/xEDfKSbF1j4vR+0ACZPSgFU7FJ+bIceqB7
dFYCkgSmflYlyanEn50tZuEAKoGiqBUrzgavooACDpJzS10y+Sng+ewDcGu7Xc9TnhAnbgQh9Mza
B91MJDEqCpVjwkQx7S9HPfWersCI4a9hsBCCTeQMLm7PSuCyJc1MIr+SUznsIX6BIgBXqnaF/abq
86xUVjUonlytp7HgzPMRrqUJEAQPCD6tTtOPhwJPzZSq5VOLnpLbExmEQRA7KZdK1RRZ6Tw4XFw/
0Oeeb58y5bFb/FdUbUYa/feNRq7mXA5HHk3AML4yHbdzipv9CB1/uPnNUg2gywdxyiE0tFYCIM9I
r2W+cWum/Cfbv0dCTJPjzgJBWlhRpde3pfxCsV94xYtjhGK3E5Dh2sTbh2NKfzfOBNbfxe2IJ2ys
DdG01/I/KVpJQVjNKQecmZBUGkVZ8sXG3XjMkC9LKHYwtZulmThyUfXWabe0CEcz2bK+UA7I2AyK
ZnK2LmqY4zw+Eyboyhg7BPL3OZHe0oPrdy6c2fCb7TF2nWrZIYj0megWooPs4vbV6M1KX9hqxFuk
CXc0M/WHydto+QI792B2ZG3Me4LA4yzBghbRgUDtUO9/7WRsyD/wwn8NoUV256QtA4X6K5Yw5mkx
uaASzgiMkC84AVeKpGXIcBUhYwkojEttxdOhxIebmJk49BlcnD5cKQYAoX1i5vZVq8NpLA+CTenM
SAR66BtpXBvhAjDuW2ZsOtxNYVC4DyJX2rn3XpsL+gS72pJMm6raSlaJ485F5kLYT1j6UnJtnF5W
fvwr3LIGSuB6aNOF5BDYerDPDsFVUtZ/NIQ4ikDf7+iQ6s9zqrmVYMOxUYQgX598X5gcqxajNFlA
cAcA7jl5NbHC30ft5k3FiIusNCtmhi2EY/KFl1mcb3o8tYl1+6VyX9E2M9pDPTvqDlZc2WzRORct
mBnt+dx9h4D/2o7gNDUCxYFPAq8a1g31xIXgBsQClcaahTcdzVUSlaE8CwsftiybPNg1Zgx5Cg9e
1ufm1dwlo1ZjCQ18C+kAWdV2+NlW7/aeuMi6Yqff24UAlWGGJq/m99W6fSXvRVndBAl9ElIUk1Kx
sQo2cHaklOHtcynNZDecoWOKCf68eRCnI0weEy7znVl6ZyYqml8zJmixLoutxB1zbRV1ODPy4rmk
tg6S+0R4f45ypxhp1JKrouUAGVojtPr2bT7rdeerfTevk6BG6IT4Xnv3AC/dlBvdur6TvOQZkh+B
VgI+Xo3J1V80e1lYnpHncc+PfAS6tz/B7cvRRQDY+BakUNIjpXMhIT3X/QhPkQiE3Qs4lfN99LbA
IemZP0xAm2jlKDuVcJoCLKj7KD4KXIgX0Ui234qBqEskrE/UI/mDhh7d7pR+tO+hxW6ISdbnCdnC
8jG/kjK1c02zt8a1Sv/69qr98Qn/cO0eCTIlzKGxKQ+nS2uboEdlI2VgvMBOXgSYrPMeoSdGJQBF
zNEYq9SdxPFU6CL37ibm9RQhe3DSK1gPSN+xkk2Su1zPzx9AuC7QH6VsTgHmA5BlELBoUeiACRbg
2Y1j9pNun8BscAnbHPh11DbWZZLbb2tUJxtDqJKfPOnXoUsf2PpfmxlW0JM3yz8fNQ1XWX9H37nb
fEPrZzIFtcP4B6KnyVu7gw7ktvbJGnqJ/f+sD/qi9zMzGzVMg9Mv2fLdtD+glUQVEH3cSC9ct0ca
AQX4XkZff3NF+UkN4Pnx1rkTm/1TKK3MvwC6j9O8/5BNetpUrqJrycpQfszvr9sW3nNjy/gjdYFK
2aq9H8JwbXc2YBs5EWMRwQJrM7SBjnfr5O3glAnca9ARjqiO+Xjw4BxZke511rR3yXgXoMoT0/Kg
8oCUVnlybgLnyT2c/GnCVpYTz9JBL0Dce/B91qfQZBy37TMIvBfhjcWIg1UT4ESS62AzU0BwJIKa
slahtfCz3/FrdAUYyitbmo6kBQofrXeSXa7xlS06oRDY8hGsT9UhOctyhHzPaPGagUjY/+rJOCNu
iA9+38UEEt7ZMzn+MYicKfc2FTAVnEtOxIk62H5EboR4J9atFGH1xx63O3V5ubbh8HbaifA97fk7
ik26tvbFElh5WV+I1by0vcjUAbht9evTWN4tPDl3m9gbH50Dynk14RcWKqGO3jee/P+ZIHmQrAko
E5eS1hUbGphPDQWq8FOwvKWCoYJDc1C63DrmqlgjI7Jmud3YKAvuMSL0uWtI/hUQvzn+j82e3EcU
pXw13cFzKkq+jLYUNNfLP0b05rybuuwvh+FEFP9o+tGNpdw6c7DDluJlB5EBBiACuyP00BE8ZoFG
6MOlLRnhflGYc8wD/JtqkAAoxO0+GV98ICeV95GBzIdMyRwoGo7pU+u2/pckiwOeIrCK71fye3B1
ESvhWVguCFYDgPoDy/49zesPa23n06F2yg8VF7Vu93Nj0Kz77A1Aj4fjYb4paPcL07Visl29rKoe
ioztJDR1TxkIcTAHJain+gSIhE5V9HwtPI75hWu249g58tOxb6nBQ+QSOa1HK/Y2L59GuuxEuxEI
NOPkHXu2Tj+1y/e/2VrTM8Yk1Ay/BIzLvukHrviNZvyM6MgXFSmpKFSLNn+ixxIHpeo/YvrhK4za
5rJbWfy2FO/YqgN8qLSghfVDMsolqP6bYACNQUrYSt/PaRQX5u5Dx81z1ioIxnbSyGTRvbVZkZRw
8vGxvqrjdjUBG7LhRejE3LZT7TS4rnW0mQS0jBX26s6YCiz1dvVVcqAjO+oLbpiToN0CmDZg5+5s
L3UpEn6Pqa4teMivjySJRi/X2pXX3mqpaXdpqfu4g4CU6F4ovUqmvtdcwqkxhzIIZPXuBoULQBEu
f5KPfEc9q52VzWa2k3Sukru+2gBvaSF/Bkzp1RY+KVlkTEVHV5ShZjY1HkFkq+QNV5E8b3xW1APr
oZYhpqjk8+2lExfWEMSiw4mAzuPJSl8JD/VGU/Fda4bOeEfSsEpsnU1up4sUAULKcPgEqkgK6ya4
Xf8xMkEyypqa1EyGfLmJZsMgErXEPRqz3DX2LAbJNriBabySna624TqyFxixl5PrIReuxn4OkMBZ
ph9As7b+Wdkn0gV40cOpXGVQbpX57333GLtFM8YGkTdFx8k5572JIsS1S3fWZK7i5S3+5MuaabuL
+MVElajhe1laIvWD6sieqRtEBCxdueLhsScxOEnXHehoEOeljF96S5jajb40lokHThh9vOVtEns6
RDyooFid9JIZ7dlIc4X2WhT6vqzx+/OteLJgPjLaTlv4LI3wlj42ZszRRzx3UNSHCfwWnSoQKLvb
K61iyiVmGlGH+NgPZXWJKkdUj9S9F4BMvk2uV4QhjOwGxKn+z4+7MYzm8Y6QosUDMya/G1SMnuKh
oFTqDr4G95U2XAsrv+a58eChIXY/rSGKqWPr/xtgrpue715QkWOFpotJ4CHk6GWxT4ka6oE/RTwU
HryhTBVI9GPjCbR+OVF+Totr8RUflCScVLHj2sf4Yvn8bSbvA6xr3bWtEoV16BuuL3BqH55nkxtY
AbQf1cbkjdYXh8Nja7YkjWTsKwgfnTH22ugmOAYexFOJmO4StC/GlCChhiwijXP/fmpQvtqICEK5
ltPAtsvbmrbYeAWGFLcfi1oORodQOq26ef2k7x3OyWJlT9DyJL7pQSDacEbEnEzq6yJFIHp6wehO
sfG9xCa9+IWIZ9nuI/S57k420JI83lM4WxCs4u9w6liXRPSmxJUKc66ds9pk6D//CLYEtyqrFN+W
7jVQcNlaSSknDyxFjl2Ir31DQTH5N0m6NS+El9wNcy7+KeM3qSy/7CXAZBQYDSHFdrtLmp+yXBP3
dkbYh6RiqSwIZfJnkdogNcZE7vMgpkbMaHLzXGyEw4g98vkBT1Leo82zJoz3kg2dzjQCbRQ31fNC
pQhDCVcfxHup6ZzO8K/8Jua6LRvhsY8GbNn7ZnCc8v6g1DxS5A4FNJVel1UX2lyUgiKejfYUvF5c
qhAAx9aFVJALnyAO/Nf7lxfAD409povCgScio4zjEsbXqjt4MyGUZ8bpiVrPtT6dKnjHMGalBVsy
WOthblT5IHqv/gMwAVAO8WoEoDNa+PPpTZZpNDmmrqdTXXkpAvZBvChQQNIg4Z1CmClK3aNJTqcV
vqCXatHp2f2yGJk0y3TDpkc/DbKGOHwlODHbU6+TL6XOPcRJq0ixfu9GCi6ENn8FjrOmmPCpfsIt
IcDo9BCDE570BB4ySaLFMqGObUKP67aCTQ/jLA3AEMIplJBteM97CBWRDRNhaONwFzxHLlMTqqQf
DgIANI5bNOixvb/E59f0A7t3ITIdKwDkTbxOgXR3EUgoPWSL7lWpebuq2dxOby0tk9eP/YG5pI9k
/+lECmdsYdDB0FtO05crvLfmUri84MGWzCp017n7/+O2jyAYKlKKcnjQNgjJwi170xGqyPCSmOOx
ezcRM9duDXHeET/4D4pd9kECBOAb3/+ZLoadN/twxa1m3CjSv5oGJQg66UuasKTcpN1yNU+gKWnl
U0ZXYSFe+sRmGc8pqyolbIsN80t3+FF95aWH5hFKxqNBXasAICb6Ol8Ct7HmOBvoc/y4MkOhN50B
X0PhGwhA0OBWrPYOVfKp5CvPL6z8KfPfHbUFzk6koiylGVmpsIOcGnAs/nHe1aeuDv2soaRmgxu3
F6vNpCDD3An1eoYsTfQa6MeW04KLGTqkkj6EEvJ4Eqnfz//V4aluD8jl9m3NeDWvDsmhuMdKbe76
dlfOaV/AUoS2Bc/Mcd6bTKonC9SjtoyFCR2i2DTTIKCEQc3/OqT7lVWJ2W1CGGw5Nuv5iKe9JKCo
MWx0+m+D8gTkxswk5NJ/aA4RnmednYhmtZ/AIsJ5IKTv3WeiUcqY38IcUT+CsSDTZK6SwiAKznTS
j/OC+fIuRr3aj22uYB0UIsScnfPSOUkBdNw0VHNuGZpYU7laa1OaSvYpA6nOVInkMeFwolfwWYiK
h2Uu8O00i3vieQ30J8+B2+xioQisfNLxuW1azFc7/Ed3+AMRNGUXcZeJG9QUcvzZMGz3DL9Afimr
38lb3E4La2uzpU+VJU7OAcMkfGeZAwA0IkgP0ppYMDPGOSCKP1BfEYGrllyWPTJdR4d/puWCWa7z
su86yS8Yf7E5VXCzED6EsWctz2C/dtgD1Y+lkXM9iwUctdxkuQdN0YqIdM7s56MRiQ0QZki3mEgi
VWnCeEEDS63DHrzvf2h80ee4bZEimBW9BBj8Py5D4Jdw3IGEkIuAUmmyR+LQozKr+zXublt7QvKL
CpojqVyPweaoiXLitHlHykbqfkOB5YsnwQiU6nP+sjBmdlpKZD3Qre9iqV4BoQsMhB5/Q+u++xEv
30ys902rdUSgoJAYPHnmw3wLEUsczsGpcTU629HIMUw+sXLokqq1jYsZeQDo+vj651ljmQSdmVKM
b5a+CljG9hBU0VBXGF1Smr3eo02W4sl7zLQXUQn+eZ7FjbjXLiwpbZuvBCNzBZ8JUlo1/3a7yXCV
OQujVvsoHw0cTFHo4yJne/rlEzmDE5TXukItDf2rJPg9h0/Yju1YQTHp/TxYcKE+6Kxi3alJjEU8
SlpYIfTNNuPvwbnY4fC4yl8fiARSNdPw68XCQJL47h0QzKLmsAHR6s080LhAFnHPxmfqn5Xt/qwT
sSgyXxCgGZ2AM52+G/o8us29cE12193GT7H8fKsb67zriMOJ5w6PlMh9Y0OmhL9QFeCySs06Rppf
LgZo1GAvucug+2OtWa5ukAG1m6z0pOiy28Je695jqT1nSA0mf60ZjKF11alAxY0GMUzykhOWGURy
oCT7tIh+knD+VqTzr7s5NSpkALUIKyln5KwiXloQsDNXhMncAPiP1KFMiIf6yZbb5LP9p+czSucF
fYZU5RuhKdXfvwMXpBAxFsQ4neYWxlyrbCcQ5Ls2sroCXnr6EIZowoiNzFCE8qseXtdZE7ig8LnZ
rQydOIazkE8MlDMISfqoX6RIjPbpyMt3nRZEaGFAk33+Eg+PWREOvzijpu472AOt1B7xfph5QASw
QG87veVVJURB/pPmWh7JZVALVviQKCWsxvZbiGH3zdjUnEvg9YPtCbOcABIFRcpmIKTmbJ/IiQof
h75s3nXSERIx4HXyQc/52MU0aU3/9tT6qrESzmuZEW9bVWLR/6/8pNq50jHtr+jdN5TvGkdyiyYL
o6sz6JC0b7q2H3E+ZROXii24k9AfYkiox4ZJ/4MtYjVj8t0Mk9/Yamm9epO0vV78Lg6dm2aSOFZ7
ei4A4abk/SO6yHraJF4WjqXFI108WRVujB6M5qBqTi0mJdD0Twj2AuzhWZQmxLI3zO+RleV03ZDV
zVKJ0jrLZ/dKLkNKV5pvJCqy1i+WeBbCsOeXkPaoG8m6Em7O6IcKHtHxz0AmP6tMyGBJ/MBfhCp/
S7aayIwoEwt11jD5PYVXcwoAYcuGJU1I8IwCpC6AQ6o5wXo6NlIrXo/ksgxPWk57UNpegO48f1Gl
HO/xvHNy2iGtTwSj66a6Ee7FdTXn0aUl/e4nvS4fy8O7akxirlJK3a7LLKv8HMzTOOI6al0Zys0H
/isMc2+zcJoFS3kGxd7LF16981DnWBP4yob3Ji52kl9Ew2HwgqgPba+VAfURAIrnsWXljsZzSJP7
9Zw1Px32haL3+bxl3yFJw9d6WwhmxaPTTI4mz8l493FmQdSCESw0QCMnxELMqzQWj6z6gSXIBXBe
laPqnkLmC5uE3NQFrj9oKzDVcO3peVIISoFf9erEPXNoSTZ+6tPOP+rVrAjLfREfQAFxBk4TG0ed
9Ul99Ge+9yEJrO7udEenejhHM4ghSytG3rxHaVOuMzR3R+cMGZZmtBeOX0w11bkMXU36tR6zjac7
nVh5zqDfjBrMPTf5YS2SoECt1WN3eUQpTRnzQOqmbst31htE0zDDm1HMgrDzSqJkwkpWLAl6wgTT
gPWHjQij64gnquUbqbSuVJPBa3vcPl/mIlOTklgbT0+4YdXjTETYyT358DWsO8B2h1rnYfZc+ECs
wWW9xClQ6YIlkgKh58JSpjocsdOzEaHZs0mSA3vVbycLcuJU6Yq8M0Qd8+6VdLB9yrCaKbsDKsKt
xYhTuLVPeGO7jDSJB3pvSIZwXGH0eEBFYRvoOkBAFKhY3GYCmYVAjUwkVM5F9UiQZTMJsLOposNa
OzVxf6mONqYzufjEiTqZadMF+qaKnhzSLWWTDotGW6NQ7zITW2BmiZiiHQK/KOs3D3tQRvn92PTc
46esVmdoGRwfELhtacoCIrjwK2dUNt5mrrTLhzYFQcr3DGCpV3wCaI6VhC3D1M0iNinL+LhElxOE
ssAmwK5ze2wKT7iz3ABl22vA3d2XpFGVe8Qk98zdTDpFyduabiFlUjbkoGlC/+NiODCbg/iS0sfC
SvQKYmxf9LF1w9vwEBamd/gbAkdStGdg85eHcUPMlonGWUPPleyfgw4J51iS7JFmGOVauM3mwg0C
vSZXjadmwd4v/91o7Wasn+jpdv2f0fn6Ai/nbj6jX49Al80a+WvaBUiWqWVHWgrToZ8PuIgvsGuT
3Lprb4zIoSqR2kg1bZvA5TgKzsoyNd3T3Tf3016KiXijwAjfXUmQuOW/neYxPD9wVxHL48bJcCfk
AEs4RmrKhdD5ZRFkWL7c5QTlQo552MBDq+JGuc7NjjP7VY9uq24WP+5ZrAkh59Qm7EfuK+/Cp9E+
FZdgp6xTZnhtludpfuwZpL3gfSDi+1SobK65PAN9KxEGxQsJOOBMxokuKdVibzKhZGMg8UV8lv+b
KPrJQKiqxf027jWIyrxEPTeSz4EJqBY+UdOlzC/UMsM5zD+s5ENmIqe/DbbGJJLAF4igGrqDWZ1O
FZdaJ40NL4lHT5ZajwPKFJXwlhV1ZVLgUNBCJ0Qp4HYicTvsIGCQRiW7E2+CforAwu3oOvYzhyN1
Pn+p7kFtsFMMqdfreC7EI717FpAMeOUE6swBoVGEtCVDR7IARAiHd1f28tnxIk451t/E2O4FehfH
vL5JDAlgWtg5P8ZB/edO1LIsA7QaVXzqCrygbnqwn24V/fFvHxIwz2q2mi3jJmGEm6jQBScaS+WO
FHodIuFB1GlKqDJXzRmiAqrJ8ldvW/sU6zTRt8/MedWUxsIiVwnKET76PvF9SZ2yZRIPUIcQMYKz
NVfCMftsk5bl1u/tM3inP8mubZzzK36IWX1O15WiCHvuIbS8Hq//hygEpw2p1Qx+Mz9ltF1wU/V+
1kCT97YbCh/u/Op+0EXoWyW0wDhzPIFUuGenfHYEYP59kwvamGjIfhLQTfrwXwYF3XLHuPfXu5sl
xJ7o51ezVYg4Jm8zhrIwpMpjAHbfQd0iXh8Ad1J2lWhEMmU96E91UNukg+Pj+9arQZ0V4QnZrXUC
kwRbKceDTa1uEH0n8r5MR9OtmfpLJnw8aQ8gKjEDb3iPek7qui27jq9L7V1fGlQofFJMqDTPKVl8
eqDT8sxEE8hyNvco0K5NIQrVwTCl17h6JyvfSWYn7b62KJn2Mw0VDBdk0zn0fDyINVO+xLKCZkPz
n3F+KDT2b7syFQite5AUJ8jwL6VXPRD38/w3srbmzTPLOHjR0La0v1zZ3baQYAH+H7llQuDvRHIH
PrF20SWXkiNfzUKTdf22Z7628scxBVHdoo/a5hhXrMlWeZuuZ9UWdropS40OlulZcTGIbVRHkjGv
eur2G9wxmEMMoBNT2gGbE+mThGRNdtDOQb+VFcXu/oiklMw33gW0sggXuv4u8zxzme7dfRUSbmwm
kPqpavxZ0zI7u8kU/lQqHeKDOjaK7PY15kFyGPEdB8eeKYEcEgC7Qlc/uH6MfK0veSj5B8aEPO47
je2Ek1iqYtYgnaEJixNV2tb1hmk9w9Vk9EaayoKQUKI2QdYA0Knf26I1vyMzDTUJKFrfmOJDVxn+
+ZI9gq/gRHwtsm/Ab818YLXQ0eoQKu3sBknQSXW1LZqW9WeVbkhCaKLL/HBS+RBT/e4XkLOiBz3O
E7NuX/9XepGzMrRqz/6RXp19ycC5MGaNxMn9IVZzfzVUbogVCgTQDMTR9KZtY2pbnC43d+7J5DN8
uPmNJjias0pdjstRBGm+6kgLnCtZqP1xXkBXG6TcY7q1noQtp/zLwZamdyQkVvRystYHh1c/KkrO
WIZwSbwXxfVAiCrtxdxoFnmpw8X+uqU9ZgtA6yReDZbDSS980IvsuH6YmQRdd4X9R0Be7iPLI+pV
opz4mhYzELVbyjA0IfMaqoyv/uu00b1OWgvZis7CnbAvnHaEpbq897Mh99a/DHh6rvxhC1iiO5aC
k9VCOUBB2zl/EzXRHj4NUAE+PI5Yx3krWFJcWt1iUdggUiVT0eixyNcQ+Uo+B1cUXTAh5JSC+hMI
FUXg90yMNq7BGKPfsKMIsJcjxY4U9o+44ALMFlr9j2z3ldS/8g/+upJsuYB5MiJ5ClFq/NGgSGri
XnOLkUfT1wyez4DDCMtea1GQFivGb/TPl5ErdBBRttvU3OCrMUre6hvf41KeS5fXx4AjFRq23YIw
saTittW2Maf+ZD6BS55n/xexVNFqC66noqiyr9Tm5taiCgh8jLNh9OzLahLIyqsLFVgWshJwvYfl
o8YQUP3UIdWegpy4d7NU5HFT85J4G8AmG0/OP/8eBEX5PDqyeeRggCeplbjDUSM+cDhhDU40c9Qg
lwUHBgkmTs0ham3PXGP5er5kodmNJnLjLpmFv1yKBQh73CuZCLMt/CamvyBCvrFNb14kV1uIJDQ+
OtmTRRXCNJT2d0+Vdl4REw9o1nOWYqzjKFGZn7dnpuwWwJHY909bXCsH0heByhFoK+GZbtwyZBEl
4KiiQNG92tr8UWEcjPZnbCZdW7dscJPs4uJ6z9U/LFiqHR6/iJC2d1/iDWCYawYyWQcjUBpRILJc
MLj7m8wlWrAq2HLdKpiFQn/J/QQ9v0RXgrgzB42AI6jIj46nQRNr+GCjS0nOr3zrB24Hdn2SjNOF
AJmtKttTOQmchT25h3l112t11HQw7m0+Z7LzshsEPFCAtDFfpz6oUnw6/OmbfFlDVNl/FlE33xD9
0EPZLpa4Ywg93gCRQNMA+8mk8EkNJkACdFHIldHs+aBkmAKWXrnorGNeqy3V/PQigY9+sRzD76KN
VK0ZSkX0pVHmKhzyjEVgDRsNbcZyAkguqI5P1zScU9742Yya1jqsNah0IkXgkacIwhaNwoyU7xDs
Ad0IZSlbVpaLbsNjp0HF6HSgr0OjZ9dKzK+WigPtAXEk7YPJrFOxoQsdHcWBNdTGT7DIwt7CRCS2
vlB5gRkrxTOjBz8d17An/COSKCMLpHy5f1JB3bc/cfUmnnf1R/gQbVsVcBuh2MUSurpJG1S5YMfA
vLxjHfTAtUAtmScJYdHAtH3mRed3+fKYUaBkZGCZ4N6EhmdmcjlyQkarHFfWSwkfhHddoSOdQsbB
9XXHKBCd1zHjlfuatup9mOfh3vuSF34BI3oFbHwlI4VjMaQBjTBajqIm73qvzoYJyKXEvenUkjQT
/Wb8tghSZ2Ehmu476x/MrnkclrOMWh4htWv8pXvHwXPekg4j+rk5dVn+WvuOu5zsS6A6U0VRljMs
rm/s8bzu349JZG9hrvfUrKhvf6nObC+wwO45WxIfBtMayTJHjik3py62dfAkJYnD2WXcKCTkSCQk
xUwQpidl5NGL34KqDzngUfnR8zfiLwHZaZ7QAmrP5v0uOncztpJ1uYtHaesDxtzUtZxDh/nxj4hQ
aQ1gj9Iu+thHRLQh0crImsgZ5yZlgbKW7/r0HuNWUyOqxlw/Gqa5rhYsl901aj0qtFgRDIzE6XA6
6m/Y+qWn9ORF8AneEPhtVO4mdBvZsg4Wnt+7PZ3rSTCjGlq/CBtbQKrxiLeXKPdL3rseKDNyTkWv
kyqjWGpYuPGwEyWAt+VAQhO7CNAU5h/B1q819SuG7TQnMEZE07MG3YszEcnKk+zavt4JTQVvFN9y
AtZ4yvUHpbDixfyQ9/AJdKA6xbIJYqb+IST87+0TAFCosnksJzvW4X3R0/iwdUT7+k/4bh87gIj3
vwAqQwqdM/cQ+ZTe8iZB8E/QHB9i7A7mqAulTwWCKGPAJFS9Tud/+7g0ujJf3fVWxR2AOcywPNYN
8jO49xBnY8Ss2xMp+pnu49EDY4ZJpLogApsvgthAm0icfbEwiBmzT/mgTP22JlM1/F4kdbtgr7Kh
9zDdWzZPKuHzD4nRusJsqP+ogVkOdtpw5Ek9uMDl+R/sHZlp/rFsvlNg8xs0+5Dn898l2UZIjido
i5aG9thcrT+JIY7ZHRd3nGnFzqClZLdvw9aV+jP4yDXGv0eqcIoT4c28XKLQZF7OxhIBENkmlBCn
BkmyaxSEp+0+jjZ8rEGtByaWkG0Ihg8NqbKKrKeUHhH8yKCG0vkYBflqm19QzFB7HuGvfksE8hQP
iKryYYiPWqh3Lfi2cyHpyKQfdjEDXpTdiGCQTpwIK3efrcbIzF4vkyGHB0sU8lq7YDMuUbfcZ/mM
W2Rygx7OJbfsyoGq9ikDffZXZSJL6Y50lIsR3BIlRs8dLaOCmvL0YpH+nffwbF89t2+ocgz5Lu7a
pYobWAIXu9HUosxQOLoJaboScRha3arGL0SFLwgD5VCyZQTv7FUey70HN7xCEb75hxQArIxJWOYd
9x4Jf/keArDDGa7IBmD1Y2m4Q0HrekAHha9SS0WMGxoP2VSVa28dNKeI3yrSS8NqIffD7yzn0j4G
yyzxwG4oR4GGQVXiFcHgzG3P9dk1uawIViabrxf5ENitm9LhhxX6opt+lAGerN62J1DAnwR1xPUz
GN8SdShLWvyimf0Api1IpSnjLye4FIUhhtLfCV5QhybhHu80pk/ljftdEgOJUtmupROLzRMEBLk8
K2E2nKGYeU4mk/1YqGp7YiddBvLDNiRg6nXYGe6iJSuJnEuC4VTQcmonL8eq8A7fKScQbfyOREVQ
A+7QRLLgXWMSQ7GxDWwNEIu/uvphOYahqu+DIxa2OaOU/nPwNMnp9Z/deolN8E5SXcxSESoNA2Ac
od6vBBgpXssw3Ibxmh9azy8soiIf7hkaJ0/8IO0aDtzZ0lFGMUAilCknXXt/en6VNBudQPZgiYmZ
kCR+Ppm5AsCTiz3QMPHHKQG4QFFivD5wrB/8Aka8RORj/yqeGC9UUz6KNWva80myOZIWXEKJRAPG
WoShcgXV+qKyINu8QDlOM/TXdrRlizvMBcxO2Isw+Y9LOr4BwzyfQ6yZrCt5ieSLUtpoMVNE2RkY
kQe/fuK+/JQkHX8RMJcCQ1h2mhyLONIDkQxZ1mZO7qO5p/o7Aa++kYBsjGO/2x22MWIalDkJGPIC
n5BWltHuc7u4khb0uSTOq55/t8sFZehx+7JCaTXzkpAHaCQJvwWjAJj7JIflQ34nwk2ezWEnud+u
SMg0zxUxUqIDpixJQ4aDr/qWVD56RAPDnO1o6YIiUUbDrnrgiaiE5aBzFvDKK5bGwZwsNxZgb1Kw
GzrZaRC5s3LzzEDAedB/Ko3me3yHPy5iqdU2qd7tNc9Rgtscwxqf+oQhKrJ8hPgAqIW7o5Y1gwAi
1i506on/cU7ExAwA6xTRiP21rVmW3sBDfQ9hiNgevYvW/tgWmVyb4fxEYysTa/v+8e9A+9s+Nztg
Qyhek4adgSaze5agrgYzg9/nTnkmjoz6ZV+LlFZVOWVT2QIQteVWZ/eO4wFJoc9waxoC/9iS3pv8
4u48YRkXaxlIobrN8sFWlKhiKyKXdQ30tK2NJ8b0BfxiaW4uO39cZBUgO6safbclq1oTIMzv1jUm
LZCPFdfiBE9PmfHzhNsX6aHfSDjSXkHosbjhRi9yS/voHW2Zggk/OfofImOly1Lcv3+XjmvWYpB0
EB/JS1qVYhJhwWQEDnTIVIFVRLgOtSKFRcQeIMFDNtTU2SCrTyE9Vi9RJ/aN6SSk+nPlE4GRr5O7
V+2hZTugabiMi8dIKDrwK1gEGRKMBJmsDFvwDrvXJ+WFigGYNcAkYFZHU3oNTO3MqhbuOVct1rZ2
L1f+eHPKgkvjgdZ1zgQl38L7w42LmxnyYe34L/Sf8FKvxhkcMKaXTEWNmJB/N9C+OcArE8WITkFt
1EGhAsvo8Sag+odjD8Pu4SFjsjCQIFCEyjwmI97TYJYiLYxLgFhlEoGKS0obogbbuxarO1NVdKug
AUlO3XXsAL4Ys592+NxOxw9UImqUMDPCLpAF+2ZVkJc3HLQtdD0Xa0PCmpST1vwf30WXj3Y9eEZq
Cl6HXEccrKgSQPPdJrGdAmdteKpYcxaXuzyFPvER8zIKfgZjw/NTw5qNCxYsap0SySayb/pJPqWY
WmPDLg3TbZnl9VYpYgz80D4hOiG+trHXdU0jfaSgGmjULT32R4WPmoMSKeM4ntLrI6eY4Jn4yFlJ
lrMbRKXOz3i+5JUD8iAkfUtJFfY1C33Zs4IeqFhZFIh3viguCJcKQFAPGq6GU4LSuXBTOY+XA2vl
T8jmXsWm5RVBhWHhh2PGRhC7AeG7FU7k6yKqVdNLyAJ3OyV9LSe8VK7Iu+uhinWMX6M2xImDVIPk
+xFgsgRbZz7XSyGvPSMCbWdh4woGDjzQxix/mirrl0KM46jsxCJlqn6aiVjsOVdtB3DZuxZ8/k5A
9sS45/KNICr8p+/9a2zYcpXjysxqWeHQK8rYlaE5yh+zW3dEjaXGQ7Ggg/Mn0w3TZVMfLVUOMv3o
f6qL2l7jpbSRfdVxZZu045YWuBGa39oSonT9d75WIT4KgZPjMyK/c66q/Avw1BWfTDEFOobQ3mDh
nRQwXWtLce5SQ8wa8HW5EC4O4HBbPEQmPxsA81zYBwteK4SBkidIt03Z3ZcN9CJ4lv30/A3R2kL0
KRRCfjxKsXR8lA0OTiy95IvMgXGY9azXmAy7/z+ZNmv4BEYebzFNo7BPNBL54JZDTXW+mOPZmXVv
5y1Lh2EJgEI+3V17J+ehueo5DrUbbMuK1hLov7zmYYPtSvczDqEfGhtDZwIwqAaGGuzlq55Ieexa
Ra8NHhjkBusMj1NsLB4yPol6Sn1raY2Hgvob1fZ73gSxVr7f7zr2urFMjNJJFZgpWBiYQm5mZRiQ
mZENlJhp8Tt7VKgqAlTS9Cq6CDEC5JIxDyCdV5GUp4Q59naYLnZpar4axuvKAZXt48j3H2Fbz1ai
weBmDKdRSsjv9IqpLiysvc8b24FesqXcLgFN3Ox0EbDket8rDKHqN/0/aRxtvKieZpGTT4IJwROv
xeo+20yQLAxM+2x9DYKBvgOuOfA0GKWNcoB7x949PT6HFzPmmtefUAaXSGHyMMXcX2s+MGU7FM3T
foK6K0eWpkm/TJN41UngVvD83akhSHKwNHWlzRcGDzWJSbQqvKsPZDjcqBdkhD9AtMDR4yp+4PWJ
TDLpSoLdIQwhaKU9BreX6e4cRcDvStg/sjHJPC/A8efaXMMoVY6vSN901UAFUR+NYgUC13QdRlO0
6pOx6sWoG+Ay/V4rxRzuJ/ls2/Ck3Mvgy+v26Iyoso0wofffUqISxv3Ud3sXtQIPw9hXcHMX091c
Rr4iX40Ol2YoTe5GdpVbkD91G+wbyNbewB72UgyTGEPpjJmjB9P7kpK/qeuP9IXDG4HWl5nMbKrp
WQ7FGC/FnPHyBD08+JlxI0dZf15OPXyb09qTvVdY/40kZOIfOR6bieH348i37DTuOrWoxp92H0Zt
dnq5BtW7MiPIXHJh2v7VfPtBS7T5m2OvjNg6I9kPzkckbbk7GAmhY1G/l6y45UKyQeEs7hdvQQxn
AaBexDdUekfLztKMnokjWjparw/o95XjUJh0h9V98GIGzl+/iH7woTntZHIGxvO9vzx3Jj5mp4fm
BDZVzj5VwaAvihaTEXHyC6hIpaKfa3ochWSId5/66sWEWxDXDxoUaIL9oHwwXr6VW2nGh3LFT6DJ
F9XUDz5MJnQByT9btItiKf2j5n94ZRnCyGQ8Be1n9F4/rGMb6MWi6uOzSYBAWfM/OwxvKeztwCtx
VZM3cNmPPM8PXvo7khTRQeBMWch0PCCUiwgqpN+vHnJq7jKjzcrIsavbiBARYaDmR1rdNkMuZkkO
gh8eLNXtFiKJR2Jqhai3MPjgAZHEho6/XoVHQzViVGa2WlucqV6/taDuNsnwk27l1gJ3jKreo5sy
FOcUj+7y86OBmVQoazb8x3xRCX5OFomV2r2oOS39s5tQ7xAryGfbfQstHliMm01Ou2t1m6xsq/da
nt7nDBkJfg7BRTG2rYFUH/dmt5s2dcTFUgB4bRw0r2mVk3sR3CAE6FTN6XVinNopJHH2guooK35c
rpxFxRLwCGy12jJvndEcN/l9CWRuI+ssBioITY/wK4ftFmjqWaTV/ZHTt3VPm2r1l/8aKilV8O68
Y/9mvk0D6Bo/QgEdsCGr1VOD0PU0ODSK97WCy1fc+Gu2/lSx8zsyi2rvT/0D1E1XeNIcDo5M+l7t
D1A01ujQTrhyUluvxZ2zEBnq3mFfdT/0rL3wfrl6d99gKUQhZuJtMRnaJ0mZnT4sNq3BnRGVRSYI
ExriUSNyjlMu8B+Id5GocDECRYDgu78AZn7KTt16vapBkOCQIP2uOdB59oKTH4hnr6RXoLtCADAP
Kx6cqgazpR/o+tnpv7EKRIDqyR8bazOeBixcL1O0MH+8rVdWC9J/Wdidt3FuD/D+NhqXkBbXSWAF
zS6iA3SZOmjl5ciktuhF5mcvWDr1hrBUDmia2Zgpnvrgv+pbrkGn+fZbVI0pJ7AKpWVCSO2XcJen
Vq1Wl1pOmC1amHPrDnjpOqCIs7CB4xLex87gmzk2vDwwcZL/hGY1joydsKRYovH7vn+iZuiBWoyK
GU1g2PYpG3t+QvsdX6mHMHOmcT8ZLQiaZeihUggSb9KuspaDH1WXO8K0PlmthsyhrM6u1QUYQXIX
gNnjQMWXgcuL34W1yMzYsepH0p0Vt7H0kkSq6RBqoDJezi325OEtwlca6+rdndUhLZp3moFJrJGw
C4lKtIiK0/XwKaZ7CGpaJxN/FbB0s1yweLSyh7sb2hu3yCHtd37eXWRs86jcXLG8dCxjq5Vn/Xd4
WzCXb596lgMFFM0X5s2xnz1WMzMEHwsntKRw4jni9JYpOgympb0LcyHpSW05Lv6573+UgHPyVCMv
NIzZXQOIIrbo/sTXYuLOgVWLGzMVM2ryT7ez722prEeRAwdvetaMW1kjMLHb98/LYLx42wszizRX
oLOBkmfnr7J/aulyq8tnpdytrxI4ZsOSP4YuCcwxVXK8d2fcG7Z7/W39xQXICik6G4Y9FdFXSj+a
5/l2sNDyewSSm2mG3l5lefmQGpxo1fmdn69TmkGiEuMFJU8uvbR4qVN3lcXW3EZGExHMq3x4dUPi
IS1jlUccvJmCEX8huuo2kpalm8pPWVS6ObDF1iUrLwqQ63YR3zlumAVAvA5+cLRvCnyIUwq1Xek8
+gat/JFKxQmJiZKD2z6hIk+hDq3JjXKdEI8DLOiEy56h0ZoPBMwvhJI3srf5YZ5pvNJ5iZccz32K
Ix1kSlCIZOe/+37yvkbbt9LvC7rHTrX5E1DlAAT5VLmvKp7xTFg4oHpxauSCN4uraCTLtAXEVbn6
DZaS2+osfjrSprXpfBrzT5F66mEsvmO6F40EN11FMcXLG/t4Kh0f13zvxd93aFbWCMs5Hq084M43
fdQ3dsodH5tbv5bvJke8RvoBj981V2mfV2l+ppRIifRfLjo13r/KNxQAKONe5kfxlyI9lPk/1c4B
mepKLtJ651sEFViZgAgNTd5J7scfDfQ109SJ6+yUHvFW0Qu7n9S73YH1OYpH0oxjYQCXgmGiK5ih
TU3MppD1qxM4BeMiv8410Nvf9Q9B7cpaSfSUkehuIjvo8N7VEQC/AlYKjWf2b6hhnaNW/iLaRJJu
giEPS9gLt15XaFNyYArpVFzQuJyHt69x7oNT2SE4C5uvWjltUPAtWk5zyRuCeTV8rjLhQJMQdGG5
LWnwK+U3/hVCmfnrtk6pWBLPrf+BusDD/K3TGEMhaAlV7RIKt1HOvyGEC/x8wSjxJfnONzG6m40G
s944x2U/dEgEWp2bU9NrELDimZkdJ/sQjseBJnV0eSOsrp/x2l5BWq3Ij4BQ9f4tBBgPsaLTKt7G
8qrR92xVGeigZz0apkmDJnAuODicxOZuDEnX0x9cj20G0qLrns1MK5o11SRCyPh9mnczqGigy/jV
WB2/uiZBGVz2LvbO2BALeyf52pTb7s3OxPkMah+v/N45aF9ALlnQ5V01d6+khv1kFDYp0HjOQ+5o
fDxhzdsNEKoTGhoPycyAzlxHxWgrikOaCHFw0rPwqk0ke1wHq8grRHXmhcgMvg15vs0YBux3sKZa
893AmO/ddcJWvA+Ig8Bi5leAXO0ag5OYfcutvpD7hHbQsihUXIIP5lPfUKd54q+GkdXCDdjjX3KW
mM5eUp8LF/+rgTVZAgEFkdj/lgrktfrIYdF3v0BH6zprZPPU9fC3nPMtOVyFQrYzmc0E7sGJ0B8B
iGHNjOZj4W+pf44m2epPUPGHCGj9/MXph8VobogCeWW25OIBrZ9k7MdaZf9OjG9eXCCESOiNFvvg
FDHsNg1zmWLbwJEAh3x+a/5w9BOaJer/KgFpivbdcKKQZc7BFN6iEr/mpcoW3wkcxEjljRORaIjV
2kEvs/UZ1ykguoJoTcWttMhiRmwr65as758G18BCe4glY9FgYyAvkjna9slLO7bdfsQHj1Ddft7m
gJatRi4yYAuJx8MPn98zfc/bhhR6aO2wIUEuJ0Y3w32ZAwt8QkoHPdbXZOHyiMkQmZPr2XJP4J0R
SSYt5b5LNVi0AK5f7h38b1HwzlomzfptD4++mc7HxRrltoyg7dTLv8YAD7IiNC+HDsI5Q9E3yq3r
YgUOiqw2y/9YEXL4t/dsvuOCUpNCv2l/4ituirPkcsSgTaJtsGZLn6CuTrt2Dn66sde8JHUWwshN
imGdwuSUckkEG6ZA1gda4knl9ixSzHMAJjOrsJnaCD9jjS8UjPvsJXQ3xijIZveh9DJWX/z0yEnD
ufWQkux98WgI6ekFed8bQM6sAfC/TORCXuzzMvBvVIP+g6IxGmVEddNxbTPWBCQ159BJxjUREzf2
wJ/tSuEaMqa/4Cp0OpK0VMHtzehbALjKY4Ql0AsarO5suXR+ZVm4mH9FxalTboLIJ96klQIzOvzp
DBCanx1zYzB6s5j+D4GfU5mZYadniEhiE+xYGSuLbomeohDI50w8tOkfAkTUmgUKd+q/GKGhAiXz
R8Dd2jGNsXM0mJYXuu8pYby6mR+NZmYHwrQaqWCEFkStk2Ji4cTzD8Wcu4fyFOcVicTWSf0muopG
sUZxe6zCt6c4v6obwC7mQ+uyOyVdiVnsBKntgU04KP5SGRc2Qp3cbGNa9eG5c4LIMeW/MpePELVC
JZLCC45qVsG40UHr8p0HTXWBySMOxJDb+24wAStkjsGIKIojjWEB/Sa0ntg1JNi/Vtl33mXCc4e8
XukGDn2AW7VPDjedTLNkONNXgNSOud2ySQiRfmzFkDkv2g7tj/GXklcEj+MSWXJyitW/ve2VgA3Z
hIWjvR+UchZbWQEX8X8PrenjTgm48BzPHAdjLIXlqM+GBykOb+vciaNTYekH3IZypwYeSsAjCvDg
oowUmSvg9/Lcpv6ToCPpOzvDIJLm1cxclu1VMQ5NyTFJGuCXSaF7U+HZsnlkr/2cxw7mE85/cee4
2POxqGFhaBMQhJdZvvawW8LHGBg60UJtc18uiLCA2iod6yOuOPWRxwNyQP9ZT7bqLDtLtZ1LyKpw
51zHmyW5YdUaIQGUT03K7m3SMD/c2E/CFc19dY0bE2NO1jtvOlrWw7F3P1vX/mLOKzTKbGV3txZg
Hi5HiKaXJunY6x3diwwqjozEK/R0B4ujw6pohwyTCeyMSL51foAnf5wLGFBYTtp2iNc+gXhFYK1E
+70UvFMeiRwsYqW6o/RWHX4fYYNsohRN2ceW/1TdGKLAu5jdx9XfpwO+EJXdZ4oWZuTM5f9YwpCD
I3VKPeGQDQ7xxzErujbQYR8enJCOc1drzBCTaHopR7zFMN1HeqITfEbsFeQvrBV/16dMm5nPE31h
mSQ444VLA3G7HzkvHwjWbSg4TRlzvCymsfU0JixzRI+xNlJISOP+/zJBLXFQnCtoo5imwevtjTdq
eIlZlf/LAvgnLr8xIcvb2Piq7hd1YQFSCMBMe6Oy7Jtn5XbMQ7YUM/t0VvApWk2jzw9qkhlE+hrS
Y+ZYrsO0sGuZgxN8nHc0ekHE/+StNDHZxuTshBn3gL/9BjQNEgHPr3z45tSBzHgicnacwkkUdF3f
1eO5a02vPoasMeuSyHEV+nN6+OvhVFSitX66v7kjpUVKSXgqumC0uLB2ar0YawYVseS8O+PuUVeB
arjK/rr7OokDDKERqp+1HVgLHWqirQBA0X1RclboJwuwTvGv9EaO21KLOXxORlSKGQzjByUCkk90
4F2P+srYOFQ8osBN3QBvEXlnHmvC1wUxVJ6emAZZ+etbAMJb5M0veRuiPEmpbKxjSUNMWoP4sdg9
UAVpFSDkgbfAk+EwPLdOh64nnUAOsiwSdV5XeUcyr4MlXxgvjlSHCmnKDYB1eE1TMOkTuukoMsnY
VbhlU1+YqHP+yGcOoyG0djjPBTOIbs8n1XPYRgTifhGK18DEBGVu9328lfBQd1bSYHSliChW58P8
nGybUYpmyHdRFWFanICpD6k5j4fJA8aNOuYIVZeTXmrFrMOLNpNzknvimSu6IXdbZS07+1weBzLQ
Rh+rpGDYE27L3/DjQjOoANYyrJvBAHAJNeWM//C0YNFA0vwGD4HDCXSo3Hf5WYJAijnZEwV9pkqp
vqxdYIAfaFwCpM4qBVyWd+w+uLZXe5aPkDXegSF35s6zQPfZuCcP7t9EGrcd71SDg1O7F7NTRFM4
Hh3PhZhcyfDiAXf3VwVP+wgHoWdCf1DoOJ+mxbd/pxt2PKkC/lY9qQPGkEjXPzxKfZfuAutEMugL
fT2c4NuOTbGhl0t7psEG996CYcy9xfoBnRf24LEG57cQffTTh7S8zOEAU/dBubEDIqney6kdSWks
ht2qxxq/ZtRwITeUfE2lCd2Zyu98nh0p5EvQXdF1bW5p3tPx5ywrYxCeeduMeWnhdOEiXREJdeke
mFmnDCbr7W6q4ftFtKYusNyNyRh4hPblLYd1dgkGhWkPT/61B4T1LPVRIwRBjALBMRHM7xXvH3i7
VUM5ySn3Psq2Itha6uzCK4Hrv5t5+wgrQJxXazjG1NWZzfwWvIOkXcyzbTtuZXJKFCbCSCVocBVc
0mQ5sg4Fkq8p2auSlaOE9ko4sL7piCSxH/K6DKKVvfZpT6FQSzGNnu2Wgon1dhLOfzSvUr8tKV7X
2ekiArsixxzqu9dgA4YcUoR7ISxE5Fa9srCNaJsXi767k10qPVI1cZlNg3Cc74hpatEakPeIVYel
04hCU6X4dz0Jl8p+5x21OlqTNwd1ACMJK6O/Jch9DC4heRYNLlrwo/CwLXSwFRTLCPkbCnKExMn8
l2Wzz8ghtM61Vu41eUMgvUqUT5ZsDhp4S4qhkaIGPZIvKKJuDDxh65YvJTj/CjPAXogjO3MAUy9G
GSQU7XOSNLxUeHTekeSlPMPNZfEvKyftEeFpwWJfAt9BHhhfBf9hWALU++SlNZjnTy1q9S/sGD47
q5PsC2wo8E3TSkwAyjRQ3/lsxz0/T7GzxDonSAVCzrfZX//uI4RSNDJ2l5Rm6HtYe7Ijdq4cAq8d
cOI1emfYiIzEVmuiriD0rcMgXS2fNLese7u0xEH2EHf2UTkqcZrTO50Vt2Qn74IPs7770xucDA2d
Mbf1rmbpZfLNjXdr7ZaOcercQbshT3Mi2YUQAxseiyogEOGuEJHhOBE96Y3UoRuqyJwLlKcz3hsX
8mq3TdwvdFlfyNc4zXLzTPnUG6RjK6ScQFeHoPBgWklSZJMZS5xvbMRviKjSLtov9Gjvz2MOZx9L
wq7V5g2dCyhQEgTaMMB6UQf9oljwR3aIiazrMh4gH0yieycSJqzBStMLZZNghTg52NpHnUfxnvnZ
cgltNDTtUHPaMtXywAWx0K17mfL/cov+hTgr5exiAdJs5VSMDnxj0eR7Ap9B5nlWsvuG7Zp8V3JN
o/YK40cegn7XhyowqNjJL2tDw+hzsBvZ2B53ZA5SbN9kbyUCnca30pF+ARfM7G8ZbwSjXIZ3ctas
dXTQeAhJ5z6KpVjfgGxaF3obu/mtL/MbFc4B+IrRJE70xNTdwei37KKlBupbGCrfQ8Rl6xwX9i56
Lcj9veyl6xCiZLQRvCFSAjv0OKmAK8rDtRdUTmj1p4eQpUaC2gdNKqg1CaZJAF+1jd5ilr+0oRZd
ZKfjGUaGd1QfHC/oDCuJuy4gWOUczocWkon6HAX4dbdvemWLQCWNYmOCPJcIkQjn2eojKQ/OejVq
vQr6yWDSfGRv+dpe3yWbpfd0ucttmqEQ7QxZtP1mcEiUl1sRpib7o9kaXhk+HZMiItB7iX93NMRM
dcttGoA8IqiSbBYyaRR27j0GlLzpVjAtbpGUcLnJG6KTSGxXplBfGXD4sdn8va2/m2e7asTyy+yr
pop9m4l2pICGpogpnwCF6h4EeDLmxGlVjPZRrIdrftC8MGaXcfIJdPKLF/0NI8lfQRvOCy5YsaA/
1hJceG3wnTcT2Y3IdKVQFzHM1766B++8i+JDOrWaTDKZMnQden4lMBd3fehB7/sEXaEUm4VR/rtW
WS9x/3QnYHxAWo3Kdc8Du2FOTY08D79GHM1QGzYMa3ofuO1JiCkzJT2JLICh/uJnKeilsI1P/O72
hhWu8H9t9HuD8ygV05rbdl+NdfzVFyqtgK5NLxamLzFwNYup8yhCx8yFed8hNbxMn39Y2yiVR0ga
VRWZqi1q7ug+p27AUfG+8Xy2fmxLpQbpD5pvxWl5gSYf5g9rrms2dyNzOJ69lXV6VFx7cp41wepK
5OMRR16NziD7RYqu/IaOQ4XYXkdIqa57bv0N7teGwlO8DF9vBh/3lAtSCGoS6e9eCMpiVBLmy8GF
fboIuJ1hAiq2qI36ZcXW0U8WdKcvc9MQt2o7QSoq99fZHZovBrfTYJMeNFUU1YU7HDOyh9MfAQeB
HPWUa0Bf54UsgBfzirpdWcXBNlW+zBBhE8rkeY35J5Nztw7OgOU2OcIxAlQnX6fYMf9ZbUSeprEO
KHIVu116xurgZX1hL5agyKmt3oUndq6PkwEeSdl2LIYc4Z8CP8oJ54ihWDWhSBVEmsF68B/uPNbm
1kjHQLxtpn8PCD88sBjNUF3WkfDH8Jxgis6pXi4fYqJOW5YObxHCbZYU97LKk81Ai2dEJVOM9ZkC
/9GTJzanUXtmuyufxDRDcQI7CsHolfkXPDn3ns8OAiVyl3hal9/zalj/JZDuLnl5GQzR/zSfed4j
RMUq7p178FOwpjZJbGA0mufmceqCnXGEzkLwxQ3XjSi01JKvUEz6G9DY0xrD6E7mv8FM9JObk1hN
7qRtBgsZvL+qT4klLv7ky3n5u3yohAgw+vCcH8a4qFO0c0e1YZlol8it9gbefg900WLmtodkK50l
YKWGuvHfklrkU6KZiuaVQdjzx1e1D7Y8lazw8lcFEi3QktVsp5Q0flYTGW2Nj2qGjTDb8xM+R0T3
xHgK+YuVcpl23ah+L5hvCfAb6xNbRXZuw/3QJs2wpV5p1VKQBDXEq5aVRbfbvznEz177xTGqK7RG
3s5kkryBVgxCct+tozYSKHBQ2bjql2N31Ly4xWltNqUv2WY0yDRvcQzEN7BcF6gy0+ZMD7GX/ced
dgSemqST1oCxfNHStGQYvcCTucwikTPPkSEoJvtD7vFmnnfu2UjwPnwSjKi2UtbLzGtB5rpYj8Bk
hN+eW0a++BKyCeIMdU/9nYbf9rwoaxDhOlwELdluMPSCMa+21msjzH2jt/tdOqAL0M7GRNAcWUtK
nXNiRwiVpRO7tSqK9mzx3OfIICwu5ltNXnnxFiJyCqvjGSlpdbR8LHvrT4P0e5CYMQHlSYZSOXIG
UOhyQJRc3HrFp2b0Y1X3/ukJkA6rB5Ho4cK6pav/y0HkE/QeA+GojNm61Jjgpl9QZUj1GuSwYL5D
1eVs8KV5EJHPo/PVym8Vw5FQ2BlvwSg+zTrQaC88708b59KVKGxII12JNeb6e6ut+oxEOTEB9bzo
NE+H2VRdsBBtp6JetzQlSA6YkmOxyfbLu2yxiUKWTFYW91P7fvQ4VpMjhZbSkxTIS6k1LHO1Hrrq
VkHLOFRIAqcEV14qsteZqTSQS21v+pKciHxA1vRTVw7GmlELC9ZixcYbJKpaXASJUfX6IFPhU4xn
xSPabnM9tz1yHIBgBGAgBBrbYlHTOQI3o9EBezXEZJSs9bHqZW/TGVHenKEOzLqXv4DDDC7EWcUr
y6Nvgyp88EBaMlZn7E141oSp2Marvc53+3yeFpZlXvzeUIsqnu4oOASWOy/14rDH6FUIKv6hzKx6
Tn502aUc8JRnATRf8+QQ38FOVwC46mhScTDaYihKYFBnuw6TK3jaGfZxDU4C3BRS3Wgu/Bf14jXw
E5KI3JQVjybZ9S0Q6Hk3lGqguvqO1lkDCGhMgwf2blNUujwANadcDITHJbh8GUVNSwyORDZZv05O
Kp5t8MPEAVy7j+KfS2lz31o/sS6sTUpIl2QvE/Z9/fclrD+9OCDCycedXCDDk0/lzYfJUMUzZV+3
byxpczEaHg81VIgaomNxZuaG8m09yjh0ddRDBJoKuREXSJqOjqI/ppEPJhR8ZKe8CbRjqXVEzteM
Ua5mR+jKBgc83jT6oq6A9Nja8d6JbEJGZyMBnYzCEducecLHwoewd58iU5Y6WrpWkof31zefEb3z
I+kztwhIjxK9FpjKZt93GuEjKoBnx9hHv6OVxFpNyGXjecyIvIznO16az/nGcYQKckw0YMq95azM
SMyL1FjidA9VCY0WuWGyH+FHrYmhmwIQ/k8d7WixYejjzuUnxfIrwb6E+PzD/6K7LQ1Rdl9I50LF
fd9S0wOy5A9yzREHZ85iMG4lnr9ziFQANV0OJIk4xHegbY2ffgrKjRo9JlW21+7DjMN9GbhqvBk0
/fBxvV8qcBMpLYTzrV7fHZ82l1FkLKM86DX/k4cumcGNsVvQzBoFMv6JkFVQs/8J3jwHJs3AbTi/
LfTo5uoKtgRkL25wES+vEaS8Ti3GC41GPYtx5/sEC0ztc32+a7B0tBzaVWMVUUHreyQcQvd1Tpl6
XojFCFSgOba8rRW8psrdfo0yNNPDnS5+/GrIjurIEElP8wWsWEN68TvMEs8v/uV2Ks+ynUsQjkta
jg5qyVdVVABHljS+NffFklakwUlWli10iRlB3DwdmxMNK9lC6chkbO7hwK68/n6x2UUG6D170bBM
SN4bXxbdsMAt05HqDlzf1Kod4FsZ19tF2S82WgoKyr8/8iYKp9FSr5m3/ISun4Tl/p3sRotmnheF
9ihruGokVdAPxeRJ1smxI2wtI4tvWQDued9fgb0YKnLX0Eaq2r0CHDvayEKcTUfEa97u3U8wwAx9
LOT6BSodAUF0ppTeRXOdmoPIARiOC+HcENEh+ZHoCBN0SOYWxS6lJauk7m8JFSi3pmRC5RUlXCJh
+YP+qp4trbFSoeZeT5MOaVnLvmf/6uwY1Y+MrTJ3bkgDN4rfj2Lm4hxrXWiyEGop9stgg9tGOKSZ
v2ag2Miy8v6hC2AqBSd5mVj2radxb8aSPZa21lxuqzCVkq28fv0rgBkTxsld6X3oP2QAJ3adAHna
+f2mw9AsyIvBJpvznOHKFVLIA4iol1Uqmcvh1CIm/y5zmhWQCWoZaL9pyVsf9L+hQAbs/fQRLVHH
M1Pc7ZlqMBrYxMvzEqGF9XJu6XE/fLdWwt/cWx2rQ6x/SSFV8SPstCYzpArtDx1X2EvXXhYVMjvn
QtqB7H6+BU1mWl5hSWX07wAAJ840T7PwqcRcBW31Nu6RsDryC+pbzvm/4tFaXhXptrG1pGeHQ4Hs
rW2gKYXHUf1mhv1kl1fISqAsfQUBtaRRKbXi96IGyNLqtx5ct7+xAs7yLGeVOZ/Wq0juMgcYKHmL
cQLs/e6dZNbHyJsKlutPZWrqaP9+iKd7dD/L5v2wP8nFeKPEVBwKfoigu0zLfvM44f7qmueBxcKX
T82RXVMpJGZCLLvGp2CHiayn5XJ4H0+TK4N6JA/vmXDT12PJRPHibZ4FuY5Rb4veC5KnNgLLoe7y
Sl3DLwfql4IatnKXLMT0fgvUFmS85FutHVJt/DkII01Q73cJNCY7MOpFTfkabLBdBhOv/NQHuTKw
NHpWihwI2Lzzo/3/FtuI4lR01uclKj6VTVbPrFgLamCr4txi22wYNN47A0k0yV4rIf5BollOFh0u
chm6DpQqJISKxrjnIoPU3CM8a860EpquSbYREAbQFHsd7tmWRpCi2n6pgSnZD/dsZUEZ1wWkFJp7
4ofIqN117wLqKdjQLJM5Jw6RzkLgLJppcB+N61bQywAAYLOjb3PuB8S3krBeUfjX6HwC7Bak14H9
09IFGkw/aa01dtKsJVfFp1gq3pp3VSvB/Ge6q2shNhdtkPP73Fa//jp8VVRQpPE3rgxy1lvBRDv6
rJP+b7HNW02LM/JbvIHuIDpyg3IA8Z/+tpY668SJpTauunblBAMdia87rz5ir1HYHZrIz2pHJWff
wlB11DTrl6h5KZhCnfrTXLF5AHsCcpqWBgVkGzh4A5q5hF59GTEzBMfvZaslKWUgbGY+ta7KZCn2
+2scFIYUhOLLKnrG5MbUcdrky7zfh8clsVDbR2h42PLmsxtUhmg+0w5ZMqmwkxKv5p0NQfsZjBqT
j5fD70LZIXNYUpb+9G87oDmibXIsluBWLFknuC2vXHvDmhnmc+anCV9qfHfQjzYcOjgU2m2lMAIp
4N6yaE4kRDQALc+PQKwoA20iMMzdiUXL+x7ccYCfborW+bQO+nfVQG0YJLMTRHm854ewVY3sHETq
MQkxZXiY+tmoL8iHhImlV0A4gH1hE49gSzxma8gIbHpD7Ji73UCXQC10LDinA532hlRZIrzStIi8
hBn2+7gP5eh3NdcwfyHzKIBfpnGm79sIKSW/xkn6ze/+u6s8KoRGxcXXD1VBMX0NATJg1lXKZ0Sz
7VSSmiO5Zieopcd2Uwom88LWpaMJySzKsiQ4GZ49oW97fBRLEb9iwuDmHEsFcPJ54CcIZaIx5Ymn
0d4zE7wl4EUYx+LzaEyLL73Wv3Y3uJ+Ibx4fA9EyIug2JPN/AVDPv/ewNNRlbbRsbfbWmTM8EUfm
ek6v664gcxS5K1jlbK8U5XlpbPIdsP2EeMD3q9V5tI4y2r+KIBU5MrMF4e+TpdWTLgrVLf5Ut8bk
SiqGlKz/KJbeAQ10RGXSdOwcDa4BDqtW400a9XP0RTel9xp5wRx3qm1vI8SEn8rPG5qNUAK2sRAG
5Nqmjx6pMeclqzNISMFiFYFuzT859wgTwkml8nIHb8nkmKgnrXtfUuP+LmgicuXL2i+w5v5zK7Bt
LyBJyW2t+wUXxHetqTO8DKfPfZex5/5BmRVh3tB9tZrk/MPMxtaVXddsv9N1BW+QpD1TGc9hh4S/
ARAen47ua+ig8KklAFq2dKjxNBXWtAS7HdoItlDaZdjpVNSBUnfTLKK5hUuZCyYyB80nLSx8TYrO
W7Y4lD55WQ8kt55gnxHM75d20O/bov0F1SmxES7y2btt2tmlzTFaPUGMgZOQM4Dx4J++KjxGzBdN
ecZxG3N6hm4sALeMVVOD9B9MY26Lku+slsENvivq3j+4DGFcRgL/q+G6wl/erD10+MPFx8cMTcaK
ODCTEwLK3/jmwyiOcqVcp5LyW+1agg6qNqCQJg05rVmvCalw1rS6pqCXbQ4zjDaTAPXqnSpiEGVI
EihOYsOy6CDwBYxUVB9io4Jauo+GI4NA8JoRH0hFUCI5GusxsRosMOXe84mFEiEuMqVRDvZGxTJU
RQ59dnVXFwwmL3TD5sRr+y+KjeAjJGy4IveSRiqzCwWQlXeT2rsODdt4tncbTM9Fy/VwCKgrn8DK
bZxYUlK1GVNIleT/uc0RKI8uiamE3ZKbRpynSalNTmjaEOkxwctpNaQPreBZpbHTiSK5oCeVZpCV
v+SRQi913EavpRKOW/eeiPoBqz2aPtV72u0wvDrnQhlTlAccB3sbO6oLO9JYIybOMQGph6N3Ews3
cgQlZKuru8EiLNMQ+pUTO7g5mAvshSYqkE3HbRjjSg8WxiNP+RZAafvjxjYGO1HYBBJtC6DOdlEd
Q0VG1TBGm0xd6j6VgdpKkkf4pUybyJ6LKCee9p0AaHyDni2ZiMqJTLJd4hLKi+G3j40SRc6+s3mp
WljMARSupslyDDr5gxySdjdxV7etRxSB8cKH1qOig0ziMuWfInb5UxEn+6scsRs/Z7p6qvJdmJlY
QOcu+v180dICAxH+eZDEof7auxgpxPPno+OmrGhXrPKSztwfBFIPDD9JMnbmWSFas35HJejORh3Q
7q2Cms1sYQYOgRWcvXRwXPV3ZCH9vvQzS5Jg3f1lBIdtBaJ/qF9tiFmqvYvztgqGs+lsny/7F6OU
eZXnpPDe539OSv1ShHODvGIwn7IWRnfaKN0yNqcfM3vaSS5mJs5CUip0IyPoEC0KePvwKaS2aMzH
gNDzuNbUvaHzijC1qVBWg3v5BGirD90pezcdR18TY8jIVoN6b9GRyKP8qBGn+OZTkH9rtZkdTgIU
HWMf/RZFaDSw8YQLWY9J5VoeT9ruKYErzpClrBAViMe6yj2cYfmZW/RiTDko4BJNxn/J+VNbW97F
ZbB41PH+fP/3lYPuKB6jdxaEWAjbqV5zLSM9/DgUoaqufSZRQoauZSM5kTl3SkiU4GCpQffJhb3o
XsIkjXbiqhoejU4s+fOAWF5hOnZSMOFhPFAxvP1mOQogBlc7ZNjoBtCaNt0Lbe+VR8jkeQkQGuxo
q1YVTPBWclFN1o0jW7FgNIbrR0xXHuIcjX1977pTGHQH2d+wQw5JbCzAj6UsQRL6bzGLqs/PadYj
BeuHBT6aOk2Ea3f2rKxEAUXSgRjiCD3G0UCH2w5841/KfqK+eTIKxZktapajaABcuOdblI6J3sMq
HAqWYW6At5uTW8siPzxOnbhi1+vr5OVJBQr9zqijjLO+AwHZc1HeRAykURSaiCS4RqsuzgcP9IJF
BaCHmmYf+CLNhtJDTFiTeQS4KACkoDNWhnmgJGmfCR1yTQs6yzejYAMWWK8T4DYc5XFRUXKXWa3u
3fIe/96yzMVHmxRDs+xJ+B+v23IRN7nWJIHZSdinjuHDDGj6eoyY5zF04i0b6DbCC2NUH/tKsSfl
N9CkZLlA5QCMo+bfJxJOLKloRdLnQYepd9BB0sDK25b5+eZOeGNp3ZN9S87eWd9T9AKek1UAQVDc
glTlykgLoFu3/beERAWOGEn1GpKD/gnV1OQ+G/M8SJNcANNYOadSFPlc0AmgiFxIBHqOixu0ra9F
RHPvliPp25v5m6o+vr4nefjcH9+LbrgJXnE6TW+4OD4v5bWYQQ2KNqjhmcULR1svnn78AmuCXkQX
JpDNEKrmInRj4lpYpCNTIyL2lGEjQL3I6BHMJdyqlWOi6oyGLYrdkIDw6FCCKXpIdzFtrx8p4V7r
W+/iRztz0AjoLhnk59tPB5BdQkgpYzm/ZZUc5M/biTbkCkxe+tq7+tQIqMCVbIdyiZaGDCl/aKZO
YqhILJKcsLLAN3lubA3B9KQWYkRZhqA9tB/pALo/gjcKbZ4pbvpNr8Am0tkTC9Zzq0uUOJfDdBBD
9gn7h3RJzq/QiA6pez3C5W0WJVrobwbZBBOt92frzfD/BGDjlQh2jSPpx1l7S8AARgUm/6kL2MBl
G8Eu8vaYU/uOkeptqsIszGbKb4/m5t07caf1DtQ4C/mQcp+tUc0iQ0BUaneqSBnfSXYSaFfELYMk
wEKG1nhhc/1eLBAtSXlBD6OQwlVzEaf7BmyEWByr+610PzaEmBjzAs203fFUoHfZGKC6/p7ihh/H
f1Xi3R1zzcylqXSV614l//wrZbuXYkoS+DLLkQeUr4qRac69DvLPJVkFRmbwvLIlok6lcUWlzUtB
40E/TE1Ma/QxaIzMy+Z+PH/tjeWNGzyJgFrN5Hg2GQ0Yw495Cv8eJP1QFdq2dkQumRjQhZsAkxUN
2BxjuALxXrDpOzQu50mTkAtDCCZC6InFYy9CrNJkyIE8TCKoIloInHM79VoFJOTKdRzrGoI9EEAJ
8n+IdA+qO4rZB/89yXnpPUW4Tui9z4KQ2CwoEaabauyXjWjxKLpmjeehbC/ZVOBemIW+WXo6+9iH
6sI01u+lMRdXC/W+hhUEqJtYV2fiklRHP70C0t7Z/0tDxfQ8ZwP37W0WEHeo1BG+Y9lN4xdRw9bq
zTo2WQYwELp2SHN0N9vqIlc/YNeLhcrSMAZDTuevpK/fBxjhifh4aRJeY63Zu8uhHdiK4cDy3pai
elwSSMuFrWCPcjzXgt5+bRroyc2zcdafVT3E1LFiIxF/0KSek3cc8Wg+bTVD9IjHTNgm9yxFWSuh
5g7RGr6zA6T4dLTXdaHKzo/rdHyX/m5NQVUqsd+xZe538dmokPuHv74IS951ln4n1MpnwCCaf3Xk
VABnyGBl+HdYY+Gff0OQoW2KaEILHPqy4+ohKRoj5xeHaTHLl+PxEjD8mg8cUPR+H5dQqBt2zVh8
Y2qdLlrAE6EI4G7BzSadqARpe+wU/sgeY28u1cDmuwkrBXrjzKLySgWG5M34EDs/hdb/+dRQaNco
VH1mZ5SOzZvcZP17xSv3ahwJZQbe2C4pq+G5TuFH1FZEwR5DRdEfR10g7Sx3unZzNWKJC4zxgijJ
DbAswKN5dI9qeOO1awrCBqvhDV/GtLSS3rnmbj/l0G+RcWffZbt82764lcpv2cnezF7VSVA44Qpi
f97f7SAqV1NLSByr3EEDUFJTnHw3qmJwTH4jP1DHGSi1CxWV6bnavsQHgC0RxMZ4FwM0OrAwDtTh
UUj7usah8ysGs3yvLVVyBHN1ioNVjFlmz7dzAVgN5/0SQ7E5qlHA/F1BAReSoja929xuQK7Mitfa
bbT+mn52sDYb0mqqFIwXihfbn5W0ufr3aMEvPigKYGBGGFOgQ5LqvnNuY+Z3/OeGtyfGQb+En8e5
Ea8cfvmtvSAsUf1KbP1O+OxNdmd9T+iE9CBDCRjceSQpFVVyeRTUH8NtFinXg72756KEXCglpdPf
hpngLmnX15XqZ5HNEtQa6QVVMHLiOQsGzbnWZbhCH+qt2s01Q6apYmQ9y0lbGJEJ7C5F0wmqd37e
6DRXBKBUjilqh1QKAFPwlnfrn3XfPzGpH5zxUmYC1txjsID0tyrSh/TjoJGT4r6zhVUcERP3YpCC
zeMN5z2fwnNqY6oIPWoKn54kourLvtRGFbBbuKkQaOaUX3LYzieNzTGzLAjrV0mcyy7qfuDPvy5E
4ssYtRlLX9UHpa3/XWQeWKK0t+mJ0/vh1R2QecixvlgCiQXH0TDTJeR93hgbIDeb5zGOpFtCjGE4
s6pzFm9eRxkeir0vuGoPx1CLaryVMWqPF2OdYFlpTmsppGuRKGdsFJBiXfxYs60IoMcEIyYus2OS
zWBgMoQQ8SvNROhJ3IdrKMiAFcYMLmXUj65Mfu8dLcPyKEUaIn8PWQ2V5HrEAts/WGqba/TKiqZZ
q2m5C4tpwCRgP78+yVWA3M8bzl0j3fvyxAfTctcaRld0qxmK6N2wWr8Tct3lbN6+l0RJdjxKWVO0
QIQHKqC3U1hNemiqM6YzuWI89lZ5JPDkHbHqf8Iz70iDdRdhOxfhQirlRzx+MuWROX+m82VupDzv
yjVD1RBmVEfoQkSHGJb+I4K8AeOotHNER7RAX5DJ+TZO+8X2Mr/W3VCIov1Suxgxiwn59f8zXzaZ
02TV7jRok9kQi8ttYnQWjhZc7gfh/9m5gu5dHrXCEVtStMi/CPw6vcL2ppHNP4egY/tXiu//mYsF
YlprtcJ5mcA/5FhAOqVTAknLm8WZN55+47ObLvB/gWmZP096v0uZCs2l2VO3+0zdA36hch5PPpab
TPlsKepFHBLszCXQM1nQ8Pc0KhloHS0sr7tafQ2MRtGadiityL3B2d2J3ctQ9xn7L2u+AVaGwEVM
SeRISquaVmYftLj/G/skOpS/2kESzIHI/UdsrZAMGb+k0OYEP6QSYY9VOKrbNyR0lB6BCGOpCYjr
Fz+Wrs7ZlGsfdWYl1eiYFvEioA2/OijsMklnYumvRfiAJmwTufRytFFIq5yPe8keyC9sHxP+zyqo
gPEm9yrda4QuNXalDXjaa26Hfv0iHIqFTHsiGfn0f33qqx05EgHV00EeA9qxQAzStHXh03lnAlYn
PsbIa3zrJuVzVpMaMTe7Rev1X3rxehL22sB1tF4C+IVPpe19ipwtViqaZ8Gu4guMlCuR3rDQa9fp
0Ires85moZIGvK55H+aUaXXBZSGL9Bgs/R0xKOkrg5QIu7oR3jmY4wzSAdmZJL/HTk+O5YsNb363
54V9tZlaeviMu49jT/LvyxZU3YbF0ueJn+lJGB8OkxTEC5am2PatNFicVvXf6v28/jpmrTIsTXM0
BZ/2fQGgja/kX0SA9yh9n2YmLPWuFDDrGnwYCVKAEgVPPi6QBF3uSL6j4WWwNtB6AGOfFurvmpOV
6dk1cX4nyFWUoRehHq5R1AxN4K4zVvoJvPQEe9uaujcV75/cdItdP9i5R3HqFFghuwEnV29jK+xo
a2ugQ9gqChmiR+Y+y00pzEdp502FuN5bILZjeQm7jyPNzw8G3KcY1WxUQAO5viPzob1yrVazyodK
D9+9thN62yTcmy4cEHg+g2mh9C3/WMYAdaeHoBoWB5ssFhErK2FbTpr6bJJsHtmCkgNb6cmqhlCn
4N/0hT4epNDQxs4yZQqSx+RAK1e1A0ZHIvi1XrjNaBRmiwyn17PLsB7vQ/bOkiTeWBC/p6cKgwvX
YhvMn0z5530N1G4RpBJo10ThLmTxcAdOLxX77JKMhm4a2MWizjUiKkXZPNyCteLq8+C+jhdfHgfn
ToKYCNYMM1KB+pgLh4SSyfS/yoXPya2Jl4NU6EyhPtrrvfK+QSdNMbQRZjVFkUl+YzP9fqQiAg/3
W0vzE8U6aCC7YJHzs/nqgvoPhZonXVH1HmasdWcf40rA2ZfTv1a1ads6bL5O9U4J3O+faQtTzWxv
W14Cww0Ct499c3VEfdd+7I7ktT9TOKhsgo19RCYJuP1AgwonXxj869slf0NvS7R6gYnDOmG0rdbD
gn7G4wCtS5WIysHHoXDF/zTWDkMVqbv/1T060o+OoM2n8RIKae/P2bXYcSEFsS0Slb7YAfQM8EOQ
xf0iATXeI0aJq1PMl6SuEMVYbx9c2NQZLKeUiSY03fGXmfj10/ogFA+riY2I7Hh8eQaQ/zh5Dwxu
ia2SWcWqqGrjKtB+I88pwluKGl+y8gh23m9Hk7jaScRlefzUVwnPnvuGrdlPlQ8AkhdT1ajdm6QI
Dj94IWLnzR4PPo49KFljfp6KKRFNXah0Ww09HXI+f2RIXe0/ynopLcqKX9iFewtQJMEOLot0xuev
qLedfHm41NfMujxOLDMTxpuF9j7HarJwueI5Yr9RCGBCFoeVhbFogVPrx67EGfhnAX2iG3VGcnbW
ioRxmBbeud/8knWIsKbStPZ8EpoQGh3X2I2wD0rm2kJsvGrHNVfdmLtWpCY45Y6rxbO/hcTB5JAR
rIC3UMNbVXgX3J/a1UnzA84NfYzHVMXjDKWyWGfLV8bNB9aj2EJbLaz/Y0vGjtpBwFAjFfTHzOtU
00o31WUUvWyibVNsAkgm6LJqxvRZHJiItiTUUf5rKCLsumoVxJerbR152Fps7cJAFZbGRlfwEu4p
fdaU4SuKEcdllQ86n7AA/6vt5kSwErMkwH0h3aIFyZxkKZhgOfHY60o7/uD17uJJfBPfW+lQNXJX
aFJurV2Z/DXVnHn8UDhy6Q1KpsiFO6Uix2YDgWECto4f+kt/In6u+8AqYocaThYTn9/42PU1zCHM
vpWD15V9zNKEmCbOEOXdt2MUA0LmvP0GszFH2LjLFJ29fz4yyaqP1cK6ZbNCynOM+Y5LHRmVK6gY
6Galqcrb44++LE21OX8wF0rzWrhYHIXrmahFfQa0O6M2x5b4Ezd6CE4yR5P9Ia7IEFJgU8+5hF18
VgVQ4xdp380Gl+v3k2YtpzFhLOJTjT7QG5LcIkpwffLKONSYeZoiRi22CrM7qFUGlZUtZkmd5Psc
5awaUFq6TbTYchye7eCetdJmwP+dXyPv8/mWiIbwcM+rEqC5vJhGCzhl+6ah9RZcejPabKEBjW5i
YskCc0/5ltw71yESrWqnKqR4S918vTDxVc9KGG4u62ugIoze0YB86BOiqPpEg0wF+zjdD55JsVvi
rPQf4hw6NFrmhI4HdiQyXjJVWCEyeviO7BDmNoL/udkExShsp/BnDsPBDq/NaUabOOfOsR/8xwFa
1tGNSIB//DtSdmLWJAXXmAKu0gUr2qw896QDpbSa9W9n9HRrQqd7qkneFNoO+QeJuoNSb/HOR2hn
qlyYQH1HA6IXDXzwWDVBN9o59czEPKSJHCl2y+AGTsZ7E78CT+xvb/1HZATEkLBNzA+1EXUVyW0f
fxPdCf+L+1K8U4/zoe0MmKfsiXeOUmBAbRO7/ruslSD56NjxlxH+t0CvfYU2xONUvBI3A35JNqF+
VBbEV/HbJmasnP/DehBTlI3mFjKd4dbGAMULvBTUIiWoKNXI2fooxHhVVYxqe7CmcmhxmYC7BH1g
0I1eLjpGwNGtB1eHiBIefS/ZnZs6Oh0aWzDEMlV2gKg5nzIJVUif7ch3P5S3W0Aycn33TC+ilqaw
mehBhbe1HWKJ9DSor8DKPs3OvlEdLaNu5ynQveoMgw4SU65F08/xdA2mYr4LGwXxvy92bl8Ihd3l
gZu0OuDunif7zF21tBzj+oOQGgwvD5BiEPG01GwEoMkWWIzcpIajhUKVeUr7Xds8gsKC+QBEFMJN
fwDqg75La0qJ1r4ekMcda8Hrq5JkfDOgvKhpFZ7/O5q0mr/XZUANzaBCuTORm/Ksx6Cc9tzmdw9p
b272CkTE+0cJYr1q7MtY8GlDfNA2I+EFLFweVMv8NrSrAQZ3Nh66nEzxLONS5KuxIFL4CJ9vK9Zy
0ori9D8WeLMT4lukVuAUKQOvAFOlcmYAPFM1OuQCSxFznbN+UI1GrgRy3OyOjZp1DreNKrWhuSO4
HDyvZ9nC8N0BaVM4XayRM1mMXQ1ISthhZSvq9D5jYHDccW2xM6Cb9ns3i6ClotY33F42G8wz5GzO
x38NJWJjhFWBfuEWxU4mQvUxslPe3rc7+MSZPWKbO0JplabCrHEztgfszU0BrU577PsGUUNWmEEq
zkER6lnBKnwrtU9IZJPKy3vgL/gU2EKg3s4EcsfhXbFLq8AXQY2krHhqeLq/ououJjEgi4+SxOGq
W1aMzgKdqiB08kL5pQGJGaOEKwTXW9d3f98mxDAy/saWMPBVn6ITvHfLd73p6Eahlsdgmgh7+gSx
mcr6S7RO31p+dRfB8mt1fMTWEWjD/EsoupoK8s3Wg61ISx9x7OlVh5qDT/ZnoDOng/pmK3Wdq3Bq
nBr+kgvdvEzEunvl/wRUhIO/++n23JjSW9SI2bLwcwVF99w0JzF5yRAGfGKf/SBfXt49h+/YP15B
bos/6WLAJmipH2Dv1o/i2SK9kuTNhs+vlULnqRORaR7fE9HoI7M9bxMEOWiPaQEcAd2QAp4+AzM9
apcjORTCAOrxpHv1GumhX02UH6bB/Wf5UYUMC/d02oRyR6NPRFvoZBJgCq63mGTCFHyt+JVqLIBP
Do1jvTbp9VjPxezV0tAJb7LyvfJorVuhyipHc7Kab89tE/wV+nHZeWYbtwQLBmQCOwgWQiUraGAB
FhpPP7dmg9fQBG4ooe9Z4MQI6pEDGOHXlPTMdDYmSqARkzSgtmHtb3qNda834dSMZR2yjnETkYac
Ok80C7iXRfGJrk1Cce6yR9W1zSLnq4iTXqdclhw80AbjGEr2lWpivCvibWZEQOlFi0fuRDFEe3Tu
jo9ngq+veYBTON6XD+xMNq7RAelNHQqap/OaQ6FTdpStxdbSqgz/ksFUpHFEYhyG/j2ygvJyW0D1
ll1OshPFKDfyVq1xGxs96Ol20B8NMTSif8CHQ4MkIHEVHKL8aJfmKFzM5x67+I1lkPoBU5DoRIKE
bIs3BQMVNizwHUnNNGSoCHZmp7QzmtoEeWKlePEH43mlwKyHD3+deyyHFUi8IvqTHC/2GGQnOpWU
GZrrB/TgmxPg9Mpx9o56yYBwgnecVkxCBFMLxzT464xMz4M+39E98yM2s+0oLxbhZEyx2CO1HTH+
SutQo1qfyjE24r3raqX4jd18BOJqM2ec53dv3rDZK/PzYC4bKUVzR2O3T7NwpeL2jPSYzhL4BVJY
DcovQqrU7qm06e1XqtGvP3UGlZ1WkxylaREg7pcY6QAbffHL0Q/SJ5I7QLINOhuLRft2T+Y+dJ5v
XXDG85EoEhGwrnZPz6grQIqKbXGFwC619lqGvGYjkAHaaH26EXhzRq4YdGpLmKBCgTauh8uGu0TN
AvlAI72dr0mBtJoI8YJa5X3vH6ata7eCWvEYXfuun+2H4CEElf66vwuG+VPyMwYyCIx1h/VeDza+
y6kwMSQr7+TfdfC/h8hqnulrbak3V7ludQ/QJcfKvrqRq+r4Nt2LR9OL6XCNu8nlYQwP8IdpmPZL
KB1OSTBU99co3S+VnZ7xbGz27gbP/wy7afk1+DH5nO+7QdOoeHKA44yR25ZydYT0eZChiFjbqdct
VEKptkHIY3Nba07s1dA7Ch3Du2vWhl5guYlSMZvf91yTmOBiEY3qBGhd3I+fThvUtltc6xT3uKO2
OlQKxKeGuI12WUj+uUVLu1kJaDutfBNcexecCJdQlSi9vukIu6prULot6HjfiYMYKJ3BCmNNBLr5
gAOhyb64fN0SquzouxsNNz6naouliOsMS2x6HUhW476b1H9wcn3ROU/I0QmVFeMscSU0RwLwe9kY
w0/H68a6MFdSVLz7+kSsXDl+ddHC40Pjgi1Gkv/CXW/QKQ23pXGQC94NyI6Sc3KDgeNAwsO4UVhH
tgmlPArbbWOEbN1t24Pn40vG9mZinUirnbOT1N01PbGMRc8s4YCIrKQ5I21XbOkYzkJryrGLm9yx
e+cEfkRUHowrdMDwFzak+t1p2Ox+d8qvbRG+kifjRxyPSzo88UZUsSPscb3/uJD7eq5t5BLq/TaD
yDpQ8ypf2EJkb3dPjXEFC+RlR3aoRmNUjX53eBDJ0zQdmcOvenMB+y9BMthMFLsMjIOQ6WuCuLmJ
zNVQ6SqmNdokwiEYfCGEXGpIeeDKRKiHBZibRF13AxkIAqK2ZiC98g4La2i3M/9O7HhWnaAPa4Zy
OamvnmnCSRtRZiNowmbPTB+xoewwaiIgLLLvThLmx4s6xsBxyckjRjpFJ1+YCxRrbUN0hKef81a0
OrOwZiiftItYpPuooMqe6fxZlKDASVZIIyZhVyk67fY84OiqEx1je6m2ODMiKC8+u07QPUzy0Tp1
AytoM28TWzdWsMyRn8eLDU/b2FDcMhCzeA6f33cLg28LIef2BLiouGhpcyvZkU7n8DHjE28srOXy
vs+pxrLbsTMykiRstUGq/uK/zXwTx5ZRjE0PByFLtfQYWKBL8BH4If0pMmzX3zzWjJW3nOCDuB/r
p9EECK7nd+nRXRsZ0rdXs/zTfzhM46jOPIj+fMGM/35GsJw0LqAmcg1y3fQg4sFTWuj/2xch6HHf
vnIh7LgqKixGRi2vhMRg6fH1aFGQeGgrDeh3LhYEHcpClOOsfSPyTP44toHOrLL2+XZncBAs6mWL
YMp3LalKE9FJpgExIT2fASHCJoYlk9HEogtaAlK/fybtnEPKtdeDwqaXFslrBAcc15qDb94MX8Ih
aOcOUeSLxz2SBjx6C0j5HVP28XHJNfo7RaimwCvOquUKiGUDhpD1xcibJqSRbrF5XJ2uiQkOZiM5
SIImscMXO4u2t7gUq/IGFoKIE93MGtk3/0GOqqQbZS64bgcaQXq9meqN/nUlGkSNxbqaKSRpFLfy
M8+OTCyusiBUv2Rfomh27eM2DLCuY2rHWpxhvar8zbDHY6x6jeQdUT3JQoUfP1Bg3awpb80K7YNL
RNyIQeFpuvN7EVHspGrRVMqhqVKXM0D4diBsP+HQTzxAIfJv2rxd0B/LaqSHGnvTrHL34w9VhQzr
A2UsBCxFDQNwxvaDUiivaKv4kYSrrVNAEnxqFwp0aUvJo1Hqhs5XmhKHf9Idn5CX32p2UIVEUqrh
+VKIKIyx7DRRnRKMrBmYXkbgjU69HEdbiLEl1Ac4NYpW7gsDpkKEvpyqKCwkMf42KGCgGFK9A4G4
TPQGauvKnmxDSPgsFEBj8TEw+jUtXERfGtfkDX15CtO6J86ggs8vzxD5eQWqAeYae3hv0EwMxqqO
WVAFPjBtz4mo4SXZ2lp7mI4vR2PfBDQsUzcZfYpHppxAtz4Zg5tACw6fLebmcd+JYmu5C8ZBjCc8
2/2HHDSbEV99x5iQoHNSVx6N8fqR0MHAQ/+TrTcy1oo/8jYqih7nAMyxc4V/A5a12tpbYlqys9jV
PdIPjAv0kAT6ePj3fGBJ/rhwTN6KhqpatNEuHa6qVk7Qvr/wHJbF1pMkaiVWjaKmiUXqOMQVqZ7D
LkQSKMxuWqIYrRrF87UxLRDpXM9/HR45TzdTujILZ2/P9nRnPTAi0J0biqKhjbS/h5n7k0xt22ZI
9o1nmI0Cdc4XIkGu/UtZwosNO8bEfkLau9WwGoGswGbvGGvzyUlujAAbgHWcRMKU3zHdchQddaT3
pYKovYqfvXaZs47dWEFM1YI1LABHd6Usphh+jJ/NxMvqfniVVRsSVvn2ZVen14o8Lbl8cbSKGr0L
3gEC3HZiqidvSVjtnDlzvXTslvMA7YkMmlws8c3165f0oxCoDqam/QiPZ86EGzyg0IMdHa/7KtjA
ZzGi5D/Pn8WFg6eQZxnMCbsxUgtlZdJWfu+/BRWobdybabA6ClXv+1FC5X5j5V8dPIo08Ur7Q+EI
Vzgw3FCeWnXXClTGmypiNVlkG9a1+848cL/rqOCIEUW6Sf8woKGtzJ+VEBnnPQzTYfJPKXhvGDfs
xefD0WVGvA0J1Oej1P130JPthIL7ump5SPNc4vb76TTnIZN0qex6Dey6WJafsnDhuHsV4JBrCmFS
KBmC39kE08rvR7ldZnUdvwVr5iGzw5WK5GqF18zSW3XUIRF4BcCBYDi8nMknixBOeYuilFlfF2tb
35FLR325vJ4lvIQMMEopM5sFtZVt9QYY26ytOEX3WDbpNVM8n9p1OBJqQ8G/etRujHqoFxye/jnG
z0jxwFQeynXsVadY39gDfjgJg1tBhPlGtUowoS32uUnVbi8weZQHm5WzALKzt8XwCjrmGKUrTbcx
e/8rToQIC46wnazYK6P+nhP5wEe3QmkKQ3IsHqpS4RsgHvEIPKMQh0eBo0WXTocZbcDd/jZdVaOL
v2SpAAKswnALD1iN4ZhhEHwhCItg2U6cPkGwoSYfeXCQQ7FcEf4hxb0cLh9heaAsjUrlD1J1Q4mQ
v1lHhY2IsUPG39ZIjnVAyiCg2e6IEX2zEqvlyec+YM7zoucbBIV01Ymyp9Rzi+jWwiRsuoa+u9RX
HH/VWj0zPAfdYRim3gHLyiQX4+p6Nl4zrtx0MXhLb6qER1ChGZfsjcdBwFhkI3J7oJPBEOWkMlMC
T5+lEBWDltJLTnRqSH/3RmimRIWr1edJqvkF5ul84OTA7pdlS7Q5kZICRGuNNvchXgC6PBrMMp6A
DVMrEuEaIhHc6U2kuYBTUJzf86BpWQps9aTPOlQEK2mBSSLUiakzzmH01VTvW8SGQ/Qwf3nMVte3
fgxXFOwNdUbKPAelW5uGskY3DbIFuRG8oVyVyKORNOj8wUCxvAy9N23FcG7PQCBCrWIM3TJZ3Ftg
gJY49t8rQNZh+L3UAzT+b6UzDVCz9uGp+eUlWYea36Vmri05o2yOnexVkCUlU0+AEtbB0mGXL8LM
ei858ICX8O2rQ98IeshATsK3HevpCJNQKjhmJvC26yIgh193FRXe0E+wOTULL3umROVUM8QASPRS
mtZ1WAs5LjN/yTLcv3FYTf7D/kpcgtZr/3YOCsI5rkm2AKRn5gNjMZUvxD+24uHmXQdSR1pGfjGH
US1AMOS1UjzWHXUEPTOoNcH/0mmhcYj3ZofUQUcPT9lrM1LhwoqLrN+d3XXFvHffQfIJJgu+HFJs
qO1yqr+vgASB1yt8SkyxxuoJXg3MjD3uZ/EitH0Bxkf6x7Ny6puesRvhxjv2f2yhD5MWrclxQ9JZ
sWX+cWjarypcu0DDIuLXj4Um3EvJCELl2qfC5Q81793k1y8UftOdLSGJ3QIo/UTAqBEbDRQw3+AU
sP5G/8zqv0wAiZOlKGIdO5xPGC9LFpaZJ4fPXPe2eq9Tvj0Sj+QmtL6Tkxx2QEa8fd9VdArUZcF/
d1fzIdBfU/G7B0mBni9kij4npInmIdfahAWrqIejZPRG+DJgZ4v3GRVswMfPky3xaphLq+Y79veV
l4l6qx+YDvEeW75SpIVM2blVI3fWL9husgwJFfsfifoqXlILdscYGkw8d0AjU6U5g2GiapZ9SJ4Y
Fp5logYsbtGGAasoQ9AhxOK1RjA750vcxHmnLaX7Nwl+eLCHPaKyUShCClsP/OcYsvauoUOcvsXb
aYfZNMW8f386Zv0js5qWLjD9O2m9b/JOI4Y5JKMHIogt99G0S4wB5y0RINml7GV+Zgv1dZEYA0jC
/tafwTSuDbsLVNK4SmNNAB1isRsF/CWlkpRxpoWAUyqdr8p3rnl6MBgNg4dY5lL17MWBzWHeqpF7
b73ZdncagIJjen4x6yABM0ZUUY/u3S8dZdnbCYr1zLlnB4GoWivBfiRH7g0ySz+doQzg04enC58J
Q5100u+jkAnMnXoefhWq+LgLCyYYB+F75QOyLHJPp6dyhYCUPubcaYUIj8q/mkS7iIQig+lpW5qw
TIMCNjYM1syxizPH8rMWi9TK05JVDyq8Rwrwdhz2IKLOVf7K36LlMs7clbtPxLDO2EFDMoa1nmqI
tCBN4bOQXpv1bpYoy3/kDVf7CHhrLWMh84EDDMotMcn7vlR1/x7zkyaLYb8MyKCavU44Nv5w+Hin
STRdn6RI2K3Hcc65cRTpvVRVbFZznuCHRERZe/6vQmy5BEhMFIU1vov6GVXNoegsivoQIGpavFMX
+D/5kslJZJaSIhmY1vWvzz+FAisDmG2kYj2KRVsyDdX7Y+9LuZzBdy4qYffL/pF2x4oPgI7gvU8R
VcBxW9F3wrjOtRgdapIp5pBtKTbKLGfpV9+DSKomnpzpxSHbChwAY2CHa1OxKY+ZcPGJ9aThfsY2
9FH3zI4EPvgwYu7yiRo7Vp8OsrOrI+IWacv+gi3IFGlrwY7YjOLh5Cjbl/wvJjUom/kcA3YfxnJA
a5Yt4c+BlmTvOgPoLJSDUHK3xxiZzi2vsIMcu9IKRaas2ZlNHj99zBR1OSWgdUkfcJVbD3MIIsad
HViRv14JzuljvGJ5gphK0J0AxGcBO80hvy5KsazoErA3QYIinfu/PfD0htUI9l8EoMTAtj6KiiGu
T8ctIPRdkN0nq0aRSietmOVvgwbONUqKkOhPuoOBDYxRdTaq2xU+rFFAdz8gNr2/oPTliRUiskAR
ZFO7W15R7dq0ZNMPKdmqkD8314Dr005lJtstihj2f7+NdMdJl/72bKrjeZfZk+MtVUYpQE4NKjt/
3UO47ac4VN2oXsj+EOGugi37Bb9HitPHEtb5OYmTbIg4Lrr+rPz9feoMazZmOyYcgZDCSO9ygAU5
p+OW1McaXHNd0EVEg44Ps4ptZkRBfMXAxojz8tEdAZH8Opavb1s4vpGeD1QR5YY9abdFUBRzNCrJ
UcpgR9HDXNmmvJv13dH583h9TLTBqOi82e9G/JxGmc0L3zE4R7tv1Vu7ndh4tMHg7ebIPTYDfQb0
Yt7mSDZvYt2LeGYZdsZ0J5YAuFqowOnyV6KVaY1HT4DQqSyMhMPcXlu0DnJ5bMUP8CzrBIua5QVB
cbBThZ2biekhq1nlhTD8/PiYOc7NSpFVUxzO8V57lRZzAlM5SVy/7jQATTnb8mEbJwOxX9fVx0N2
leNGzUpdj4pK8+Sssh3rRyJClMh566O4iZwJaCAM2Jgl37aHrqYgXIMphyvlIFcxdS957K0nUjQU
s4PN3/fdmWD+85mdIt8Ck0NE3+cvUEBLW0Vx3vHFBM5QUqyqF64xeakUgeuaPXmcmyw5elQthVBG
XBrW2tTpNQaf6KDYU7oT6X5FiHC318zCMyYJ7nbNheBxocIyS4FR6WxPhkYwB8EpXxeXZfsLDFj9
0gnwMnaTEGgj0eyimbZjEE0AEgES74OBMnSY03E9Au96d3dg2em8HdOHc5RL35frOHc7vcFFJgpA
9UoX276rWxkkUHMNo9tBOBDHF63tZQLnfbyYltzlyyOa8uQWGDdj6/pqIlbADH4mgmnTHgPRq9Ru
0shvXKbKdijSGDdmNENGrWXEC65zKnk2qj2g0j69x/2GiXo0lQtgEcntVRiUti9GefzmtyANoB3f
VkXtlJsxLvJTRMiJzCnBkuJnPvXLAvoxVLCr4kd5MYyNowG613558s205DdtHAcGpbkBOaRxQcY+
/aYUP5Kifx2v3LNcMI0gSSWEbIpzxmjXzahNnVli8MLrPu0Mld0mG6xqgtf2FhbnQ8LjZU26XTN6
APVQrT9sMYixbW/xyq73U1CjOiuflD6jR6XhAUTpJCQbUJRlWbQaorjWgJI0o7zWuBjUY1WMKalJ
zqKzqtE7IzbNBb7CrOnMNhGxQVtPHfUy9JJzZ5lXi/TYjHoYMCop2kHUPShZ7l4d7mR6mKwc9MRX
uVsr+iUFIMys+rqctiWB3Rz2bSCOODPnRFjbtsTrGnMjlWRfqybVtTHYl0aCv0Wi6fFr+/E6i1XI
gDrlsKyFvS6irkifqRytMWFNDi61zrkxV2cXMfTkfNDxaSMQ6Y0x7Qt3gRXtVv0k5a3fS2IuwkUB
uu8gCyNvfAZrLBHUuN3BAkD6Vsygg9jtKBkYVIv+bmnzFt21tXxlAmO1Z3bJfPvrI/77NOLYEsVk
w6owVOAqYkTHhgR/zXVogG3mCVC5/8dLkg+I/CEM+/xTp8bWHXGOcxKYQLGIwDz7/7cMHj6mPvze
TnakiWo5YmQLPtJlwRiuY84i7oiKBbUiMzE2DJEi0BClefHXsniCY0/lr/dDzo8ETbfD+oHKIwZR
O3f+oyXeLOFjqmJhwB2ls3JHiSDPB0pQjDXweGOfRflaXiAweEno2+flolJc79mDxLJj2+rHiNZK
/Hb1WmQzElysXengKpXUh2spArOePezRGbTgrgtVvloimpnrGAZ/T4lPg3IdY1A6R9iwdaitMcKg
XNkrU4nilEMVTJLiei0Aks3K0bzk1Xz4TucWO0bC715sMU8moiASR0oTSFZHzxKtgPyDpL1/SE3F
vZvdaSwpFW5xt4jCfdeegU7/6dBwVfEZCZGp7jyeJNYj6TBsmnsIWXMiojFG8x67bCTGdvGCqIgO
PAa5uVUPOIYuK5cVB0OfXsexHMyxU7L4g7f5p/aifmjnc5rSSpyUdx3dqmMU/ybN6It7CU20rjsW
NY85McKGj+/I2kq4OPsZv4M8snJnn9EFDByoRuu3GEJimC1lwuHYWZ9O/VM/2DPBZrGAGS8//+Tg
lAQCItnOzPv5JAAp56CMAdvdFK6Rah/elJuJTjmFKsQCFN3eAu4Wq/tY35OVoHbOF6UzCAU10Zim
kk2L+pKpQUvqYhwncn77L2uUdjnn3rKfdTEVqpcx8U9Y8mvHNDiBNUZg68uGlCmHzZonxMSfzCLP
Jks2AcSgcLjopbemorym8VidvNXw0bK0dinLA79nlv4NxHVQslWhJ6gSXukrudMqf+L3cr8H/beD
qO9vRjBak3jZGrZb+AUSY/QMFeU1rpQYSyRBsxdsk+59CJ61GgE1gKfCUEo1PhmdI7+oTY3w1bbi
6bAu6x5KP+4Na+R83cWVGke1BDD7K7OF9vWZeR7MDTH+nvEnNO1yDEQO/Fl1PPWlF53+vXVMXc4d
lPqFS1tPGuXqohDS5eIFzBQx6p3eG64NuUUGHC8YgDCpO68rSP2xsb4umtjmm1ZZWKVdNe3ptVp5
ID4saYAOvoqnfYlErorA0aSS1S0NCanf76db8Z53Gefjw3kV9T30NKL6bF0YiEyuO/TwCo2YR+tK
pku/E234TkMwQCvRh9eh4VeweA4fFOwTa0FWp4tSklL13L6Dk2BG1UHPsPNKFKZQtoiacASf6Kzv
d9Os2GE/Cp1urVE2+KaZnMAYerAN733TP+b169DmtZGumuELfkcKxOTi7RK4fHT4Jq0s2Hx58wAF
xAckQthM4FvU/b2zXD0cqflMpQyWnN8Eez5jPjo86NI4+9LzrfKfa7XkVGj/iHG34b6HWt/sR8Oj
NFswmlpobEGEf7FfJw21Yl8MWGfbmNjQ0bG57VrVm4tPrEW9j6QaCsINrbKq28oENGMfQIlaHWrn
j0BBDNYnqjkGBziNfuFyLpwHRUYnbZVlzF9sfB+XR2T7tRUUMkBnOekjYL4/ob11KYKZ4L1mG+7p
jb7KOBj3bBC6fHHgrlxHtIe23em3WOSFbLUeG9pMBAuEfEhxcImofZ427qCRMj275X2N2zgBYaki
W6N5AlaDvX8vpyNyYzs+t7DrlU41lhtYEIL3rmpUEJ9T7PmKAEJLhqXVEzRQOrrG03A7qLnSCRHD
ck4gz6d4uVUv0nDgYOsAl3XWA1DK/PXwCLnwy8sQbJ1wIpRJPd390ow16VqTk3jNmxXQAUmhbaOr
41AciI+bRRA3/XRptq5g0Qh7JGETC286/RFRXAW/piKLnnwVWHt/WmsUyiiuF7dQWUEBpCn5vDjp
yNQd98JaqrTpN62lKGdM4OBU7GFXzFEyOQjjPVXvoZy4KhJOqgeauqh1jJAWxpUR5/DQuHpDP59M
z//38lt1WfnRGV3gX1zSyZJotb+V/0yk+O3ffWeaK5sfwCx3n3ksXtEJBTp0tNwqF4gizkAbDubW
lpDwNgBESvvpxXUtzNBR/i3BgjumBYVRad+sor8rvMbjSf+qtnVKlrKqClUBi6UQKutlNfEqYrWt
GywYqSh2aNW7RYMm6uYwBzVAAaZ0h5Q/nD91fXxIj4Eao4144BUjX2TwxjHIHFCwD23gAyXYNgdU
W/FOVYCThjmDNWg+Eul99mEwivx7FF58k4jX42M0skjIxFb7kFPri3DuZLT1pgGqwdQeHko1ius4
42r/ENfsxStNJLjfGP+24NBA8XCYGZdmUkUu7YW5bmUXoShsC9VJ2glMkiDQUQmGNTnPRq0+FhxM
+6xwFxGzp9rdh/dCC9NkESzePJljjKLEqmnu8HVSrd5HBhJqRm0j1izYbdR1ktbbt/ORSHan9ZEJ
POaQwEIBiAxl5ss7YTrZGSRLI5ibaq+qiEKl/md9Rg+D2NyhkhWYLbYnjUmxniC+RbxodI04+o5n
bw757lJh3rMBr1IjbCTIXDf3/Cm138Jfdk96tMoDLm5KTUKm5wNdITE2xp4qWJx0O7Kkqb3TJtbX
uR8Fylm200B8Trww+rkSCloXZHiwTQoxosH5sVoiwRRNEU5IIeSuOzpmTSE84QZrjemXc8j8KWVK
euHt7SR8m8i6ocF71JaS2Ys5oGFQ8azSCes6F/XcKzbHgmGTqMKHaZKB1EZIjSmqG7fVKscvTvHg
N4cRiuYpBN1pVV7GgYJd7/VkLjl1HkqJytmrt1PgXiHRZZUgbjAC0KCZF5imLUqdxGE78pH9G2uW
t6mTiGUpa04Q0+fXKG5mDj/kKrc9t+SvdAPUjC3bbG2uj6U1lxISI8jBHcKj3yoLiD26TqjIx4Q4
oP+n6Q3yxR6ArW0z/jJu3lYefFJZHDs5T040H8ZR5RL5blX9o/iN3ryho8eQbc2vQqv6tCf8xOrr
wKHc6Fm7MbZf2+ro6jrxRq3ktj6vLkUhSyz+oQ1Khl/K+gzCLXdNPUCV9x/Ak+jdk7gn9w+lK5rD
We6UJwvCzVc/wpatnWdyGvwROa2WLbwCZod9QzqbGOE/3+EtMoLMNCHpNim0160QEede0jNNGWoO
n/52KEw4xAicKXFfI/jR+wfZEta2QLg1+ZNJgCb/jqS7HaBHKGxMisVyBeG/psuISvXEo08RwAkw
N5sY83IjjV1flk1FITmHOV8YVWuL32/5DkBYX7gZFvUEC+Cx/LbZOtDcp3jd/LW5C9AOSDtgeIxj
AmkrPdcVZCYoCll5A7SHRTYnqVHx2OjiSTtsr6+Ng57PzuoQYYUquAiIJSEv70joHo9F4KnUK9Pg
3rs3bwZFFlBXrOrRlHBGCvqtNQ3v4olOgbZ+K4WgZiy8wZnhC9UPRCJA2YJL8Lw2q6Jd7Xwl87UG
6yataqCCLEO+mFAPoTVcMDW7T8aW5c34mqCf5BRrWN0W5holYoCzAugKoGmsdJQ0AoYIYpagzgUD
Pc5pfQ8vBYqQ5RZCgip8oTBp8jML28fAVKXHTmCz+nPivev0BJIPTnmj3ityjYdp0v4IPpQYP0HN
2Sz+pGj0X2UE/dLSRNc59CyqosX4XJQRrad8m235iE3YsllZ+CuY/qpiWUU3ey3Or3zTS5diX/Go
Y79q13WhZTdjtGfZOE6oj2E+owYQaqrhXizyVRfDdl50IqQZpqNu+I9cgN5nCWKRY3kgUa6zJwCu
r2qFOWdKwV+23+KuC7Hd6F47mnt7YIGFW3CNXx5D0VIpbImv+9POBRA6NafZt4w/5M4SoHVwyknd
7R4gegHvC1rw97nn792cdtItineU12+p3uOryl1uvHF/SIgxhenWGxTpkiKaJ5nmtOpe6DYAYEwM
xA1a+Vka6ulBem1S/EopP2G89Ghl1OGqkL9opXu0ZR6VYzWP69LEF8BZvEuE4hvFoOhJ6vRVuF/G
gihEimBTbEWivn9Y6INZvgIvL+MwKeXKd4StSnhbmiFPTeMgwGuWQLW4CLQjrkIyVzyxd/ivpxl4
gmTpZlM71Frq76UDF/vLC40RcQZ/dl5DkXPEuhht/1oyfsjeT5sZyOs2wGFcQ6eGQUcbdCL/s1RX
JWhPDziG5PaVL1FRK4qBTbP2YDdfY7roy49RV88aTx0uDNQe+yiCdMQPseZ48aKr68p3VhWuMAtj
MPL8vFQ/VO/FaqHxC9y43fnlTM29kwgg8FHn3ScKZU+GCsWPrrhb7A+jF+c1qjhrnmlZOYcTgOT7
Ofph+/gpmwK1RJK7EUGZFnVznmj4DJDQxnkYI5B8+uzLaK0bFzYNqedih00o+mnL0cKaJ9Noyr8d
C8IlcXA8S+YujV0aabV+rmjDRguc+RppS/6oJcnK7xDbLZAUav145aMBbprJZaYNegsozUIeN1xp
9yss6VOE1GBx2YQhbCtfppA7ekiWrz98gjek9miJ9PelATNqPARxhOmSaQea7NEMsR8EGM0zQXjy
JwlMf5t5wClu7UXybMAm69aPmKQWbj+9EMV26v5D2aEHuasTSX0Gej1aDGnA/wtnW0WoiPuWRLAl
OmCFCO/SUDvJGh6SJM1/yFZdSZRq0junosbLI7rV0Jmi0/KxS3TjYKRUTMUTFU+4wW6b9iAXS0CX
ehkRs2PBtbRQVIX1moYTndr1PCKWmOIlKKUHKkHhVLQMQ60BXEgIYpFKoRUIOHQuyyEuoMljdfeE
jBvsnp6f9EixV1hBpNjWKKe+lSSKBkGCM2kYp7Fdu+PSmNTFLwi7KArWwloXXfdkbolV2O1BccdP
2CmlhA5RZGtAFu0Kg50U5DoGMmfDrkeQZ3ovkXCQTm5COp3Dy+D5zQgz5hTDT7czlItY2WSuNB8p
Tbu70eGx/l44U0EMdFn8HdcbFLi64hLChNQ2Jf57lYxJaknvI94gpRE03DlQ7BfScvib61NZaZo3
Hqyar/lTBWAUUdLSOuoFO68k0tBreOjo9eTMxswv6mItYWgDEbgiNlpNn+EwVs35I2F/jJZ/RKbg
kaVp5Zid8gAQd0I0nU61+cAGwvMZdB6Qrz3M5B6AiuNG62Puge4OBcpBKCKVwSoPiUzIf1WtyPV5
wH1AKXBv0vQzgY+zzx0/vzcMnVswUm+c8p1EO3KeXM6bAZLu5wCBKK24oetJ9d+E0Haek+jadWTX
MkBTvGpdpfA0wtUSozGQ7VY4eWFuiC2rHoxV5Mdnzlr3zuuXi5VyTk2B8bH/sL3RxWAuqKHSyFWX
sBIju6TZBozjpOLll9Do1UWRnXXBWG4h1WtNoK8pit/Bnko83wlu/XLrLTF51XfoA5aqD1LoxKWe
5VRT4Nf46ZPKk9S2rS7jlsiU1sxX+siEk7Dn7r7k2EeZt16mKq/p6pSBVbQ4JbS6e54UVJiRfCQk
vqStMCo559RPts4s2xeMX3zNoNsgOjigZmpJMBAg3DT2MGjH9dKLrO79hCM0FodFvQlLZO1H0Tmw
kQ3lHBVwv+WVfIlR6WSzaKFvzhZZ5mdVqqJVb9CsHIlUcaZRwg5t2pp9TjYAnsZg8WuPDo/pJpho
SS+pgDt8/zaV/+0ppAdG5HdFQ1bOJSYdYet279FQ952XmX/pULifMcsIajQl0zxyyNJCWXW7WKa9
61EO9omT3DGx8deJvBCpemKZNBU2BwkyJiMw+dVft/D0Nic9Bs95yq9hv5/Budu9ML1BSY2zrEqx
wCl0Rse84qLKxPik98raym7wm5Ky/IFiqYe5//922M5bsUEJppVjGPQYeRSEupXh3Sgtr9U9ajVS
PGD7JMgqStqbjClH3g18GbMF7OkJUiiH7Czf9DVKqTmAZCO4m2yUsRlF9BlfU+vWG0T4Y6NplbFs
56z9A3rPq+I0YKXhFK4Q+jElbT43ZadEhogIMbGHOgBSYV/rIKDoXiKstNfjEmF75OC03EnPJAyZ
HLO9FNiFFVIKPFo0rYgxkkEawxaKXV7PQ+W0pTxgKrqPFCyMjUMy41vWLBdgEkp/pIxPY0ZXL979
I29KINfE69joQRZsLj71ELe1zOtnwnAZqDTKOivttQhL4rjzeYG5JKHH7ez8DrRLZLFaUoYN+aXe
sdiNwbYxl195hsejRmiC4nioegTSKIOTBShW/N7yYPe1w8nhfaxNuWh9p5XWLPAZ/VPyMl0DDtN9
vL/NFOaWvb3c0a/krPKBGRualDEclsH72ZyftmdzGxhmPvws3wf1M4TCs3y/0ye+XRq3vfPGRUD5
NRSznjU70Vv10fS/Q9UP7k1Cdo7FoNHZpdGS9RBG5Y1SnksbbTpko5MpV30cE9yMjKTDPZVo02Yu
I/tabd2ivkW7X9fNBfmoFg77ozGnRz4Qmzg95XkAiuxN1Dgo41+P++QGZK4wSDwlpAtkwQl7xJZ+
G+vuJb5Us8bab4ue0Ew4hYKO0YRRTUXLGcsaTORtCyAb0IV1jUDXv71AhaC9lgyNWe0V7cnA/qoi
DRkbLdSVzGEEhnwurcRDtLcJp2e2j+j1Ua/4O/crn5y9jxEZrKZz0Q7b15Vru/FD7fPf1ECQq+Na
G2EaZ5WJJRxEAlNqK+D6JfjiEnO7qUAAcljBSp5rotXo5zCtg1tdMqUt6LOlLzN7lw6KWmSlQChw
FT8fXRKh4XFG4Vv0Ry1Z9Twu4HUo1SAuu2Pr1WgnqTW5XSML2pSN25K52YzGyvF9bK3E7nqFPiKC
gdZhd2ao48s5+5PrxdrOEt8DJfPRmAgR0/y2wm5Q2sUXGh31WjFI+MLJwZ9XFb6qfUu5AnG7kLBU
ndQ/9V9i8ZB0QAwadv2ZdGv7gJtPbcf8uaX3PO59MsbUeZVcXXjsr20cCUVmI0j+UB9w2ncg2cge
s8gUjxjFL77GVBT2x0jgebAP1JhgfK8nN0Q2T2GINahqVrTHljOMZyGmPCTJDVkiwx2bNxdobDYZ
Qm9NPCQ2by6CKhAptYDB15MliQ7rhh5Kvfpq2h9Adui356z+xOkzRNip7mzjl8o9DXYkM//jraI2
GAsR4C0USKcrS/p/2P8LP52POWFtowuCDQVWM/W1sMMxgyXYSVSVLQctrsQ4u4Wdc1E+MJ65g9Qz
1IQUOtwj+/cVEjpbcl5TA4m0sGXzvSzaAfQ1m/88lrJNeDA/Q1XrGMM7WAkvXVmMTR1N7uwkjqS9
05Fel9qmWhBSaCgaqYCBKrHHNmrK0UDlVoD7bWuYFGyxU0YN4lHAvMQLTO+yOjb5XSjQOVUEe1Bw
RZ9hKzq0BRWYuAyW8ylIOEnN9dOH9tIDT46yuGkWAR3m+u1+8ebtg7pfkK/lEvY9nQChuf/lYnVq
XJOOKrkWMvBYni0WNXieDD+PQXJ8LQSpwePkwGj0A6U1UXoCkzewUE9z3KJ6Dc/3XEEqHtGcrfmt
Gpdbfq8J/1HZX76OAjU7ZO484tUpQA1/5bptRISV8yhVDS5ua3JyfhDLTFEXetIxbF6sI/uWXTW+
IMXOoNloZi6RJXEMcfbBYInd7aDhzCdadAfeAiRdTr+U9dLoegfh/HQvBvjndnCoW8H/SfYmLzaF
XDlG3RDtqQkvQXprebNdOKcG6Gz9/17H+w7hkq6N6YDDrAGKYebU7jlmv4ncVK/PCAal9rakE5bL
4qMU6gr2w9AtRR9B3i6dQj9/l8v0pkq+tkK5Kph1efSjv6pqpOTFMKnlNGbqka9LMIaY5I8nuyTo
sqb/5w0EYH+8Bd3k4hVOBVrhN5I89xeFKP97iXodWBtlPzMZBnB4na4SV2jiVKJn29MO92xExmUJ
dLXNN8LySSh8HVwIPVtC9IiH/0NfXZdrSilGGIml9yKNNDanwRcN2LI5HSCGW060jm2Db5XlUZJo
uQJXX+xqDDeuhPH/Y6M5r6vbLfvC8WcLdEvJjYa+H5TDN0qwJzevEYMKPvs9bVRPHAhm4mcpfHt0
MpjGVDU1FW0bEEFXbOZn5aJMiv5J/RS7t74m7AXTbSr9hAL8Ingu1gZwm8swQWXi6wqoGFtp6PxL
frmOOpMRFH5J2N8iJOmUHDVXSiGv4mZJG3p2MyAaxkDkVZKddNK0NmePk8yyCXzE3453xZ4jtTsN
h7bVYrNoaF4/qXe4bUXL+gWVEfKmlJvdHXDWvMkpes9bFPFN6IneI6KFjG/rWxrrJH1/bUV6vtuD
oYfMHiUaGEwLJQur7fXjlxVmP9WowtEcA/SPK/fPTFZJm3xJnMAxNqE8uGaqWMaVoLiL3aZW2Jca
5UpqFCFRP98vJ1CMHhzOw+pKpLql4f/YV9diwTdHIg2Q8hb728Hv8mKeDkwhtb52hpzUlpQ4odrL
MH/1umQBN9WF4knXSENWs0IeWuFZQKOVk7RGF8+gMazb7pMzmuyCBkarCrNp5bZpXt2oGtZhPDze
817Vep6lI17DJqgiJA+Lxvv/CO5awFd6p0KexvCL5fv8pc6ZUszCU7p7VPsZh1kdhvOSzoP5hldH
kzZWZ5k2/P3kQcvA0BTg8AY/SL0+fTaIj6LqlvtLmBD1FKL7msI9jyh8Sdyye9SHWK/qoNjlK2q1
yaSN99DJqk0vxDokC9AF2UNqRtQ+JC+GPESsSh/qkArIFIjwBzeqQ+5yVoXHyaCHZoUYo/F1diOP
btOh6S8anOyA7R3EetgJKy6zRBus81GFjmYHGjTCJ6G49HmWTaxXq3A2oks64t3+Z98ZNwi1SBps
bpP00cLC8cCuCFCnE+SHEZynVehTEuO6JuI+NdE+Vl+/TJXh91UxNP0Gn0wC7jRYhSuEgdjhd/T7
lkglUdEK9TkzjKEdp88AD5FBl9db6XGTGTu5UyCYSC/0WWinVc4+u8PDWwK6xrJYOyKA0HCFsl0S
BnIJAoVJSQEVx4XPpWLVZliBl8ntcVUYXLCBgNv5mOdJn1Bw5Vt22WbURvylQh7CXE3EsW4uGYGR
NLm/LBr/smk6W6p19472vEPotPSG+aiC3PQgRsqJHkgzKvfDi67Rx10WjBJObgG1Ln1KEA02Ciel
SjZi/S90ZCb/UKiV+tgbSbnxRcUR/jNRrsZGVFP6R4h2pDajkO5CbdCJ7EKIYQXjA+thKuI3IN6W
yC5du1fXPnYGhDLncr41jGbygaTyD97LdokMlYvsBh9E+NVTYaH/g5+VKwt4Hl1nEacUeoV2PfRz
FqOtjipBfL7plwUAciNpu/juk6GjZjFfZfEqfdicXdMM+dCav6FObYNudQKFE9rtC16Bm4jVXVwZ
wqjV38lacmH+fIbOGsCuJpqu+DSaFCcZPT7EPRwkQacIc5YUJAxc1GtdRZHgObGNGe2kF9jZXhpr
qBmEniWpQqWGqswYzVrDHr89WdqxGG85eGcZd0f0eFvbn838p05yZFFTdxQ0CGDmfMRxy1riZjuy
IcGLldGmOYMX7gIBnyGhvfl8GKo0YjhGwbzCct2hx610vOXYokZoB2/kgqpRFyr6acIogyW3UagJ
qypuoa3eOQmU6886qcRimw9f8Nw/BTh9Xc/2yL/KxLStjnHX6z7GU4VuLdtxw0S3S9K4Q9Dq9Pnb
c00nyq7aCDCrC0wOulEkiQY+Y5jn+g7DobpP0B+xuDK9+wEZoL4iTOffloUhHqNkB/Z2WWAg3vFg
b3IL1Z9kAXl3JYPL8GDmlX7DwHUz4+tlWd8wOJ4zZJxqrBNslDYyRKGhEvrrPKNW+2lfQ/ggp+it
zvCvQ7uzrQbrKVCV2dwtxUgeC38TOzzxPXR09nDevonKpY3lhJjW78nSikMcMaIAaM2oHwWhxULW
y0K8s81iiilcPy7Er0LCYcxVWSKMLcXijJY5cOB7yWXOPUnO7snpyqYyNDWyGbkXrpZ4kkYDXKcb
5xsu2b7OHFsbQntsE2XL/VVyW2//xM1h8/mAuKNeIcueHBpdc88vFwZLZBmwVIjBdVkR9+nTFLd0
mvrZ0oPS5Vvh4YtV2MqHtKBmHwAURjPQHS7Y4/6V0ZnGA62Kwsos4a0NAn+n2c/UpAto9YVPopPw
a0PhuJ6UyY0a1JjQThFi5KiA3NTUt5bHc9qfIJJxbiNgjaWGXVH1piccjFve+FvA0CIXRaeauG4U
K2pPuFjxDbcdeOKa0MWC/YslgVrT3tBPWE9Nm/FOWwQ2mw1MMS/ZTnVBofJsAODXh+yMp3c7cnzQ
Qt4GJKUm5AfV6hJ9ghkdJ4682TBCSBPVP7b+LTJFpZH7m4NqzRR3xkk94j1L24QknpHrbAnqbWD6
v4l0Crtd0sIEI7Zb4KNx8mQcVh0M4FLWG+te4trm8Hg7MmS6F4XBD1Q1x6Y50IfaOL2fH0vyNmAd
HyyDEriUp5KZE8aKz8xBdGGeZqZQD3p+vvIP0oY7+4EOyDwZ83/y+MkvKSHkuoA47VpMLEDVbgtw
mDdIKOjHaheiGtz26+6XUiMS1KHd0snvbt7RkmG/xJ2bQ0YrMU1NaIlu8JSp0Lxfbfeaqi820D3H
+Vt7rDFXnOChux8GC9muNCRr0jntyc3Pn7lhI4uoG7dXlf+/hWfQcSATUybH01EMfhQp3hvWhzdu
Davlx5jzK4NqNwxWkCeJz1+Ugdhr2mr+y5GrfcH15ct/0rzhcp8ZhK76fHfSRPPCgqfGJ6VFe5hT
kPvhTCebr3c/6GW+ywxfrion7XdKMMNr7RDq910dWLw4iudWE0j30HdVSM7yGA11vG8LdJFMp2/G
U8PK3Xiw6KLuLfJpvsW/vHNfs1ZBV77C+LORndGHiIWMcOBSQHc6uFpG4Z26WbNy/X+to4OAU0aq
3+meh5SSym3hl6CRhm6bHpdjJP1BHPBCg1meTMryx5BpE3QSRgyKv0gBJN3jTqvwMe8hArg0Ku+N
+PZKwtvsQ13bo9R9w/YDGpuHrjunMY9JqHMRLxHSHdcxcwDudcPGyFBc5weTjOI6ezdyeFHfrdwY
MLMCyMAgx4cSHUnoKzKMdlETP009JP/1d3xuV75TGu0PzABrPh7giwRiCH5BWOlmgzbPaqySJJ4B
tuJ7KkzxtwVDtveFLGj8ErhF55apKMzvPshtTHlvWWOVGT4d3WAY5KTGL1TJKEg1OKmfv0CW0wom
gkWtFdrPIvxNpLQkT5Xj3k+W1cdqojeC6Bbq5YFWEKMIoU3Jys3W8GxTPw6RHVja5wNTvzHN0ZEf
6n8b7cEz1kE4rmtqRUvOeYhEO+rdlBCJ+k1RggES3V64BTZbaogJ0d/gDaokvBrA3ZDbYElQw2Hy
ZOY0A5IxCHuCuOBviFc5BHIu3ubQ0ZkjPyMUVfzDaHu11P8whjdDTifkK0jGVi9PljeLIkhJmVO5
CZrmUbEXyNJF/Zqbx8YyV9KfKMD/U4znl5gOXNpj+CzZqE3lI/YReba2B0IKyvghpZWWE3c9r1Nv
bB34N9CxsJUOZvaXqL1Wa+0AIBQQBj5fMxzgRZVm7TgdYIU2Kf05NaECko1gfQnD/JpyRkbeTMac
VxYCfeoqmctJFLOp7fmnQxvNhrvGGf+XYl3vAJRb2ZHHgvVC2lJGH1ALvVNHfx65JbP7Kalf46JN
XCQMR7Jx7l3wm7uwq8r+ubEicLjoSBIAsgbyleJvZcIcqoY4ZoDKtRBAlLflZkZv8CvKYoRHF+Ku
NXOYJpLJBcu8/7xPyJ9pEBdRsEt+ResHxd0uxDPkKiEthDu3IVvfreFTaA+y6c4cQi4HFz8LOpqc
B/Pu9QYn6HyR7Tkyfq14epq/QiAG5mkax6RA05H1MnwqfxHSwoU7tFy4Zj5lryxugg0Pc3kPOW/o
Y+ri3D1yjjH1qRB2v8oWNagKknwBqQtellQwTJ3MQPURL7jNCW9EAW6dtt3TYn97xHrFEm1iKOj9
hPK5md9yvc0jYvOWGBmiURspnOQlQnzXUqfH3Qku/StNxxRNHEOlLnCOAJbbdCVT3CMnGAe+4bZa
vjrT4yS0XO2P+sU+BcJyMMMUR6HkMwTw/gjbd3lC+TCTdJkRT05/MBrMOMJMat4r0ntyr2EF662u
+oai2tBJubeJVGWwKlPvN6y74fdHZKHpi5SkMyH5x+TqiWzKsgfWY6+s7MFINHgDCnyyAb7+GXYb
U+faBJ4m0VlUmhg1WvpfIYzZlhc/uuNyNiF8gHYEUe3DFG3CWZTTKjTEJLQUg7mwWVUhJuu4pO3H
KyjwGLBGOLDSXOoIZPFNKQwsyZhYzjGHkHuptY6u3oNjsMun105NqS0RPbyqcx179Zz0RSjsQXgR
OsfJWJesd2FeOovJDstccw0hYf/0YX8k9BtbBl+W8qDhLmC+Ngk0Rw7XYS65/u/2jhtpj20SFvTQ
wdWtIv4q20tK5wgjssAR+5jjoM0Xf0I32Ke+CE66iqLtOg6utF1OqsSPhMRGpr+7ajzOsw/64n3l
YvOblqUDdI/Cx7g0Eakb+4lb4HImmyEH/uZyXEL+dKwYIWhxzN26Sj/UIXnDVK/ORyZp8Xjj/F+A
MkYrpFHKU8vddEVyYS3q6HuIJVfxzCnVkHBhXHH8adTxK7m2W5D55omfKGUBITIe+6nL9OhlgjJl
hQ0UuljfejhogQByaunVMiB2X67uZdIomhmwJEFeBZiJJd5xV+VtlKwcnbqRA4U94sXbTe9MhTYK
qx5z6XanbcrZh9woVeYMCoRjZSmt9r+n7Lms2G0TgODr5XdQ/xtlOQ+OWfqE+apRN24XcvfgItyF
o8R1ZUNMMi05aOdRH6qCq08fnPqmCuRizC3lekIWT/9cVz3+xHppsgRE3cX9mM+Ow60ZzcEIKGX1
y4cB++xR1LF8Qhy0TzFkNj/Q0nSAfg31GCuEpa0M155AG1AJlqnNOXKhNAiGEC3MtxXN8998oUix
+bq4vpmP18tcxBqICNjnP4sMHk41I90W8TUIvov2hFGmwiZrRzumO/zVjNQxty9GCQU65ezfStgW
eQ2M+zyt5Hfn+gC1Lvt0Nc9fDj+FmaDSBzYXp9TC/Bb48y2f/6Z1NBqd0naFamLqWEuRNHnUMlVj
WUgXJhJXxrYeJOr5fYTZfIeyEuwTQ/MBNd02Jhuz9yPSbw4KZTMKO+9R+b+aeqaRxgTahRrn5jJG
nZS5kjhCBqkI1m18mwNHEzj4BUOpSbpMUsEHhaX+nHcXuETKd9eQIM7qgThLLjxPz/2PH9Y4G416
xAwKmNZMjLmoAOsxfC0aTPbxxutbi6vIvoYzu5/xm6BSUA7Dl1vE9Aq6zPlK2AYq6q+mCbFKedtz
ylY+G3PvyKIbQkeu8Qt+STzl8EAHWeho6no+h6gmskDpmUw56F73q56ZIrhDxksUCzbGhpDYGPBB
qmWsULjFHbHVEyzXO+EfqVtCyCZow7sE/f+DIeG8xUBfMvnTnWzFr4B3QtiZKjYykoDwowYEMHYE
GkOlhZL1cMLXgcIPxpOVvAub5YZdpbS48PM2sWgInmFHsvZfNuLVv4xf5HitoVqItWWoYSsURkWz
MFFq1wPXeli8cub9EsXatMzv4rtJ7p5wtZsaf/eSooTZ7UIHXCSWpRkFkCFjZHWBBm7vqV3xYG0/
flWq6wEWHmWQN+F8gYP1NxrLzqrM06KyIsN3cioHJuCVOD7Mmb9e67KxZD+vFlJLdT3uIr57OtoG
Jv/kl0ZU4HBfTNrC1KsNAQb5Lp+szBClbhlajp/Lt1/ebPCcr4kDSZ3O4kQDOaMCiK3sYAC7PAbK
6ewGHAtYgXjGBg8z1p/nGU/9PGCOSj6SikHMtIiILj9iJUmJXMBLEiu4Et0WWeke+fWOlqZT7nbZ
LLkWv10cSA+6QF5l86hdcvxd6XbWmbbvVvy9kzLJlUPSqMwHsLsBWBiVyLlMUW4iryguh04Hs5M3
cxoagQLfeSSJ1bLImDDxjEqjUggB9IXRrb1RjE91NkBaSBPwXEidqRHCDxkZg8Ym2tZ+LUEhKNCm
tQL6C9XJw3JHDj8BDi4hHm9dQpwpI4Pl33Z22XX61/alm4ZkXxBnl4e2unhPbVRdSXGEAH5zBbTq
jlkyDaZYFsJHCpH/mwrAPgHDRLskbwQJmlQYuxqkwt7pv9RooYRUGmIBoR5MzQ90Qlo9EhahJtZp
HHWnuOHVWZPhxOlit5IHXRbumIMg32i7lqld6QIJ+LklpcGD0yxbQsudaoa/vtQggPbQ2l0hrqAT
Ga3FRl2kjVTiE0+IQWhAW9WP+90dcX864OoZKbDpyzFTUqE5FALFFXHnVeOnMMlhzRTpOoM6XMYu
P800jb7WU177IrIoywOEnaVYYlWbyggH61o35VsKHLGAmnUVOZFzCfs4QWQbGty74vxsNe7fnETv
MZGzA3Mx+SuVzytdkVzzSOyvcW2MtW+K/bGSM1c59IvklrUABMyj2ojGIP3M4bGrp58dPBZkBT7J
FOywalZBIoHxpRVc95bFQcBvgj9w6+vCutwK+gYyrGR9PrMMnJkPtYAUeJ1wXBy+yALHujqVEL3k
B5LvI+HMIR23n4sbXTc+lh5F6S2Dm9xLT6xcc6/aRSuYIstBxetXA0kaFtK7OxPF/kx6fFuz9arH
u/U5SXdm8H6AwgaFgeWtMWyFLnRoQVPqm81MOVeaUPDo7fE6H6ixc9rnx1ngObU67gkLepkK2nZY
kA90RGjX1kIf8GDWdOeH5N/Rr3CCAIcqgnIru9O2oG9d1WlQA4NRQa9InAZAnPX0oi4MtqZ7CmGr
blUEhBfgxWH80Y/p28LtCIlhDg6ib/YijgpzSOaB4MRSMKVlCi/gIdNzKmmiAl3uhmhO6uOQG5kk
QLQMoIkdc6rWvdD8zz7TSsyasONp5oFLTjYkTK1vQg+LNMMgeUenA/5E4l2hOOF1gJHXSQ/AE9LD
xYPQVbiAhNzoiHfCTSsCOgsxV2E47k/65FzyKrXnNRKN57APtJf917SsQprCCmJ+VDWdPoAD3qP0
n2Syds/pWUnQ45p+C/hifuMxQ1fMgXgLH8FRFB1sSKo7ZkJrgUKYQeIfaRtDutK7t60TQHPssVnd
/yakv/JYC5AAX35SIbF9TtYNFP7+pXwSu10lWsHXdtlJZKbgCB/n0/mMzcIDSSf7TrOb8eTh235d
FFKXBktOZ/BBGoWN0HLnke+hjgg8Lqo3eqfyy8DdksYpjbyXRqX+UBQrnHrCMzURdq0YxKdVbMcm
cOMIN4kcIZtzw9DErYo2vO2P+px0cTDO2wUn25fZTZWZ4m3QjrTB9QF+f8A0Bj59gIZVIBNjMyzg
GyMNC8D5Q06Qda3PyZkrCXg+MiR4Ys2I1sg97FzJpPfXktz8+rj5RYPUNZlzDhFdI0Nlj5v+iN3a
qgJmCnCfa5T+z/HnqXVGOJsn64P17BqpsU/lB0PKpShOtP6OevX23F1jlk2a/9ICua24zZdYtqLu
kopORWAWxXnRQqQFNIXyOcUxDL8JqExKqs7J1lBVow+RcV82GpUIK15Ug8JwUhqQHs0qqx4WH9zS
xGjHN3HXu49ekCTdHJmFAcYeqUMz98K7wFytVXVRmPLEE0KoPJrf2HGp1CHynVatZMKkr2rI4gbM
dA8fjZBgB5EXV58OaPJdYgdfsVUGp1kaXxXtgN2Yhz+YExlSvOymkH0+2Cw8luTJx5ah6VU/Efen
HzbJMeMeD8DESUHbXj9TqBOLbOosFouC9FNN2BbIopU3K3rzzDrqR5i8QgXZGZoMxP4bxJUxEpet
/eIDAeawbAStlTvXGiZ2LCuiR166HYiVvH/7wXSGBuVyWDD8rE33sildAl5mypJJUzby+zNoCrar
Ccz+hfRPB6z+OOdPPCNeJZ5oOHSzaTmt1u0+1eLLkmhFW0rzUyRWIHSzFFnB+wKtcdw4tsCirRiD
COL3GQDCzGaxKDYK6qPnFu9EA2LvxnznMy8UVplSN8dADTkxJRJ0Vqe9evWoQ6rcd9jEb3Q52al3
cGBe5wNZJYV3byhkz6EUNztaKWLVAAH2oekJcG4L6A2GPKEc234bAsQfZsZqYOSdpmV6vNb8v7Dv
Bsf7XYHuK1FP12+ZgzD/IdjME700aXvKM+ApaQs/cCArsJxzDG/4MeqtSyXXBYiLmtDmoRVn/n5S
Sf3+FU1jHJZWkeC38GKZ03Dt5mKv6jDUY7hAixaVnakKDRAbTAWPTQeG4cOJiQ4+lLwyZ1c0T85d
TMgNUbzK4YTYxLfbFhqi+Z0ZkZBkxwnTmTjr1n0JT45fSKYXhkzKDLGmjEHbz1zTdrR8/iXGXe8w
dVT4P0Y4QDZXg4G1VEOelBthffQISuBlhJj3gFBITXqr2xebVGkG0xRyJIRkXYOSTYOjuetcNwr+
sidZgKf6cKv6GwH7C2MTfxb+vIXXr+tsm1zTaCrmVeXG+Cl49gkpoe3hi0l1W1dcKI0KuKok5TP2
OGEVP+MkopmIOAjL7vwQlS+ow5ZeMQQ0S83syXO0x9WBfyKRpaRX7NOW/AdGGAFOX7VP4qZsqB8z
myRLU1+LmnVHaUpd7Zg9AvLhLxaR9idPXaFg2cPvn3zHllSfRj9sDhiTAdhOQIgikuy1dkZgIbE2
/W0ohD+0lbfyHrqa4eTfmTgXWXiv4MoZ5xHHkLwEhiW4JrIFOzBWOl1gFa2p3TPQ8F4R+yogrfIo
AWGmdHZwLGMa1b8fAs9H6s8HURA60WchdwtKRKyGL4mWcfjcqa/P15w77qpg9ISZfkHAOJCXzxZL
vXKNP2DHwDZUvZtkQ60IQjF3mullnKZGAlTYyyqIHMN4Ao4R6Qq3c1HTuEn6upeHpxDJHgWAt82E
2NjoAnWJTNrcrbCBeNj1NokX9p7e06K0MI6862ZBxgyIc3cmQjjJZBQ3R0/Hn36ScvXpdtri1KEq
/xuf+Wd9s+FBdC2ciLUKCPpzIUYAG80Rexq/0jPOWKmYSJkU4ctHKNhsr7C4B1dJ9Mn3idO00hRh
wU7V/+pVVcqTkzz4P1V6jH0fqNxWOibpZ7Euife2a/wKFJ5Vy8vAtwDdg6U7nE49VJTMm9W/pw26
XN7dAX7ZyfTpDTtOLV6JOZ1JKXxgI5lLvkDE3QLUVUQnbvXA5/WcQ9RQ5ALU1u/wwH5nk1OP+H5b
dlRxo5TW8zn9V6CgIENXRIlxKYWrl+N5lED4uZ4RrSSny5IqJtHyyCBkVdWdnL2YVTJT1GmJQ6uw
1Uz6Giry6P+QVPNZIf2MTu6lZlT0D96nKjyTRxP6SRJAfzHZHvqmmANwJYcW/xFQafdlAW+6Nw3H
KfdJ9baNlG70qf7lXRj0mZvGK9XCFxDp/PnFImX4l3dSF/98o5bIZNjE5fL7COitjaDD+iMCd1q/
Hsl6gylc2/TOG26ucMMzlk4DqhdgXkOdT5g+FO40yjz42H4lAueMPGST0/KtgZyXVcGlkesgQdsH
Ho50ImOLD7hCzFknkdzd/5qQwqvBWdcq8T9fH500CsKp3PGASnNYXTEAoUPFHI4UEieyzthzCgvC
F20pcp2q2tRA8lpjb8UafyxXoF9PMUWRl7aS2e6E3z7kPJ5wQhhVbwcnLz0hUjZie9K1cJ2TIT+y
kWmiQk7dr4iEz7lpYb3kdmfaI0WKo/cUjYRn+BtlF/FydRbYY6m9N+xdtOisG+Pf0iqmSBaffZDE
fvO3WcSTTnwcsHHK1cYs7OTk1SAfh256UrTkM8Kh8wywCg9UlzsSSt1AeQq65KWz2YN6TYe95OBV
HwqH6dNzWM8gVhlk8fwx7+x5hLF6gOU4Nn960LKuPM8uxDnLaaqJ8h3XRivBEk93QM3OSRlKUNSZ
1C9seE1v4LI6ENZFklrKF7gfC36f0/ljYrNWJisVlXmXCtlC+vM8ET4TOWBoYsFuyOW9jPcpx1U7
9WHsB6HEjF8AabbzqHg/tyHMsxF9szEI93/WKSGc+hUzp9NI7cbKGq8jV8VU+49OKBXI0qKUTTF9
MBOy8rBIkCD09p1xAbD+rYOmAWdDDZ+Srzllys7O2KULQjiCTvlEtyrpF2V5F0DgCpkvdFoaHpds
04iZe58h17+2CrDZzZTyA1VdXLEH5idO1JRGH6L0KgydLjHHUD4ZO4gNxBYVlNTiirYv5GZ7N01n
F/g2CX3gxls+ZbQ6bqF9zhK3n4O5ohM+1zuybYvxDmTFaDVEgsj0OcqJIzYtsZJQs1TghuaMdQvo
hmj2vGcpI20k1PMvhiwHwHReb/KJz7dmPJx74zff+354Roud0JzSMqlRaF2VMBH48CZ193mPM7Zq
Hij3WfC0l7y/vCcKWZN2gLcwRJF2rm8JeH6hbf7fd9Lw1kaY628oxxY6+FJq1ijcYIUVHjVZTt5u
JhQhB7Alfh+yNEuim24dywl2wD5AshHZJewYIQ/QSDltSCUkNQGrJF1rQpOBfHH459thEWhkbfAZ
DvSyghOkfRfZJbmD+Y7Bt45jHEEzr/fguQ0w5on4xmP9p9N44t2/au3HhpYEkdO6C8HdYgFBs+mS
FB6ajavH4irKG6UzFowxnL+gZNruCox669Ih6B5/7uK6LyWdKqIzKjgmLn365pKYrcQnRhfp0EU9
jEyngJQmQ7zmfpoj1TeCrs13UwVbCGgh8FDg9n0Wivk4NPjRVLFed8hGV2pmt0tDqwp++IfdICqP
6jLTEt8Ry+REg4PoQoPcBNWAo2MwkpGPQDV1Ch2gsZ+rfK4dAwqidHvYM37+rNidjoi57EcWEgqT
AA+Ho2GgKbahT+LvY18jlfSguYwfuqUELmP7Yi3LQ2e9wdQ0ZTRTU8Ah6RG6bkaxe8LQpDl5uify
8VhNOjQpkMcbE1Cd0DnBHyDi/GgwQrf6eX0PkcP+xYxLY8VaON2z9elEhSldK1fK0MTffWavtgvO
URtf6C9eFB9lrMcECgnfw9N0fVB8xtsS7CtUMFlDVPOhuIVPsMj/4CEEX6DLbooZ8sFjKVjiCQ4r
RGp915GAqsP9S4wlX672czOh1uDOz/yGT0sV9bkavs9DLhi9KT5wsy5xgSbgNR/M3mA5OJgSB1rJ
V6Cq1kdaTVu4wLRuS/NBAnUS1vtgM/8y8qoz1OUOkipdU6PER0KxuH8TJ9bx/aax3/FDgjw2eR1y
la1Pes7cV6Qy/RHAEJL4cl3gPu/DvHbtX4eFcAzcq2MIy74eEzfws+d9Djpd0koNvjhjdcITvJzD
DW7BY/t/homnhmhPmZmrsOAvKnBuqgaLN616IU0KI9d/Vumvno4mDfGZjGZSspJufLTQY5c0R14B
9PzaOoOoAUgCRbA+TPytiUB/vWtjx4ChzP3p4TslbJq8Yf8dDT6+PsJubM+s+zQpa9CygxlK7cNE
kG0zmXo0Q5MEeizWsz/QHx1x/G2ZMq//2QHfTr6eA4wJ+t9/ipspDOwBGXxdULnQGgjXlpQQOTil
CIkvqFQ7wB/7DzWjlejYaArVL0AJF9WTZBwxpKzdnce2geBYqke16bdwyNPwPmm1q7vqP1OBii7m
9Q2ldGTNQpkfjmmnDdOGArcWj3LohuzNi43ARFmp3qIOYp9TT+lqoDTn7dwMULRj5hyE8nkcNSZp
ZgN3EBxvkag8j6SFCzyeIm90Ky0tJfZJ2JJP5fVIBiAyZFvZAwDyn5RjOViBVmMjQjxEkkw5HfKM
vPbB4fYWdGF10N5+dND7TciKRc5AdruN0Aw3mHWlNahplLeuFGh4jcIj5U4F+tJHw4ZpcRsM2hy+
Z87q1gLdKiQsItNfpVyoyRHZpgtMlQs6ljSQzRILrxgIz+WnT612pYM1ynLABnFyC2m3uNrZ3xdO
40hJ8VobQ4pzgGUGM3FWGWis4Mmhb7l3M1uaTwUT6LDQrzNmbYaJrOfes82FhnBMx8Kg6wNLaaRy
Ll+MuH4oK2SnBscpAmFES9KoK4/95a+5WLRCKb7Ir5O6xQrcSj8bqcuKgkp5zgVfFeygtDJSpQhq
JvgzM0FsRdOxp9pZDYcOjQA9cPR2ZbUSB/ZgsF0Q4aIGrZqsUCkST7t6X6oIJc5TB2lLwOgWZy1+
2OtOjGHLyRdn33/wHZNfjFMSir01o3NSuXtNQdW6X11j/HnNUa7ALbi+8c0peNCkhIth0YLi50oS
fUI924pLHOfCaE+jp56YwYF34BV9MArpIuVmLQXa6+dEXKWhYu6dpKTEAuszauuTAcBjIdI6gnBK
zTZ30G05swA68rNzXoN6Mmq5DXW63alC0ZBWtRMNfz+4mypMb7XwEzMnFcQULQfmdAntfDUDJDoq
KbRrgfRbiLfrlNSD84vVoQd5Vz1dVPOt2Sxb3U7p1dW9J5tcVMHz2Q9aI3vbpN1nYouMAqtQjcSt
vy7fg4gzhvU+IPaGHr+F9BXzRHtZzbKCRZuGRn3NF8guCFqVRZsUS9eYEHS2kCV5YEDsVTQuOhh7
gPBVPzUnhMeOe0Vkc81WiFiXGeUGoaRryIO305fS1sGkh1zzULP1ByuDsjHqaHtMl3p//thG8stK
NfN4OsEwJc9TCr/QeYmZfB/bflPeN3EVR+O+KLNfzFRtKxs5iugS9IFEIfCoCeo0/rjWMnrnWLZh
fpGoaTcn+nT5Nx85zr6wxeO/PNsGsD735YskQ5NI7ObN8e/0mAPvr6GO4fw/lLtF0ywoAAuK6f5G
CbasLTVjDUtKX4+7KkNCXboe0PWb2JuO69YF+9thX0/53smB6WJIWdUt24D8XfTxSa3fi6OSCLWw
SJ4gbGtDgJo9RobWAHEaWHnDLk7Os1FWoAFB2o72FxFGXuiUeurQAnNEJlvCKQt+SihtiIab1N5I
6jiUdiDIad3RCtdVn2l7sTBBdwL64UQWoEY21BBFS4+mZyCghxOSMxaMTPhZbvazNaxHt69A7LeD
VAdXtswEB9p7XFJmXUgAWXWuH/pD3PiAHjR91ZOKtYWLSAcViKQuiSndsB9xpLd+G54ZYWq10rpg
BZ3qSyXtY/wuJFxyvm8vug1cWzQD1RKHfHLhU9Laa9ewl5U1sKqVht1pDNYqbcJWVOjDlgYtyAwa
hBM8NAjHiyz0jgdJ575b8u3UTSO1FQlByjfYQphA5lm7ESZgNB33PVHxdeH5AOh8F1KzD9Gy5Tn0
kXGPY58zCyOIW6XaXFEKFeOiDcteryiHpWun1sqLZMiG0D2kE6dqicctSFpiG5RHBSWZ4amRau5K
JVVwJ+/TyrbiJytv6135nogkkmHk9pHhDe4ShuXaQgBn7lPElQkUAEuslM7hrA4SwpjwekP6Br7p
1Feeo2e2zE29E7kSzRXzNmKQBv0mvDpwJ4iFhOzCiX/POwMUUJe1AFEbLTcwta49PV6iSjleHSEa
MJ9aF/TuE3LJ/MFuFXTYTtThRc8Ekl6sVh5ZlfksgT2cyB8YF/1hTcoDz7MNd8PF/9GA44HVPzKf
2OY2y8gTETQh0lgXNpWg/1LQL9TvYQ1lwGGSLgVFyfTz9F0LEYXmWBtDrnUiNiWNmwg+Ty+6WMYs
mEX63wZz2Hynz91To+7ZwejPZGt5QBM+Ry2HaWuNE8RnNZ+9wjrSWzW5Oe6f+R0S16aAaXdE7Fnf
lW40PyGE0Wgk/+cWL38bCXnwfuX68j4VBw0jrRWJx/GAMisOxRCL84ZjK+RAo0P1KfGrERxzGuaZ
Hc9vRSbFXu+7iYXgXqSiwdHItup0eVtSx9ux+T384F/23UP54xwHDDFOvkwIkuzIpD7wp91wZd23
XoKqfdlDL/g2cg2e4X3Yep0XK8SkgHfVkVH4jZpPqSTtfGE9qj76VoVEdWBaeYSEHaSfeO9SlY/F
FKDOrmqz2112Ants+yfNjNPlxDky1vl/0CyyTsyj9LCVsq39Ws23RgmKz4iZYDtjabjk37VdDf26
FZ4SRSGqHtq6pFvpK6LZn9pyw8cjLe6NaNRFFshVcQ3NizFB4QnAXal03fNxxHIce4b4tUq8c/cd
r9+b8NmPPtKTx5UZDkuD587Q8UL/pAdaU1F2+OEmTYLGc5Xr+yFW8f/4IcBsdw1/RXD170OhwVxf
P7gXj/RpD3zDKD8j4zZQG+3Wb6XJu2+uBb/o96k2Ca305kMArSVwn83rHof/DnSj0qOmtyUDrhPM
2UUZPPcRrvG657mvtxvLsl9E0QURysieOy9pQ9Oxq+Hsyp+LRu0BLm1jgpC1jECTIVw1aitycvv9
q/DqhqpeCaAV0tmlV9pA1xBX5mtRGPML2syYnu85/1ZFr8h9VjpncRdUa3/J5nN1c+a2o1cbv9RY
M9aXdqF6uG0zxz0C5uONoMpMOrbpN9Wtk6BLx0Xq/hJIb5GqzQKcDvkA/+7TyPEx0EOQPQO3FcxZ
CnwmLrVfQO74YsnKDrI4dv1h4r5HwK2dzVAvIP+3v2zhiL2oUO6PIRKep5QmSXoPBEKDsqxr9Mel
qVrM30bhSxVvS5DI9Jf1+cEzE4aBURIMGIbRBepxS74y+5cUg5RA3Jq7awtM2BdHi04veUB3bCQj
8CfS+ihOJKnCh5udltuwWgvU4WyPbTzqqfNX8qOrdert4xLVc9Y2ZE8TDmMAoTo5iV48K+IFeWZH
7Mr+BDNljcIHMPOEGRIOgsf1vJ4Sy6q/MYzMVWhxSfFBmaSaEV5QxNJwkNqjJlUWVs8Vw2xllFRM
IL3At8ZriDJ9ahggRhOSDhKPMUV+UYz+W8UDDrIJCI4pSMt2CSL4zLkzsQ5fRZauv8IUvcEbLs4E
s5b12d2US06T20J9fcx41Cz9gEtNv7ECmlsdJRcABTdOOjAAtja1Wq/9ol9CNm0JyXBTgd3VWhRm
y6yRyV1kVZTk2vq5yOrAZC/cGptgf2H9fcpKh6HZJNxhIjjI7aU702nKWRfhR2j9+lPDdrQHCn9M
Him9y3PMRyW+nZ7ZCFydPRPhyfs901/WwvDnU4XWXzyyhsAqj3k7wV1FXXdeHhCJwVhKnYhtCCei
iVSZIOKOw/IT68V502kstR35tWqvpEj0269xKCFKEprfeBInCtt4AtztSAyAnIeygxyvWv7j5fP6
hczWpB1s3dB+K7dHo6wNIZ8eQR6gwGyUazMBCvS3VwVbHETHfLK6eM98pQSgkEl+HhRcOgUjEWs5
xPeOzzNVJ5MfyM7KWsF2UDxfcOT2ifLetYY8Wns8LD1wO9O32x9OhOWB2ndq1gmyGNuQwW4Z+Id5
KORxevFH8PkmHigF3dVwbB0QosrWDI48u1t6YFVhO5ANS6/WbnL5JUp4hrXMprP6G9++50mVXm55
LMEJRJyExk1V8gR9sV3izi1ODIlG51JTbedpBYG4/nj9VM8Qn3QtWmwZsdjC6f42/mWjSKjUq1Mm
OeFB9HMKUOQR4qj3kWoaFy4Pu/RM9aMEmAHtb7rpLiTeBKX3ClQ3tr9kkPiyfU7PfNBTpn4MlC5L
nhAsG9J7I1RqWEglR0AgFiTeyJlKx/Mv+gIx9/pZxyH6XlaH4Ap/84AMXek+QdnaO+dawfoECsul
EDZbR50FLpywCc2VI8dBaJTehvqc8gm99jMPnQrGUhGG3hvw+VvxfjsehBaWQU39fpRdeRcfHcQQ
xL323pJJMmkhwTKjbv77XzdRdB9uT6NKmKDwgayxrlZGfQoB4GuN8yMAdp2CwT4LSz+vjMkJeeGX
Z5Sb+NI9WKNm9hDbsdd+0ExHP+iEuq8q8/ir4w7m+AS4UJ/mKyoaqtqKWCY5yKixYRjV1agQ/SSV
UJZc4uZntY234CFnam1Nmg0rqbJC0+f7Hs/X+ZH4C5Vm769Jpwfsd7Ooia+yBamFn9t6ErgRESdC
j7K7ZrLqT+jGGdM4Vvo0RSnj7b3jUooesJnLNTG2vi2GtBl6N5I27eyC14828PtJu9pq5lZsIYCp
WFkTbS0545SunIxev1O4q/DT+KPWCcoTh92U7rw/HbHapu6CvY599/0o7OKsblRfWTBR/uIBhbN2
hqO+JGo3+Ok0SwavLRd+eCZ4u9K2cbrMsviC1iMdVEblZ6h2PEPj4wOLNCxnFDJbX0GIy5j5I6I1
fk/6bD+kT0AFruOCeWHVwRktL0pGbK1BEbDfNxGP2m7a79X4V4ZpdryQeXzpdMhlpSrKQZlKtmbY
cvTBNRiCnBRfWcgTMlSlm56vjTl4L6VPSY+vbzf+/Pq5yiA20A3vmcxcVBrlSdwmVWBroERAlShz
J3qGah2phRC25veldxsDi4wZvnNThpW0wrf5qbh+NOq0wMBoHYjQf5FItdBzO40eGFBwO/quFoYK
xRnM9lRbVwcxQIlfhmmjNR13Iyfc4ZSZOSWbxtByGspBREpI9sjxLj/skjSqhTmpxYPDpXypLJFp
SN2tn7+LvrSC4e0vvL7YrY8eQ5yQmy/YuY72s8JtX2D55CpGoK9a2DsFpi+42vSUM4lGZfLh9tJ/
1MMvmo1V44GvCiWTh9VgPv7mdBIQFRf2WFiT3doJRbj6TP/dd1YHoYRbuZ0IVAFsWq77woL6f9Uy
0WgryFCgkI5B71EkGcUqro6BNSpesh9S35nAbAWlFHcMGh89MwX/u8I1n5NlU8PTmw1T5mWHIRZ3
erWPe832vkmvOHmbCJsG6Pu8kBRDvhOg1a38dRdanRyUjV/KXTLtKc95hUt6n9ZI65uqoOqCb/Es
6b2sD09K1C+GOqfrjlKcu1JFpnCdEO1bmTm8W0jeJfRwlcZIwpqERW1cY/d9SSh9wNLwhJfF+vUp
OMZpzCo2O/E5dtkR5XdTg8DPoe5lshlFqNXQO6g2LofZOcivcFs3rD+5lHaaZ9LFsbL77PEoYmOg
LJvPby5k6EUtEaqflQHlJD0F45fXQvoghuLNyVup1W5Qt455k+CXs9R5N53yeF2O6kZkoy88/+nn
HXHteKtks33RAWNQQ4lzLg5Vynd7W65bzTGkVqY6HaPg5T0keYRWQ/iY5MF4kSdfPqXAhvrA2Ib3
ZGbr+q+/WBXfkMGe2UvDiXpHj9jXQO/j3eMj3PqwkCa6DISiLFfko4ldn04tYBuZXG8VpFAM0l58
l7z7lhxbyUT0+hOHf7Mp1l2PAkUuztYqqXfGmRIccu4U20gh85md0p1BtJ3KeNLlUpmthXYo5iHn
+TTeqOoJH2GSUztLo7+fwsyezQzC4d//PS47eXQsrczHUIYa7AiwwoLH62EvsN10L1fuGuwjwHbx
CWHv+7RgfYax14o82XZMlRyWAOka0o5Mx6T49lYlMYZnwX3uFPliRo6awSya7QeOmBPpAZUtfvmm
svvS1LCEdC72h+ZaiaC4aTwvaZLCFylXexN65itbTKsJlqd2JhtdRK4bk+nNStSItMkTv8PV2mu+
vjHCgpwmOjEuumUq3AZp4ohGamEbT6mMRn+1Q2/tb3C3k+VmZO5G81h2pK78bJ07lBjKJkiWtPMr
yH5bkXkdtPgfwH1M8MbQKLkKif9RRPcN0OzFz+DwSdDTkoZ+fBTCqj/NdX0l/G+spggtG/wr3AQP
PpDLThLi3jWn+oZ+qZgjVadeqtmyPYWCbhmMm++ovYPLyqBjPL/x0SYabvl3Ur0Z/T6fUJSnOR9o
4NnteUPuINzP68z3oB3YL6izSLzNUSUnOvANxGkf3U6/vEt8InwdqrSCvfjR4dNncSf+zWExPL5W
20Xhg8Ul613R0K4MVsMN5z6XP7lgjBjy4kTMah0MKxhBqkQEsYqmHiB8spjWbSmHK8TtEQRKeqWh
g/jeTSEg4xpNfFtL4VkavTPneh/CQezsX4kQUaP2a1dJExOZTwdcIzg/RRlU2rn7WQSosrn0IeYM
CmZqM9W37Vvi7TFPMZ+6xJRr8N6NRBoDD0jXAzARiVu8VUK1Nh2hhppD0s2M7J4OU6dlVQ5EKBMJ
ZgF+vKvkZxDBCQQgyjRMUOgUzHkFFlfoLnSLhol6jgAH1Pqv0yODWEQKulgveoI400S+XzVuv/BX
g7mmaoOsVuZcWC/JDbsqmd3//C+Cfcc4obe3PDSJA1dFh06LKSq/lF4/tLXWt6jqqPGeWK8avEEH
wa7+YRqbK85ixcHE0M/hqBCzEINb+LQbTAYLcYTfFCU74UySf+FIqP9vaht2msUAk6k/jZlV2nsi
zjwlx6vBH+U2hZxG9r5MubgGbOjixclx7xkzVJJDH9rpC/OfkMnh5aYTDVl18Sx/Q/O0TLb3fY+s
ZMf/MIogjqT1M2wYHZ+0ry1Lk7qGXVRUjxcEKJKwo3TtZNiteACU7ZgW9GBUspdInYjYkF534PGC
lQMcz5GA6gkQARjVdx3XKtt05JB+zdntJ9jP1Gbe4Y+tb1atDezThNlS2Ed1giKOnG8NxeO8mS6f
P0rrDDyG4MdJrSzw/FeftKImK3+AJQjjSFUQ3fVzJHbh1KmSalQtg7gUcgcadg5Tsozbn1hCnwZ3
g7EnU/SF5y6hqmZUMTRo2EvdXLBWNQ1xk7pnLeVXhlXS7/0cITbrtBeS4GCmOV+lFjOIG2Wl2crw
3A7hglfi/O4aMKn8gZ9Fw1wbxxC7h62t1ZVqmMrr/c3DnORg/HceHUuc5tuINgb0Qn+bkf5rgmwo
/zefpx8fiNdj1TCw4BMGiqmU9N6FFAUOgTUPv/e0gNJt5qsSg6eJA+HplEXDiIchst7ekCqvJsJS
ujZjSElWrqUv96zNNpzFSi1KMkrKHmTzA6rJOwX2IsESdeYDpGe+OE9aQQA1We/4GBu1s8bDY6/1
3mzIfX4g+o+2Iy4J6aAolaDSTUhbRrmj1MfXs/3RIGsvG/vQCQIejX5rHWVjjquHlQV3dAmkK2ql
ONA4q9qRhdU1hE+xOA7s2buV6/cxogIzAEFuS3Pyv73CnBf+haEvbsyVNXvCLQ/CQVfmX5rWOlsE
010uMwzvSiNbqG387MdGXLYhp3UR4dhc+A5j8JmhhUv6t6FZmLq9ScbGFuO2H+VFgS6YxfyM5vvE
V2j44c8DhpXd3kXA2+E4MgEoI3X1da+dailvKIOZbCUQUobMEDu98Lz3kMoXA5xj+khegdCaJ70b
BxgM6GxUP1RucXzLga2ZLg7z2CLcwSBjYYkWFxJzitPZycIZAkWEPvlS+CbyYqs5IvteDCGHBOFH
xMC/zN8mYMNOlNtWedW+6CSdJFVYzq2oCqhWcMiRIap9tUGyTY+ZzXfjlVRgVrg9qvjzuHarO4qr
ThJfL4ARlHcKJWOzoY5+7Ej3al2de7J7o6jF86SsxSMkJECNFNuXq8ljragr8H61rpKcLJlZXq+k
4rOuyDY4gUwcL8ow0ivtobh3+nhEIf0mKW0a9DOpqILQevLN2zp+ujtZ5KkFIV6uBiZuC20fYnP0
cJuxQxkhtK3BU6RDiRTCcus7dGJiE33N2/HuWGeBVZRDstaqJVsPJ0YtqtpLQjjM5Qj3g8tDwnfl
nmkVBu2HspN1lcRFcM1nb9C1meOooRbITuFp1vp6yvHtuCGXgAb5w9Gi6nyzZDVwanHjOUqbtZyM
bsigDetWrWacWkTDkyHDS/fc/0MdZq/xSyEk60XiUm4qO/muhATJEQRAg9EyoT4aAbOODshIgp2g
uaXFb6bB4J2vdPNM5G92+VdF+H6Ws8O1l61tfsDq3jyyCoSd001KjXO3Q72VNVoKmEiT3JhiGLon
rlxSYdCOAuYqcIBKqBOcXxEtcQguwfeBjotLN0+WgnFnJBBiQ70MUvETRqUetqn0L3cjzq8i4vrO
SLehkkcv3114YxbcborurnZW9pUGUruM+ZB3KfJCDgyuOrTI1mRuPwvkFRuVcdrx8pLLdjQ86+ot
eDVvL+pg7fgEHC8zGVowkUwVSuY+t3ghguXQfiLcl+R39jkOhDAe2aFu7S2+tFscLYbDd6FTybO2
h4jxd+VbQtQm74MwNAvwSnF+NOOZv1HmXQi67ZvdT9ggoHhDw72H90qi36ci76HoxFiGeks5AcG2
yvo17Al0znzX/+zuRfPFu6hHEJrm1v35HbHhnUD6LhTMJoD8Bv/MJ63vKg/2syG8ZX/uyt4ppLb3
Qi9srkwWYEOnmrqS6BJoW7GN6+g2NcwhI/HkNguSVqZKFwHSY7TZgaAvKWfA4IX0jG6ASVOPgUhV
VJa7oZea9hrfOUOL4KdSb1ZyFrDOy6PHqC50J4IiYgMXX9Cwll9vb9xokAVTpCeV0F6Pt6Zste4l
+yZoP3hV6xOVnRy8wf6KNp11CYWosyYj9QqgSiNSE3DLvzifg/Hp5D0oeJGTLOa/s/MVrGNGGDkZ
D2L9lFEz49Nt0XooH19GdgHOKq1iL4SS9Ml4BeKZ4E3C6mnO40McXZZ8RDHCLkCY/WrlWG9tlPPW
aAbsvStiJ0hThqnODTlv2uGhgZlNval1UMqcNeXlWgA/NzkoptIuSj1HFQWbPv0cgOTqu2jQ9Jt6
ZVrzGmO43mhQ6yz6c5dZFxBgy5Nfj228slSKF9mD09HWUnCed/dZzkeY0PA5KL/BBZh8+ewqEEZl
jQaNXlSRu9xgjJRiyFpZnD4xLMklsSP5EgYPMbHUVWOVkDX/zpgaIWawlrMljWAodfM5jiqAdMKq
Q7+5IE2LpjVSqnUVDIs608kRBgmMPes3dy1ZJvF5JhUEF++2mSM0rxGeBL+mS/iFJOPEpokc4Nee
ISupxdjRS0MrXmFgM1GEJ8gVuLH8z/6+8Fvt2eDgp8IxFBhPt5MUQP6kGAgV7nZuYn0VO4xB2HHi
tKqxb5Tuwqw2LHArBbRyYExRBYl4yvyktAdXnik9CKZe3gFAyYOGAfQvEF2t+SdQyA4FcHw6VtIH
Il1LG1X9llRxMzjxZ52QgC1zSE+yLmmAYItlIj0fBzkxlJI2t+Qdlo+nhz+kpdTo5DaiR6RYWj2x
GfJ5M4zNlLh1T5fhQWOwlTOevvU94ZbA7DT6vcwHFDWVbrS58C4mpVLByeOZeKbBEb7x75w6gOpj
HByXGnBIOlOe13USfUzG8oiCOrdmR6qUqfZArQCr0cnoR/tMw2uAh0l41+xjJixRzz6N/wXadcCx
j//CMwUZx555s/zTvALF5ysqbqAmRWFkX3JeVW0jh4KjUz7nYN7zX0NCF04cTIQZNU/MDB6qAifu
MtjEvEK/B57vOqr/PoAf7akcw/goFmBsqf9B3l3XcNnORSc7/ArYReBz3HPcvExa4rAHD1EHHRJP
+X46N9bcB86ndBA5YKUIissngHmrQ4lJ4hyOw4FgP1nWMRGFG72PVTbQ31VDvtNUyw+2L51XbDdL
vKoo9FCLz6g4WKyR7NZ5d9DdBs7WW5qyodzAc7mEC96NRB2XEVNXrDlVbBVWrapCG2ZW1FJAgPIy
LcuSs9GvVZqjZRwnp3mVz4H1OAlIKUV67vRoELB5702mpTzxxXwkLdtzbCO/kXOBWsPWoOKVSH2F
o/H6rRMvN3XmfFy0WU6BW9v1vCKf8nOq6fk2s3hrtMHlWQ1nYTUbk5RNyEvuePNDvAvdWIElNWQG
X4RZN22+rpex5HUoipMzPht1ymkUfvHbemE+3WL2bn3AJai5yMhKWzMr5WkE0TFQ9Ndm5yCe8JQZ
hzFWQc9tAHJlLNg8tKH6C3R1/18bOY3zDqGIHZCcIgSQw30w+LihADTk1+htU8mwKePcoM8t+W+A
eBHVf+c1XrRpF1V3mQZxEBFkgW8Lb+iCXDPpbB95nF8TVJvzveTdVbYON6gYF1ZrMx+bWeyFtjyC
gWf5sL5c1u10oy1PMPkDrc6z6L59csjVOPkRpU2sgXdikVB4d8EKqD10wj0AIh6t44F1foM7lKPj
LHaBh9/Og3Pz9H88pJxfApuAADvV4Nsahf2sHT+2MzAr3OFvHAHvchCmWMY6gFnrrCZkHwk5Apvr
T04+dvPN8qSZtzVUx6gZ3IhjZd2UW7Zd6cBCYrfu4l6UVJ0xQL45yHk7FVciMaUdJYdDt1fr/BIM
DTND24RagAi/Hl7mrkXUVczumHDIWluVu5nrQBbfOxQ2LjqKoXUNYkjNtJmIza1uvn6FPdwjMGHw
Cgz5L+w7zv4quh90yx+T7Mrgdl5updjnwPeYHu08vVmaMuIMg+j6b6Khu4C77DrPKlUSIvYEuifv
93JgZTwt3zBHuwTZ1N/PDMrPGe8+/yXDSDzz71wkOU3VPSK6REkwVcpLRDQl1MykDhCbCI3jVxeR
PMCQW2//QmeCN+yvxcDXPqJFB6cvCDoNoFMIV5VF90lXJ/Q/m9572zGRXninGVTAJDymPXttPext
4ceHCBeOto4iMqHHf8LvN2bLePqEx7n3qqcXx4k7eiWwbmTpgrGN9L+ElPUzStwN2gGabhz01UEG
uvLxZE3vrV0IgnhUrZcWekvz/tFlw3nE+/djCNVdWJ1+QdhfCq33Vw9txBQoS/syHDg9xBRqZyCP
U0Qt8g9DOVZ77G3TnYxz3kJKXESUDZDLstcDPgocYZIBQl8s39O+h4yBpJ8kk8d45k5M4PK3orDf
+2bxiou/1d6Zr7KGn0Q/h1XGIf02BXEuzQZQktteiayus9LhPUAfrBhlAx1hHmCkZoAakTKCPL0a
zWNB6vlS5HIdkvvJz6q58ZPON0L+PFVoTKVm3Fdo7Fyv87A/jmc8bCpilmgnfjymxVLHjgLPFs5R
lGYJxlTM+uJLnn3I9Y5GXBuJgwFeVsJ7fcLpDtrkElwHHThTvPvINEGPPmiJVdm0ziB9YfE+nBKC
78ultTNnUSnmrqIJ8k/j4x4nnLk0AMirF5NXfB249LRhqOkQRraMSOHX55qZLm0REQsK4dYCaoJ+
bS+Pf9yiaJLvNkt3b/gx43GzC4hPK8S4lNV8BEc6hxDarkVQkmZzFbl4diui26jVI+tJnharhrFY
U/ozB/waesNqiwx5hDhS3blBk3PiUOMy9RH0o+0F4o2x34tSu0UQFy7rT2QtWRdORuyhZnhqq4Yi
M59qsSCrlNFtYYddQ6B5vfgJf4NSl+Awi1EFrznphAxn9MU8GkUJPWM0PeCAEWklmChYxaJkg3Bv
LK1W4Bpq0Mk7fRQqaxYB43a+Si0oN4JsnGIjROOMBJHjZTOmas0391lxEVbvebC+lU0v9rVs2Tj8
vNt0P2SdsNO+9dbXglLipOTo65Zvi+bQnSMLMJnWf8h9fMuHWN9SdUMbXeaXrHvsG4Jxk9A977vT
cq8sLFhAd2GlReNVWzb/87OKHqK27ToSkMOcqmQCg+3qLnEuuCuS6ny4pp5akjeFQGquAsCtUUcm
ClhzIwkB7E7oLntrQ0r0B/Wzf6wKAQRdsjQVcD4bg4WsbzW7LEigaOmnOhdhvIXZhkHl7gBjC3uQ
zsuMeEP6abLcdjEOpRY+r4O2s6f4Rv51Nz0BWnFlsu198OUloHOqnMjjJtyFty+Db5bWYdNHfPMv
Mz11p+joAd/OiL3/YZCo6H3hrL/9i3Y+gynbm0DJYUk8GRAMwDTmMRly6IiyXgFU+L+KjZQLly+N
r4YPYrMlsQdQgjl+BftkucqAUWnIAMVW27kTSEcieq8W0Jwamt6nJakISi8UehUMWFAD8GKL+y5n
lqHd0S6k2YzOD80h1BA9cOo6U0yhI2Lxa6sCYF7RWBAsaEOfsMWIJtDPm8+CrvzC14YCKptJKWOd
7ICRk6Fg5MSLy+2o4jRKJp6aK75SqES22CKoPueB34czAXh+e1jbLdtBB1QcufWqW5VWt2T9ippP
qFPXOmFUCt9JYYFuQTd9P1aUj8CNozHKQwBwqe8CfmqqXqy5iLS9rqvuzwYeFUpQ0tZaeOeinCFk
0zSl5Ng0pZjU8ROh7ygWHUgna/T6WuRDmTJWRMWpMMtJvKsd5veDtSzTsuzhI7Md1GKvA7hvHn8Z
L4rU1OnxXbWbTABUfF1GfbEqVbvwwn9eejHZ/CnXfj2kuKko0rIiwAP4MeGzygBSU3PEm8ba45gR
NTunzcFa1pkpenkFAO/GDsdZkdQJc74pZaLJiHg2dZdPFcPQXgOjYD7bky1OXM7t4rFYd3gc4FAN
CoMvelyUKsyFRnFafaCkbzSuPmSKc6LugNfmhKkg1g/W+nERN4DOighTYmAlEx2C7d2kQgDxC+VX
JlDr/fdY4zGBn7ZqPCpqiB8T33Fsi3j6ylNPEhIV5HBxHJrdNADtdc56In2DnnXhA9QE7kGkjj/m
Hrzi6mCyeQT/ClzlibUlZAA38xHZ9zyczlqINN6M+/jqRtlAC/ZFrSHaQQeNw4fQ9dwKI/N8Gnkz
Vm6PRdlsXf8H77MUhocdOBuN2NhiJ3LadXup2xlh/4FMyH2o0lZ08LJ5avRSdRiUsHmhJUKaAJ50
CMb2vub7gvzbC+E8NfeP/DfdJJxzsP4IW9MLKapBD6vd+8Gn82G0iLNGNUv8Cpkn0k+jHN8a6nvb
wENmJs8FnCT9W8vwPP7MvqCyURX+/OI2dvw17AT+r850UTQCqTZ8T2dDxrdvkt67ZX7xRGrTvRHk
8g5sQ4+pAibdm2Jv+Ux1zBzWCxeeu/bBgA6opDH2m2eGbvgaZ3gj5VSQA9qVSpv4tkzx3Cp7MV0g
unyjoE97cvudMlqx6iIKiTGoZJslZEeiDR2ImRghg7E0qj5IV+2RSd3PxVPN/X4XPU3H59rVTawG
ieDuH3K4oJnrLywPZnYe3YVPHabnZ6t/TWJzzwFy7kHyDxULZNVZZmmmZLnGq4rMvB6K69eKZD4J
aIEk9KUnnDGVEZ7nstEUltB9kOJveNuGtt00fRKzOtgdfiEtizqHPxydQWIFNbNy7ujsIQw+QYzd
mSiHjPxnXBDLwONfIM2HiADcHoUY7RjaWvssyFDtl7o1uM+W9j4aKbNC4RISx8p1pBYG0Rz8jvT2
TBufhEuBKyEZQJL4xkL8vh1kn7gQCBpsXVE7hAN3Es4RcnONc5X6ln7Qba9nRZ2e+1fyXX1I1ZWu
w9oHdTGMhNKLsh//OItUicJjpqbujzv4uSoGJLiCVZWmZd0rm7Huh0EqMKsU4c+2NLuZ5VpBe9+G
seGLMGb6hkUZpu/3ogbhT0HMn6LjSG6XGoJ57eDCEIWLZYzZqEKrLOBTKeioWOXXPOenS/PqbDfu
vyU9Yj1dWczGkWKlCQe9PEVR/m1e0hmgmnTNc1sVD3nEN9YIyCxnLjgRZcmg+8Plf6NFDr+FPl5Q
qG/ya+aqAYwaYCiFKB4oen8/5c4RGZZNFqW+E2fnfVkv3fZBWN+7Qk/H+3gXZrJAyRAlgghj7qKy
3zXnTyRNDUKBuKddwIgbQBmUa9li8jaS7gldgtf2+WAO0CjiVa8MtA/G8u4BIblFtmGy+OE0SeDC
dIEW+p9ZU3ycWx/84XDA3VYOcA+fkMUgoRBQduIfqbpFw8vzBb4aN3tlWQchmRg0FWTRzNWJ74xr
nTDiBXZfOTH2PNkGmDjnAwt54+JjqDEACqO1ZA2L/APif28gcXtYfcHcE/mFwgh4Fm0EIfEV6hoK
CLXhUzvJSJcdjAtJwQzl0TLKnkZSxf3mdkiLOGmtUXkb03CfvDNeciESFfw8Vx8g6S5JNmCz7Tpn
qWnZgSd+cr0BzThWsdLeLq6Y5n8GtatXgno3xrUeIH7uA434+jPRR/JfYcUx0swYc1KZBxkciphM
2dcclg1ca4GfCQy2WZ2VASppbT6Fl04chROroDncTxba/ashe6+7wLa+Vk9f98a1Eay6c6QwFfGJ
naxF2FRYioLbBshQYcybA2N0VYhj60CklJJLZkorc60L4eJTwjIFb2CkcU39kQNluIOVIY2QsMrt
t93iPGaUV+cw9NhqcO0qBnYjVAePRoNZe817TqW+gv7N2Tq0QMsSCQZDQ3wZHrCOU95KYRhrm8+H
4JBvKOBoT9vlc/lhpWBUa8HUI2yGssKEDHvXKu/9YuO1f8bNvrF+ukXVpIrDHGNTM+inObUBH8cX
hUuc/cCyrn3zEp2kOCRrVmqim1vFKH/TooVM53J0Z201bEsqcCR3AJabR4N4QYkSvY1b8H41bmO3
GMnRLQZD5BJBvbo2kS19KDJRBu/IL+IyucphtL07cHh5+54Q332vNkdwCPq69tuzfGcgUEYiEHH+
DnbE/LbkB3zOm36fLwtSkFKzrVJaXezeJpSvsBOwf+79tAAkmrEXE0Mk5Uyz6dGywyJeYBNelkny
aI9w1hB/PDV44AnfzLIOMru4Vt7rN8ozGanyGEVxMus1GtOO5Megsynx9k0y03mAjf2FI4TfCyPC
RlQfmb7l1FA+rcGbe2bzNAkREzGPQlglCZ7m7IPaHTgrCKP1O/qYxvVHejg4f4fYd8UIN+KgSTbR
M+eP9SFITACmRIY9khsZRYGNapIGyS5skAx3qa6QBDGt9DIdOY6kUJIDODUPYKiQF6mXynhP3aCg
nNOA7MibvEWFzZP4g3XaSF2enMioGwMjqSwI/vsJbLjxNbnbOeXbR3WuDHdge2h4akSIealI0OFs
oI4goD50SvDS76DX12WniByCMesG5mGbgdqixLLiNewPiLmtl4SsKOr8jLtGA6KYBuVNoBPbisRP
1ZynOwOC7g4yXY9+/Llyc7gvIb/myUUZK18Sa11rx5s0yH2KbXC5Crzzai5wvT5uOgdw+RPNtJuB
i69Hn5Dj0jjVcuigwdXo2QnVl/HQZ/PH4GvS/CneR/AjdwcYujZ9K94vDXDCVQBvob2bvxn3iB9u
W9LjJS9eSHbzzXUuggtRMxzYmIz/ePBmd1EJ9zM6T644Fp61tBSBwuYnJRIxIEtiUg6gHXz2+r0c
ll+lBx6LZBHLZ8b3ayHLvG/NTae/OS6bD1UUO1CCB+Zt4yy+P2OxfWnYgFl5EVAp8Buzz/v2jKP0
8kVDvo7Oi8M/vJnCIippeYQmqQ71GQ4tk/0YX10bFgkZGx8yyd3iqRyol1dW3pyUnZjkCitpdD4i
NXxHEiDr+xnHsmbd+3StJKJSvzBBYdmaV/sgnwS9aCoY7mov1NK8cLrYdTa06dnYDsUmC1/9tln6
2C3Hgk9Kr0mIpRJjWcZDSlrsb7QNI7it9m2P1goX4PQUKRJmDA2mZE/4eYbDypq6NiCIygDXYEMg
y8nOyPhb35h0VtH3zvmtIH9WJbyx4mBp9TJ1hrI24zvW8dT+N+qDdHq30Ltm+VBbQOY7kqQXvn/a
nPxYqC+9Eaqv1iyyg+h52tYIC8pETYoH8NCSbFf+77B2Ne8Us4XD2nrvmwbv+NDQialh9qfJdQVY
JHU4iVLyP9erKKkYbYfCck1TiBz7PSTQP1Dka+DqOEX72j3dtDbvDM8pWk947a/JVphZ42mUdv1v
jHQLUACrgo79S34HGUtQhiU14Qe63ofSvsQGJ7jn75gcVOJnaq5lPKMALtN1jnZqHWX6Xq59Xn/+
XLtoxWGbcmQ8kJ7GE10j0sEnEKLHbumVvodf1w9/N3W7qEHrwjI0mB1pslSMXy7NSbVQRHwQZcOD
37IzQh26EJaPwsk7PvdyAP33D35FD5KSlR/5aanV42/Yz+zcCICnzqI8seXygeePesL8tp9KxRO3
a5U8pIJyBkJNBNTVRc81al7CjK6oOAteNpx0rpgYr5QUbaq29MeQvj3ZCces5b8EmpjPH59lCdFT
D1jVZVbDIoPKWn+3pLgfE4UJws2JKOwWyrKLsSbQvEB6Q6/jflnuBuo8WhoNTwh2vBHTtfYXrtvU
AVNQhESv/O00jYLXGgE570vfevd8BPnIm3P7KgrYierq1JXv1GmpoO/1+38oYzKey6dODItCFiIy
SMjAMxcfZ9ohMIA8ZYnTDxBe33fWefZsEg9Ja3XFmsXAcWeO8PrMsCDtpxp12C6x+2XH7sFTHE/Q
M7BgamyTEVy1N9OvxDtutd2BuveOE2Pi3zWeg6MTW4DiWtyHDekRbHqsPpYLtcA84lXdqeW+uBO8
U+yiBk/QzpdLLMSYPsiRq0emHShUwMkZJge6ZfocPLWfdHZ+RrPduoYdbTbV4Jn/khoTdWLeTDSB
Sy0H3GND4pN4zE/1ud/eJmp6SkQP8ztqaOcKRCja48cWJ+k4/Y0pjivlkQ+kx1UN89j1vDO9uc/y
PcK1It4Zg1sjacTtI1eDo0vKY5HbOvNXkiE9j4s3/HlTgDtWWUUXSUH8UkO4kkBG52NQgbvScRpn
Xf/mBJlByZreQS4fDP2HCerTLXpfhMWQL41/pQpBWE2M1vOLW8yWr8XQO5ZSk4Gow8qbsK87gOLn
tYYbiNGf4UXWefBdFGhYefDNsjlX2jYi4vNTUuFtVxpjr7XaZsKP2KiMxyxMUtl9CcFfqywIMhIH
NoEScRdBQFopHhPbmu5DCmckZRFDq/U/sUjH3e+d3O087Fby/3/wtP3dmkn8+1Q54yCadL5dJZoL
UDTal/LvOGV/LEl7U5Fwz0U6gj2vho+daxg0/of6remW0PD74ADJkEVkG+v6i8AUcA+mFdTR846w
s8O2YdF27lXbX6aL7QycmMr383OP/lILcpc555ThWFpOg7hTIQt3nrwzBCz3hSKmX+bHCqt4m4r5
S/mMeO2kQ6B11fWRg+aAMA2+CPwp+xY0Yy6y1qJrbxlOoBMgeMpzA4hhc2UEenSOIJ4ei3wJSjT+
ZADCVAabCGrApHX4m7RmVBxhzRIRg+BP7QM9qsnxhsDhmhf051PzWTpPXiNgcTryWCAFIMOn4Pxt
zvH0ulSsWfr73E0PIUErjYSH01nY7O1hoVojDp/D6GPQ1/fJ9UOdU7B0cIwF7YsNX62syzLXJTw6
9fsx3jVKaf2fcuiq1gYB+wgov44Sa2JsEaTWPbJdfOf7ASH5q+/SgkCiVzCZH4RnIqLscPdDtR6H
FcoLHJlCmzL7c1Xr3fHxX/hqItqfmGVEmBiVZBuwddISQWJmnwqSqWB73vOTbk0iRWPTHcYi5K4I
jJUOJJZ38z6JpVqvghQ7sTxtG3/fcDkpscmis5imJIqCv55gQep04u6SfgBrQPr4TNFRHOyTW0iI
nVatzLaAfLprzsnqblqNHOcOwXls20PFcB1py1QuiDfJuYqISLGL0RK5PnZHgqCMY2qgvPeu1wNb
3PPq04DZoYD4hRC3akyrf7PFmFlQ2Y1L1hu6c9bOff3ziudLRwES+F2XcXzOhT/XAqKGBe90B2Jp
OBc97NdsRPrU4Vy0EtIvue3ok8cmmiIrSF2vP2cpJuVlSN46zb56kYPjv/r6tcrPJQjnaofHyQMn
xQ7ODvSVX8VLT1lS8wfP/uwL814bHe7Q6UnHw0d/NpzNsUctf5EjL8SJCQMFTd0fNr6pe+O9rz75
8YSXOWt851wVcJ7YPG4lGXGGSqAHHJexZ3vgW0VkmO5bpIzmwNnyS/Egtwc/2Flllw3D3G5aivyy
nQfrM84cA+L3r5q9eDG+8fvEhBLGzxDvTPZlyWBnRVyXkFC2RRLxSNKS+3rrq4jZwXfLm8j1DTqt
8uvqDOXabzI1h65x00sJcHVm6qKxRCHhrAfmu/zlINLMeudB+sr5OwS00v1VGxDybQA5kGFVXleb
PumKQKLIjUjq/yRv6JOhOJqPs1LDVo032a4lXKNF67fR91R8JOYHE56b1kTC2yLtFeCwSzFm9e2u
aXR8ykSGVlAnAFV1YVF/me0ZAy1Hqdsphl9PthhpZ1TLW/JrMw06ZBncmaLuRq4di3yHW8wVXujI
xmYhk3N/IoQuoPZoZ3SVqnkBL3jEvqvplSnN57QdyUgJC9MVTvDiR9L62uwh3bIcjXMpIcLOFvkb
06+cFNjcCAchIaZLxJNFWzVy3RZNuxN2eRlFdpIQ+gPq874EQnheKwBx16oJDHshFLX4ubRm3pU1
/Dv2sKqsm/WjiEvc3TX4lsWUAefc6joIo4u9eNfRIcQVvMZdNbe9n4//wWVViXQv5i2+oinaSTt0
mX5MtLkjs66zpV+D3hL8JGn1vafQBFcjD1zCUMRSD/bvkPk0kfrP4IZ/O6LoZRfzKt5DqlBMedVx
jDfDn+flcFa9xRq9ADIHfjBopnPDz+4Jx1+b8AQ9ALpArFkw59xUbv0UvVbrzG0MJfIVn2Xk7D2Q
MO3gVb6IrnFJI64Z7DPV8ipLvKU74637bdGBsnwJRxRGYJ60uWK+sbXzN9Q8CZPPTjWHy0soDZm7
K3lWUu8jdSvLSFfF0ee+OpnoAe8D0oS9Bjacq3QQsVcIMrdZzHmpqaFVEgLeYstFvRXs4YzVjZyv
sLw5IsD1Ldo6N+9fmU75eBXz/YK/GOG6CmdbBqFCrb396KhWMrinGxk4jqYP737cRjFUokbG9jOE
LSjjkmLMaVN0VX+BlM1TMgk18jrigJbJlxa2lG4qbFBvJ+sKAX+jwM2LasAZaq5hvP6tlKxzr9nT
hWhUUVjNlrxJip65Zqn7S+/NLY0YY8dGYJgs7iPbiOFQUYzXyXJj4eWiuLZvJHh+HLiMMFy6w4f1
8nmWdyEau5sFhVprfrc8oJ0bxqU21Au8i5zQ8dC5RmTWll2Vpkle0asJmVceyCK1uQ1mKQEiAOBb
Dn5H9kYgr0YLW1hudH5ZEX5yEfQpcNt9imWoW3pQcJbWRnGKn/N/V1TtrTLPNoqMKAQaQizoI1Rv
HV4whwZminDoZm6ouoPT+EsfXbLaP/+Ln3WlSTYKx26dKvOCvryCRgOpdGkaw+qRsfpdcJQOK2da
vanzj9DoD2GE1u+h6L3yE7zrAFc0XQaRLWbgYD/LjfxXC+OJwXvD33cu2QYipyyNrc2oURx6g/I4
dKU24AVt5CsAqnQkTpwGN6ndW/KP53j+Hz2VisRBoOk4H5j9ZwxQ9zxRzKdsGY9XMgb6VGGmiGcA
4Z1qzB+fcZkSiiTtQkwlfxXvjIu/uIfmQ0thVpjT6Nd+up6INDpD74NiALyr8RKuOTRzf5DBWGLW
QLohZn+hXegTDnbWcWye/5s+x7280viHEUhU9MBxJsFb1BmY0+++EPUMbQ3wbSGhtxemUGdoTRSN
FtwGG8lTMbAwI2N8t6LlJcPQJeeH+oZikwfAacEzEHNrmToNI4rwItwA7cNa50qjVjmhm7yx9vLW
n5MdsYfwkOnC5BqjvV5ZQspw6wg4Z9Ef2RiwKdu2Q71SgC6a58ync8BSi65zCYWtctumKREWEHKu
5T4Op1c0Lqn4V3CI7Q/gpC54M7/5B+6kaQM4sf1oREOxCEvubdBOTbUUpBrd4DzluD7SLtjEtk0Z
h0bLEK7HE60VxlgYSbonVAmpb/j9hQ0SUNBYUzWv5zbJJ0MXrrb8xYNx5GFn2IY0DmE0LmbZuYyP
x7EX6VdPYCBcQI5EGe7BACYcWCo8hlwGBRb4DLS8rb7uVGSdfLO+i7Oeh464D+boTQRh3hZyEJWL
TlM2sHnFTttgSTovqlIqOnSZUaMocr4taPryjqRAWTX/N5EuVVL+x/aJHb3ab4Lza/2bCLJmPSL9
SSsaNL/O6Z4kAOH4BG0q4Y9beNkmNLiLCjAzFv+AmM07jEdhWNU5rJezLsh5z9SqYTMpHqDZYssF
9S3yb1bWG5kP9wfqM5oZfZXTWjaRF819oa4rdClrAOiS0Yc0rBLpq+l1xh6h7zIaps9Gu15yTDzK
3IW8qVyIly1Q0GOUXV/TUI0AtNLbVPI1jxVNr6Jw1Z5ptw2Q16IVcfM7tZg2kXKAwuhNMzNqzoiS
pKF+bMhjEldjMJsOxTNkpGS9enmJK1NC98VZocV32z4xgFY+WlHWX9VvzhrPUAYCmgW1oTge2e0/
munwISpEF14rbUwfFWAGp5ds/sjOMNxYixPmkJd9psC3MkZzYbPYvQwIquqAMOs43cxa4Dh7rzCE
6wA3qRFkLHZWi8loegJAY1igN3zo9a4ztLRN7VUlZWLwZdZf+9FX3MSFUnV/K8O3s4Svv4zSmYJo
zvyiPdD9v5SELmlUCZSFICzyUnNX29bW9r0wGXEJkIls5paFElorlOTeHisseba7jPJlcuv/zH++
vJr52PiSd7lY8deqMeYmGfr32LDuNwkZBB2hB6zavw6rns3ZKz5G+YGTtfolVOTTBvBHcNwh3tmH
ofwTdPlqCCC7AuQ6R0Nn04THJDmvLcwj95G3+vbklpgsXXOxYvDuAP/J/QfCgU6S32WgC4qjmwcj
/gABYwSlN0I+mtx0NgX4rgQNrWEO8UWBhsRDCatO+/GhOh5vpnwOsjVLeN4pXuzjaAOZPfbdmdbl
QltvErOWFCv6mdHFfsJcNj/FUE8RiCbdtYSxC8L8mlZws7LviNmcFUdOnZYeIFMJVWdWn8so2qdY
XvflpKr1fQeA/A9sThcBZ36fgZ2AZnfJ76uTY5x5fMQzyNyTaMczEAE94tnovU+bHRS6gXE9EfDz
6pIe5cc6JGtJQsOvW6sY4e7B7fu4VYEPybmUOYEbm1C8a9poeSywpXiT4vJu/n11UtBK1rU8smC7
zb7W3gGOxvfc36lQFqNRnGEvcpKdwEX0KrE/aE8mn9yOAFffY/RC+vg0HjxqDwUMrTrLnZLVGCEx
z26lNpgbNZIYbepom174xzmbS1yLpYuflMPmLeCW43hslAu9tz8RTES8QjkhXPkpMFq8C1mrq9DN
coGSJmdeK2721cXB4EOOH1gtufegv3Cv0Pem8ePl9SXmoNWV/ryRyDtEQSxxsmISNCij1KscWkY9
z6lAWRhaiSKAcqRNTysHUWfcuwtAvCCqDtp7NWxnn1/cOwvJlQtAbDvSsKYWoofzwqghyh9wEl89
FPlLwQuUIeRrV6D+a3yHcv0apIcsSZrdmOwnqdjdD01GSETXRc58hsg5IZj3aTCZ8l0bLt1gKpoh
hVo3Wf2IpLiU67wWy+gnP5kIbSwfeV6DMyka0qrAJbpVFPr/Bueqik/FCg2ArPcRS2F+vWjmrpQW
s/gijyC8/QMAwGiEGxYWQOxuVv2r7hiY/hQddC0TbNy1WvX2iyPtRe9EclXLOFWcdf1n8X4tZ/KO
SrlN7bqAesIMdrQhsPAZf2yvcVMo4DHK+T29YCLkt3wMgLo5qo6+yBYVaDbCHzCVJmkH2WeZBirN
wPftjRarPsnmSlY1S6wzS0LPujZqO1lFxMtKeZ5xaqVNa0LXwkxLtneZfLJumc5cDNpEzkaPb9Wm
GIW1uZIXkXqU03mEAW/nEzO5pjl5OWUqIjE29Dkf3F591PS8DGMFj00zf+9XkOwH/CA+iIwHZN7J
k9eX553/ssDbvKXpaOtsn94Icg1b8gNDj64eZBWbsHfa+g5kvVQbuOZOVIiBkp25F+ojYm4fSbwp
4FVZjZVrxXCijrx2sjt5R00SLU9bbkXpuzx6A8D4ECj6P9kXck9AnXGID/ks96qu0mW0+CPPC2sq
qJ79IS/bIGVWVTl3F9LRxokBKVAPAL/d+Df9cKAx78G2HARe/SXPu9JZD4f/CgSH9i7OxitZggrw
+z01Li13apCdsXqk+p0NGhnSZPQdLcLVGpclazXtd5O2NYP+qI3V+7zVtWCMKPGmDhWTpmmfQYUC
FtTnLyeogowE/fM7gyPkOjHasAPSDW+6iJTjfax+/OH72pOPMXKwy5SqKsRW3ltCARIixCYAGHWG
qtnJbym93F5RnzOaG/p2MHjBwwOc4JpTeH9nHTRNejkGi1J+1h2bSeHkV2cJJp4w4HN/PHiaMyVU
lqIngoSPIDdPeEuNalTh17HrbxfaVJSoZ/F0K9ZBW+ep86UCCnZd28oEYrIAYr93074anDsx6Xj8
e7Jk0ctATJgqCwClNUphviqfqqcOLRyG3okxjg8j+E5QDIoX8HVjQ/fuBv9UXxAAIQd6zwHMkzW+
yXoUiTXtPKb31aYzhBIwe9Hw9XaNsMCyhr1xx33AIf75tCPbPBb8xP+FkhAcJt2v9mdTpGmAebDs
vmfV5nbeMU6MF6tc8yIbZyn6qvfJlMa/OTDuAnBatdiOcz5/q+vRb1nB28Y/AuGZ9FL230CBiuIb
JUtWqYWSuqKOLRMwbMD/StdroT7XWNmUkWzWc0wyTIUjdGQVV7Ts2UCQ0kXl6r7g3tEzzmdCcC/C
vS+f41Gq+870/L+wA9Zux/sxVTNBfjch1NoPChdBChbf8ngbKp6Fbe1MPNUjEcDd/Rl7hpPFcrc7
QH+5BwkwBifh0ems3uVPjMPz9Pc44Nek1eVX9Y0XpckuJgA/+63vxyL6H8zLd/QC4FRyaJLtO+1C
9BRNmNKH3/7pNP8mpt9dnChjyGS5ExUogxgWJTEt2B/DlU4PH2+FoENGEaLEoOf34cxrJqYnzErH
9Ciinr/MSMHVMiiwObE+rzPoDM6XQT6LNDmQUeG1Wb/uxRiizDtoCU8FOWKVHe6XP6Ikt/YWMZYB
wlA0UOd6r8h3ruqeH9ky5iAn7WDm1QfSbbHbhivVhtmZRBoMYjx37H9IcBc4tj2Ho15ZPE2BbiSG
UhiX07tXKOXRiOXGNewCZwY7+1BwqCozcFM6TDEKYUBxVpj3FAxgeSUn3n3I3dxg+xI673b9pyb9
YwPF05O/r0EvHP8zvjQRapmyXTU++pLXpWqwqMeuclFypavArPeHttP4IsdObfmbFlyYl5bhZYr2
+lSNv7Inwg933PssPjNC2/Vtt5EgKZ0Yju/aKKahiDWeIY99YL3psMhGfltW/dp68N77bNNQ0s5r
RQvYLnlIJrSyGJEBup7Z7gfYMlsvukwO10KJPe+dZxo0C29gkEbg8eEoUoC+a4Z8mZm0IRQP8R7C
sAAWlmFi6zSpL4/hx3bNlyqTHWMUQ7AUL4j6KhZot4uj4gU0xf33oqToLGny7WY3RVSG5m6AzqKw
Aptd8NQ2kvifVnaUK4L0a4wJnXHDGYhfnAGc/oWuAbNsmpQnxRUYHqIJVw61Q8++Yw4TXRjCcp6t
hBM9EryCHv9OV+qTl0nlVpwzwAwReipt3+dNeZztBK5QLWsr0q9shpO7HARzXZ+A2b+pF8432w7b
Ez7rgY/uDOgztDUa8yfF3ZheR5G1DsQwaITdy9W1X3Cn1zdZ8u4lhUc9/Dx6l5X9lqKhFCQCe1UH
Xm2+gSCesGrjPaYDj2fYYq2gcNFz/7HNykCDK3o6g0ir7GRj8pB8ZxntMIGVMzrEHCZUCq5jfyvH
WwPQ1rTRhH+hUzXn2FSKcaM62e6GDhHUSQBQlg+tLlofXW7xwOba/i7G4jxFuoo4r0MUH9iZukIP
q2yWuUzZr0Apx94Im3so5g08B9eCjksK7N3W+giJATygDdsFYAtxtN5dLZPPWD/sSLJTgSZngZEq
4LbCL5XK2lprrub2g9Br9UDoy2PlYtamwerbJrq17QPxJb2wVI1lAjl60BdI2J3h0svYSZzBwMUV
T9Fw+CUFM3kvPj5KW4jipQrzTfwNQAYOmoRKUpFy+HkDd4SmUnlTmCExzUMinNdNF3MxUOLNZW42
nRHF5RQtbWU2bUWwWuUioappEky+IcN0b/MM3TCCc1ZwyCx88SyBwanRbeAN5sJViyKF6645ruXp
3v95OSZ93kDmX8842tn4cg9ttuivHy/sYslaqq2noBXUA+UpGropsQUWcrYJkw4mT+CLWGVw3Uvh
cuZ7OrKb5WcGkyKdSxZJJ4lRxqFHc0N4LdpUy6LwGXBWAf21KjExXWPLc8RluGSftlenCndB+KYA
RASL8dK2KFDnzHG56VW8x2aBdjSRnQrwVUMrGLKsqYwDPFja7zKHKmk6gzFnmPgPmdQ5sYu6zOPJ
WxLZGBegGKLlhJkX5ahsRJ8ZJhf4pezFmi/aWi5BmnyfiT3w8wl7uhxZy+3WZMcuHbHvFBPpfZfs
0mAIAIVYl+e4vKoPTcaYYkaMga1gWECCyxjilnxz9HcWsHonlTvZTnq4y0Ch2oT1o14s4Tw6somr
BRei8hxh49w72xNGbeKnPNZaHJIyh6s4jZsArf5+5hc6K8CS8aB+5uS1JYyO2bXziI8SvKEH5/zz
J8iHxdnczIuL4Xacrt5Vj2xEfREiIDVMkF4nQO4/BFE7QgyhH55NNEtq4kj4q5NxylprJfwmfriX
Wu/G54eEScahar36KRPBNvQS+0HlNCFF0z0stEKRy0A1gPppF+pioNccRDE5wfqdax+c3pURBIIg
mxqdZ5BRNEyVNW6Vpjkk1NiEME3OE7RZavJrjNQGrXTkCXyTM0Y88/jfvMiNLGAD3tLyZtOcLtTh
Hb02D1BuMxE0juXojLqELwJY0YQ89m+b7Y9R8vKMcq1QTWUMzBVD9NyFW1zK/1PNQXum90cSM2rQ
L0Oypa+AH+FY9wE0Jd8EBDhPIpwPPv55RG7W3WokZwzk95l5gbLzQJtGS1qPYg3W4JLWzClvVWkO
AJwOfQtaaE2O2Ppb62JmFgiWI4nlj8XMe/vZTkBoLPg92KMSnhP5TdblAm03H70br2c2epDVFTC3
yu7GTUXpk9hD1AP9ynDak9MBgniM88lkt0sDYBXgNVRuRQy+LhNVhS/RIMLuo9f4C+Ef+IHoU1aL
KiDbSPUTe85eleinuE8Q9f/nznVyWFETCZ1GKN6s26gZDTrQ3ZiJcRHFWiPjwAqrkA0GaESelxT2
7mfYBPjKcxGVKh2fWQ/5hbcQuLDUwYOWnOpTMoTC252Wl4qPadr5uPea4s9GyefGCK6eVLQg3oFI
Hh/whd9zsRlM87vFlRWfSV6hL4hQ+7wVAPiCU4nDy5bvXCQk083cjGov7XVlv6BhBKaJ5aUnX2pJ
Sw/NSfjBLT/2cVMyGJMURhjN9BF1yRiUyNo2HcQIKHlNS3WAToeif+x7xcCz8O+xYlGhYU9QHG6m
H+hwutHW75U0mT9qMMdFXhpo1BmrA76Jim7vhS2/bWT8jmPK1SPSoDzHV1tBXjllsBEOOXWhGqXZ
Z229Ar4FOU7tkSTKjSzAPNN6xykwh/wyJg8H/qsn/NuyNjD5jLP7wJHUENWqoxDC1Z2GhFHhOs3v
glnjzZ6mvkv3OsmC6fUwDaqyMfl0BRTAOtd9xmqtfHTLqQkn5a2xeV+yhl1VPX/KuL5Km7SWyw8e
W1aBA1CpCMgbahHQIbuh9k7D5cfQOt2Pk3bqmjlJt4onlmyeAjcRDjAl1bxa9g1shBN12XVGzztj
aVXkhZ1jY50/HuldgdFGefh81xj6sAgZbOGKMF/kLJCK+MqUFbQ2X6yL5gFX5USbLVMCR1Llc2g6
CqI/pLAeC0U5hIyCCHUG9X4mt4MPCufZ9FsWIUdJumqyZszY2LZy3WcexHU5HXuiEskJXCVrFN37
6r7Fq1j31SF/Ylseyfy4KDvzJRJl3b87KUQF9/JlmIQHR+46QVIaVmTPJ6YK6fOhp5uWRdv4a9kG
u9sDbukYE05QAR122oktEOGOX37uoCxOy6bMLeygGiSVyJN3pfXdWRIdFFxhkEmnjFww4Tw2Ui0L
HdVJZSzI7symv6TfDWegpyCb0Xa+cY5GqLtj/5CuASM2khrz8/R4uN/VXLVDmRwziS1YuP6i+WUH
Fw99hLBcFD85S3j+Gicqdv9d/OBZMmHXrAbTY3H9PXUFQ1xLU+NOl87aILuNeMRHse/WmEoyEpiG
XyjIB13a0LFN3ABFxeUXE2evXaQKYez5SiTsDe/uB81Q0y3XQiSe1OODM7qmpro8Vam7HbJy230d
5SPMnf6N4rCBifkdYKoJKOfLHnu6+xCt1HnYDOsDpSxtAlpS0eDzkTA0kruVPe0zgPGx61oDlzL8
/4Errrj5IYO1p2g5Am9i5ZisGm2cu68h+qekIHiwovU2h0A0mZp4xqUaohcUbFkUvOct8iwXH8P1
k08DnFS//Hq6mtlzRfiJUPOYrSWnMs7B1Pzd4Ow6Q9IJMlfz31OUqyfbKd8Jku/EpgyobQ/d7JUt
yhfZQqv363RFZez5jT6QqTQK/XQlnD8Fiv/2LcXjN1vwJZIhYHSpILQ+R3rnfKc8RltrIJZlw2YB
CBUpOqoqf4E35cYzbCyVP6iSEnjAAkp2tRjBHxlIEf6cGvSx9sBAOgJzQokXC/HJthIs9ojzIEMn
/K5MahWnrG70UEJhSVvGhbm8G9BZd/1rF11AXQAcpPw8Eb40Ki0EULOSVWoGdwcywBVMZYMi6h+N
gkxSGWXnnM1IDLCcx6lFbX/fMoU76raOp653KRDtjf8Km1+abuThWi55lPY3qlwyd7VJ4OIW/mBy
de/xgy40c4uNm29bMPjbWVjWs8sbgiuUmU0GgSBAHEETHwAbWAEDINwMKQHPb2SUrArtUDfG4h1G
fN5w+4AYTmV8eAsyMOJr2Cld60A1sl88CEt6ZHjSq6lSF4c1LgME2q2TG3Mr57Vn5sqadZE14uIs
8pC+330nZBTvdjZyW/06fkSHLQPiGRPAhbF8vQTGyou+iA5TrzRhm9NgH+4WTWljh/nSRu9wFSd/
Ef9RaemsMRxa87FO++I1OyVOyG9EU1aZ22oJmxLm2wYYXj+hHHIIvZ77r8KDkfXdP5lt6uALJOov
n9f67j2dqeKG/7pjx2m3NOTlOpGTWBq//ZnxsoOXyQubauIzCo6khtKEpePJKuvx88URtY98D2Ew
FG3OVhqt3rDWG37ljr2MYfHYVAxF0ujjLyZN+JvNFep12b8+5BgczvZ/niE3i3GEbiJpG4XQhHl7
MzisgnaKJSz+bDjjXRFS0l3gnADY6y93mICXqGycwGcMNZCqP75S8rNWcyBu/Dszp5d7AAw1PIbA
lUS2J5mR9Ik4UjIsTKt75yjdhOJk/ZfXQVfC9lAfkxVHNsdxBUQcO+SiN3HbsY45DpoZ7o5fjJ/H
0q64sqvCIqeTdYDXMWGtTiSNJgZM9zNyw4sVlXgCa1Q/wT3jPFL53HaGwbdQCT5utLYYvKlGo4KO
jAJuaKgwUh3/fMtymyphJb6tdGJ9CLsAlJfP6qUEQjOYiZCP70IksCCIoIPd5+Tcs+E0A01BZpzG
+8SOE75KjVt9VdobsMODMusb/3m+PkcY4E2Rc6kv8qI9RYsjjoqX9fkCNT4CrEavpL0oWYFW2lww
MvehGK+U7Ji67BGuXWaOROJ9q+XJzRBTvRKOP7txGLJ5EEJWYvGkRXf31zdv9qvpiL2wDchEJ8FL
J8GhfE560poKfndv5VcRFhGEugbSmF0BLuxxU7G4AUAmL8CS6q5a2s/S2ZIM5JIYtUsRbDmSmUJW
Wbqp6PVTcIznJ3pJ7FMEzfO2Odu8bylIoiImllDPSgJmBGrg/uE2oS3Yv8ioyy6qgmZH34lZNmyt
j0npaXinv2Fi21eNEd6m5CscE7S6JOcHHdhEJgOyYpbj8qk350b7b4WqsQ8v64oL9JeVPLtT/hdR
YQtOVPxMiinMV9GGBPdWvThp4QMlNvXu1U7Ff8MCocrOWmuoYfSjeFfx1lPEESPaJLJWplTD1esz
KIZ5t1AmE1Zvhb0f/7Z8H2ZPk2N5oZC7TgF1flMZaxfI8bGktH1PGLtbwwP6G4Thf8Xw4fVBdLkY
44xEIvyhrIalbv7yTnb2PxeMG9h5MRoWhqqb0eVNmGXiyx7WhJBa1wyw6ZXYjIDSIfb10uzfubRB
6hfaJOGN3MwBHP/XUBLeo0Sz37ks5hl2I5ieJJNDuPBG7AfEO01DHA4CcfVpDCWj3mr2iuc/rtmm
muMJJdrZTYUbkSiZ8okpfI8GmVhdk7LovAXM+cShZCCeM72oLL1V9xMKlVQ3DsE3Zo9nzcdVYcaW
zvcmc6ii7wHTlkjYqadg4yZmuvdo9tD9eYlYh4kfpqBnoB76/AVDlAMb6d0cQAINdnCD+pgtlduh
piBiyUyaMAXoQycXfwH7M0n7nSRWmUUHPS1mDI12vHIobeaSSXQt8cH4dK5U2GwaKNWt4cDjKNdO
zj+8UkUbNI8L3SP/WEMr8V4jbYlgokwpRpK3yqiqqY/PIubjm9AnQG/CCM6LZ5IbRBao11MD3nxi
JWrGn5qVC2XbcPGtKUy8tBGZ33tzNtRzKNCfBSF0EJIkKZXinrETtaWc8UnB6IBzm5cSJhMEg1mC
WdLqlEoKrI26d+Wip+H6MtauHRPiakZ/dlPkVhJqKf9QmUzWRU6ZummohIE+Oye3oEDt/aEY1615
AMTMpRHviE65r5ieYQtyJ1oW2NZr/Mq9cgKv6DAQmeVwlT/AdKZqAn7cgUJwlK1S5/CKTd9Goe9v
YGHAFt/7RLnQuOHm+LbhlTWbQBJd1b8qZLZXvcavy7MiPaUHeZWFCdllbZbJ8eZ41guUw44SWJXq
kcm4E1nbVabvDBWemdLKQevw9dKeykMF/qLgMBxWww73AD9NeML9atoRpHNOVugCcbo85CvpWMd4
gcXWEHu+RzXvQv8OgjZZjjKYfiz+3rpezBgRCGEJ8PUbofvVBcHlKOivXn1Zi49RKho0hATuuyky
BDTpoe560iwWm1EtC45nDnCdMjwtaPzsK98YJKeBvpRxA61cOKbYT7349cLBfTgaqirqYkSplntQ
9rQ8DVM72T09nkvlw3r/mRD2HFBpRrO5aIsrlXDh1yXxdBDCu3E1DUrvU+Pm83NNqVevg8snSygJ
4PWWII8HnX48vF09LH0XN+9H8Msa0cs6ci9tTfShgg/zwMIZEk13916muLyFEoQiImJLN0Y3MMRR
DoxBWWP1ykdIJJL9apbDjNTTnpqxW7yLuW6ZddX7v2We6kJAHbYAyc6hUm42TxhQaBBkr2dCIqjd
PC/nYr9+lSZIu6MdV1ewoP0qfRbgyj32cm0M7DjP5luG967/81AWABU+Jwvk5TUQmN/OiZ+yLzNY
1C7B8Y2mJ1N4xTq3RuIx/+8JQKRi9Dnh2N2R6pBcwXy+GZROA/x0V4Xg0MNLqO1iLoSzxbxOsNN1
jDIyoxZd8DAORY4QX/GzPLtt6g2n9ms9+MXC/tAD3XV67cFZiwwUpjTc45eafScotlWEtCtyCpEa
Eb2vDgBlodELioCEgS2LoqVZunCxL2j7gpEhKo6Yn9QaOiPqAXMzBxGP7td/tQA1DSYF84Zw+3th
fSiTHZ30sdPxIM9hp6uW/1qwX/sSbiKvnZ5VMfu4sFkN2M9jGDLxfTqWtdC9UrJ3rYA7x+4r1wRK
UC2864RKNPVActNR4/nM0IbaepwTPfTip/pTVMbnib2ORMHXlgFeCI2uYJkYj/YU2ZtGuxhHXxrV
LDaiEFEreF4kti/4RDLl/gc02PlNaTUOW0G5p46PP1IKIFxxk4Sqg/J2LeTMG2WeQcj1WZEnIHlo
Zne3Exhe4v4TwdE6qWpmB+C1p1p+Re5wgyTWw3+Ik9zrKayhYiW7gczP9WLFPQu9w2m+9cMXBmVX
tpui/geRnUcuOyzTMpkPN7vTkVFCXGi+0S0TdCew927FuDLH/ZW51X6mGhmqKQoIC9HP1qSTUz6k
h8cZcdm9X9dN8k2XQzKJtqmf4o4lm5lKEiBylEW232kac9oTw40qN1f67JzkujlBnbrY6Gp8Mnvz
UHhnVP7xNBXBT9CPx3/oGXyLXkOA1Rz+69ymTvXAyzRpLrkyiFgVxgeSduKnr8o9tuX//btfd18P
zRGmY3xs/XEfcmrRlEOQNQWysKhHVLGJXQkZyXfeipiOAb0HLsh5+HWio/7Ba/h2phMxX+zVjz1t
8EMUveOA5x+x2U8viqJplHLC8L6+sT43kSB0AbEgjxNqcV/ecXPBEyqtckmvmPduaqC3IVF5tihj
t31DlWe6NKjNHVTDxsKrism3jENXZsV6tTJMbP8MX2QopDUu7nkpKyjaIJBB18QOj+KVvXNr8t+4
BNKXyw+QOXuXE8o//gq2gWHzJYk/gg9iEuNgCjgr0xwcIhPJafc+BHoVSkPiAanJXhJoKBQ4dT43
yIsn8LONGgGaLnmwRNhObOpKRN3F9AJ0waKVnkkh5LsK0SIoMpocEzmrXozF9VVIz5ELhpRRGDRs
lGrVzzDXM4lYKalh2RyAbeI7z/teBHQ1rsDGJywP7n+nrkB/KCw2FbpeKJM6qd/3kzRWa31jchTM
RmmK8rOh94V8Yodk4C1HQSlpnufC8EYmR7FjVuNrRIIx0w/QTV+2fe1na5NQYz+arZ4jemnvxI7f
LAjYxStkRTfBKMrOw6ELFqyW8ro1cZ2ZZIAnsWsWQ72fTz5lzU+DaXnqjRBgGGl3fSGP759dUdSZ
6mhkpdPM/yzthZzqBlIkUeAdKc6Z/LAm+sGwTRpufJ7GrApOKbrMmSiVXSOJd1LDp30ga6DLVHqk
a2Cxc+10f5++f0wXy1nC1XGDCbz5uPIJPQS5h8dftWtf1ucjrBfhr2JchTBmSfOlpPnnNdT6QHkV
0gwX9oRyG7u+xADoctVO+zDW4tC5NiNPfvsjztX1zr99jOcctBwkiCU25Mr0EJ6B6a/gqo9B8P7f
KXv96U8SsD/dtqxrd0kkQoFnRppTTDA8UADA4jrL49cOrPbi39lGp3uLTQIk93HMQpjOoZiDKKku
KlO33oJlF0HuchYkuHz9PvUsQHX/ZcILXL5P8cOJGoFYViGIginIeNR9OGenMGvunVBSNLn18HVr
nLl9IAVSV8ca/jGdwkbBIDVT+36MH9vsXcgxkiI1ipORgDwQQZq/bk6Gi9VNp38yQLLDi2VztUsp
iy4qXuY7cfqXeVmO4ssYglM4rXd/rsiZJN6IrU0k3hKkgcPNT3+M7EgSrtRyP7caLtiYZu5Ijyna
pKy6U2fICtYhvTma1s8IPfT+LfBkBF0B67oWw7wvOmlyswG2JsnCua3pJu0JQWA4mScSigUEEsFO
lY1s8b89AjdkS/3G0wb109Xau2MEcyLpu2prIoiWar6nuqgShPzBImpUyxxCRRFM/VnUheFVeJZ6
ls4eODOMtSViPjg71/PGblPB87eH6A7d7lGsVIswMLHI2t+VmLEYeoMwY5Uh4hRwsoFCPyyEf09l
5twElXpzMX02G3Ozie4rNN/FspLYY/HyyvO1AtmHP5f8qRqbXrpTHQli7BIWzjOuv22tvDZRuCFh
IGznmRlC4jJQddnmytS9YMDgRl77bs/OZ2pQKqy76GPpY3Cn20nWKL4ch35JAyKWSDQVr5uXrHc7
/EAgPnxpXGMFZ42qsjJvqefuGIlvREbzPMkihWMy7XiB9DLI0oqMf2Oonsms569BC+gC3cK/I3EV
yRRMgtyPHHDSdHzW8QFCvT/HBKdHtsVzlIbw8Wg2L9MHlVVHXyzyGdVvMJ+XxUcOfTaIVu8bdiNM
pBhIO6OZ5ZK3CDYsyt9+K9EJiInLNl3XIxssbJHk5LiscpxWMAG/H5iQ6Pe23G+7tft7rBzpYhdX
eOVHzp27i+Hzd4T3v26YSoxtMK/UpEYESWhI8zPyLOLUbyfI3c1/SydPD75+ufIbI266jgaZMOzJ
lAEO5svtcatyRHucTc9Cz9wXGHF54swz/lDvrxYE2KD8HqvyBaOXJ3+otjdd9yFvznf2j2zBEnLb
VWSjNIzibp2YZdsUYhjrwWecXsWIgXUOOGHBJ2HaWwcMzsSdembalLiEzLGKwtUHe2/vxGuXuLU0
VvUKxaTKQlEAPqg4a6yWsl0YsRQByxmguqv2yW1WMtzOMNY+t/GuvAG8MTnKgJEPeqHHXDEAiEZ/
Pp57iGTwfrDY9Vw588W8GuJ7VMYQtd5UyYsJMNGyBPifhuPmB7ieJwEBbIhkk0qedQA61fO4yvPA
VQb1nECKoVm5XVPrr190gexpMHi9TC/jKkjcBeNsrriwm0jUrX1cDDptFnBVwGeoRF5gElst0MQL
pWCtBQj/yszLWe31FscsOQDqHaxMFHzGLSzN19HzyHOoNv3421qfXLyn7+1DsAQON3R1MackjwHP
wgHYf5awOkZR6Lichcf+SKaVvAoA7wdlD23sqEmSjyaFRUWBzNVfHo/fasBgssj2kHTsUkDvTgjP
ODcW6FXMHqxyf65hnDAC4LDrSusB8o6Cqpnf/xA3p0gVHU17I2f/QOW+DhePKc8eT2claOcz5mNU
kjtZl6B02LFG1HQGUwUpuMElapztfiVDwz+Z0cSwCBycD8gDwksMWW2O6X+WiexY2PpnCUrXpthz
gvza+tFG6AWp0q1g0vgApEZGL/yyooG3bkoToWAyI2S1E+yf4n+SQEeZyHTNys2aNXm3IEy8fOKD
6oIKqO6vFfMZgEadk/AsUZKflJZtuoZ2atPlHDlJbdEmxXRE2TcdOm4FKCwhtPznKFs0GI+/KlNR
oMA1ioLWpzpnjutmwj38zY8FV980JUgp2LhyJzY1vWTdzvEuU8Du9RcUK43uOqgVQt80XCjwLg3h
wKMCjbc0//DU3SiJRFp9veaHMreahGrh6C0eR8pCrs93IT3/6JE55rZEJ8McfBCDchVZklZJYIGh
dTFnjGUYGGdrQGZw85VVQ3M21zgh8DzX9NlFZy9suNrhvH0ZScZUo+/ixeFALW8Aw4JG6kJXdzr1
hYgGWjjCzBYtfsjxe1CcH45vTbvWNHEidK+YlvRzGkU+AQLIGmHx0TNbPqmnPjtAkR747kYXbb+F
ZKQlNQOom8pGo/Y+F0rVWVHD5qi9cX+Ipsf/uArnZiuWrInFinhPHrST1Eqaq7jQ/9E8S0A0ZWWw
7LJreVJL+nbb7DqECh+FQapiYmWGaYW66GkXHMBm5g18Dx56sy1h/j4rMw0Z45VIh6PR9IfMrUDX
ZFesQ/ag/gUesKKkVJBMpnXdRTrj6a+R7lseUe00cjdAWlWerNuGNEGBH1jgx49ybJ2x5iv857xm
NEoV4dIA+KbkqHTi016rDocER5IqbqaV8eej75qgrJCd2SjUvmFB5FdzKf6/Phr0YgP3A4xFhHDt
dMnRfA1eOSiswNyg2CazQ8SwbRvQFuSkCOqt5TJ1DOPu45l9upmItX0/qU4MfjyMLdqCrjOR1OJf
167bEXvZNAlcUNhgYQJK2vMn/WBYRkDL6GtqfO8dYaYuuBdBIBtFPiz4ylAUshX+98/6nAzkq+He
rc1r1/jwuyc8PiCrcgIBFfbgJy0jIEuTP4PBI40s5dexY576t7VNbNNoRRbkXTXSwRmVkoIyBlyv
18+T9HSCHnrJy2YFppl9EeLHTJ29bgDuWTkHzGJXdfNJqw46oXr6yuNwp5pTX51WXqwDefw3efoq
LSt+TtO+lt1CleYTnaSxnTGSVbzDd+ZLkd4XezdJupaL/UdWOA7LK7T7ctNQ8PpiC+X9bmRjQPlR
N+SDEWKsE4kh2gDgN0gkZ5cZpbkvNfk9CZLKfTgI0HihN3Ad4d2OPpC0zwYUowS+tXk0m3LqBHVu
NgRGBg/pNneJhu6OIpP8gczGwx2gkGBUKCKGv+LGqCMyO99ZytKDJgtsB2lFo2iN2WMTh51fxeQ1
WWR/wNFqPme3IvPRnq323wTPuFRqNMbHe57qZ2cP5dbZl0tgjaxrHvFSdkDkG7epJSPqeHBL6/08
Kp9uKShsboTPSe8tQwTz1wg1at+MwvS1XmnNgUtEe8zAvZlU1wMKNoOBssbRtYi8AbkhQr9NGPbh
AiNjwnxidirAMjc33C4iqW42ccE9ytpcvISE/HS+6EpbqAzb4Fb3v6aYqy/movCkFxsnYLoYYGRj
IdhLGZJhrrH135JlV0IGX7YM51nxE3OrGtpV1Uk983RkovDLmv/H3o8w/I5Gbl2NYAwANAgMe6yM
IlGVb0fpnah7KnuMdXvsbI2lakyt2eW6vxYBRUkwsS2apLJ5Ts43+tMWmeFbd5NKXjB2BR7frwsK
yeSffBM9a8FWvUlkTlRijqLJ8Opb/lGtRXWmTS0UytyJWwrgaSjHe0ZUjsNZ2BT4YSRpRv14zSQ5
Jc2e2Jv2ZMQqlWFXRG66VvAz6qpMd0J6eiFou+FaDhDq6/c5TVWm/u/ZDdznqBhsIwbguzMeZLO2
7dwyqBy6n+VTeMBdkQ5VaSlSw9voSAN79BYY+o1tGl12XeidDJw6kbuK6VdrRu+TpR3pyPY6pigG
W1D+D58SLOgcjClX9ekFEJhH3sXrXzTjKZv/BKVTKmLWGX84NmPGSxN4TS5xPMCWoq+293rYghRa
yi5D2d8CTtWQkIuunrqPVtxUViydNaUgGOnaFjdvpu7PIZ+UwIkmNMPWLk0tfpCNzNyZfmOrNw7K
+CYtMdu+/8x/Z/B5p7cq9r8tvlz5GWopD00LKX3wQY/RBzJyji4GYAmzkICiX7XvfNvG617P8Q5A
e1x0GP6sNR5qqF3q4hdPz67chHfkA9g9+jMw59/xlqr0IjDgF44JMpyz4Qw6ZhwDiNz9t+Z+hqGy
dAcqIQ9iaXqukBFymnAFgCStWOtMtIej72xgoFwiP1y2t1xxjHryr0i2tu3IQ9axv/QtaUfkDTmf
vduMBfFoGkwQWNnlcONmRBDFvN6d4FmIpmivd3//LmHmSme0PoQqbx5EfV1IzISN3Z8o2lPUc58B
6tP8RClSSRr8nSJiH2GNXfS0DEknqbpt5VwCdIkj2JYGtiXuw82wZja15pXHXDkZhe4aM9jsbyAE
rnnncmNuWda12yFnWxzizTRxoUuk+qqnoGbSYZ7eaSWA56rHnj0/PrzBI27NKO5OK5j6nEVYTEru
YNyunaBaHMQVtUm1Eq7H4VSOeV7/Ar17vtfLTugajyNiFq87ONjeXkSHW9ZGbZHeQeVhPuHwqgMQ
qZTjfKYFPb+ZTO3nzM8Z+7ztoLMwCpNiHrW6KDehi5M8SiXF9cCYu/HcSP7XAtTMIW+GEzAIS4qb
YR/3OvPapt0xEeEOnwNgfCCxAihTuPRI/BgiEbiYYUMwzhcHu6w4C3XvkVarfrehwmJwx1deXx5x
RrVzlghfFg1IofEVfGQAzMMX9xONlGoKuwT+DYDDKdcM2laRSeix+Ay1pqSUssY9UF+u+Tkqv2jB
lpCqcSU6Auh8S6pCwtwsPA33pld11qgdD3Rzz6O7dbMayqduAJb/97kdzR/Nr7bAi5NQeMtVeAZR
SqkrisQj5UZs4KbGiLeCcStOPozwBahgojKTXS9fH2NnHq9bGzfWZQHPPEi+VWriY32dK0VMkeTZ
bORa1okWCJdTQ+UX0KDbR5yNYsTXDIRqIh7mFC9xBlJTO+8NxsdyYM3N92mvkx9m2+J7FQzaUx7S
29mwdMKWKGc4WiLNvxVYLmLiuECC6InP2ek6OOTWwTxpFMIbdSUecrqitUhGmdlX+VXHOmZkl3DH
5XBDiVa4zVi9ZyXLpByo3vUHy8dOwcEcrsqwePsRyRnR+QwpV4zNhQZJF37Mj7ShlqLq8kRU52Bu
H9oKjprMEdsHZuRdGWtvuu/ykAXn42mx9TOd0B2WhO8oVXvzOniYkpn6duAg2zx5iNDEL6+fFvtY
kRVouZM/WmlN2hEuqk2ha7Qwl49aUxFLzHtHzKx9haoeXCGgkCDV31QgMj5N31yr+O/m2AqySVZj
lVBRG+BxVhED08ZFn/EbmwZwUBIPA1WXS8EmmWW9Q5hmhqctgG8OqQXLiLEEbrbLokJ7iZLcnaUV
5Xqy051AQBTNfxavoiglq1jyLYkCezHIs4syxmsq+KF/MQ4QzPUbbJmdOVA4LMQ6Jj7R7cq2ALtu
cJ0Jb45eaJuFY7cp7JTN47145bvZkM/uMYf8CvTlPrkDyLCN8PaKbtkdnRN8kuiiBagHjGxFOH8P
Rdo6MxIFDiUCv+gVON+anV+OlsauTWSj1JmP0u5yvr6obcuVpp3XUPlCbRvqVsNiU5yhe27DxZb8
ksIzj0HHe3icFuPBgz6x3hfS+eHTr+wnyuia6uIN/ZAhW1vfRNKWQnk8CtxCwfXcdWjAJBmBEWHR
5AorEArWkbPPHAUFAnZPT5gdWVknxTThEFywLTqKhr1iyyZ45QVqNsCH93m1nweCWg8i3w1QeHy6
VaUGUYfbsd1bTFN4x9khnhbayVVCf3a+hjEOH9qyL/8v7iaa6aLnXI/1QKtMm5ddqlRe/IM4c2xc
FXz9C8ruSy8t6gyJqnpZ4kK+ZAEvLJJNQudwmblas5Na2/c64Hd/lj2LMRbQTj8huo5fihMzIuui
TKgVG8/O5XcDYdvp4xahzti7nqbpSgkveV3uBTpmqYYYH3XJxBjFE20InZ4ty2yis+Cu4OJvMiK/
H2GF+rsfU7Qa/duw0GG3lpfmxvIZVXlXShXDVjM1IbiT6Iw3VmHB2Ndu/sjb0r8gPyQJ/KQ3wqZz
DHFIV+Wt3OtkNZLlni/RA6HPc9LWkq3XKM9mP6RsP+AI8wj18PqLdI/iyVbEoSyGW/VeEG4U05Si
gqK36oLSnWIMfgfEyVO8FMoStXFl2gEGvRLllSclqqY+NDX5P2uCoVua/c76VoT/nht9CTObvA+k
tMaZCDlos8WZypUv0pExEd+GLmeNQhSQoJ0lcom1azfT72fPrtupZHhbEDNm0TyZCCR0AX8obJrA
5lX2/OU93OtrJ/bgjlWOPzHPn6gUtq7K3N/B89NaADHLeS5t8epcDszuyQ+XT5o1cDMyIxga+Miy
h5o9kDlZ6G9kL+SHqG4cTmcdfNiYhxroiJ1YMFyj4JA7RNLHapgfNN8pCV2+i1OQelpPZ6bRvto/
hja7xwMWIcy5iSE6oQd3Q2LEIIb2EorWuEVYFtbAQj6+aeKR4/PJy0uCcJA9Gg877EuAgfnTKAX2
i0j2PVS8MsDIzB5oHdSJsoa/GtB62qiz+Zzc6haVsCmw9rWff9U1YwOUijzF2AzIzwM0eETSLMOC
5XmoJxn6VIL9rFA/hMGGKmQZVRvxNm7hmmA59n+/d7QUbmaKw6MhmjyyyoeLe6w+m63NRqnD22XE
M3TCnXKtCQmSnTgGUC3B0smfBHrU66VVMzNuCtx9WId2sKBy2GQryoO3BFGsckmXh3PuzqgEiasp
/IlNhsjxtFjwIDgFb6gh//9OYrqDSa2yCBNds4iBGX6Ibj+3GLyV3gkUn6QUNTIqanP1tFr0PZgH
cjoAkqsELmlxzsWgEdv3gmW7791dj9GDLKYk2P1FzrLQ8FOHbKEyQdueGHdZagrgcvAgtcIE6b+v
MdcZG2DGYdjRlH5qtl/hDcJ9t/KyQbMUebfe7ElmSkV2eHjE/yI5P20OX/dnh6TNKnBbvS789JBi
amuKKyfqS+C7L8t41hFHPmRxLkctJ0Agta5rr7Hu+sUg1V8kKwuXxJX/4IdfmvuJrXXLG3w1jIKE
TXSLJlnYeAPbuTNM+2HLcdpAIXKRe+/G4pdGCmFKm6tzYIFVbovCpTjq6rnWuosZK4GGP9BlicRj
WGBbUlmeYF2c+zbftKM8KOJeJ5ZS8bSU7Oe0e6OLCnkvVQJsiPeeHDTH896229cDcCgSRoeV6dJ8
gpG/E+iAJzzIMh8wXk9QNwgs/ll9OFthBbyoculHX7hCHa5PHsIvF3iYYV4mtRibzzW9s8XeRb66
Tpy+wAGpRgQ9xQYnifjLsmUl7cI+Z4KrrVNs9zCyzN6NF51/xx54CJiqdgo4FLynPokRGh87rj8m
z91JbWnFbv88hNYBO44ag3CCcvjFtSgMGRPJopEGqL8qdCQdxpWA61Q7A7My+gDvAPCqbe4vBoDJ
BUiZqTBTAmAKgRwWZ9Goabs2+QvxXou/DCihoCpx/xX9O1gTHDBVWWLh+E3yXpoKusurvAJqlb0x
u2DZH5TbBpCcI0prSJ24buhtJMclOGWof5w3eDnvX19aJzjHqr3Q8VsqioDtntxNrkwf4POz7lnr
G81UllXn/0m9T/cmPuHQNRa2J0x0SPYTp9mvPzU33ENL89l+ffqSY3AG5qpAfFpFP9OdrlZsGWAp
h2oXwDFvqmLPW3OcYQWEh//hBvccRCbgiLvbE64LQoL6rrY7/gt0O06aNFdShtRHmMl+MVvUPgnx
8vaUgcsa6mCyFU+2sef+MLxd3yjApkO/v828lbImz8fmjjfC6Sh+BWJX4ywKLsterNMn/LDLQZ33
mgQ8fIACArRXA37xPVb/HNbfg2R3AXyJnCGvh+EySk1u7lDhOJafTeVs3kayGh3hbfZC2avhgHBS
Cvo4ozL0aSz97RP5wqxz74M1cuqzCgUQ1IIvFDFfKTWgVkKmpVsHmjfU0qTzkHWjXPpMfColE12c
RHpsDLfEdl3K+jXfM9Kr+QllbdJwiCvSR1mXlDcdlv3GKokvkdNw+t5pdoOK+q7YS8D4JFhrUOw5
9FuQMlcEFD7265YA1j8LETE8oGG1RMqNfzbLMZ6jLOtyfHQsM3sDvMATuUvk8ud9Xl7FqO2A9QPz
oUUI6WkA54bPjC5uopbXstfEAI4s6RJjD2SDzmARWbuZUQHdjEmDQFGvgApRt2G627jWruvJjGGj
qCBjQjrXo9cD+m+UJIDsnGCyq7pJins8wBAU9NNS7xD/dg1/Idy98wAUpNQxw+Kg45LXDaptoj7r
VwxTP8sOgMb0g2P3Ze/slbXDojHeRpn0hsok2i+gpzX6KqO0ZnNpXnHEyTenokBOuknYuZ/gxkb2
rwLjiNBZ0JqasjmMUSOMIy2/5TO8VH7Qep/l+7+ph4AblWLkPVzm58KTjvlA3AtTlal4JWTLr5lv
RFu4Bh7FtfUd8vDuWA3E2HTTnjCSLRDRsuNqIasldicQGKehBRF01h8a4AYqdD2vEo3gp5T5+uhP
XH0cnvcj3I6roPIsWcRoJGHd+yk3mM7ZA7S1nltXeg9zhNgQEYxk5Z16olDahAmz70SAdTRvqOXA
U21pXv1Rb5UobgqtSYg0fB8UhjcgAO1NRQGl62USdEXAmRYL8+2brYG3yDbVsUH0qpIlGNVKOymI
jQEpJScScGfrmuK5zhWNSG9gktzc0IvWucZ4TK0pAYEQWq1jZ3R+0/yRBiCjSei7SWsbmb31mBo5
vXDfuesw5lTy3wyxkzkouyjGCiSnROWxRRpe8ARpiRcjuEA7vYKzZsPv4HWEx1HXBDJuwfluCC5x
EUQq/Kn39b+PxX2twBgk/4ueTA+ImPAo61ZQkx3lXuMUzQZkLkPnFapi3tTLMxcMLAdG1I8pCatP
+JVqTHmDEJQLA1B524/aeheZeAnGUax0HrdJjv202myHubbkU9b6CiFkBdbEQkhPRSOonatNUgCk
9fexVHVlQbILGfGB8OQ+LzSv5COqCywDGa5t/gsqqBJ1RCWEWj0PJX7Gjl5GtEVOLERhX3nysaGf
IXvyc8pNxPhXWpk7i51c8mx1T61XhvDzhRgIkWNgjKsF8mAgOOV0Kn4qqc/s5znu+mXV9APu8m2s
1MayaTQRrg0IrHMHSIbM6yP3Lg0HDhg99S8ewU3kxuYUfPYnlWgVJ2AqMnhv3ATu7xGID1v7mHMB
3F+LvUmJThf7vqKxJM49niZvtW7WEy8Um4St0x1AUUTIuaIkyWzlc6s7eOnfbI6YunwezrcP2Cj/
ihXI6gO60+o0UeDP7Y5Ac6AKtM2l8x2lF+SxFvw/eMjRDmTCYg1k7zuSt9iuIrJbkyPx0SdU74t1
keCzAIniixFDZ2bc4hHqdm6Ls8VhyFFtK3P24D5UsQju4munXLI1OIGcIsmSrXnMegw+U9KuDCi6
1FOpqw0bV/+8v/hsVYFti610pnNZwKe05k2cPAl0UVh29uDNrMa6l6bEaFKkzzutnUnHbk+iQhTi
HizTfE1RT8/ktD4kyfkufXTjRBRtU4xAfdYXIMFbwcTSnb756rQ7HClZ+GcWky5ViYYzllRu0Ha7
WwH7jCuJmSb6MGdqxCBu97wUEUcPZaB+XBGEfY/zUrBJZ5w5Wb7EXVWyVFCojmOpTjTzCBK/6QMx
ecZxsp4AgZ/hDI3gWWx+ocr6W1Co21gAQaDbyxKuYowK5Ak8gHn2SfRc4Xv2H/kWMob+kTBRCBIk
cf/kvNgOhudysid6AGuT0041CRUG8LNBK+/az3WDiKHWdoc2TgvR6q1KREq0L6ztErmP3PxokAlN
hjlEe4+kmBR97NQLI4rIesbI5j3bRVw9+Ahg6v/Xy25k2FZhL4urdyHY+5HzANL+l+lsrxEM4Nlx
3dOc7R8eBB3aBTwxEmG4rnUgbvo/12PzyVi1mfXmmAgBFuh1t/vMToOqDRWkf1k0m2NSZBP+ke8H
HFSiUzZ/Poxl71kOeP0xDtPDonQG1ByyOaTC7sQYeHtf9IZNrdwJQIYdUJpDmjfBxtMTs5b7Gmoc
rqF5WSxNmnU9nqUHAoZ0sv5B6TsgTHlHpTdLpTLXXTlenJMt8I3pAd+NNP/cnN7WaKg8uaRrX1P+
eQc3XXtae0bcYMOR6+KKAecrpZn2l3t3/LsC0xI7Oqa7nUuDxEpeWmil8w48xJWN5Hb0IFjtzAV9
CP0dXY9lqnHtDRVOBRUknN/Hh4Zna9CinEGlxZH1u9aB/ZT2bUvETb/HjRpmT2DhTn1Aqa9jgyY6
G1YfO4jcRAyIAzdLB5HUIe1wvZeCw2iiH4J95AROVx5bkBCfATKARIFspc56HssLgJjziTw4XNL6
Tj5OypNypfJ7Z1G6dhjiGN278VY/tYYMsypJCuwFNDvCnEU9p44YXExh22qIAnPHKnS8k/wgRT0A
xheWbPhfpYSy6tilsJgUqcY4KITjriPk2RCYDDciF9QyrpkWdFs9RdcRPEWRmss8hvL0i9DtnLff
/wcK0tt890ycrCIhgomBC9Xty7k0bzgMbdJEBDQ5oJRtY5QCYcqbHIdz6CX9jC/1xANw+TINlzk3
u6ohrvOLPuhplBS6vQKfpBvLq2BlgjZwOwFyFsqZVgLEdlZxDGPO+J5cOLAplY8E/1rG6YViWx5N
U97n4AkqvzFFfZeSxdPnE1PbA2WxZb+C66OPTFv+vZg6Z+sl4Fwhq+2FuvRCCsbNsyllreBmMnrF
s53UDwI21h2RFm0wPl0ipoC4pBuU8Rl2D6ALPJNHFlt9yxO8xGR/C/AfrfciyQ6MUF1/qBC1tFbR
PPKdGvHjdDArH5YmlyhG7wx3BPTNiOJZ1CQ29U77qViNMDSiwmkwHaHXpXanLGvx0NU4uWG5RMXK
7qEBz0jK11PjXeSRThp8y9hLz0c6oIvP6uqn249al2P5Wkvnvq9UOHIUiSjnxWyzRJMma5ju7xEd
b+z99oA4YrHK8J74b0cgMwdu2w1zci5xs6rgcBtZPtnmw8o2zxOzwnlxuHtdAGAeh8e2It9smsYT
SRkzqtdLGsTQXvfKWE8mjUIic/cB7xb2mDL0MAOajkI0UBMry05XLH36XievU1U7x14nVpVnmihR
N1xvVAUA5xPkqQMWiyldgvOj05LFFEVYqeCDh4s5DbK1zf3Fa6ryuQEI/BqOGHp+PgH5V12EE+a4
WCXf6lJjT9BWwxqQLLzQltOqXSgw8fcABq0gxi/kqsSI63rxdrKM4Hi//HF8YgmDAPZPfl8BGUFW
rFaleRd/YORqxSeaKCvASnUct9W7nEdle7lW3e4t0t55mQ7wJ7uSc8VoeYr6Lv4+d0XEMz44Ot/4
UgJaJBtrJSKjZdGbN44YKucHZnM99VD02wNwytau8/In+53zy0mQ4x3h8b8rC6WcNxdnLKQodicc
RFi26TVrNQXVINWVV8Lk/IHYIOHlkJmE6GDDLU30yu6ts46BCrWLGGMRFdG9I/X/af7+buD3r1Me
efO+H3V+kXS6NCG0KXVxYye506COSSSCiV88jJBtoIW0UCqjy2xLgFT3ZXnDoWYk/kJtvX49apc8
ORE6hAV06QdRF7Ga9iuHibtwK+wP2sNmmLf9tQyBTTv8NghfefpwDcC4V3AJH4vPNtauQZZFcrJ7
7swEv3UTXR1UbYQmQ0hZ22qPxl/KTNbOzsS8WJDVB+wSq608u9RC+wPvM+TeGcTWpgazq84yaHfw
dMn6+xJg2PQGauj2dd0XWhIYNxI6160+E8YMPg1b5/zZr7vVO2EqArO1qgMgBffZRnsHKqglee37
Xc3xnK83bObZtrD940ydhkMe+b7zOXmzHdsFDpQHLGLRnkHBcFRvjpk+t7sbyuO5JqVlvnbh2b0W
Scc8nYIxW1pEainVWmB1iGWs5C2L05sx2GD9NKcFPjoZOt0D+bi5frvmaUFtt1v3wbCoJlNXm+4t
0Yy2NM1qO0cUqPDImiYvpUMYzU1+I+IUkgitXM/5eMvD3e7B9KHxVxr8Ied3+dHfSwlFHXGmwkRS
APa9IxlJRLod+/RAJhtw+cMm3Z5NB/BkthwL/FjtYbLlFEE1mHmhSPkMcCXHYRjiXfcNSh2Dp5ZU
XmQqV01bxkBtRs3tXEyt3GOiGKd0vjhGoOBPIwt4td09/P+qZvBbbPDgAG65nDTVHwa15ipdIKww
p+5hN21T9KEz7iDyBkFubnVtwo7iMk4OXcZ1OqA+oh3uNthcSjIecqkdiwMYD8COGZz5YLxlvPWM
delZpY2dJA407VYn7gMhwGmMwMlYv2b2rIBt6Qck6L7UqL0ASXVFacf4lDlNb1f2Akit+/nK6/A/
KBSO6wBKf4py74nhtjIuwobV/xOL9+cBBsXkxvzcrOPHiVWVLBGUgyC7xxfU2WOlBaq7xe6rKybi
SkFY6oND+jQypIUTPo2Tju+bzhguhLgzsFwYhRc/N5yYE1Ml+1YR3I6dvkG79hMdW8VFQGfJ/DKr
RE2G19+XOJ03hV9VbBXIDEGKuCgdgZFien0oZK3KXfnCoxKJClRMKYnn6u9w9ixN3Q4VVspZzk1/
svoW1EsIB9J1ZN8nEMJ9fYuGeGbKM33XKuxhTzkYywVDgqXzBYu+nEIZGRnx0Ux+Lt9RPtSf0QQq
zPCVwRXfgX/mB7b7pRDeDAVy5ZDG3DtHIP3ck0QjIqNBp7bmXVv9ZxqIKV1zEhN2+K2PmQR6Pb88
Ib9T2so+YNcemJgvWnhHpGDi6u9NcoL2BBnZ0TfwexxZf4+jKx2O22Kh58aMJe/o5jASJFhLylSW
ufYbHCuHjnzfEff5eHK+HEs6W6TOQ8VR1zKr9uO21GQqyMw8Rj7GK/ACJaBmxZl1ZuP49BYwI4Yw
Se6JuOpGXIe89LoE0BCwCjz8e1W3WQbRIED1umOnnkdHDOvaHQf5oyr18DpyY5MHkinQ7DHDz2r2
NpVK8W1P6H1aLVgm/RvF2TohiFN9tJFfEjaYqFJsOql50EkMBQJ/dZB30zKkogLL6FvdkOLEbkxN
UIkM6WMxHyyy8HGCjYBAUf4UgWenemveBInYn3NAKIMoEy9vgPd1VsyZcbOrKb8ja3J4OosJG1gy
2XGZXUuE3eL2XwW16vXkkZXOaLxoNWppmvgK/20CvZQ77OgcC05y8HnqJ3Y/86RN2zo3IaP3NkYd
vadsXRBbSuxMabGeQulZf4hmJufpcciM4c2U7N5/6O8HWAAGvlKkiNdZcUYAmqX5IGcCdNsVLR2L
J+157khhzV+R9wFuIBip1+n3v8g1twE0yG767urJTyq/s87eq8kjnz4SuSsqbkAr4YMXEs7mPHdk
CEpB2vyT3lyzb7BMiMnbhVJeMCgu0W0QRFGGgooRoBwfRtfvm6xeKFK3Ipo5wchDSKtWZP3kXm3R
vp59A8bmYSgyBtazoFv243RR0TlhWdrLZaro7C/DUkmmkE3iW5rclNfaenculg6yZJaGpl5PhmlT
LzxH9Q0FJr9RR4JVl5ljdNHQrvZSSdrFbUv9qHO3KcZAeimYawbMCBWsQw8mYD5wyL5VilQMM8QO
8cL8cfnuYTHy95QhZVaCZhCiq46BaJJzZJ+6LKD7vEsqj9d0UN/TCiK7rm69igJpB8Uyz0vcf0Ly
1EkJMkBimHtrJbZ/HyF/YPSVwYJYRq5DIxxxzlYIS+TpKFTbWWaelip6ucju10nKLSW1nfkMHYhY
VUrrDZUomkKfjJJEapRZexjsy6HPkiDIlyHleSVQsTf1Bwy7iwzlk6yPFtezkv9jI0g2r9fXlt1x
K7OpsoQPRksEGUw1J0Lq3X2vRumU46+wqAz51svNxZ8UqmgcfrhK3G2PUtAh4Y8cumI+H9BExpKj
HK/wkOdeIwBZ5vtPQHU1HNEABxl0DLAbETXr+OpQ1zWKnDzmXd6JvT4nn0oYP3kwe3T4XcWua0+l
+kBP1eIGvWgxFahJ2wY0aM0YdLRnxqcTx/HB4pCyjgC38AVDxdV3OdICuJfgbf/FFtXkO+qZ4McT
+Ctn26TJU7fdoZyxyhz5dJA1gdQ+4afoL11UkyqtMg8UtXulhWjpuL6IwkE6aT8cPRstBSx9AEOg
Wh6q/50ZWqcR4zeJoGrXtTzxjLMxRHTShDKTjfW5hQO+Hi/3eilymVgneV44gm/toRiwPm9790n8
yMiqVYdQt/mZUPswApMQuRjyPSzA7G/6dKTuIoHnnIlTtjUXlQf1cH167X+4nkR9YREyqDwPie9s
maW5eMOvdHybAITftU+lA5K0/ZyvCezm8WmN2R128OPtwkkn8FQYHQ3xio1kUvmiGc385Zduv+3T
9WDi2kCELQ79yxhTzLST4bf925wTzl5hq2ev84OgKZawi8OGgrfVAjYes3Xojcc2m6/2ONCxLEMP
e257P9dBeW6bXrqDXjQks/xYy1+ek6sQEJKYOFFyE+BvV5I4PUn8ZHsjq1wcqdYCBc6xsufig92c
nb+9OVygLJDXKamyyI64qKuQ+bdU/cO1Ee14mFsQJcdmkn3CX0xIIYZNd26gnl3NesEoDB948B0t
e4icATAipzcEKPjaqlNR0So50Tywiic7OT4tNY3ziB1P0DsP1B95fcW8xWHSlVVzQZgOH2B6wYYl
iYaW9ZK/5bcv8JqW+0E1dCDciVLNr5UJyLULAGdS9dmr/tCO/V6NwnW4tAWylkS9Bx1fwpy5RuSm
qhhanX+HQmaT+6VDb1ScKm//rSc4VM4MFedcdSqr++BU7g5936vV7Ng0p1fILxy6C5Rnpobtr6L/
y3YbAv3FrbPUwKg0Kcwl1YkjoD+bPndo/wb8RNLk6HlaskgYRGOUiO6vBzs6OgK4ynuXawkumQC7
CQWOaOGjHgLi0QgVHSR9Rp3MDaFpEDc099ZI84HNzq1vvXqLYriv/Os8adGyMwUyc3I6R0UTaBYr
wWj1tjja5T4iKBO/uLmcQEiRgRB/cqvllSBqSqu8ecpRsvxx4Tx2ydl4J0/qxpi1tKO5+XEKwvKg
OZZHL0j7LraPEuYZLglGjof5i0GZcUba8P42lDbz8KjarnCdmXT4DGp9wxXudt0Vs/kdtkHopi4x
ts8ARj8KQ0Ms5q3E1N8Mb76b58pWyQSPn3A4jvDYTrSgtWFVU1B0HWMy/HxBGEQigubVwf0gRlRx
JArjLEfSB4QKF89QG1Umd2kD3XIADS45nTFNJs+ZPRyc1Q4OSx50eeW8lMPVcQ9fC5wLW6D5uV2x
7EYgHM3h/KyLg2m6hTxsM7kDiNETnU+YcMlhqb4koUmkM2WIc1XXlvlZDiyRTgee9kG1SgoUqYV6
I2UTVX6NolUwHLLr8mI6mj8A1ApmaZtqNU2byAtSFslS0vaO9RkKcW4Qs7oG+nrlqqj9jAqJzexi
dh/k9DvnrU3n6WUX1yAKK0eIlBixk84GzsCaG5H+YHuSTtmUZ/GuGEmCFsI+5Tz4zFZIuGqlikzT
X8tI0VTtkTkB5jZ3soBVJ5MNUKfAgYzhYHetZ2fRmGZvB4iJG7LoT4kqGMIcMGPtbj0yRxaUPH3t
V4Pv1xHJZWeqxIdsMuDVVpH4NSu8NVq50YC+yF0s8KQYuXqcviBedEdibrKeyYcI3qBDPwyNVe8R
qA1sotvybgImItRCNNjiwFN3/byiJ2xENqxsKmrdbu/xG4fyqvtprV06ZFzGheavziqnAyJ+ZfFO
DIGtmJ7bek8vTdiYUw4I9TC7pnjhxy3wievHpeoC2owji+VxSydz+sw2norX2aD0+wzK2NwyG42D
W1AmY41Ie8nVjSbQxGnjA46Is7/qMDW3fdZ8Fedh/vga3vA3KssCDrdTj8Dn1JqrbksWLW8KwWzU
8VW4HZMbqZ0J2FKE/KGISzqLkjqHMRrgVlND2rD5FfgOFQFwsBYVBMvC9E5LFecH2fHT5+gToLdJ
hXMC6GkgPXEOePHR+Q1BNg21OomKfb987t74u5lR2T1b4STUDfSIvoLM2eleWS5PTJwc3Vz9KQQ9
fItY5d5gTOotyZKVya8r9+WYoKkVQud19GPazAKyWyG1l7IQ1Xq3tfLq49bAjXmJpIocGyPZ7aNs
vK2OHgIZoEENuurZqg506z5SJnN3AXnkOX0RoatbOh4XKMrCYCpZxk1/G8PGovtZiaeBsufri7zB
tBNqn7j0AD2KikUxSQX7zmjDBC/XGu3arYUDODobKb8yfs0N6cC2ySDG1MOMb0Zt2U7Ziwh8WoFN
3f2YbtdTaAKTJB+OVOyL75q0u/5g8hd8zmpIIOULotyTthO6QFn92bNH1OL7+dRFLaj3CDA4ZvN0
5/ZzZCNjMSk6s8O1w1g4eblQ+DbPGPPbiFkubgH4z5KI74k54teAH/2sV++TFGu0pjKgk83T54zA
smCCXegkshfe95zGp4AhTn2DaNSMIMPkzuD0mOwlo8a39EpQDaso8MCXSL2zNvlqfOrb7JZg/icL
5aoCnBtgluCEedJLAWVXSCr5HcAmnQMrr/gEBdtvPquVFTGQiBxP3mZAU0ngpnhQsttLx2i6dyDg
zSOKmix3yK6zL1eJrwEGuWojOm4yyqt2NsITHWJRmKyJbxLD1sqi9dy7o3hUeqsl+F6lTeQbRIjd
K5KxYxSs4tgCPe5Vz0VE2gAD+fKjIxAO/yPvHnbO13fjYN0yAzVnbqB2oMOyUOSzKMV/D6D32OtI
gAONTEMnfb9JJvJ+nBwo+6tbot6etKnaytTo8NWD01KtLE7J9HrfBzP9RrKOP5WUj/CtVmkpmdPI
AeY5hR0zl5RY2Lobk9bi2PzqvFEXgaQG7WR/sp1qSVQGN4DfQvMB0NXSKsOzkc+flVQWQ/bw0mkj
ld2xT94+GplxpSNRPqg+wYd4IcOHjDC9ag2gOKP/iK/GUO7pcX4yhy0GnsgnLTs/yj594c3+7b9m
x1gv33ZUO+2ExrfJ613s35bizEv93bP6KRTlBdB/kmBK2vZUQTgzcpuxtEY8CbXEDhncdemyazA1
bhYBmHUxZzHCWSHKA9NvFOw7M+HO/k3upYZa5msuUO+4xKh9Bh3uKrt4w0dYhupVrnVBZ9g0mvuH
jTJPYZlnMPFnT1io8jsJJx7PBXLxQvlbHoBoNNE0Jnzgsf/fgwz6PtLGO4apFLnxyNjemyYpx+lW
+0XpwdpFLWuUzzaZGbud7r1wcyCehvI3Vgg7JJlDeOaDlIv+oHETJkK60GWeSCj5/0sgXmksrOHn
Jp9kEJ5wNzqNJSg8uxEsAIadrGkaGNztqTaf0D0KRjpy3zQpM7W0exjt7CeXwOF0Rf66vVASns9b
5NhGlZcL3bxAkOl5uO9laF5hV8SmpmXhVLzfqTFv7QYK4G7SjNe/X+9ZPRRzgFE+E/4N7XVi4HPw
lbH9n/ZRTl+b7Qg6CTOjrf7x2LiVmMAKCm8LWHMwMAroUcd8+rHjS3bxQAOFEr1aMW8YyHhboHNj
4chhAY3+018N7jmqOJntAX7/HBVe+EUg/hkp8e3VsumbDOUA+G5AIWS8F5AN2zgcY0pAjF3XfghD
IAag73JdWk6Ev3xJr1H7eKj/YZNUxo2lwlpWUGUNt2u2rOoEqRXa0DhKw0sIF75hgExIYuy7TLDe
/6OQWaOkdxLLdz2xDLCc4TGkyWlGUD5VAGotgrEz1s0xfkFDnILJva+A1nWv33hp71Rwmi4epnaB
Tz5ozK8C3WWQIkdKSGU+rXd1ZOgH2AA5npPlcPzCTqBqx6cJJ5hNFxzl1wNbprE8CxyGHX6w2G/p
iz2JpB7qDFxspIOsyJ7NjAkrOWbXf870usbG2/VnrdaLbbs3VzTGy2ZvK473vSu+4oX08IL2sh/J
faMAD/te5AY3nPMjyxbBsysp5cmKwUM+vnUKtOzqL3VT/ebErbK0SN1n01yiMqC3KVIZsvWvCDsJ
eiDCUk8t4ghkXs9o9ZOxP3CQViG/VvVzKqZ2weY+heQwDlOKLk4dzx0zDH3oy8oIIBdUYMzohYI5
QoVhOsHT9+nTinvS1gSIZjSjfz/9nBsMOQxkwiRXhFgi8eRuAgyKKdL2ALqd9Q6Zj55fc0wy7JZ4
iJuI+sij5oHRuRxA8hKw53EFBDas85ImiFxYIpduNfUd4ff/+tCkG/Iz4utdo/aNQLKluPV3/hU9
xmBv1rOi6Qxl1cjMaYiWlxPVsbRsSAM9F4xv04i8/+6QhKEqiQ3P5ovOw2Yow1XdqQLYCqewB0jR
YwwAnmI8AxRFK3p/JrW0PHkJFcKb/hXoZ8KuTfh9O6tEADL+qqdZDr0oz7y1caitPQqPdMp1jF/k
Saglp/y0ZA+fsbwQQU5l21UQSpFvuXVFrWpg4QNd2yEl2eqiNcF4Aq0rPGWFtwG+NNObAHNth9nK
qTulJezJl2DnKeRLu8nhrrPPOIol2jnATMJQZQWrU51nLniU2svSb6/L3IE6aD4Y4a687hm1wQQ9
gFTebNOXMOvCWFsnJ75VwC2vEXBgf860or75fUn/qX822jm9dnwJtn+qegHyqSIZDb542PF5gIIx
ASs5Tpu8NeQ/L0LJqkilEtKqoMd29xNQDTeVYhpVBkUw760atnDlZzYgNGi9u/PbzDaE7ay+5Y1d
XyPxT5rRABpJ+55tPh1gX3uA7KOF6qdrzEzP7kOThaoewiVqOUhUgn2KiLYAxI/FLr8ExBFXwnfA
SIQer/E5D2b5FLBOZP+kcpzD7VewiHlbpMrOtcL7iSNV2wh10JtXdBPZLvGUYarkZH+8pyeWfCkP
9oWm6rnUKkMEgV8oE/deVyzn6XNUn9BPYw73qdWKf0YeKYgZ9GNSqGOxTVMiDZFMs8PVrOdJWs9q
wJpAjtJSt/PwtvyDWct7a9/bLsCygwfgZaXinXXCyDM42doiPyJK3i7wfvY895dbNjbCXUtYFFiY
3rlpsPY7wiLuEcmuAHQbf5KrBrV2zyXprmO2BJA7n79tMQsF3XqSnQzTTmIGrVBFKn1gpn2qZ1OU
AHTywcNrx6dWUcdR8DFA0KtOj5YinKWPJjCT9O3RMsp+AoDU156lIWvADT9KV33T5SkQwHw/hBt3
2seruSS0hvYkkWTgUBTG0cw+uOVkQIGBizmFH7e3eSyFuLMY+fFBkm3Ytg9c2VEma0veTJT9Zz+c
QK5HoV/B2/H0mzRjIaMAl6s9kI+edAFV5yQ5LRLaG7fP2qO6aYrkAMsVAOZoz/306E7t2jfNUNq/
QvGZc7ryA+gao9LUW3uGgwtrf5RcY/kHPXHJ4mXgKi38bewT3M0fhOsNMesboHYEG+l/97TItkpD
rWqzjJIB9cESxOOIZiHd5nfywShtk1vnZVyfdqN+/K0DRwn+pEMyZjbP9kNaHh703xUNXJRMlQKR
Fgr6xbe/lLrCnBY+zjqCB8dc4PzkerbKCfplwAPqMcWaGLnV6tpdHo+9FkYP32hQvnkzsAKkIqGC
cxB45h1PcNWBQ6XIz1qX9IWu1EMdSnFnPSoQLWN06iuqksy2MfbUpVX0x/9eloyy/j54AIgbXq5+
04eD9LJz9ZPf+0oqCuuZZ5bYo6gEtfjIW/1WIc7onuYR3gVsDRPbAee7s6E2V5sR23DYg5Gfia7k
hzYl6IJ+NMdb9dXA3BB37XllGRLqbNBVHjDDsZk2tjzrLUS70NCPwrq8zqI8SoRezNxAkf2YIAPU
LaoBSq+GKTGEU0j/EHLhUByIZXdGjsk2pOK6rWfjy/EiuQo1D3mnCB6pkls2w3TIS9BciRa2fKga
LDjUPmekNWcDlDmsInCxozoH5advklxcuSzz1QQroaqnUQPr7u6/Xyk/EAEisEOivKnyduCw12hh
BKiEWz6aDPXasP0+RLg+TspPE5dzAEekyxt4/fs8HOWyg7L3iblB2O8AzW4SuJhR0k93ghzm1DWO
uS6Iswqwm2uc0fWrMjBojEbWqGVbQsMi2CjkoG8su03a9TwC3gQ99uR4e9Ot4/9TReovtgLbTgqh
rZ1qxFLLnax/AHOG7cyFq0Wgz132bQAldSD+rejE2wdgWTizZFayzwt4UxNIMitkhQ5+LBdyklDd
hWyKOjsoj21vK1M6xRICrvon8ar5mKzTcNN3GF+IloCT32ckw8IT0aKLLIRpVjReQe2uNUXpSo12
0qSGNvnzd4W17RJF4GEhH97mIKThamgN/Qmm/uNAGCBPzjcaRLx4T8imsoSQ0RLmwZGtT/9blO0c
TpWcII63yqDPWw4POt0e42qD7NI7jw8po3n95trsRtmLwF17wTAEZDPMy508v2adFYa8Il3xrqpJ
AQPDX+8EPlheg/jbgpjaMsYe8X06Au+e8LNQm2mEJm/fKunhgU6jDlQewtr9tD6dNKHGfM2CnTyn
OWuULj7uZF4C0cwRGD1FUNzovZEZDoyDlXMs8usz99P1wBIFPEG8LiWEzHuhrxVqizf1oTUFk7lc
fgVfUPQ7wQrNHRUuECXLbkfDfpO220QTiL1O0kBk0PrpxZya0AQJ3pe1TlSz5jY0f+Favr5NCHZ0
lin8wcbEkLJ5+wG1YiMbt/UA2ttqCEomogsxbvSjcXCgX59vOWzutJW5ZZEGNlXXpQzvkQgxQDAv
z/1WgtiRCtPSmGKYeMi2EzbO8sR7lpRmG40gSkW+IdZ8Y717B3hnIuTvIcQ95OA4Cwtdz5FaAOky
Uq6uhuRojlz3z/PzoBBm7iVRdALZqFVm9nxYrtF8aFJGVj0Am8DjG8AJKxiM/t5hs35VqwnG8z3b
rYgwPlzgzHufboJY1PUKEBlaVnWpPK1mrHU6ADrqyQ7U+fQwWsaVYLxhjFaTmJQDSv4KqlQ9Pkjq
3G7HSgx0tbewb2SGQKMKgUiUZFSmQmTOgiyJpLRNURgeeYGn4sIZ+jc6dudzK5nESy7lyqbQmeFg
5vnDcJWpH97TVQaggPqyTNuW8bQ2NJMCpBI31IbeQnscfSJ0C32JeN65HfyX9GN5bY47sP3NHSie
yt1wOrbgxr2PcGCcSzSowfN8F3nnGRJ394mxcoUcIw4VbyL2xY0egDi14TSGCfym07f6C6YD7Vi8
z8Qf92haw3JZ51P1F+j2PsPo2ZJT29HxN4P9Ch1MD/zda1Du0T2g4qlXrJ8LS9eDq9rKaUBbWQlu
HWhmyMSBNdMX35oogU1yLwYr8rLCxMGotLO64dN2dfSZFy3bLwkJm762041VOESec/rZyjeqrcO4
Ba5JmdjbnKf1gCyehSnpIAX3u4oedM25Z9UzS+xbe9Eux9qu3riSJqHh5DvJktjQgS94UUY4VLS4
EvK7iTZFKuuZrMFFg2odaUNV1mWOb6jEjW6ONqcafEh7SufN47ho3ulbA2HEBN1dEnri8jYr2jik
tZs1ETqrcPGRfaFF0Ok2cJUEZ7CL0DLmdbmnfjB1Y9DAXylAs+wBiAbH2VHuEIZ92jgi2yPefqPe
xQd1I4p1WJkd9TYH0/P2W0lXXzy7Pl13eZ+qb/j8DvAUW2pnmT/bsO5bpvREA+/hHGOciTjwN02g
XgRTl02TJIeMbmmiIxUZ+/r8rnIW4AbAiL6RuYumnOxEh7S0F/ROUvvXOjl9psa1ku7R6Bolv/ID
wk2rbSzuaiYUDyOr+NgHEDC8vE321WhEaJ4PSAbiUmgNHTTotQC2X51kHtVcDbbhMG3jULzcNi8W
c8mQY8t6fYkcxAQ0bBK50dqiUuA5N6AlzgDPMBacTdZFZ/P6WIq2XRGUpSFYrKywhz1Uaz4LSm2D
yvvOiANGNNSqQw+tjU4rMMOqEByBVL1IJ94oRQemDDBZPFr/WxlPrmMX0nP5gS0Yn174U7lX6nWX
6pWy1bGmSLEzI51RuKXSE4T2iYk+5fFAHMgqqq3LTPrjTM8Jb5erM2fKlIT011Os4htJ98cLp0rt
7y3Q8SgclZkkzoV3EHPg/UaofDznoibmgEDhNeAfxvnrhiOuHkcEt9hNAq/8I6bThYc73lA5Ir90
JdbNiYBdnAkADH+xrcypGF6sggG99dJfCkwOsIziGUNrQbkZGe5PXPR6RrFR2+BfFKtZbgYE9Z/1
utOfElELhVeArVA26nH0vo4+DSCMyPXWVW3I30Fdp55YLmjAgmt0WochrlRzSFgX9wJu7qx3qamO
v5mm1T5lNaQaHfbWqAThCq3T0Nso4GndD9EWNwEz1J4mKJPSbZ7buT9IVPj5AjZELFPPmVQJSob7
WpONXMNiGF376aNJQlMKGIzQQJYHPPDSI1pBgjmWSS2cUCU2+yK7XUHzVKKXWRyUP4/3NZjDJ/Wv
eX6+AEvHr/VXNZWbN9mvLeEzBhjETeYY6eYIA4u8L4o/7bc8J88UYw3KMmaUAqGP6CWnsLtOEkxE
oPdP+OZM2dDKH1Rom0TtfD0HKXOKd/e+Q4mlfPyE8YbmotWwjNnM/zS2R2sRyqNU2f6STdJZxU1T
WyBneFQhrCnIknvivVLhN3oHADbEfMYSLBtKMAuCyEXUZJV9mPZexH6hBLs3Ys0XSF3Q7BlCvkIu
jGYfLzE3vQvOCtIGVEriq7GESbMU0PduW28QyZfoOwEp6AH38eHYmS8S09mPMpreNoIQm1sUHeyf
M5tZqQNFBPNaOYcafPv0b8zvJo57rX15nm73kwcPDRvSJpyg4Q5n8uZgWAqVTLZnzPjF/iD//PVz
/4cpmAA38v8oX9H5t0s9FoyJ2To+DX913+AClHDdl8C+bIQnH8kWqME3kVwqDirFvyUCxxjlmrXh
a2APYzAGqIEZNUGUEAFZFzv6oYjH0KyvokOWssXSmCdOJeyEPhmdW0KaQ9vauFn7qM2cKMpg0ias
Npx3Xos4KSEwmSiQ8SRv9ChzcDxzBrZDJKYhWgCJ3y1dwb/u6z2CjADxFWuzkcHR3lNYPvon+x31
GgL8Gmdy68KH9lVKgaYgaYCG3JMKlxUTPq27BP/u2zXgiXCY1KeMAl1HVGyuQD3VEdwzdkCbsdu6
sraLFnmYHJS3jY4oKBY6b+SBpxIyk6vU++9zLTEZBVwYw4C+2LYpIKHbLnA7bpY5a++PtWmEquzK
c6GSpkC+6TzLg0mE2pxK5x330XiLXX8w09N+vTX2HFJeC2reP2D6ujRLtaoGzQ1CzYnGFIU0q5gg
Du5lhktx5EPXxde+ngKMvS3Da3z6cOXo6/30w3CM2TcNUgoW2ueGitjTN7Z0AV5IOL1xE/fdn5tH
/6I9k915l2TMT6qsBY3cDOLQ59CaCoQOMiAxDJHmCwpCRJ0oBhcFhvK8FeGjoOXGn29ctdqv0a1N
yzER0BryoKKY6lwT+WrKI8K6uY2B7FYZeQd2buXYgHvlT157zATEAVfpmHfyXDXrN0ki0xRKvnPr
oJAzL+chauSoXjIpdFJcPZtsKfsWhP0FOIg6L3kR7pKj07zNdBEsP77HOSqSkc6VvVw3o6r+uuVo
2Ja7OMv8bYzeRtIKwxkY3JIbXobeHohDfuBF61IeMkXAeaxIQga2v+DcM2B0cL49H+EDr9r7ooLL
B3SzoNIgaQ+hKNwfUc1Md8r/Gnk6u3fEgKIby43eh6rXEIHJoYGbMLdG9XVU1d/7mRbFq4wro6VB
EyPpF5rjz//a6ai/qoIz20J06uzZLQyvZMlczBH/VlyaD/xTWKbMW/cDcDDebExkQ3SCdCyeYLt5
DMxWjEJRpuxjn7/KuAKmyIuxDrue5/zm8BF8YHTZm2JC4xQLCDesa5U4zplLYPR82Cl+9gLkNRcH
3dbzaJspw3v6oEFzftfnIxk8PLkTnYLQUZy+d9fJ7NLeY4nEkGuEOZEXaKZdeOULf/wS9jiaII9u
7hTkX/mEcZrKfSWH1/UR1o76xPIIrypPRvLvonQQMx8wjtLotHab9uTOaKEgjsapg6kKV/XhOzjW
Z9WFJiScN8iohlokBcEMvqwvuZ8DMBuRZJwpTiZ9HSibybzGrTnisAcrb45Pw9goV7CoSqq1SqSL
Jwqp/F1g6IH6nJnFsDkaBopTPJyoH70uVD9sAq4oC4lElfk3wdlvinBiPQ1G1It3U/DvZyyMmmlE
zt1c8MUVRZIG0LqipQ2ABaYBVkGzIj8JxxQj9VcpqTYv9FiKll0Qp0OGGDgONjRnqTHbC8SxoZlN
t7dl2eUMA8Y7aBO75FsL6BTLoIKLOyRJJmxHY7nb2xV4Y6vapNq+QABEyO4SwPxSEPb71jANSVx4
ex574vBrTfRBhPMeHZFm+AkzA8rrIj0xpcfCLIaOP6EZzMXPGaX1Hgqa+5JS3bs4GzIybF5D4v0G
VMvCTg83jaG31cSZzsu2zzeyAvMAhO9NdI4RehV03sA/rEvvwtavWBCwppYJ9fFduYP9APUHAhwL
bj8T32P0rnWN7cMaLqhbiqdQNKdLRXipn8UcKle6l9L0GsU2R3/tPkWCiiiMXeUp1/Mq6Fd/axDb
GBvR4+9JjxiaY7YRxjNxepGFLUv+foMj8gphYvf0vxYZjt4mDgvu0vQcssLiCyTMz6395IMO09sF
g2dOzzytgqLUHC3PCwpnxAYmC8+kAf6chEOVU9zodq/BOxxF6ZoRICj3vGYmepBUU286pTXRCOlw
bfh6F/t/CRwjOLMdepgJcskQNWxhosnr5aaFiWdGUbjN7iLIk6ovlKI8jeBcpk0wXAF/bKM7tkkQ
hFozbCRquxHv9zP5Y4LLvi9G0BSucBtIt1KXWSvHp4w/NZptU8wMI9P/wsnm92sgVCVwkauOjVjU
by57xMbAEFEFEzbgl2tbBPrKXcYd2NzUT4cXMco33c0yX+HmYPzNitpuzh3rQoEPJyKwXGYwCdLo
l2/GRRaqODLZAOwNhbz7sNMQTpyp7cS6nHPHCwIgdKVCyerkTKfqQsv4JmmOKGHonJHgbXmCH6wQ
XxJL4O1ZYvzTCqW3lGA2nEsCsrtAj7Seh70HGRzYZar4A914VtFisH2osAF+5HWWLkhYXs/nqNMQ
cdh6Dgr3JJQTcC40SGMLdbn6xv2Fi2Fd3FQuWBqnVv15MugOxqs8S8Kox+AlOKe9dX8Q+yvq1j67
IdzOVJq9kKTzoR/KtN0ldIgpLJVNN6ZEw/GyxSokz33vzIoI3ZWJXOWTrWA8H/5ZFPzie2OtaG1+
FrosNC2Kn/P0xbERj1hv7T2DK91XkxZl48SEdVhVJL5dDPy1zfu+omTUy7OHRgmtZYyOfexEUTc+
VMw0oFzfi/r4twFfwgDECfguiXo9xI7yTF/jGH8L0hqzcZJ3dOkui1KZFfQzZ001Vpi6taAwiwdo
aT45W+z3ScsuYLLW8tq6MoRNkZF4gN8pcWZ7zN/Fz1V0J5Z2nCmMWChejinliqEFm/Pqc4BsUDzv
UBKOyQFE+LwtcZAbNJSHZU5+r6LpwcAtpx/exwD0XvZTjQ7BWo6vSpPhj5OjC2gJxxr+k6BEJY9Z
jJHEC4pAFtB/7rLkNBx5b7M988NSarNwauZ5qeNS/TnVV79nXdAsox2cN0yF1EOSYwcf6Ie8OYIf
cfmIf+Dl9eoOwIEsDgUnqD8qmTyr8m5WTo7Oev3HRYqmZrjUZO4VHVaMfH7c4zMSxK/5E+VpAhaw
sZQeUFZfsm0h6jE+RpYmbb1tj9V+vwECrzS2ws0JDF46rCEE72gjKRsPU2NRsmSivCHfM2KmfoE4
5UZeDUMeYxwUHkstz0L+zKGEToB4Egmkvov4D+pvtJCNxvAOi/y62L/Fs/GYryl72U8WwJpzKny4
T3N8M031uysebkThKS/it9ta8we45ebC3JCH+W/EAi1FJ2s7fcer4pH1rgjviGDm8ptk3rGopnlx
v2a4NHs/4gNgD10AU4Z9vGlgzF7f8JqSn0EJ6sWhJG5OJUUPrxEmWb2RxrPz+PQ7KKZadQkAtQmV
gkZPWVRb4prD9KdFypd2wZopIN8CBXL+Kd0JJf+QBMU6bW79mW3IycmH8MDhA5fLAtA4Ra1asJlq
lXxBqyifJMSfbQROmUcEUoDc92SqA4og6INelfV3u/u/jDyPB3L2d5gNG+AH/5UeKNHdHpNzYthw
Cly+/DgrZouLihmMSiFnhsnWbGxhurj7O5+nxNsSlQA2Q3hZOdPTXSI38mVskeaHWyJVvrgnH7P4
BPJPeppENTWB1bBs0XfhqaufPfuU2rrgyZTh3cykLxU4dl0Xlwk1bqAyQPYEVPNQqlMp61R1hDeY
NEOHRCtCkdARj/Wz0Aq6cbx/XyRdACCH2wHkXX32Q9wfQVxh1xBT52ZPYQ4hZ63yXg7P7vnY2MoJ
A8LcCWxs63esbWq9HqFV6UPLqXJzM30+P0zAaPX/2Q5BzCmyn667V5L7TEgBRwmNouWO0mVd+8Xl
80fm/w/zwQM2+UjjuDvbEGNHitLZeRYGpRVM2P8mhagVtPV0UdnFe1sKwpK3/ui1mQoMlT4TxnDp
YVefsytM8p52RRpSM7KGAnU6jNByv9+vobP8uKfMNRc/BPxw95jWmqwxSGG5qbtMySxgUpG2ejt6
lZELyRbdczqOSERcpg4lk7l9Tc9KM8B+FWdBWyMBvbJ6XyVMH/FqZM+4gIGTPfUlhIj+Pw1OqJLd
Sj+HwBLyEGwLh66fKR5mcdhunBmwNMyeixD6DXNRpgou1Izk+6DJfLN1N6aygISkI5OFkjH0o02N
Dh3F+H4eHJOI4E+FqJMcaVAOBuofGcS6KuxcjZiJ96LTPFXaeYlNj/xNlKOLiL+KLVN+C8m5LvPa
ku4NSqJUI2NynUMpJecpafbGrUDgzMgXaLo8bPp0P08qHnKj0Bd7o+j5x6/sjsOIGNAWr4LQn2Kt
rhWxTDSd6w7VJ6TT8xXh7jvTqjB1jm7HkZYTuqz6ATR/mlJQwH+jqDuv8GSdYtDoP6Q1W/+RNp2g
qGdNotONQOcRfUc60/CA/GmFfpeMagYRuR6YWZg1URb0mx3DAEh8MgHxIJn7sfq9GdO7NFnTynAI
9fuiSfeG2lowq/8N9bxkDnyT3RWIGoodX7TnRMzCclU8ES3Fn1WxzmiVmX8aAcSX44C9R5jqg3D+
gY3WIHZELbZyNj+zzuterBt+syz4ukg5lvlWbbbI24u+fOpMaTZjg0vmuOTqmOz6kR+vWJnkp9u3
9x4Pj5K78efjZS8/ufMsKbAoekuE9kEjhb8SOqq8U26GpQsHtNUsRXji4xSWfGm067gW2nHZtlC8
GVXV8dc64FddG5KIgl7Pjt/BYlJ5LrGlJcQgSWwuPWrMC6NgWFPRrx0yWXOTZSu/yo9pkRwZMEJ5
qkOLqTDWcdgNCS5KHi1i3v53ldbDJZcYHsOsMxsR6hMtkQ/dlZDNdijPNy22tN4QsK1I0IoTeO8L
m4YVZEADKSLva5MDbGeK48QVAREGiuNd5X18+zOFaK9ebsfHz1A33JUeN77CrWKOFEmOf/1mq4cv
3Wqhai6xx5p5FlwyiCOJNXG4FDYt+a4YdFU4BCEkrzqrPSt49j4gTXAM86zDfQA0Q9lG6XMHEMJ3
xSPjF1pdl9DiRgqiG/NiMWAJljoY0pNc9AWDGuQexzliJmoBhPU4gGEb14Oa0NJeiwLhVeRBn6GI
1d/u8np3v8f6gqBYx+IY4vjLfRNdbeawi1Yf8QaO3A/cBKYAyHs+VVgFwAq7MtvAneMvF1KpXiCc
i5DMWmBl/D3Xxtquyn7mMLXucbh0ljPYUQkX5ObLHJiYei+UozAEpNB91Yl09NOBIdfGsZBb5Yf6
eZJx9GSzlna8OoklaV/CTNtTbRlULqf61JUkpGOVdXHo6vfPUxXsg8yINovwKlaLbXU2L5fwASlJ
dlBpegBV3c4ewgeU9arHWOWB6GjAdGts8LZC8+9cQgGnJV/XfOd7TkGvfj3CYw/40puU6UT+V6p2
eh1SIEioGE0gjFbUYHcW6GpkA3pTC8wBwBjdcku8DlxeZnNId+r7s5E9hjuIvdefyFicgI+HK1aY
AAWtE/WbzhTALriGoyaEaOn7njQaGmeVP3gKUu4T2QcmTuvEiQdH5iBtB/RCCu2hTYZ/+KfVDZKB
LBKjI1ugKd8Yv1jrCeVIKLNt4sV9ZcqBGTRqTx/2F+BE5WrzXINPjf10sxVr6G1E0mjArqGOgmUL
5SQdX5L/GkxjYIWBiwGGtu1BvcLoruXMpB5Aj9xBb1VDQ8fOiCF+VLXziGuXU+/suaaGcFuaqoG3
GZOMDemh2IOitCgjB/EOtiUNQjFYGzLos66WGuuHeCiAm0zjzlYwwKLASxBpWjFmX7HJioX0V0j0
drECoE+BPo/4a87O7mMO87VOsJQ4WvzDmLDdvVKukx/IKfahJ9S4ITdKAk2SB1TnxIU9fzTk2Eos
HblBSUf9rlrcMtAn20247oqMR2Fxd/yVqNDo080PyZJrqjXeQLop5i7ZKSeNwreG8yJ2ObyBPIz3
kVN4PVIbnooVY2727W82gV0MdXfaqm3aziYSIW9TtCBLkPh+EeeMVMTpgWfyfxWkGNLmf7PxL4xI
fiF/UwTU55SMME4rTleVLp1XcIkU/OallXqcJuHmCTk95qIYoVCewK+AI66lUSaOGVmFVNbypSXN
4yFiXqVqB/YSQor7gogU1yafEhtldYbFegLtYjJ0DoWi0Co7PAqduOZJmvSPYDmRmRV+VhkHBnX4
EWQNmdt68IwC/DZwdhcahl64SBS5/QaHBPMy0DmJ+zHL3a57XYCt+J8kmTfQz8KIiMME3ZhRjWCd
1Yx6VakQjLNhDVbSynVrsV/sizWQnQQaxMi6ZkNHXyrYDIeuGEwJqoSx1lr96Iviz8nSf4LagjPi
hOXlC7KXISmQabbD9ZXbS72n9mU+YjibypB1ak5RUFOilyW8mMtQ6NRSBDBIzokgwged9n6X3ZQ9
jRaZvbIJ4k+9AQl2iP+oK38gr5IlxguqEE6Y7H2N8G4sn4FGSz/SDXz+1NguiQai1+DTLljWcmiM
kc4H3qnwPgA/p8NWrHj3nr1i1rVmM1jRNgTSX8Fjl6DTTIN7DUinxITT7iSk1IkWgn/Q86gG6bi3
YgHcIte6eKtZNt+yM62RnFqNAPXum3xR+5b+scdtAXAj/BSHtPY1oCzA+WEyYNrvHcuAbyctWyU5
goEk8kIe8DRaytTlrFBVS6O5owBY/PNFquLvoqHBhfN7V/MM+ooFKgNGDaVi0/KUJuldjvxkkGZZ
753/CNBbq/8PYTb6nnyMKKHx8pFa7XxCQmK+bT0zXzR9TkcVsin03CHCmLy8yAE1URugMOapTmtx
yg04RMXxDYN20TuuI72B38Cepa/gjhyqN1hjEee0MXGDubDI4lK2er+DoKw/AF5Qs+qSbuBtR4iv
93NlGnVJfQvfhMnfz5sPWfI9cKV3xL0glAofbgxKda/Xsz4+LYLFEAvQPvw90bOMHNhEgnGig5aC
DePw5HjI57vy2da5sQ8sv3OJbFFgvD5krd+P+NeyA3vk7+zQxktU3fTU95aRlaOCJXYWkTzIkgsl
qiRPuxW012pttw4Nv0S/b29SbbeMq3t8sMEwWGRgF1SVmT461pRxbgRiAR/sm40Ez+w/SBwSYl90
j2sxxBLaZrYuHVascj3zAMtk2wx444OZvVUe8rAZE38PYPgfqAw841x6imOlaj0q9IbuRhViYr/r
8X6rJk0zZrroMUmqreNIthdi7PEzxDaSzT4OdGFBZni/OQLZ3O78WUICOoZzQgU9TkD5eLavhPhO
SX4UXFnBpjZ9NDdL5Ea3voE1f+t+HfibqN4DCAVGqM8aybysU4SNJEvA3cmSIMtkzpjvtUQUpQBK
sdv9Ch7koFGmMFT5CsgmBSjxqqy1lBTaXPpb0a3ThMB7En8uwIMpNk6z8wqnEAvfcM02ArxG8R0c
mVI/Z/kkk2nXbQUtRNrInsVH3PdLU4O+o1lbqkIzA1o6B1DG22OZkToUCC9/P0XacXjnNFCX1ldr
2P4+HwDtCzueScoH5ZGtjoPMuEk4owG6EcXf1+5Nmps+wRq1Z/iV+31W4hDH79PIlxFMoCv57+DQ
MGhPwzp/X8TMxo8szBHADZ9QGi0P2w6BciScK2yQiameTpHmP2EK2jr8ZHVfWXkTrh78zjgfu4kq
PCnO6vJu17/5bv3g81iXww3911MIcRmcxU7ZaGQusBqEOhUTXqRomFhICqPk6qkMtxpT1GcX7xt6
O1709Et8zLVZclNXoFAJJEI6siwms5UsaClb2rO+tiHnQDQ0SBC0kUeBWyVSV+lrsfOd9sOErF5f
WEcFOowdYN4a5jUwmimRTYAD7xU+6DNfolqB1nwl/9ht/PyuidIklLBOwIhRVoY2lvtvaVfEN/BJ
l/K9ZeFHAt6jGgmS8jGmJ2pvIT00Jja60Vunq1XadyjSIGfS4J0hzarvjU46LqKgQbFFCfON/RQA
mfauoL7dY9RUxoP2pNIgNmCWtbFvpYbkXhgYUrkOd26xNveKYmfg/i932WJbWNm/L89suqFmjgbO
DGpZXSutgTtwxFvIwuTfytWBDEAWX4xYoNk3SM0TnFhVGObyKRitbMBkNNUoFx31cs3Ob1flD2iA
hS78kZ9ef2MeqDg4G1nR/9f8ApgkZ7uR64BXc0t9lL8i7Da66b97SpJtw6Dav21Al5xIU+2RwkA8
mb7Msz6ponKwGdPq16z/pR7vAIZJ0vPgzyzO3KT2raNZ0J7FO2Tuj5zesVI+WDj942ZDc/q5RMGg
PqRsxCgIqC8IZfqMtqjdjlzc83asxo35BfAITcDjYpytulcP/xM15fWO5Emrin1/5dUU7BajvOZj
HAjFHHwyE3yZ5EY61+pHEftWvJ000yFQd0VGvENkONsnMkrcOV0Z8rnrIAnzp13OJ1joFIbW/tX/
pSE2DKoVyTKu6tOZwt8/YaFsZkFsPhojahH+g7RYvCiDcPe865xu0qgFJVWj08jS/ZLKg0oLhAVz
sc/yMdJiGWW2ICMuaQJLssNd6fi5tgC5DUrUJXRLtXg2lit7EFhmFraurnjZ8QvnxY6uamAWxZMB
MRT48jTXYNAz2JOZerhl4Y81IWyH/YWruXbYIiAkqdxpzSFIPitf4dXaTDbXYQJEhJkQqSyY0AX/
pkPPZqLwMmyPBd9fdp15lCyx6cr2y+00+NJ0Wy3FEgTtvP+jf2BGHydSnzTOdYfHjCjHV9vjNn6b
2Gfno7u7mNbKY/0eLIQZBixzFqDGf9Gr5yAdOF3XvUTow2PTbERupZ6PA6esJfUyw3H4XOKEGMDo
b+yg1QP8DxJiHM+Db+o7dBGmyCyo4J16JUrPa6HlZVzAFq5r1u0bND8zb9fyzph6NsJGD5q1mXtc
BT2uwA9uRxmJnD4PyPZVAxFnM+hyAwhcxrqeumuLSxntbLHYH+3jaj6wOTbD4z37PTLJogWPDKzq
MIcw33rKv1U5PXkGnpjBC+5jgwaViEmhzaEXmzQ6xamfNDUIz226hSwtq3ZtXZpfJSRMYxga+35I
zxmQv446GR+DLLrajHfjnQ3aQKK2S8D2Wxlfc1HtEr6eveGiDuNSzdTGLLNaVcAYMtmqHRS21rjp
7tt1f4d0zxS0pDGvhxYYSqPnHdBsKKuIyzwVFzNeSvPNwGvQz7FhS5irRebiC2TqPQi++j8Tdxja
RdF9HpeafegWP8YhVdpHK+oT1BKFMiZxXKOhDb4vRYDjdnMXL8sI3T4aTAI/HMyvXl9oAW6AuY0i
lVZw5QkrZTOVG5WnDhCwytYXzuR4m2tk04hyEj+dwiW1kOg7TtDCId1BZk4doP/0V21RBFNzL/4d
AcOue2cuOPoeyK2r57jm7RB6PYv9AEbbev1ciaKOZgFq8W5l2jnTtPLTMwXHFrQAHKFTlykv4xrX
GfZ+xJTyzg+AC+SMqulljwlP1RzeQI67XV7GdXVvFtd/7AdUshmzixcyRBCTHz0Acyk0JiAR2XJe
OBvePdNev/uBZF/3bb3VGzWIG0C7gGyBZzLC0A17OldAC/apBV3Y+llP/agzi2Pz/nrigNP0C+cZ
AjamaSCPB5q1PzasMm5HvWFvv+52IYA5D0nscbB09lMcm1KsBnx+FjapPCkPS5M37plfR+LNxLrP
f9N6EbbGF8SroyJKXccplJvprqVexjAvAb7pgpC6EkYb3KcLfjpBcHRFak4Jkj0vEuPzpg72tJY+
ZqSWEgjDMpEJmDrA+MwHvMc7slwDANurUPmaJaEJY2ooOoehblHiV2WyAk3zFOKywL2QLVb/OEtN
UNollP3RHXMKkApHnchGlX28x1Ubx1HtX6ulDp9Y9QR2T4A/rwtuREJPFJjSnrbvKuA38z8msx1u
5q9aC8T2ZNf2/LPKFhWLiFFiKuizsGI1ee0gA4hlbXR+6rzrmUSIeqCKqMtMkA9uvEIaqAPDVlaF
EQDN25u66n+vNu8FcJPyYOIbBIQld8dZS9AGZb5odZZeWEkYqe0qEINpndIeRaqqrG2pH1WNdP/7
FzZujGn6uXiYvAYvSKEU7UxjeX4roZiFtEKQXda7V2sxXEmPWG+CJ22Fx2msxZrv0N00YeFSAaza
xY4GiW1nxLKDEbIlzXaKCy1crMl3//GEZzXGeGJ7xZx1nRX9V6kDtKeeWNSSZ8uW3E3diSOHI4wq
ZHX+b0wH2+Mxu1kRfbY//TUT7XwSN90+DwyraZkgsIDFNC/5yRd5jqenGJ4c0WNqL7jGXUrwMaHl
sVsi4j+t6+TtmImlzemiy12NBDNF+EopoqYs86OLlSwtUJiPjeCwa6ZsKma2KlpaXZxI7w872Vnn
zLdWhJen+pJtu+T48SmI+eEh/lE4CrBzTTHRocX9M26v06w7oUNEK+PEaD5AStRz6EtHxyW7UkM6
PmofWAgsnYKrxD2yZdZf5twhVdH0Lc2VHVK9uz40ip3iRRNmL7z3cY7Jz0uCA3+B7rdvSMtN5xV7
NDdPGgtkvqQLgdFzItN8FcFSVcN0rXFg1NTi07GjTGg1fV0f4aahaD4QO5Io3UtsNyqF6G4muAg6
r2BhBRslUaRSNtWp1o1Ck3Jb4D85ltufYPwKylOddj4hOG6HdWZqmETpQ9FzkTm18w378egQxWVN
Vy9pbCUpesMM6iMutwCuqSA8COBHxVyfLL+L5HUFF+uqfuae8D8rZzDMOu361Frf1j6ndO5oZ+kt
cY6yYokziKiDaJK5jxPcIRiy55UyaprhScM5/Mc7IXAMy5mK5cgPM8d3LkgIlUlOZ6MnElGQ2Z+N
jaEkf3JpwlFxQLJDn1FU5cCQj66kXIb+E557w0F8JZBmM665WztGLpXx1iLpC/kl62YO0SJSVWv4
nv7GpISKFskfAJxAomg2PuDqCGDkqDgRrgfjLmXsd4BdxJp8ntOfDh0oqGCt7nQVwY3fIwvnDjwb
y4umgvU5fkfYW8fHe67Y/JBOG4vWXVzg6T5JeUVNROFKtgwEirg+Rh+ENXKibIStwbellZrIxwFe
ysbmH+aLfPMVf1KlSqyfhy0mQTZzmPGaUN8/JpQQuNJkUiSQcDHjJYWMsZu21KUurtEwfjWFSkzZ
CEXMtQCcdCKsIyb6bopGlnxNxJVCWpHg+F1MuYO0m9aXRuBrCbBloYXMdKwzOsPLvUne9nlZ7CiC
C2Tr7XtDjgvXvo9HNdIM5zKb+e6P3gpOJgV2D/jj3IE6OBH3OPgJyFngz8yOO7wThh1ndTBZl5V6
EFtAdFJNvGLKrfktYvz7jocXjvX4dox36IKNhwZDF0GfHdE/fXFTctENQXxwazKd8XN7fT45w8O2
AiZbdEJPW+r+NptMos6ZXnyPJml/J1NNJI80mmAkLK0bbLQFSgM3BdcFJ2cNZHhJQUcTUxC7MIHh
sUK90vaP2GLIIUUnTI1Yk9zGKEIuR0Vi9gaqdwAaOyVQs1C4bgOCuWk+twAYu2F1rJmp7unhJu0B
JsSzOwa5CB1n/3zacVMWTuwqDMdJT6Y2pcEx4QSIHmj1Ix5yR/XKQ8obYPY+Xf+/UP8c8qyaKUhK
s3ldsWiGyV/5IzwVz8PoN3ecP1UFZsZKbXHmOlZSPwmuxQObQKOBKLs0UIXodQGSrW/j6HvO9iqS
qCpSFr3ZztLdeer3fOnHLkhIHrxrlgRKAfFdTcEvf4hIDDEy/7uhIGwkpLC9mdT78aRQSg0unDqb
ppER/um5+U0S47XdQD/Onk4GbhEewVDq/OqUqmKMH/Rqi13dFpCt/N6Xe6owjoVr0YatsJAJh9u0
8u41ZbFnTQJd7JUv2QqPtAdVX9CBw+UBCMPYV/R6opGe72DtiDrIYhEER53Ww2B66EkVWOlupUMq
U+uFxxuFQoqOSPgysJCwVcQ8x0rQTiCax0rWSN6VA1FndCKTGYW86BJ7inSGqCVCXFT9HUUuL2pV
Lh3tqUToJNznwVSC2xneCux7KCnLwLhbpPHH1adE5n+oXr2nnKOqlYgAPb+10v7sNrhCDCLBBVAH
aI/4rf21HvQDsf3eJFJyOfX0w/iuPacnf7AwX0jVqr8aZBNfAKS5SdrOegslpBEgXDprtOiYP72q
pnzk83ZxXmbx53IfXSna+zKVy1QcP7YXiWaGwdoDv+n5G7ac7ak2SIxHp2MUs/TmeLOmlWH/IOlr
m1WBYjvCjlvs85O6xVKzW6ERaQj1L7znM/dExvazg25VBRfb20nv4E8/LRG5UqDfHKPosPlj1c4I
7v8iarlWzsvS8EEsJa8D2+MaJ7ELbshGSRd4IuukPLixLmGOxO79sgfYCuvYnU2zbqeQ8F3WPtBo
fTfkxUDhfHcj+ueSdZX2nJYmhVHjJNziMAVLXDC9AXj8ipI1Pi3bRntfGFQsnJeC1okFg1cYzrvg
TTz7wwAk01cPafsFFbSfaTvre5GjqKz7vK4Ahavoy7nMlwv35lilGxn3S12/Te9LKKyZcNULaqbz
uMh2bjACJfHoUKAF/vJUiVGKpWyzXyrDYrz17giYazo2xIZW9EQtqQeVU2LXrr6GbNopQeqBw5xZ
QJd/v6abA9EwcJGmEBctZV1rCU0rEQUEPB2dhGyRJEniD1P/Iz3Q/K/5JlZqcWqTMgeun7DwAR7n
otn1rkE2ZfP0b0GAV11FcQQR3776xJFsza1foY7fcVfawUcmDSMSJfckOBqNxvziPUpH3biDbpKi
Wnftn2tXXQFuubaoRfV5T8icnQyEqXAUzbJGi+F8eNqGDi6rP87BgE+1sgKzdME3hWdJPQrRFvCN
bkFiXbOoRZAHJISmKQi/mARwQPeb+dbE67RN5askAzTq2wNQZUZ+IRBtSRZWs94i6GpRyOES7BhI
DXssPYXtLO1ostnbtrUu0nn2tteJAonT5XaOwoJL31H6teBIp6nuX0SvAAWsbsnq0szHtGUgyRpE
wl5txgTbO60Y2ExY79FkpSFMVyKzpbf2e4l9d8n1vTtJgDW2MLgIK8fhvTz3pVRMe5uKnZzgzRV/
lSJW4cbYxiFVvtZYn3NEeYLkpLDZ3uatrPLtZhLNCNLByncLHGrVs2CBSvodl9VJILIBTc42cpsC
QdbmvgoSiMbq4rThTONa6aR6EG/aPa/MZeDfYcobHdgUAsAKWiBH/blM1TMptpkXBKRr+SdBp4AD
JKNGLLeDLyVL6Duv47lQjAIyfp/I6QN5emyMZmNCWBIfpxhCMRKskYICxDuv+WnbTlkAudBIq8+E
cZlPJqBclWFGqQh/tG283t/B3OTEAR2mvgpMJWE41P9v8OgToJkYlHMrrEi4ynn5/8tSGONd3SeZ
pXMUloFoiE1NZ9jSVpNm6WQpRA8kg0rh1t0muYTlLfb7UVxxnnSQvaNE8YhMvwJbPwxwN3o69Pk2
4wMDO6Lrm4B9ZXeXsL5iVroxeFQKFxGyFKjxeZfBeBV/zszoSOMFyjJxUa+UC2f6aEGo28aTVgCx
4Co/rNji+ejVCz6azNTqjryBzSobZqbuzIzCWiOz2+Uc7pH6SMHCVngRHXzNjAm5FIPzeV22t37I
AlbZmO4vUiXre7gaQqLGQWOVkq7fAfF1Kw6eoOYddF+M7fYqSAyw7OedWCpBnoV8EybB/89MHJ7L
KWdVhIEZJbAaG5Vu79ZSCfQM70wQ9VrvziBqnNIN/QGHNZ+A/3eYbHTZoCzuOou1b0lQkJDJ6jXB
HhsaYNA18RVFV4IhaRYE5r++vyyDiXomkRlJXf0MK7aV8v3qQPLQ8op1WT7WvTJKqVMRpdtK4h2L
rd/38aXEyA9lhKmJFDUQx25A0Ry9BoZZDin1fblHn3U4xsYP04S3ZcDaI6JDN+ORY2U0V+CMWXeS
fSn/HfrpKSGp2GOLP0wy309gt9QL8D2iZv4+mnaDEDzK3lQrzZ7bwtDQ0Gu8wWf8bYKGLuYFOBbM
pK55/Pr1L3gfvmc6bWdIxGL3jkq3Gjx0HkN+BlJIYfg/H8jQLVakTtJpdW5njCa+6+rHraEJGhZ2
VzmClFkFYJpzkF7Ke5XUPRx5KJqqXwC2g69mP8+pLryhpGQEZxKROa+uenMVOnHvDCcAjscZf+1f
YkzMNqk0Me2KfFY/vQV8nMs1JP9bNY6YERfa7KqbqckhLBYXmvGYfApqftZ1eTJLvb8ZL20PllDC
behTTk0KXRwa+3utnSrMJcVYsEKiAaWQylwN1aemEOhf5ViAFEbjmi6JEPHTnw5KRS0dWXvP2cRf
UWkia9cPiZjXtVYT81QNQkqO9ldi9FQZt6vqDyWFGOJbWmD9hVUZyL07xJl6I59qoZwEROXkw3qq
pQiEuFgtrJI6rDzP2QqlKadmenkUgu2gBd5fZ0hO+UjYvnFaxW6CxDsUUGDE5lgL5sQVUfkmasMW
han25FXEN96bTLo10BFFsm23Rxn1ECde9Ct/EgCu2JtRMmrUFtyiLQj3Krjic1pwrQWkfhJB7QK/
YgTBaLiRBuaUylpZQFdfd2w2nSE7gxgaNPn/ecCH0zDFAhOd/fBfPA9pU5fXPjNSs+LRVMnEwuPs
yG96U2Buenqb9Qb45JuHrNWWcMP7/lf/ozfrqf6koEETzQk46X1mMVJk6WxVo9wO2aSl3x3Hj+aC
77XeJXmB4/Z42DeN3bkeLcRTX8axUybErHSXBSTv/IzX8+kqaqkKuFTnVX6nogiQGmuw33ml7BW+
CjuK8Rn8I+lociInUAaL6/mE7GTa1I8ueiaOvQvjR7ZMFX40SlEK9gjgD3QWyRcCQCOwym/WURAo
BOVrNjxypez4AXncmTB/A3ROKx1Sm5hWOq+XreGliDWsiarO0IG7/muuDKEr8rKnzBZRehyUBXdP
jhcCquNbUwKo+2nspqS5ZB3jV3LxMRwChVzSrLVJLA0jdqWEEwGYaAudu0QjlCEBAbOHZIAYyurE
PSaKvbeTHu9whroPGXEuNcKqUlNS6+va2cvewhBYSimPpWsllvgZrCAqBCvbWAp2DHeR8OVcpv4h
2DNSILz6v1QDnwGBUxd7BHQd91D76AnydG4obTgwufLcXXGUljvQMv9mHIXM4/IHyDNi8Pyoob/F
7xBa/6BurFTa/ew7jiV+2b69tMLpNQaCPJMnhyTpvuwqEK2UkkJx/NgANdGS02e161JwH8PU4LLK
yqiWkghJfsaKmJvK2DKXLr2HRRqDTJ5iTdURChpOmr8Ray71jFj4L7iNxxDt0WP/K3siM3o4oHTG
UbjaJBSBPN4234NoDEAvWA2qcWyj/B60cYifDhX5qEDaQJI1+5Ll0LjU6HEfYZS14MYCmiRArw4U
bIqtjiR21qp2IySnzTPlArf+0YNeFXTRLtZmHq8wT84qlC4Re6yb3t2u0lal+dUb/XwRHFfZ65Pn
qQrHX0eD0nvoNprcXz6cJTvCHwBPopZqbyxoefKXmJboTOX8J5UWW/4pZhq2BDg7gqsW/kzxKUNp
VqFG5za732qpps+Al5ZyAujw9nAjzgENbY0wH0WmCeHFy9rjqoU+2ykO67S2ojzqNXxrRw8FBBrK
XWnJ4H6cdY7xUcaPQV61g/Wuzb3DajJIkCKFgNwiTdVJ73CSmQC7atkUk2lkOoPBY1GGF+htXB0b
M3953OvuSn2vwrSpUwA+xBdFqaQRYnUseM9OaRjom+MC+eY8Fue2AwLYEyLroTp3Ya0B+UCAJ/z8
czjMx12AIGwbwaCQckZPrigdM/16ZITcrtAdiO3S0W2PJ6rvxzBw5ZgsEugCjJ1+QGYEn1QrDbH3
pWwnh7LcOr/r8sm2YaG1cNduHquoJ53cGyE8Jw0p6iHTlnI+hXFYQSSvTBY43TJHGWXX5iS8KrlD
8vzaA/vWH0bIo4E6W0TX94todCDJjmQa3XyKDT94c7A3eFXWwj+v1i828dijawUgxXwqB/Ai4X1x
lvQFJvMql5zbgJ/kj0shG+J6OhhaZvc+SUVWs0lveWxbdf4ZX/CPKROq8nl+9LV9iLxX/k5o51ro
gS1Euf70IMFaBefWBRdr6X3FYQ4k7TVbc0F71TJSLRcW00BmDuSxhP/I1yxMNruOSZv5gRJ+zyir
hliCXG97VG893GaFJffPnI18BSNGkYHCA+EWWhcFTHQa4Fol8jX/NkNko1biG9WaDRz6/TYpB5RL
pGV6mW+k+uA93SjecwN5F24fQ3CEm75GWvMpc5yPODr4io1mnMekWrJZrzsEbOa7rExpCMIQiDIX
Qtn8QPNw5jk11x11dqapv+J5wMpXlXwOLrlZLj7TBpC8irBD3zEKeCpQbe6asGe0qsYHkspJpBmY
SoeKEKkPdc1jBSxwAVtFoUdVMXmP2f6xNTPCqDNqO4ESNf4f+eCM6s7LF4Q7wt8DNWsWLCnRhUT2
xf4/NceoIEyhY346I21Mum3oav30yVOm5pKza6Aac0+GLdeTmfncL4g5Cea6Xp8hiHUOPzSTCjnM
PqSbPO0GestvLn9qpKQ2UHfx+EPyx1EkMgAUao4yEsTPU4SJdHJVwTPeJyJUnuVQlZus9QX+SMsp
vBXV+5FUmMMC5RZ4GAobQS/i+0oQLgqM++N+rxS/KAHATnHRQsJ7e2CxQ7FXj0qqJWWa5E11t5Xv
O5JPPo8c5bpoMBIpQcinMAnQ4uOJlNIx7tkPmZwV7edft9p6dco6qkYQrgXRE20tClUGe9Zc7mQf
SwepPYGX/Ae291x7PHkvnHHubSXx2fQmPVN0o8WzoBpyj7kArKXlRXwaet8hQwLF8Z1ktfDo8gsg
TB8VrAFVQ4Gc6Kkpon7TxX74TB6RGLT5idTSp2HYAvpmksovgoqZAvJWVMwd9sbVBS5QPvpLXpwL
U/9dPZuuYuKQ/xXcXsvlne8iThrvx4LxW1kxLf07ofpcHs7CMNWZPmAyG8d6phfYgZInIwmiIh4a
hjb6WHul1SgGhtz/kwdRhqAj5yq+M2wTPqBDCp4uMjVsdLoHMc914ac89GpCLqAaMx9FSA75Re2u
RJJi4MooGkyT2hXcznjWv84n+VQeXNyRqb9zaD6C1ySeptEp5JhsYRxJgv5rE3/SsefRby+Z4/JA
yfxqM5y2H1c8+TRYBkg/HFrbAqNi261nUXmWZx9YTRUhuKgrBw9aAj+BcVhvR9EHTQsjr6JHrO3b
K0JNoxRbU3bpNKFaXHh+oUEgDAyVpAHiyi2u4ITLpw7G5uKNCnzuTgcKFmNtHTcGZnKm7jlMDI6Y
SBC7Hnl/oeeh0TkDz7cbO0k41Bzy/xwztirRUP4DgTNV9koMF2dhT+EMKRkXXctg1UzEB3bPYPyH
DdsoFSvmp7Tgi7rnv2ESJYYS4Coan/6OtpblTrgDUMeVyOMWLsCNnGq20CfUMtVwizsLtIh+zGh5
jUwdrV9Ew6u1HUPZ+83SfjLgyBdYFe14A/RgzBQv03n8QVWHoKKpz4ilDFrFo5vkJj08Eumnt5x+
J1NOqZKY9v8I4am1PaGb+a212lZZlkbJhVs9Q/Nf6qLiLXuWSKQe17dkky7NV6QDY0jRpyMQkb57
DGywHZXr2fkpWZ1LpKf+pVPon9JR99onFk3b4/QGHhRO46N317aZiZ1uI649Hq0mxgsSlyWDJ8Mq
StJ1pI9ENPgLZ5X0mBk+0IIoMxgaZlAqCc5XTORYBWGnexNfcTveF7qAvhVYLBcTHfxfa3EgYtMr
gzkMCr4TUyfCb9OzYWnA+nZA3NXoKcilpE5joxAimtkpsZAA4kLvUfuHxknemNH0GxXoXB0A2Z2c
J1o1zyUtoKQuWroLLlGM3lE4kxsa78mT4P4Yv4hPxBFeXQs27Z/HXQl8UjDsh9xJUoqEHiQSGHg/
PSLGpsQ0qp860Ls+ZZPB0mltdHK+BFaYKH59uxsHsL2WQ4/yxkcpvrsqzx04b5is53luOnEi6GqC
T7dYHRq3RWxTLcpyQ7ZpwT3zGaYZ6/KjIrtFSk7fx/gKgal0Z1HGWdLVwpJxCiKUApz9NaVaK49e
VFK7FQRPalXMG4d0kQ9uds72zxle41C1q6a5q/BPYfcPabtT9oFUsqkmL4cbZANbiJRZj8F0Hcbt
b+Kat/z0yRRD0hzFuUN8VmEN2HBzmGLWFmOvFsq7VmvtIn2hM3Wyb0c5pO0xifmJyqzr+3ra2M0T
IKxTtrO585zcSUfNukkFpHS6iar6SiI3On6GFAcW2OWQaPwJr7wQronCFZtecQJYxLjZirvu+94H
YqPPsMmrGtwb3caxczXbPz0JRpjY9qzaKhdFei5W89ZzJtonKbfTQGtBrBoQ8+rHRdXoadIpg4ln
0dgbMOArHlXRnhvBdnbxk+eZq8v8Nk4L6wOM8ExXlLpavV5DpW3G/wxzfFAX32WvCnYk6Alwn0sv
2pWvbxPllgdb/F2QXDc5Qj3gmzdgLhyl2+GzSyRheSF77OX8BNwUmqaESLVY8S8iQw7P7GAd1qFS
Nmb1lHUU2o50O3Y6HjBiYBvoT0tt/g1jl5TSAqEwSKEsmK0ISbZYhNIkSImne947A71kXfTnLs9/
mJ42BzpXUwVddCIwzl52+9+wfi++RtiTUBn7M8p7/q8wwqHRoOGoGQieSA4kzv3XecVoHcixCrqf
ZLIdqL6u4LL0/LIPy8zdH9D5FC+XcGLmk+yeUlnD85wU+myL6CVq9d0l6JEEUZ6NdMwwWkwG2nMr
dKmigVlnJ9AU5qL9qtpQpeQA6kqwmEEu9LeQFBtIoyVHb5S39UjJyv7pesvySDfyhtdPm4kDbCX4
lEwzK620HDBp3O1PgP89hlIim01quVxNr0U3Pvq3orCUDZcG0UlR8sfo+MZhV5SDEN7rpyKfury3
S1zGiUCgFjrJXFDLtf01bJYMpMn21Gjv5Lcb3UmjvucaXaG42zxaYcbPaoHF9AIoeEwcqzmPwPZ4
dN7BGKo1RBf/DY8TXM2X5kGd88QE/0ywovrQ/1Afjl8J0Nl2+HhDrzLvx1TVbFkm7xKoLxQuXEgV
7ymtKENLnG6rO/ya/DOh1eI+IKi8VHc8CXDjIMChaYG+YV2NRWDPzo6kGGSLC6obSpheleLxQ3XH
Fs05wqyVsLl09QB1pPmHN7+iJJNwD2Earfjk8DQDbKZAsAAuEaJkk6WOik5bsY7Hy0YxEynbpMUC
8Y/LwvyK6kdp1A1MEfyJt5OFtQxUKg9uldeVPvMXU1gAFGMnSuCGytGHQBi2p+0Mvxd4l3JfBvlc
xqiUHjQj8FwpYCsSBcECsenhZAsSE4o0h4O4qQv1IK8UKVA9pqi4FSUg7dhYhdBUwXGkkYmLYlp3
1dloPNthfU4qVVjyYhlgXtcZY5LNeZkOrRku6T3bPyM2ZgkmmrNTsnbBjJRhvvWrZy2EaSI0dwjA
5XVc4vcLtxjQN3XBXmXd/LYTWeC/psO9L/QvvZc750ubAuPHZFm/28IjOfaUegktcLNzEfnLIKmT
/FKCJtm7INXqZfCVl1s7ertvmvgjkLQOn3wCYnI1AnEU8kSSM0+3C8ZzOVhJKZ6UbRGb/RHeKsK7
QUVgrYdOi/s/losBLO3rfPWFGG11wLOMjU93Bm5n2WqyII84SIlp2Ri2VEAibY1TVt/aRbE5RUP1
mtOeQxp282torHDhK1X/qgWGLVyeoglUDmDP04gIZMQEai0b2uC8WJIf2FpnfuG7y2OVats6vPVp
Ti0BXa8sITUX6sSapOdFNNvDi2J7bk0xSsGecprda1SzEywUJ05trpBu1QYFF9pRYmoIetrP/R/I
p5ENgG73zGsg/4JlN6tJPpXwDytf75SBL4J+tKDSo8Any1dLzpDl69mwyiLySc7DvonIitufOtwY
2+pHU7MOmzTuXp3TR6uURpALpIgcwvRdryxqYBBlPzAkGHrmecAuSmbnygQ/eCp8cxpXsdURftnX
NK4y01Xb1nXmRnCoc5ftikogEFw7s5YuRlwGltMBXqXepfavNinZdkq9D6Y+16JCe3nLDOxXJaKf
wmqVqiTZkddzcAhPMmw8HtEqru0C/LkSY0i+xJJTuym4ziQFj07NPzAJShfVzmrXwvGaeC7lFLyi
JQQn7WOHv1lLOjGyAz2WBHgFF0BGCCKmjrbmljXmeo2xe1afhjHz01F7z3/lIlT0+KvQkTBmf8x3
hY8IzXaDGt/0REKBGsCgHYi7jZ4ZLikYbeiRp4+f+/Vs8e8w/qCeN/7nCILWP8skMYAwxRZQLBlB
c+s7cxA2BMAkB0pKZ7sSvPs/unSvOtzH4w7L4KKHfmnF0DSvYBInXcwRFtFTL9tm12Pjhtt9ZpPN
tVkUfEshbbVTxhzQPPjjCOKaI4KAmHmgHahAWBVWwXTZBjAluRVlJtXDgePz/j2Aba3SuEwEmIVm
Jf7VpE6dVWfLftqThOhoQtE0UB1Fbuf5l5sw4l28pDsn3OHTe1so1/Zi1jt1XbX2SBLhaQSlQoq/
FMKkpsgdhlIv0JGNGouBhCCAKQiNu6Vh5lAuF4px6jt9MgAEEU7UTzwlH/0x/Zg6hMb+8kCc6F/F
JaMeGNseIIi6/pgzndOWfgI94l7ojW72G9VAv2QcNWmbWzG6HsLxvkn/maeV5W5Q0BXy3uzP3miF
61t9854iTgNbgHdIV1sD1SuNAgVs+cC8dmrL2WABD4IycOu/lG1X6LKOBIicofsh9CtaICAl7GJw
234LJ2dZpKP5+Taoe08P9AqQFfeB5L545Kb890RmZsP4a9cFC1zq6/tYOI0fhptg6prEc6HFjPPV
zKrk7whbWQrKNZ0S2GgwEcp+5K0r4zgTuW/gnLSTzThOVYhWn3Rj0DbKa1S/mj/YZJB7R4nVcEdv
0hxFAYoIh7HYiPvBUvTFsgHBVHq04sezIqQyuhDLDR44oHTbXfm7bx+E8Pd3rt1VjKt/xLCC3S2Y
pIYd0EB7vc5Ka5ZokwJwG96CkUBoTKeJqqN4GbaIsE3wplxVI2RgJqVUdLlrbmQApQ9VjdieecOJ
fZev6u8vPwI/22p/z0W+IodzgzaYuLTZENRV4I99UQyJPjAaSIRmRfnEcw94VzB30EpxqOFCSQrx
kT81jSF5h8cuuhlQaWOJRt3+AXPfNFbakOIDa0oU8NUVHA1sAIKL5VY0FgdJoVB963W5RbqlV2mH
IMSyfozAaiZFyvlDMlZis7kX+oixazZo5DjpnKWWV0zsvY63Yf+/n15x+HeCWoUppaBZy6mz10sW
I2s5rVT+H8oH21Z0CmfAx1Uy6BQaeBrorIPlWuCoDXLLcN7o1gr/jji7hzcCcRxh7kXKyT1isLqJ
g2zs1nb6Hqa9Z9RFfWFbMA4krvRpGm95ai7Uj8UILU4rvjNTASeK6OGZb9lwNTMU13Mm8Fbw0dlS
UwhAV64nigaK7+AINcuCIjRO56XKg7uMDZmXyflcQQsqO+a2nyasYaVpXFHd0xPTsQSrAkghrFTU
TD5UsFsIZagptgbMyRx3gIEcVWlMha2kT0ip8tI4rGHlLpwm1y9lyU/N/Zy3ve4K+71bmak1+V9U
oMvP34IepntJv5/XjdE44OCgkrIq674EIU/gmpz/cGMz+xhvv6gdthT91pE474cssqCkgGxHcaVT
O0us1H76R/pURvNFbbIoFI0hOEkcZwho0qno+l7/ohQp6TEgOFTCOofHztXV6Tiv6eYdEXGx8vAa
HPkMzcCzUjTqZKAW3le10ZyS5uuaq/YSsRVMW6NEmxUDTh7dl8xpwVt2/PQKkbmP2i0ksVqpCavT
gjHSYH5WFoxcME9FwrkQHBTmgXidIUupicnA88+ZXAN+98WqOz7nu4rIkCOxLAHq3rYv0jVBGOYA
cD2HJDaT4hh5CluTWLgMZ5FnMn0FRR5GsIkAdnEP5/ajMuvqC/GKZhoKDDmXDKFNGvfbTZlz50r8
G2agcCwt0MSQi1rGJljwajY47vQnMMZZAOXMq4Xxd4CoVOUHxnhPb3SGLfbDsYV4yIKZN/oftybb
iUhm1RUAMGvIADACoxLUhXHjmypdg9JZoVx7HvtoCsPmJ5qhoGb27qbHxqYU56yPf9vTlojz/PVn
5GiU+WdRVtPuH/UWYxFvOas/7NJCZbEB6xOs7U0hmPMXQGwVdUSltKUMSPsHfmEJs7LEZA4ASVl6
/3hvIhmBE8dCuR8yZXM1Q5moEnhqGVmpUKP3MRd0Nqkp/jBwvOLj44FOEdy5gpWfNnfUZC1yunfE
dvfqSCKipnXGaQkiHHl6dPWYIn0yThBq8KQ+H7C7+bga5a7qnnyawa+DRgMj3wR9ZOVEKhbyJqzZ
Eq9uq3f/tR3fECENN/6FItOUTmPSnwdM+KUmSOTCRXlAAi+hegcYuQFUEwMpjPRF9e+vMdOQo7of
/zOmkcSLksCdM8vShCIFprzberQVVYvv248/QBA6+iIE5Hy7uyKbAvZbkF838M92du7uDcz9hqTC
hHRVCu32ST6xdM+eTKQZbKzFofosAn8M+Wqvndud/oEeaXmQuyZh4QmeJs9yyyfTOlG2t9Nk393x
ZkQQlfjyrgW5lhd+yEov/XOzB6oWmVPPJ3gTZQK3zrbEuK5VU4ft5/2/f/byYgJtSgUBoDi6RfYl
SI0KF4+9tRH9Iij7N/eYhzhHzO0P+JDTg42BCrWjuBgxGf2HZi4dXLPAQjgglf702NUqTSxaFGnX
FzuJEjU4GKYAyM6rj6Bf8byI9s7Q2RQvznodZfDLjJ/gW69B5L45JN2KLqsw1sQiwSe90wSQCq2z
lndlDq/xIwzJm0qJlf5PFucFZk9NwnzERlQNeJj2WZmkMowzkznG3ZmcvlbrNw2QeHwSJ2kJPF3J
NTgMSJAKswKn+bSAsAcb3D/UwW5RxREN9Eda03ujHk1j0bIouSknMHqCZKBnsL5r2J/GRFny6ue5
j0J/Mvswzvx4MnCXVM4G/4F/IWqlMwoIYNCVY2q4ZRw6dWytHFk0mbvAXoqHkXJc2dI0gGEVTmMG
w1TDL9Hk9jvg/xfv8/6tJwv3PcyAJzuQKncO4GZEAqE38dQV18z3+wrFuVrSpDgfbJ9g+UnRQwKc
xdSgpTcHP35ktNohSpb69CXg1huiCIJgd9ROe4i2g0Jc/3bCYn7XMUMZ+gq4f2veCr1rxOBkzrWN
yD7C9UlN6F4JXuMwuaFxRJ0orlnklxPGPouLoFnfpQBdZB+b5gWndRW69pFSqA85qwGX0PQCUVqR
klqCKrdMgWBaFIJPrY9YQkTxdFC07sq0yHA900Xnpbe3QsfHTqDg3njG6KJMH4tk2lQYQapH2kqy
O7mYZhWuNWYPq6T8x73e511vzo1KpqJOXZIyaKFnT3nr0V6Y5Te5R80a3+DxUcN1Yt5fu81pfuC4
0JMKhFklX1fn5rVeX3AbTrnXotalm/xnXu9SLC365TQPHVJvmvKDivHec3M4Ah9EsmwtT/Zdu0cG
v/a0zzksOwEMwAWiWaCjjTFI45tieqSZG7Jng2ZgBthBxxcVFNBrNeu5zj/Pm9l3wB4VYhcx/rNW
nWZtbBVvYBuiiaDr3zNAi/osl04w0dJAFPFE+L7rmUGBsJlTkkNyeW8aQRgzaO99PvtEQNflk2t9
1pnhXOg5/uBLkJ9qdSrUovPAreBx1WTIzp2eXpmDhK8VY/hnMuLbcgVc9Z+kgCUBByfI74is3/1f
R8Mn89rtkBrH5HCK9FFr0RPtEBMr6f8lxdsoO46yDBmDJCtG5XkIWi7HNxrMK2gU49NzWGBS3fGu
sOgx6ADhUR4eD6L9e0PB+SbnyKcYSxsAJ4O5Rmuty6zApooihMp5APtTdFhSeO4wBqGS5GtEFDtW
+vP1WrAc8iwG5zkwfIYvoATHb371zlWhKlTXEXqrYJZkKv7dfJKRxaJKSkyBYta8bPmKUCmGNWQ9
CJNYOW8kUcTgxN0EozgsIj01/6Wkg/nZfCWBSiweSn+3RdVG6NSsX5rUE7COe+XHlxmwM9RjugeD
HoFWyC8bhtnLhWnZplFUwdgHOybCoumesO8o1umwjynCIyaRp4bk0YREOEap5AW8SXOFK4Sfdf4d
J6BTObyhc1b1ncR+mu9x6Hmx8OHeGOFig8zLVuMD5+Y014JoXO/lNE6rxCTFm8D7O6S/PyEedXcT
t+4fktzkQeXwvjdDjSVnGHAs5qx/TXeQUmskVlCl+NI0Cr4ckX79vmEO48LKHFwjPWyK/tRZJUDg
caaL40GPpkz0f1W6m+VSaGi0/Wv94WtnM3AaB12c1O+4AFec6MRTYgjYlxNQERP4x5D0H9CevkwY
cfHWvJrpd2FdboDSrZcrLpjQeW0cvAOkMEZkW0KT5tnlzWca0G3FAn6zD+3ha2zUbPWHdyr9BvoZ
2Ot0aNycBzOZMcFFHaBRgY8cmfVQlgqcxenjlPhVCUBNFmCBg6IUlm2bWi4IV/lfYXXOxhuhSneq
32uzBleMDKD2rY1Z6tWwo0DYGMGtSqxc+NVPfrNl/vV7PiVphvT1pIfZs6a2b0/t7eSSsXxh+xwN
9w+qcFUGPdjkIQh8okSNxhzgiupKGCyN/BvKTlSFNTWECHlWPDHH2ILMlgS0n7fZfJpynrUtBh0/
NhcX3eSYGU0sCIOyishV7/HY6cRh2qQh76skRGufp2EJjGtGnvEJmWsDw7zsxFcnr4zf/RAdsjpv
EkU9IMZv2PgIMk5/UsgKP6vVzsGqYeDLyWF1LNWrohxVXj9WIT3fSiPVTBk6CpciQ1pFBS/TA69i
W4lJkUXvuocrvUkL7dIDly9aPjtrqP5ucLOZEUvXAuxXQVOrbTNeI4+dsqstBsWj5P07laQ+QmYA
7CSJ0ntDnCGqsunf7eKt15uijV4MqatRC9PkY92GDVRUwwO9h2DXppAqdLGR8lw2MAOVuWkR/da6
WZznt+vHz0w9UNjFAAmXdd56ObM5IZZCxbNBc/OeUGTGJpklWWDBCSuGZwYzyYHPWagOUijHYrIr
zEEJ8mEL/JBuiIcus9lJZYauW8CEnjK+2Yjy0gA99rN7CzWx9Zi8FhpJckDysH/LiVuzTOiyERLj
47ITFDaBp1wj7bRnafBiJzCcT0Y/69hYp9tof/rKGBXCk7YdIi31GcGAAeawvw1fwPiGaU4Z34Ep
BOPHOjnSiE27TDUVWteFcGqZXCXW+s2Q5MGtS+Iy2BHSOxPLi1nk4Y0BF1NJHxNj1WnPSxdIKpFM
rrRp5k+4YjvxLMQRAUJIkxU5Mep6b0R8r54Iud79Idq1A7t39jpnUI1BofBySy1NBqmnZLf9ZXdd
k96BgskSKXXeL62RTS4C/+r7qPDhTLQxMTNjWBsx1EbqhSrtxNJSaGsF82z96jmCkQWwhL+k0K0O
H9TAEWF19p8n6MqDZdb7CSQhFTDT8r8KM+BQ1M0kf5juUV2TekQi96hMHaP5DzfRQD5ZxnEuWl1n
fIxismtSl3WIOR25qIDig4PjlOddms04HFMEdvn089S4HfPHZqHMHNic7FWSNId2v5ta9PataeJQ
Iu+yzk0WYMzwHV9TlHBc4ZAOBNkdhjzpyR1vLtWhmVEY1AoLZp2zq/2i/+uTA1HeHA7m8oaOJlZ1
Y+VEzFO5K+wTBkr8klgOU8yiSu055+81rZZNwnb+82BDWYUjiSO+LBvgdaY5PAGoCtjzq050ggUI
vuCWxUGiHjukamisKmAFYHs3J4Tq9EVhkGVSSe/18WI9aW62lbxTUvgQzElU05FmaAUCUz82k+q+
+NApydmipJZz8P9BtItUWHKTcQ6hetJ4Uc3xhS876q5MWwN/cooiONRwxYkXQ0CXkzxI3OC4Y74A
orruVQHrKX7Rsjb2LkFY7UvPUCR9q6E5Vs88Gk287F8YYO1mQuldiw3CBLiIPQbmSjI1vhCJ0Xwx
nce4BE5VnOYWt4HHvy+xyWIuGHLUFUae8wX0JjswGAUtC9/H7NVLqKH/jWTdWm8TrhsByM47B2sA
Z9LnANz1TpgrpWggT2iBFm3XQUtngtpicHkNJdnMfOxbb1/HELEq8T9jwzeH5F/Z2Tb1KQYOqKhq
PGOr6erFtqZwmaBvo+2Z1kh2uk5QwVhI5XrDJxfojG3LQmpr9HY5Ivr89W72eKqpocNe96Soo77P
rKSE0jUXJx63gZ+1EAFEOp1X5607Rp+tR61g5B2WUGCSYpLcUQOjrxIMHs/OtD+Lg33GFXxj/jVO
QiF+p4h/wtpBQKSCn85Kxtya8bU37f7R0eoj6t5peIjre7dmFSbZBZYqkIlHS2m4xHPymlskSB8b
mt+NE96pnOb4lJH3mRFDmRqvA7N2HU6XzJpM0QzubTPm5dMBvC1OayUIPqdNhwEfVRUzsrs6Vmws
fEDJbyhajsI+Xk4yONLo/nxsjf9pufhlJ1nVI0wbME5dpi/NgsLbtsXH7vgOv/c0q+bKRnP4hVSL
rOMabYotxgNGSlTbMrvFkYa+4u8Ka2xpYofiwM2Zj7k+6mjY8YXIEn/wMiyqjEnbEOoKvMFU+H+U
h2qY3DHbJvZcomubYvvOiai+5R0jiiTNnwBIl3jkuEtfZopsd45XPkzk/t0ScudrDkUd4JUwcGCd
Y/24yRHrYTl486BedwEm8pxvT85pB2LzCnc5JooksWnL2D7RotlBlEoiW2/q+46UdYIXByztGgIr
EhRQbFfw47sdZxUFvoAo4oR0wySX9UEu/jcp92PY7KcRxJyFUAjl7jYXmMLdbIlM4oat/lBrlNca
I2gScOGVcVuyG2kQn9QK9f82M3jCXNKFW76vg65MssdbTuDVi6SCkrePjIAFBXSNzAAaevU6KYuI
AOPZDup2ggu3V6njE7oTa7i0u9mrPU0fuOI7rO9Zfi8Y7PtH92kXLqKJJeYE1EMfmL0mMBv29RJF
MF0DcGJoB44kkUy1d+JM6XDO5ajPSpKHS+n8iWQdSzMgWQgPWjZtrFUV0fN6rxEQ5fIuR3jBSny8
0AKxKYmCdA4W69Z2CvajZQ5S4bhsDk0m22ubUlTfx+O+Wj3MNhpAgXmGMLZrrslBjHChnUAR40pR
/QCaSyJ3S/Vxaxz3ck5DhcMDe+faTu5YPy/lL31aJW+IIJD+RmSM0ZBx0IDBEFNRUAPlbTm5f4GI
ntX2E5TMHhEhD2ofT3PzypTlySXE2S6fulyfVTLfBOEZVDpSeL7JZRUkdFWvBrvi2YkIxFMyf/g2
PlC+cm8RniISRfg1GvwwKi2zws1hYY5h5yqiVxxbkKBABw5SP+BhgtlkA3nSj7eufL2NOAC7t6me
L0xxQvtqlDTj6uHg4iub19AV+0OmpqVRJblF8+EX+7UHn2Ck0HoxKNv/tENDqG/+YMIAUk2BiO3T
0gyX9L1aZChfJRdYk1hxqTWrgoQwAcRFFe5ypC5yk6jYdPlsFou1D4C6P/wXYggKsAcWqD/icEBU
/9Vpb95d8ErFDAEWTXUqdFxtRGahDB70n+WmEEecLQaJZfgPJADNnbtHV0HzGepNuKQ7t8gziAVQ
wn6RSwQ1oy9ezwNq14s69ie2YwCvD/02ZbmJvaxaSaBzR2UxkiyaxIDoy0uJfQTysqK2k8TavmBK
9d9BW9nnlHCawZz+HS92i1NO7PIJkwUrU2vjgL4oaURP1psLRg/l/sqkv5WX4mxPDWsLQsAlH22Z
xNUisfX3rRbdrsm1g2nDU5VWTwnZ21reBm/NK+dh4o3qYSZNYKvrv7qspuUu3bLNh5xNZ4Nsk184
3OzdKBTU2hcJ/e05uKtLJ4SamB9WauaEK8+yQXHCVtXeVxCEBf88A+huagIoC4HpHAfB6OTNUVdE
vEP3prEFB+mhEK9DLVi9GoKbPyUJE8FoFWlzWlJHmQKYcRJp9pw3l1Odh2aV1rF3ODzDj1u9n554
NTe5fxKzi2rhipIGsGirScM6nE3tcZ5criqmp80i5TXS2SPRelnLW2EDRUY07BW8D+7oO/O/NF2V
glUcnqxycJFldjcz8lOfl7rXd6rpBrFKNJNpQj3I30HoSE8Z1sIpq4V8Yox06BmtLHhk8zKrW9t1
nB9CK5cwKp/7PRmo2SvXnzuAt75REkmBHwgeZAdoW9BfHyeewjjvmak1eP+GlIvf17DId0tOjmzW
2CQk5mJEpm8FAqXPLBg05LiwmqZGkwEIclfgLXcok3q8mxaXE774TDroF3muPn1dklj9f4BX1BvH
87qhjW6SfL1JKi8KdsGlEbnZdlTn6qwDbp7J1QVyp7/jnFAIl9H1HmgXx5HMJ1V6LM4T1RDSQaa8
bQ2vPpi6WIaQvXHZ/Nu3wYMhK9Z3fYFVu5NfmhSO/AH2VgjmW7zphp799r4xw5H+rwbnDhGRC4S4
iYlfwDXZUUayNMSp07974bpc1iPhxMGTrfzQRexammbNodnSSyER7K93qtHh2P/o/0ujq1U+e5FH
xxPZE+AiadQi2RLY96jCuGyvQBHsdyluoJld02xI0GF38zsoXOmozSyOBhearICUt0xyb7XOJJjA
+ZdSLPpV665M1ez2dlcGi1BFK0unZb0JbJGKswnJeageXTvP+vIRNfBzt6C8+xQheqbzH8kxe1ei
kK/R4JKfCpNf8re9zrRc0dANCZ0mBbe8OVefLwH3ceiv+/7U49m1A1as/bBGmwf83uRDGCZ2dmqT
BGYIZIBcJvmplnwSuONhbTluyQLSttBHVkFO7tokRgJdmqTVYfWPkgien15NDVv1JDP6KRAVrAzX
f74vq6eK3KPFUfjdCZd6QNbg7pqDOCJZAbzAMm37fWIZbzXBQAaDmdbtdPzLnuy34yyG2X+jwiez
0i7OODnMVgZSQgnNJEWZ6cU3NyKaMGiXzctVnESRe+v8ar9X6CtYDB8MekCqaGgTFRCwjNpxmJkp
zG8kJ6Bm4JdYHSl/GDHIS/L0QV0+911VI4uAVjJgRlgS7dZFsvSVOKZVbjjyguvnb9sqsDp4RhOm
td8V8X08ilQEgisYb3ZPBwSgFLkdlMaBplng39fc4TsKj62YHX/iwuASEpfSrTdB2SeOmwdfEmQl
4kHCkXeHMcwLwFvB2THn9Y38LG2+v4O8H5n6k4oEgW8ztKljE8S8GBIZ5QXKgKcxhqXX+/fathQY
i9Fl+Rt/hgKkpmt37tLxrAbLgY2/364IlZrslhmckzU6IEks2i9wEpfvms7/bc8EZbFnXplSykS1
rF7z8KfdKRYZLHwA3jzLaehAbITK2LrpPdP5BgXJs31/jYg2U107z/y2JLiJAgjK+nbqR/vh86/A
OKFwzBBHzDv/EFntu3LqDAZCSB13kNPI7CdyT7CpkXd6+w0XHUWc1NDdQ3ghRyg3c3XgUDQG2vr+
Nltv9Yr3Iqdho0uU+C9EJBpvRx2h/IS/WtODuqaqQDWOJtDuoTKHmUnC+PNIHnXgrDWFotIK9iAa
67TKbQS3Ln82kI+s8IviHxWz/00M+57kSC11YVE0DUertqrWBuxLcwxcekhHcTW4TKeuI51t3fcd
1hqFasvSn3Jz3A04cVXxZi8dckbClZkMiQ/CCVu9WOxiXjgbJ10CQNdUinXwRhkgJWFLjjfgxg1D
S2qmQx0WST234cKc4jl1bK7xOV0j6eRDebFyKbmbCz0YiHiINps5Di5ZmojKt9vkIURRY92rPb1D
YFsWggQMgCIxu+7HiNEq9Rj7bCTR08ODAkSUTyp1HwINcnGfgMnxRCU/9zgmwpfPttM4eFaoHrRt
vUf7piVQdMTDqTb3fTWzFEtPzbiZ/LKFJcr/3fGue+nR2/Zvgi6FV9NFDRIFVxzj0y8WKhmLUPym
bU2VViuSs9co8L5P3BkgA+0voGsIeTls9RgF8MFUp9QVsrFekHFBi/MnAUX3XpZM7d9nkv1ztDYg
Iclcx1pp94F8ESoKNugWNclYX/nfoTrUfWBMawc09pT1n3q2ymPSxUmh8V8sr8QieJRmsqJucuJ2
PN6u3fHGZLSp5dNf5hTfzIRFIlc8ZllKauBpmWQHeQYHmoIZP8nUdG9voFyQMYYDhS4ICwJIZayj
bpFibnZNi+IeWMCaWi927xwv5VXFdCLsGiJZPsSOteHG415X1RS2ly+LZitCmh4/SdxC90R+jYZL
3mL2WvmE6ZS6QzNjMNL5opg38VXVVU20j9aMDOvSmVdCfUOkAEgZb7z1ooCR0kNko3Bfpts8LHIi
sSSt85w44TqGMmv6YHE9ZhvQ5W/sZVt5XcOYviIRjF7TDnI77POPOA/8V7dS3BZCZuhw3RDf7Rki
mSHQR3Ct0CBQ0TRKAbGevujJvDXyHH21E7KwQAqkR7o1W4G4GDCLx8e7VfpqL6lmEXhxogiUoT+c
beBNXTfgLInn+yLI5A+c+Vjnyv8r1tQBulqatwLKtE7gOB5Qpu/ddeXfrWxV9O0R1y926U5W1QRD
nF4E7TmMrvBTDkA+33LzJvsN6mbDppi+eFn/rYl42zFDXhhXYW3d8ZaLAGo2Y/fjyksyQ8MEMW7u
x2rBo/jBY+zFKGDK/dCoqHm6mugWJgbuxSnjQ3y6NUCeKjtnjUCYOmFpq8hKqqjjjgRsRgn797zh
mpWh221SMCv9IBu47xY4enOb/deee1wLhRODrBbEvMTLaP64jcDl5+z25aOKB7nWx4mSsRwkdbV1
ss2JzFzFLHzXyF2gy8D1H1onIbSqIIcb0nKHR9vBhECqMgBv3US0O3Wqtz1n+ColA/VazFm68yl1
4fm6svjMMoKrIj6erSXKtY6vvMuXszcrFcztetBPyR1e5RSm1LlfO4bvEZQcsw4tOtOwwyg8A6Jt
XFCTAqHD3LeOJt14PzM2csB9kgBKDX3+yPrkEnI0YH5B3kym3XtCrzizR2UEfc2uudJg3SCWP4Yp
TZTTwkRv9SPSAyBiaqt1qmKLcxUY7ufBX4udMMEbGZsxpcicZhDRneFwX3y4q8fL4Uehcea9hJTA
WWV7BFVUvVsVzdn6/IbnVu7HMOtXMuU9r17u3AaDrp87BdKumTnhovQe0v6VsQZqyuLBhdYdN5/2
nMl/mTYr1phkvtdOJn+vdu3QEqz0RJ1oMS3SVE4ukjXj89eBjyREtvM6Li5zeT3iFagIVTwkowG7
FZeQ3qvO2f9W9RCv+S/Hbo0i8UxMlfEQr0i4DUkbKabY162qTjf9GAXjTsTXuooOHTJCAnt2e5RT
g/lthbkod5ky25rQIHPxnvzMZ9K3MkpY9aj9Lw/QcvhCi8IklxyWp0Euif4ZyDwy/Mb36vm+/LTS
/XczsrJWo1FFS+IbRGUyWoTcHePpF0FAANumAPt+XVLslF0oOmWAvw7kCjsw7oz3TpRfqbP7dVYa
5yDjz40Vt2Jgwlc5cAqJnSK5ksQ5YoAsN6x2UFUhu1dK6ILeMaFBk4ZhjWpVcCNN8wvJp8bxw34j
o1pEDZjMg3s2+MzPyXWwSpXYmk6K9IGgN1e930RZ4ZRk1i7lhJ70gyMegPR5Y0sLGL3NChVw3/8B
Zcc7xt7T6Hqaz2JaiJOvS2P4lJK/y6DUh5aXlpkRtdx4zQrZWVAZ45kE4qZCXHiry01W6tfHY52S
r60x+/lVmdNjITZ/uXOBmymuW8qSdzZswy2Q4Jd86/FVh4AofArNzcP4MrJvedTa1+LPndcVk7n6
7zs/60thGGfRT2vTQglSAFCFP/ED6MKgRURRXIE7PJZTTcoW2tmW60NXZlpJVTGpjUgCQ6hM+XxY
UP5JdDkw6bx++H0z0cp5QF5UBvXOa3aILwr6KNbvKeQz7F5CO7nft+PpinlcrBQpLxP1JfH1VkwQ
ppWYLNpsEof+DW88IPnTpYTgzAhm7ryX/8CN1zTpmqK9v/2QdKZexrG7zs0L4e64lWPEKEtlPvn0
45Gnq7iASI9XY6mALTgIRUM0ECk9VRC0WBLZX+WdRB33Iu5MNMMmqrPGsAVH2DMcMjJaj67OAVyt
4H+vHiyRPOgj2dbfksZeMDXoLYsFYMIRzayOInvDl88m4ntP+Sl75jCZDlzSQuJ/Xr4oSewDde0E
Q4jv/gn73JNubOzCKfgT53ebLxh7QUqSqciA9CsbAj0FH68PFxXlsIRsXgj+1upV6N8jSeviA28E
qqzplTwLtHoLBa9+iY7DL0WOR92TYrbuKjDSnogW74GAcn4ecw62Sbl4MuZOEZqBUNfESqgIZ+a9
LOaotdx9CxoR/UNsotDX1fKcwWQ5P/INEHXpRKak/rsZGeFIvdKgZr9fA5kUdGCEBkFXMgyqUa9E
6DGa+N6cY62KMDgvdJfzWGRnIohXQXttlKCRX9oJvbLViv/7T+G6WjEIq2Fsds6ur34Hb2wx92Od
ruj5/WY5nPiOChSZ6CHd7QC4tHbc909srsxTurN7FDSTsK3S+8BtmuWJhsYHSjI01j6us4i8smfS
FUSPbg1IBvg3pXAfOojKIwh8GQ/dfw3WPdqh2CZ8/gh7McR0iiiuwacP/X0nYjWiG1JJvXX2BKD2
H2qm0ph73hf73TkfpJzxkZ7AMtRmmpvOuhRciNO4KovdMeDyLTY7QX0t50lpVfqrrP83ePyeSKw+
g+TNEceTLw+PT1Y9sUJehbGoMA5BWaVOFfGHplYCPOdVnHWxTo8TVF2LsiLczIZsRyGUCt/gXBtC
AhInflx+qoUy+HAkkX1szLuN2TQ6OTUY8gf9JTupcdOOPaiqpXcNpmIfqQVNLxg8r5fWHXrFSbWJ
eZZUthxtA+sB3Nc9kzqQ4/6sZgsSS3C3bzSjqSERsQY8GhFHOlcuoQoaW+cIPFOt01dzUSk/Qpcd
+b/szED2cLmeDWQ3w2O+uTdt+7GN+GcXn/XNj7ITDeGGPUFdtKMri4wnpt7DKUXO8PVZBXhfBGQ4
8CofvpQX/QLHXT0t6R8lgyKfR5ZYANeLYScZ4i6RZ00O4y4A+tbpQNAS1hOykxXoLISGhWan4Ztk
586ZQpsno/T+pxjP1hFmk114lRCg0TMBM9e66chsmH1C3rCEKk7WgXK5dfTRwD//XXIqpt84/ZV1
bcFX8c4YJsXLSG68qTh6J3raQ14WkyjVg1fq1k6rQybk3r3A9Y2/M3KHI0IzgMW0rVEvZIr59NCt
NF6lfNrTT3LZ9OeHM1igMSqt917RoHd+uJVytFhox4pmz4tsrZTPyGnLwc+2o2+KC1YTYyhkk7UK
FixBfLIqBvjEIa/cGNnAluclfZfHRPQHnTldFUrs40Q00DmLte/jKKmKZIa/Dmg85qnGhvoKcRCH
TMdEyGhkEeaBd2C601SD1jOmNHFYXc1TmQ4i5/p2Grk36zln82hjzVYmMOqmYL8dEf0jBDGzn1LL
8o+QmzLN2s5cPHB6PJv1R1aUT32ItwE/TzdpINPc64GIWez4Dqc8QinZz+Fs3pr4iVu+xxsIudl4
EwkwwRkjb5yxyARiOdaO0hQfe2D179ru5ZEyDImiraTLN7U2B2X80A6sI63O0DR67xTX1JDIQem5
Nk5unLLZmC+ad7xsN/sb4RqGYt5Hgm9oolIM9/CW9q9POSWZ9cXvkAvPFz8xeQpVMrdOBP182QxX
PG3hiYCO0x5lZ5iuIoJBvLOZ+O0z6hv9je+mCO/Z2gLvOSRtpglWDffd/8tVwWNAATmvaKdbRUzd
BpuEmpApflAz3ux3vpj/6pRCZ8Xo5TvgclCS1ITDk6doDRdFEWpsoMCL7j/lwkPnjzZBBpQEHOMK
sLQ88BvCygvNT0cyKp5MT/iNverMvEdL5kVYP6u23Qur6XiFIXgWjlwWeg7Ut3K1w8F4zRHNO6/H
w9gWjbXiDZYtsyw1gEm7IreYaC/krADZRYgPNW8dEyK1/tfzes+bBrUqyYnRfQ3YWLexGWJwfm4a
WUsAizJtCcdDFItyXzNya16ZUjO3quxBakHYA8i13XttRPYlEHevF/RQrDAEIz/2+tdg/ouEI5Sq
C1QkayH66eT9Vg+i+F6hjd3v0MByKvbWXz6JnmFBCZ2c55sfIa9Yv7X8qBustdMYjAbJRBKSsF9U
bLmA1YUXCk+uk046bFsq0jspMGCjfXGZTwo3WbzEFv8ulMc9yZinrBbkV7ilMNH9dY+eTD+JOZNB
ZmPDktbcBiK4zXa/zmWl8r72MrW0AJWn7Za5QAFktlSWTCg+CqGmN5SHv7OMk5vc5Rl5y8MQavU9
2btywE353e+eZcmYGZ1gW/1Zt0++1ffDerM7FoL7EjOqXRPhZKdqaQ3qRiqzPrVZR8gwxV4LWbsU
5X2FrIDOAwfzwGgOhGn2E1q2o482ssGkZwPV3VgF7zo6Cg1Z3pvYAOSFai0shfM0shKohbDOmizD
lEtJHAiCNPklIImylE6IdzhzO2VzLLGC7iYtR1j7YPOcFrcGkDeAl1ddQ+3yZJGlBCb0nNr6IzLU
LgZK6HPnovfp2aL/eGW0JPkis9IauHtck2ddUD/XeDpmEuPicwI0OfYKbjH8OnGFMJBtE2HNjloK
M9JrZghz0rIRbWIAgbyYNPtohMihcsNDUJ4QV6rEvpBOoZQZrNNfh89Tg+mJoYfkxXIMvKVE7Wmp
nBoOCZOfGJnn0weOV4et8oAZ4+iwmIyRXg4WJNqDQ3yuAY9Vhg1v3DgmlfEuxVeH78+EvN2xH+oc
MEF/sZ/jF0wdNCXrRp6hEftWCIC83/lDqRQR+gjKipsA/bEeNPE+2yU7G6Cbr8wEouirWn1GoyIE
WBgyflusNe1spogwNcJ8RjYgtopu/6+jMiFrGoEeSDnYakiboYYwVy0bo41qZEK94QewT7xH42pc
EUpn0Wraz/93fPbmUveT4azhIlH+Q+E4PIxEhU2u6pqfd2EVCCch7MV1TqynlSzO5YS7o6wa39Kl
O8dZwNPrMeG/BHCXIf+LweLkEnSfKQ8uzFR48Wr6qpvd8jy8xaD+PTWNzOZnkDf3H9UTTQg7EgjI
cj94pRqt5Bmf3uTUdYGpmV5XXsJ33tSz7t/g8W8LPuKBHbn9MRoPQfyH4hZMdsPrYggg2L2Z7Jy3
qcxHQMuGaXYP3FNiDuNxCof+iYVH7RyVExEO1ltujBAkGjg8OINKet45uUhgSMVRTCDUqK2O6gxQ
Pi6z0gDRBjp6Wbn5M5YlqSWm/j1xI1j64nm4yXxgYfiNQVtbfo0uwKyJZAtvgeeShPv2tPYRLEul
/LJQopxPGjqpQaGSiaktmzuXkzfVPU7jyIOHt7U6Us3mJTslM7+XnVamj480XosX/++lGZ8ix0PB
UCwE8n1AOeXQs2eAZFhJ5sE2slBaWM7tb/Iei8Tg3NIpRzm+vdgRg1Vg4elvLer/AVN9iJ4xWm9G
BKuJ7SU34IcVpUgwhVlXg2EvMjEIpZqPhdAu6bND89Njfaw29vEP4Y1cylKJkUBKM7wppeJLkZJh
NZyjrGfj6fiua11nWSp+tkEdYafO8ehpLy05mSCpY8ziDamSl/D5WD6fzxeMRJMubBTWS77pLcpA
gnIaU8mojxheVPDPqVBYvUoNbmUXIQWgWze0ntwnPQQ/iCFqTNkdyiZ8dteuf2gTshSl5N18QBzs
0hskffys45L3PlHQuOTG0ZGJlVxkNpQfQRfsGXNZwx9Pv3vP6Xgm0XxgMGZLOn8kmASppz190y2G
v1fK07B5nQZX0/8oGdsHYa3RWiyrnD1uvuaqw6jYKo9uBk2WofqDEiA5l9+BLRTbIsb8GeXQrw8b
twdfvT/qpE5W95u0eMzOp36DulUzSN4PVw2AcRCcJPQK1kYuO3AR4nO3frhzb79/JvwvULdHuilX
h5+6zIt1bhjf5XoWillklL5fvkx3xPyJk/Gj2DwCDE0SxQtRdmtNa+mrPCzEXH1wDXm0fgguSODC
ol69BBVXHYiwl9B/Oq7oFlJS2ZmqVlFvEh8plhVzzbdylT3NMoN3TvRyIQ/xB6Nb82ZPog1iPiQa
eSYsWVkLmAYEj04axxboIUN8OaK8w6LI1fc2fMZh74IAC0rJorflA8XH0yz9gC7jZ3O2fIs8dpXf
i9yzVTU7lVE5DeKnvLRU2m82Z5hTzkZwpGWEQgAJkNf1GNKFrlRmMtS/G35063c/2I2IrTQ05Q9z
IBGQegH0/FGK9aK4UpXlEhmRoLpkzObvvwlCHc2LSuhELKc/fSVIYSOBlzeNmJR4ftu6rVARoBBd
5UNJmfGXJRCeib7wN2mnjIsRLjxi9gZVVU7p3EwDaWKEqCG0MJAYrE+sm2UriXs6kCNtPCLGnyZB
0aM6elP6JUG5F3z3cqw2gOOjD+M2NS+LM+lJyYVbDp1i6q5wuiuz44ZOdLLR//L/4S9HdbHxDX+w
N0YmVJ0p/CXTaHmISTpXxq9585Xa3PtAB5kAO9Kkh88CZFrbhpnJ4q/YpJwHG159MlQ/b2pVhPpX
TeJh5WpEPI4gODwrUrUyGNIQYM/pwypPFyNJovaOGeXklfm2/MKGTV7n9pSyHkkdRgwAtYx4PK1l
ZFFJEpJ+JO8WRc4WpHJhlJ5vvvDeyoySTG+nK/2kJ/MoVIwg3f7Bst4F404t6sYh1b7yohUOett8
ESHZ46s5VQlUiUZVNXcmqfA9e5ArJK99Lc9ULGKRcDKlRGhXaHVzQ/58hbSFVGRjeh94fFLEgjA1
xFPEOi9R90LmJP047Ds3D/v8eOQ7nbKasrluBIRFWuAL6JWGEXQoL6a9l58ml1qhpeIda7FuWGKx
CKprOtFtMAw0nxC5KBmygGq5v+WrLg+S3w9xkHmn655QmTb7RXOyaecfvl0Imcbj1749LvXmJ9Ax
+VAqRGaA3bmvp6ovZ+TXCt/RIHKOzDypYL3aDWDj695Cwlq3dGPq7/ovYjRoT9K8B0C2DqT+bBN6
+Sv+UwqBrAD+8BNtpTsIn3flQDo3fxGPWhyO45KMG+kUzAjsXBhzWP4cCCu3gWQNNNZjDxGaQFQ0
JoNM/vOWd8eR4ToiEH9Fz28Tl/rLwPxVfBK5OgnZNk0QziVG4vahynUJ4FLjvnIMBDLlGGJt0ULO
TLbrPOiH+U+28L8uqnLVr70cz6dom06q4E/O4Vy7wITHAR69mrEXsNkN+IrR19DzWAEkArTPmgwJ
XWocM8faAObArw9gYK0B3CkmVzeQ0QuAJX0vD2cZOcGfd/CP+QWyBVvZEhv9lWDEy0a0p09vc2+5
GpR8qdqu9sTOo+/nJR7SDPifhsnggdEWRmjc+buR1+u+5ui7dAOMe6xTabpc6fGK3kPNVUy75ZMa
+IpVL/yT62c6tVQO1pRp9Dnzuej4fTiHfhg0fojJlwiwyJIXxGsBUXz7dqn/N5kqHfBKq23bXfc1
MqXb9W3NnUR3pD0xg6bcbOZq4SyCvZO3sPUoTBR803o4rOYm9oM+uLnGJxpiJFMdNZy/FxHCwsoy
87gd4mlPI+xkhOvM/O+CKtt/tUWnEN+/EDRHeKnYHqp052mG4GrIgPt+nhn4vXZPys3LHqEjV5zE
OlrNalRCyikczxflGxNXIZ+Wd9ht1S3K78fXgL5e8Vng+mI5LeMJWtUO/4gwmnnFF0r6LNvAGFV2
vMDry7OkVBkA/36yTsoRwThUH+1BN8UXOdPapPpZK0EYaGxUsITi6ywt48omE+/KQ4CIBOy7rmVO
8Jdu0+cDFs2gnnQLrvuRnimEnIYqfO8CdIcfUDzliI8ffaBVcpiadBCr/bM6UBSGEcJAILSavc+O
NLKZcPTFAXOz2WftEctwfJdDZ2ONoeWF7C3F6JkkxBHQtGPlNKZSaUP2a7wfLaotNvvxaL0QkjC2
5/+uCdZTRFCtwU0QNPpi8D7/gsVdH9VEEgtc7xDxNBekJkZ6DYLV080VqLd1p/GvbpWocUi8YKO/
qiwj8rBKiVzubjPrAbcUQ195Ahf7SUoMDz4ehCBVWZfnzJAN3q5pzBDIXHj1Geb0zJhepCzPTjgP
Igl94xUqY4obSmsn+mXHVwtYAerN2fTT/4hCeXPekLFDJqnNW/a3FgAitVkwnqKcmtXRoDnLf38h
RWdg6SvtVSVG0XhZ+Kaqa/2PnqexPybhhQajpd0AE3sOvjsCSLxSYPGSTQh3bFwcy2iNSCRq+FlR
N3bO0LuQXFrzJx3PfYWiEuFbvwu+1Tfp/4dBdsNkpDSKrGQ6a9NYR6sS+UehintY/JxrtTTGbGtl
TlI0Yq19Bj84LGgCRab2IdlXVwAwtmzEaNbGF/9unQVvBpXJsSj+BTvnOF7tEZrRnTcLLzz48sNX
VklaT4LzATUPP97XWL9ogLvFmRDT0ahY2cJvoQu3LFJrm5WozPTzXT1qfbtNyReySL7yFOFgB6gz
/BGhBmr8ErSwYLu4H+lFvO+6P+8vciiviqAu9ovGfq9Nh8iFVU/hV2sxHAHNnB2aqZR2gD4ShcM4
mZTJdQbmJhWedFGyA/JU+LdVEpPJYp45UlJ2himP1WcjSBJEwgJmycJKkW3G11vwGFzvbuD8IcYk
wUZtnWesa5gDJw5Hl5+QKdj5Qto9mLKXNOyzuSxfPbFUMnpgU+jyc90O3K7eeCcRlCMNvHMmbqiD
xHfl7cjFzfpX0D6CON4q+X7CsXVWI32gIC7dPv/Wglw5m2ghDw0xfiHmtlt7aefudPvqqBwkCiKs
THz69TIQConJT6wBGMR1LzMMhu8ImLnA0dsjULk8AR8pim+uN9ZpGxYJAlsVgUfejS6T8vLUXJLX
JAJb6QPtltwdukxB+N6C68X7tVnTrMnCdlyzb/jzSl23fAM75XUuJy9dPYo5csA+sU10vvxdqZdg
ITuRerwngvmnUsdXffnn+1bfuzAbxiczgSZfr8GJ7TkLew3n3PWgCYKkBOL18lOTV2N9DDIISE95
FKAtbDDTC8/MWb4TsIFNRWdaTdQQJVtR4ZmFUa2LFnbr7Uai22R0vFGRrF+taIcoRkuaRVRJLn7T
6QrCdV8btVm6L5SiMGN0JdD0V7JkxQoLkphrqnnJ+A5XiyzunNGAHqzjr6By+bQ32huzWwxpy7xo
lsNlvUCLjuYfF9jRqrFDgQ0CdaTqDGt41aEfJG5z2Mub5pPXB1KiaFqa1TVa2iQXTIHuO1/1fqzE
MqPRXCzm4Ap8Vbyx9xp/dH7N8kbvCKZll+8UHpEKxOGg50PpuXXfqhALilRTsjWpngSJfoLgb7Qo
wkwHXAjg+CjrrCzXemg4RvMZY9BKq3XzSSCLCENeY2yrEN7IwFk6wa3gzss9QGm9VEX8UJGQ82c4
Bp3RNl7CSL1Dqg2yy0j9FNvONlEcwY6H+7aCF8GXI/8wp0BkRAbwmVFZB7HZitvO0dcj/K3SVhIz
0k/z3Gir4t8nDR8oQVsr1N0koLwnU8/22ABQI6ulgbg4NeM08BGqMyl6WxGjWduBRrT6b15yVz4b
jMEhW79qF2Nb1S+J5I4AOE4mlat3ACsTl1sCqeWSdNwhRe6yyxBVHbyf6AU0zJJROGGxv91Kyuxr
c6cPdrGrkvm+V1CkNoYq6laRU7R6zDgoDz3zSpIxpP2PmVzFxJ2pcyFJ5YX6N+9TUFSQNlGueo0j
fmEai2vHThJdr4d++vp17LEJwRmCnNNfSKi2a2jJ0WAcUtiwDhG4ELCztC72DWN1pccCah7Ja8FZ
9cBDTdDR8t12lMXcCtNDnPACYUuHDem1Lh2I8Zz4hIl2LA7svS5kRzQWVrhvnDSSNQMDwVYg+v2p
0Yi8rPJ8H0ORanxBALttfuPv/NEP6V3o+ytxP/k9uPZdogmUjo9YyNadqNtEmGElAghvYDrkFPE0
I1UER4Vp1EMbh8qyfWLwMkeKR4XRHeq1Nn4LGTHW/YeZqidVBWXbQiQjZ3Hf3GKAZ4nJ3Y7lsYyO
1JSZUKhBFnS7m436nQrqFHuxLFS3SxQCGMD3+CKM9QVBllh/AL2QqCom0TQaNlf8aSSuUwsFsyIb
1SEn6lAjTNq/tkbPRLYGDKUIlXQCo2J0lI8gPvVMo4Ebq5f1Y4wVjOr9a8Cyhrm+tX1uRAMzMVaW
L8yxpuO8ZEJKd+R1HpambHgxYKPB0yQTmJaZitU03+4TgT1g1wMmeSlWCP87/E7pTOXLvxqdXJtR
amQqxNI2suyYTzWVUPlQFKgqECnliD83oYjGTWR0oRQIPZ1IHXbr+8o8fD4FPJNgpjFr3p99C/46
75n9NXHM3GX2K6R96Dp9B/9BUT5Nlh2ZB4W+aQJgmWPvNs1y1gsAGN82fUtm4xMCJiusaqu3ccrv
2CI35RSqVcYrDT8CIE1Em38WlY9siZvwaru8Gq1zRF0mIZua9M9oye4TMGOmokpA/G8X+hWV1bR2
0TB9rY4VEt+mknzCYh27Y1B6JNrcQeigtuSa6wZ5cWqx0El605v1fEWWFQTrBnt0Vg9YOP12Tmdu
ZdZCsiCjFo7qk2JhC3Kkjh52k5BEp3QcNZ7EP9pPZKVlzuCa7s1X7u7AJzF1o+HOGLzrlHRVgPQ0
7bxgcCtOIq6oEd1XyK/BgnflWIrNM9zdqxO2+x+Sz2IFNtfC5MguqSDj+zbq83npAMEvPfZcTu5U
aZJHrcqCw/fMWeS6HSJbhHC7sCYeoOK7IlELEF3gop0pvgPjUvre3SXaQO2ZL1u7BzdTbDeVOY4Y
wwyTBIMVpgFJwGhWX/FoQyOtp83OobMhlhfvb++yNgoPyIvAEyv3FUHE8adFVwxaYFHTiyPongGp
41CDl8CyuB3g4lEPfDewklCkaKefSX67TyZFQ4yl2/D1pP+4hu5z2882zSfTc+T2z5meQag9XSX6
/y3iNYN9r9VDhZOdrIdDYLQSBTFSHWWIZE4Vyoz147vCUFTJaE+XwTQdZrIHMpoW5aGZPvL36gha
sJh/mk5tV6baFTM2eOKMBpic9ol/9t7gyXEdlccPCCR4gEgVCLD4kMX4LL8PQOaxweXrAJQLCqLL
f4R9V1SR8OsqUNAp6qWVVXmUwmbVJoAZIfwJF5rmYXNRCiizy+DALIxCc4F8JUMWj5XjpYekkWiq
EehlfbKMznDytdgW097KQ6dQWqN3EKzQdC/HS3bvGQNYy+e48HPQJdY+H8yKPL6Ai8UJVz0bJ1Jw
yHhlt8D7pE6W0KOG19ChxheQHGAdWoQwPeErSnM6Yf0jaEtL8FVpw9NpOY333J86PwJmBYKMdk42
SbZN7WngckX3aO0hC2Dtbbj5JkLoGnx5Enc6ko53m/HDTAje3WNegS/cFOOY46E9vLVrCpuYTIES
hcIV1BoppBJh4Y66efifF/LBU+xGTkU5U3xQfNmOu/2FEvryKk8TcrS4NQQSMyFhUw+2mGOcndAm
Ay5/JtNj99HgcaLM3Ag/My13ORYQF+8Y3jOqyA0uar5jxb4Uaqu66NFr8OKDlxW1Z2jM1heVltFg
rzZy8Vitb+QXqtDS2isc/SPv5kxDccQ/4DypfiEy5DwbEDuIKJSxxw+A6HhG9k5pnQuZDAEvNgg8
rgM4inou5/g0AsFwuAsaGObxYiBxTXjek6wpqd7FmNK31DHx8Y/gLbgBIkABiBGnt2flIAWapDQ2
7LBiQUKCp51KIklgBYVbtNKHt2L2GT3PKezGZ7vPfJXz/epGXpZvKmFbkZsC3641OZMCjBuG2Tpg
42oZ/VLYKmrsnEWj8jo8uLy0sRG6i+GpHLMhDjsHSKcye1n1MHw6NfXGms1ExO0Zvn0TWIrW2k+E
V/cgh4+Nwv2UJEBsVh8i1GCzegbqogWAy1eG2ZA0EwLR+L554fQCh+Yj0KXLlQwrN6OQJqrPBKQ4
LtRPif2QqixmISt6E0T5LtWAaJn07c4edxG8mFod9vXAa6rVifzSILDywhnuelHQh7L7yA49pb+V
WedcENmRjcCd28wFuBb28Hj/9XyU4LtaVLXIyN9RafukmYAnCdlWj1FamTZKsJDsvgazSVPMvymS
+imsmKib0k5ZbkySM/XR5O+3KKhF525nNvzOJ8mBkTjd0cVES6PfeejYcS3So9GJ1RuUlotuMul1
OZDOFzi+B+P3s3IvLZEff1noaEWPoyP6/kCIhPKvrwJWnL0Thl4/VkUAxoGZuQQgGANjmAR86xm2
xa1aPkg8ab0TZ5gcfVS345DkJUnDVxEn9qiLN2BycmVVK4TMon4mNX3LZiryhBfEsKK/LUeXVDOs
uSgko1FQo/3yWWwEDrgtvpl293eeAqxAFcaEOe9lYxa36DmIkjDRQQpZVcN8csgnhQ4YNWh4wtHP
JwFFLOxa1KR1/UMMSuF/cUSUuND5XZnTHH4jcEbZYH9vFQzdSKtqw3EmZX/KBvMwiVHEAwCM4hPJ
ONlikoE/j233ENlUtc3ootW2q9s+U+was7TNjKcLsRNtVq11GdNS7xY6iSszS8kLhFVju1brpmkH
PL0EMOn4msI5Rvw6l1juTBdpv0jbhtIJYojq4dzXENmH4XNMZwPjUpYsD+S4sMeagoNkY56cwOJb
CC1mQnkMTgmRMmzAW/HR1VuUxmA+GmKlP8PfeZpu2LugGLs6Ob2sbQ7oVlFqbftslLMJIWkZCXT+
gx1qc1om50T6kRqekFVyWpzPCCofhzHlt3qKyY09NcxQQT/RdCIyUFREA6HrEOj1MST5sFKotwQO
hFAUkyHf3jb0T+WH/KzR+HDWQDb2jsByWTAkHtDBVuBCxpZn+VtT1Hs3g7CIpy8Jr7psGV4LCIgT
HHbh7FMg9TsQDm0SfdaqoZSjCmPghLh8pHuVJNzKYHkxR0+3Yi5s7Q2XKSAmwVppzjCgflyeDSp5
Q8B2Qrg4p4idIj2Wa8Y5RPF+Jfwdb3zDxjVF7sDftOUNYHVNm/O5BGcjMycQ7jHfHmQRf7NzuWAy
fn6+pN5GLibOwDrbNTHxDaVYyzVhBAa+WXpzG9tUd1GooBsPTv8pLxUsIPm95XLdYmaIoMgPoqgX
hFN6ApgdJrYdKWVvSB0BqfLailjs1pezecXfsYEn+VLK8zZ6Nx68KWzrL0Hd5uw14KEGWBjEeseQ
YstOonwiiv2w5+p4QeUHhFXQ3ZWopRwez3kvxYydpiDroFSbtXhrZ0IkZ1aSMMXmL2stAkc9kjmm
SeWxjjaAabG3D8ge9D5BCr9KM+8jkuQ1EFb+h7pxpUHR1TKludz+36bVkSXc6wsZMrE5IABSJDse
/KkgCJgqSQQTf9wGzlYl+R4PBO++UZAW7x8O9+CPOD7ZQAZESo3+w4GHuVrWJvev0KkRGnJvMR5K
54y/VosRw/6UWe4U5xKBwzzjI51VVBby2LTPg6suFH6pKs+1Hrpsh/tnF7cZSfTFdqIvkdExfuPz
zeNdoUHYuIdBpAIIqni3B8N5LqeW4uASePJ+Ly6AeeRJQu/Sb5Oja3UBxJA+x8jdM5P+A10PUVei
BFY+XkOkZA5Rwi5gQCr3x2dFNKoyMkeGb4F2/hDat88vZrET9YsguGcxXR3i7Y+/iIqLHGWzuggE
yZp+JRsKbkf1p95ViK1gl6Bx3AivVWiiXO2F4atq9SDrhcaVXoM/nYkv22B/ltZ5I02IFtbULFFa
qpGHpUExYeAfcOk6VHnzbnrA8Jujr1/IdIg04Z7PCUBJ03pyeNvIijnfPTEojNWFcVtE28dmPW1J
vPromvXwuLIvuImXfGWO5Mf6/6EoU7ELgXp++nYM/ySJ9w+gW+KGX6YHFutpFH8guBMHN8LWXVSp
L5E82h4Zw74vruOSj676/trz8ikDR4bOGGsbYgKYPX4wziyZFdz2wed7DsL40WUcjyDo0T0PKAv5
RJgg4eDWKq1M9S7civ8V+mn8yJdtv/2Ei6bhrAicOP8OiBan21KXGPp+aX2IU56qxRsALYE7A9jx
ejW7pNzVgcQLchhxAlNehT9JOtSnQ8M00p3L34uMyi3NxguDW3EEfxK9SsKD7i/OHGTYzTs0PzL3
iT3cF0IFmrh6T+QoNzRF7EGkz3jSXibXbIfns6VRD9D+463V38emqKHD/s/+okWzucDDyuzkD6UG
QT4q2r7TErSSR/5Pc5c/3K76ddZWI37Evll64d/0acy/lAQ+AA8uMN8K3SgHR4KdEvFr9kU9ydNE
LReI7t/+8GMt57tKa4LXAg1H6nU11yAeuxfT3/en3MJ+G9naRv7nWHsR5zp06TcL/wtlw9+iEF2h
701RoA8zsgz+B/JqCGvEviXtdnGCdl6uUnj/rz2xGiB4EJ+ODnIeuQnStRE+GDBbLFfZex09mCp+
D8WFuIRu76xVbM/MBPtszYiUIh+QRKtcbepzytXV6xQ715JwVyWPsA4H0joEsBdRiVK1VDV5L1V7
AwCv8L2OKscGPSdDp3iXHFAYF0Te3BFAVHVxOkHaqGZ8mea3rrHFdLd9qlELedHMAviCgu9osrqe
Xz8lt4TDNhx/fFcoHxU0QJ1D+tdtAAvaStJhhi74i1pj0wAm7Ws44g4yelOiahEsm6nc1jxjngHL
vikrtbJmqrgXpQ/oZMq2DppKi0rtK6jJyEnf23Pj8rcRp0A50UxDPTHhPqlEIaF+onTLuVqXonZR
xNCIxibr2TsxCNAiEd9zkfo6dNOETKGg9teuNcT9T2ZD++Xry7rrKAbQ8RB4HXeOraa/tJmTvB4R
EJTSoKbgxQUjkvBkSbO0FRm8SSCD82fcKABIwajyJ5WqlCFhx0YwJl4AiQkmJiQNvYCFs2RgOERi
8dL6txttSS9Xlt/gOSw8+YOBeZfFwHypeSuF5lsbyAAktNQ9fXmXpjZD2HgWXVVegbgbjBLRsZqm
9tfRWNYbs4iRsWu5EiJRW4DeOdvBnHyc2bAAd9XpJxwQL5vHKW1rlhHXnoMwJKICi9zh/c5DD1RQ
GQq0dzsVvX3/HKLSCLrrJWSk4aisAUNKUtQsp/n+MxSOm+4umh7LBd1CXsBCMlsy3xRaFbxomGqY
6MU+fHzPNfVHfPHvYRO1GfR9SabfK+RFqoPjmd46kHJYUN+njhEENUEKuTX77jPGBOCcHjhuWXfs
4Y8hkgG+Ef9UwwD8ughZ1eVO4wi675hfHfY7yt2na4plGAWiglUE+LGl8n7MU8uHv+qGPuJ6cTHJ
y+bHNoupKtXxZftFpS/Km4cNvBVCXOFbKyxf6wlDTU1oMNyQCnVW7nlN9cXBLy/bqQ7gJLimvuxz
qOphg5FvU489Xh9dkJbl47735aU8MkRwgBA/6lYiK0jtXn9tXD0GDSEWa7onZvGXTj6fO4ymY43I
Y9ifBOgpvkFEk/pu94MIDOLMqEjpgfN6ngUW7GXEEgymwvnWm6QcSVCIwohSXiukuGePvhZMuAQx
V1eA+G0JQIp/2ouGFIYnB/9m/Yjb3D/TpQh6ow7jZ00ALLTj0+o/q9Bgi/nJpTlr45IIM/n6Qsmx
wTLWHtNn4ciXXoxBBGwE3lb5Vd8wZqWtGP9RG66D05Uv0E05v6l2TWB6QArHqsFtRN3gNmmTbsky
vKxLh2N3sltyAlLBolD9uLibY0dh7gH4uRpsvgaQaPntbx6eBAQzVkGYfo6TssckOMlgO3fa5RAR
ggxNJMRcvB14EtLZE4pfCfcpfUWEXoBc58eDdjyCITnwlIMRa17ujDy1ScNPef2nZ0k+IRT1Iibf
cInssZYLFZubKb2BbjqhNQdufZ5gPRaB0ICun1XJ3STcjcCi1e4U119Y8m8qvyUTGZXr/IVjkw5G
I1rGaxGJ5qdjuM4cMPVSnFwKqSMN1CfLYX1a/PnH6GgGH+iKRejrX5gxPxwRUIvF2zoK5wz3B532
lIln8coCqlFOsBzY92HHwBn8orZRJBQIaJ0Y5jpNOrmArWQgpWgtaIXmaITzieM5K+kMHBl2o/HG
wxJcPoAvU5EjziUiRjqOFu/05M8nJ0Tn1IVi0LexsxxMIoETuxZH0+QuvZq9FXJxjYKcpM3UQ5hv
klBFaQuzhjIpcaS04KVrxQ8E6bowI1yOcERF9EY3W39w7B/IsPUq9kGJApzzihsDqdalcqkGaxRp
/alZFKd1tZzkOPRtTSvuRgi6zB+SF8zvVjuqvXtMembvKjzvHEp7T7cw7sBBRIByHRDJ9uPN0Fln
blXqngCoZ//3U/K6LzFXIYOAptZxdP1rFX80fBzf12LVo6HZdDjZoG3R6Zmc56d+aMsoHcIHerKc
7F8pmtYorsQjhZs9V8S0x05NGCrD4lJNpF9b64m/Vdqs0CoAF7jF8nYSMlQ4JjYN8cNHmweLnQqO
ZTLM4gWy3eDGFihg5inlBJWONWIbQijcYermTQvvKoTguoAgrqUISq46azUW9CiLqEHNKnJUxByY
GY1sIZuiQMbrJhkhPXojijJ+fVRC1Y8nJ0Dve5aNHUDVbEkSwt072cT+0Ba9pTB2Wb649A3NgDbi
9Y1Ldk3so9/Jr/PMHSZ70AdI3iKBjFW0er1F3I6nJITRFUDzZD5f2V/Bcfw1+CYt8JP4q4fKrUIo
NlcyIYNYeIUBb0vKrwTKkTIoF5T4MPOTFL0hY7rc7dm8p24kctkSHmiIFkTzMB1q4un7qj93BWBy
Y+ERPEaO+qNWjCfRvgaV0SmQqkl4OrJO3pAqBaJ6hD1epjTJmSZWvNNEnCdbaWCnjIMJC0hnhKSw
DYx3hwjHLfDr/zDze+CTxIebfYPXBud1Bb4AOYkkgtBE61E0H9LAjQ06gVbLFqHYyvczDVd5du37
RVApnitv2f8UUXE2rR0YEyg3vsrZTUotty3zX6VGuoMELc/L0fA1o8glqTB16OKlaYuOjdu7A5G+
CAooks0Y4fl0mKu9xopfkt/dgSMSAmpw6putXEES4woy/GnV1VSaZngc3LnrAkQminQk1khsrg3K
uCIYWKdfLHewXeytqZQ0njFlYmnoA1w/KCtJhDk1QKt+FaYcBrKj3ojYbE/1zlFNxMI+/IuYZ8FP
JE12W2F0RpRAeaiuVC3+bxjVpe/clGoRPV7IQT4y4bdJyPlBUjJuJeyUANqGtkcbkk4Y8Es5idiy
j/mq5sgI+wsL3O2aE17IBNAP2kBmXkp0TMMOGXK0Qa2gyGS05NRnjZyGK2bSgYSyi8Gy+veLDfJl
4qsOa61t6Eq2XA0fOnZUkfVIUDVY9BKb8o8CqBl17t56ppMVyeDP3LTPtH53c0/uo4pNbnSg77xa
RQtz3v0rQT2aj8bm7RlExaEFnSLou7znfwvQCS7HP4ONMnYqMF1xLP/Fmj5oJzFE0ll0i5ju3aN4
B4drMzJ8w/TAYlNQybmc8wlYVztBSRQcz9pNi4DkG2TrNK+sRUeC7NAnE8hC54FCMh9KIZdbmPi6
5L/eQgRS6SQnFsjUB2q6uBHbPlqY/u2rxe9VgS0YfbQziaz7B4fdqlmv5CdVH+d8jyTfdLNEYPVT
yxD0EWqxn/+haa8z5GgGd2llG2oKuNCpDz81xmNqf+JfrNkYeBoZXngW2xUyDcJAK9wXDD0eJwfZ
NUxPnNkuu6s/LY6GCT2px4mwO1PEb9/lIE27mlIi0vL0TCihuaJ0ZBD+/D1QJFrfE3f8vyl3TGQu
Ny/2lLi/CKl5M/7T/Oqir5JP/dVAWG7YVX7EA4zhV7lsYRcwOjZ5LwhGl5K4jIyPlwWX6f4RNd99
3aXNdlU0pj8B64UYtHZpGdIG+RTUeJu5rfWCe+LcPQ+AHzSUxz3eKW7HEVPQmiFWn0eMypoPMC3h
wp1DJQML6BZ22KUoshJxKqVBpwHmSIeUd+F8qeYGTe2j1sF9Ih/AOYCxkRKiL9CotpKpKmGeJkbn
oHQyubZ61lmYrr2mjkjStFFLm7y3B3qh7VROaRKUihfQbYJL9iWj4pJeWOMibhYs7uha5361qqmI
ZXJ+0Ntz78jd+gvtebrwz9IKcEmdT9Yd480WyskMiZ7k2S+AnEAlNbxh6kvgm5NjD03nk+TEyjkF
3cdBCbZ61zqJgxM/NIXO2/SJp5TcSEC6AIH30iEpeeMgM4JHcyRfQ/A2IEWOPzOoCnE/Z++REzul
5UqfIZwwqv3+VZnXzpewgw4pvlv8v+HxWrmeUOI5V7aqnpptUUALP74hVHymaCEeNsHGovpE8ifI
MFrYsTq3QOqBh7HuWfycbybcb8qQiBs4UrVlES7o5b2wHsJLZgaGWhlJjiUdFtblVOKUJwOBwJqb
KUhs4DVC7bGjON6LOXLbm6APEhrxlmQK5oHrT6geT5xyxYhUqA2Q/sfEGmmE2FGmiBx8DK0NOfVF
nef6Uule3jAXuNkEqqXrowOOVbmYVt8BWbcbh260rQYVEl2V3Welv+c5TEUoRGFr25Qm2ptYjRlP
6JnCwXcY/ePx7QCnz/omNJbt+4MADrjW0JnCOfEcBjnYUnhGKT5wFZSRFiHfIuX7DuFdiSeG0Nax
X4fcPa2hr6U2yGke0QWXKAxSLCoME034vTd3ArIIgz/X5rGuwkLW6v8wxKC5K5IpZO1gdsFOfEmz
uNd1p07bwA1AyTDz5Ly/lWWCwTMJ033t1nQlx4kRNP+zF+cF1X59ojtFdslkiRV4Arz9GpB243o1
g6HAFSxRsdCpqZeqCUokRv/zJYka4NC5nkeolhimX2FfQSYLaQ6KwdfdkZriiSFMLjjjWweRxkHX
refLZNO4cIhbPMFuw2SwtbHgbpyWqbzYgQ2TFGFsVsRHccbkMzSOX+UyQ4D8opkHvDQdwbdrwJn+
Q1vqrtPqoO2FEcDCs0tK+mQiWO268sfKCpAnQoeR/VoTLjTqhMXA/C3rMp9KVA1jEgilwypdi3sH
WZxGiFZi06ls26ZP3WDfuMVokSj7t7H6g9h9bmS1N6wzxAP14IG7XwJTMKIkMvcqxjLZaqySTB9x
qLQFFZ+AWZ5ITJ1meYsejGqdpZV853MNS5N3na1X/T15GC5EUkHYkcIhAjFu+H1Kqtf2Ea7qeheq
DHGtH69V5yx81cvt7ffX2KU6xqKSsIYjy6NDqlLj/CvZsHt2WeWRs1LGIAFRTSBRQj4xi9T67E2L
/RxlruWYHzv7+wxNkAhgrXUqJRQeAczsIrmxUPFB3mk0SEQY+lAIata9U8ZzlvnpEDBn53cMP4GO
j4Gpn5JGs8HhMFWsmq5neMJH9cGz00stK8VeFz4teHVlR8hNjcN3+P80EWaOFufT9oOgRqSYeyij
QuobSnvX2ukjY6oRk6hWoACIG90bFXGPNIqgDscA6X/29KDrlAZgS6Trs1g5Wj1aX5DzjsnjKORE
LTC8PTWQiBreqMgFFeuw/s2akLgkpLvrjqYBWnAoIXTO2HNjkRnCOG2Vm7Ug5PzXg6O1I2m3Hi58
4FDeof31EPgJ/+ntkVX8YZPAzybFc+PZjqNhIHO/ArxZHA5togQoR8WThfNBJ8vtKJctPZQisQm5
srR/SpiEGHri1bh5N2EhVMoRFutJybEDHlOhu+yexDjgBZSDMDlJNn/x1soqaaBUnSfuxa8WDWg/
1cUxrxbz2po5yzAlQtCGYtrgQ7KyvXcj1O0WKNGEU+PvCnrjbtVVpenvmGnmmcXgdDP0/eSfOi/O
QLVNLp1NK8K8PYEKCIvniYdDTthiAlpO4WBpTXeh5z5tVmoujpYYG3VQdgaQhHi/WCqclYT01byS
PZAA9Fs5kyOTsDNwPi297mGI6PcnSGO8ofCakJtGzRKAlxuqVBY6h/2lMMAIPY1QrKVr9D5vbF6Y
ZL0TRFhxgNHsYhFLQO4UP8i9y+tH74NR/LJym26UFWPDcs5hZ6mQk0ji/B2mQL3FZXKZlKEtXBiS
FXX/11hR4mcq8/PzT+OmQXb431y4aeG/IpSu8W93t6LoDA+MT5c0nqAIBNC56UvF40nXYNng6gP+
NMyqJiMY7HBPs37G9PHsg9+p3KMI/Hq8Ildnfr2Sg45DjcGB1NgtKjrXI7eI2qX6Ml+nalXdhobE
2QhQM1fhztZBYU108Q1lzlLREQ9D/OXR2hZTyp1BoA4PDbii4DdwGL6rUdsDXkN5HNE3uJbVc/1k
FStk1ImGiyUN6ucSGaxjh4gzNJAkNoxt/Wz4L7a+UagD4b/C6cUm+4Y3fIBZIh6Bn7sYLUV5LEVg
0LsLXUrU9Daiimako3/xziU/nDuGv5TZd3pVgSaOMYiqYLesNSdJf25pll5xRUIR7oyDl2Bk4cWC
lOOsttgUHvrzyftCjoygA1itNquSR/cz5dIEeuX2GsPJTH2MmIG5zf5XfkhE/rMVNndodPoC/2Rf
fwv9XyorV4fFmtmb+fIDUvHK+z9CiC1zzFsIkZG7yJixKEPeOB4w9fOkdHh+2bq+lzZClC9Ri1K2
R/TL6YDh27VEEOU6sfBxS0ijlJuSqHLMWB+Ej9Hvv3fYzJEzWJzq5GJeXJZqCiddzZH2Et3nnhq0
kqho1tVe5FW3crcgpINAgH+v7XYQql0+f+CxXEQnHNNwYOrxz4UBSIHSJSSVss/cCvk2SA+JjKXy
JCAHsrV1GI3YK9dHDyA93uQUSUhPQOG+V/hlARuILb/rzQuSiTlKUHwztmF5FgMt6l+BZaxd/z+h
fBEAm/e5bua2tnDM1ZSBg2Bevh+3Nbds+ZuuqxGi5eIErgxmoprLSVEw40IVzcK84D/Lp3Y+tXtf
agW8qIcZM2KGFJclkAoMJaGOxQg8a57wFHUSpZSuEpAKEQED5lv4B73xNk2tdsL7bShtZQymUHyp
9M7ArMUtKy+t77FgKI96JGw71zBG0nRkY8oPJKEXm9MT578/S1PXbggwBA7BYG3/up7ngTEvJHE3
YrsgdlPaVRD8unr4SONcpsoYaVwv92TsprRRYd1o9ckIa+8Tu3bNfsoGPl9Vv8RfxSFPlgZupcQw
WiNOKETmad2lMXSqbqQfAPC1WIkmGro+0dv/5ypldS1gvOU267mRlnx/DI4cubyibv58ja95ee6c
MUcwG620gWni9DIIjuuTBS7QeTmwnosYqzGV+ATvuwPugwQGWaab1d45bc7q6tVx+XKO4pbBCeGa
2W/3EXSZJYIzcpSNEBxfeT5+g2WMYvlXPVEY8BBOTXjfIFIndp5hqRGaVUR2XlC2zRIw6aTfX/LM
tRbFJPJ5Aofm7BcR4GZjAJvWCcX1cvQ6JY189Q1PpjeSQhdL09TsQMF1nTjZ+c+vzPXMQgHplVTR
SY7UGFuEBgdeMKkiTJttDpAEsGMwYHj7l3/86aa/8n281exXm/8NO0VnMs/Iury03c5o2YHmFpno
XZu1tiqLwX6LBeovCifG7y4sOArrBBXbfCg/dqWJAipVJfkwFRWW+XMdHo9CU+9oLSAd6vyy6TYx
1kwfjwigEOHQsKl+qas3T10QaY7CrYbf4S27TqcRKAX0E9iJIS+d7My4aE3cugvLoBBbdN6UDySp
tGOjfswvjuumAz9cJUDA6DlSSh0bU9QhRSsTrmCxh+jhEoxuzDmF66klRETTuEt3mDVP268/y5wn
EWhefmsP1rc3onhKI6j4YRbyGlljmt5JNZ8UPWOq8U90VVj1nR4KJUKkkXDHr/IqsGwxYgexcisb
I6yLukRkoghaeJZJtEKaNf3Kb7GTNykQQAzpMozbJzPp+/6YH8srerBoa9Wr8T+DZ9y8CZxkSnEN
KSY3EJIrzKUvqeWtxZ4UVOaPkq1cMPIPoR9o2Fj0ey3uD/KfsQW2rcQMmVxM0Bcl5Q2GtwJgE5Zz
83qT1hZj+pdv1JjqN2rvUnPdYhmDw+wRMx/EJkaCDG0rdhEpsSjJkYYLDEHCaa+kJFMudrXLx/T/
wf8O3mzZbwwJN0QfhMYdpyr1XsmYWmrGdhMa+QfciUoVcqWubtWmq4VQbA7L+HknCBbyjHG5DlSu
0aDjUdRJSpN97+j/sQchWE/nguAZW5RmPTPTgrGYE0RKCj7qXQKtZSY0FHcXlHdj2jqLnJNcmg/k
bfpLGiCjRzGW/2uCrNS1OiQ8QZYmhBoWhh4vL5Wac3Dd/1tdESNckKKZphhvKZ02EX9NdTN1crU/
3Qv38dIF+xgVsnXDaEo+CHRGX8nXWvmk9nBxTEtl5d2JfxeUusS2TJ5UzrS5Hmw4o73g1GtIWeO1
5yPYXfC6UvTJbdxcp2OF+uwMCZfHYsduYOWkIiSWiaiNBMLXNhgPJrWVE2BjxxuAC6wnXnid6igO
4KPHpeP2Swv2WoJnSCM59Zw4Z7450tyDrfPtrcSxPeSLNqhcDG4drlQhdz6fPE77Do11UmY90J1z
yI3Ugh6X8/mo8yvqemUHnJHk3WFz+6uKzDBKDGbGgfouOJdoAtPuKvbGK2j9PR597187D8VUyZ1+
pAluLnFiMkV2ZGZvUZevu4F6NI0ns24ATFhsSQVS/wM9senoPlZW9DEbPgC2kI8muX37cR+hr/zh
cyzA01rqsd3oXdVsBX3RWPteQlGi/qYahrTJGT/5vTp8W/P17zLR8V6olL+kbKyG6u9c7ZmsI/bz
al7RyR2FN3ldE2OJ+HUBSIcZ5DIV+uBb1iTPPQVQC2jhCqTs7MeD+MaWryzcX9wKxYVs8iWpzCwk
XGG3/Gz94kMwfDq/T6ui4bvzBiEZURo2wfcgtRzwFS2ngXyfOrq2t91QcU1hIKzItu3iKUw2qF3L
SshbH2QL/tH4Mm5pnf0YGxiWBj1A2tz+P7S1UkLErsWEOqDS9bwcu1UW6AB8C+1YdOKAFropxh6I
mdWimwAQi2sjUc+zyo9IpqSYuS4ygXKcO4dpCcR1W5KLJXaWZLlHOiaGy35w6kjgzKVPUemt8AJT
x2iF/fJtD6lF3pyPvR3nfuKKZPy1+eyEJiD/97TfVhuf7QnB9el+Z4ff32m81W715Qhu75K1onEb
CadEsyv1bU2O63iFxsfE9I1+HPkZ/4JGNphO/FIzMJwjmDHaN+3scutm/KPryakFNybHIA99vU9Z
/t0cGAPMKd0+N8vW//w31q+0iiuuWJuXH/dPxWdWzsxnPf0yDbcBGKPzmzLcbZ7mVhbl/xOL1nqu
h2X2Syh6niaJD59mgGLBZXfEvG8+0PyMe1aKy5DOL/oZn8Mw/Hm0FVq77y5v0gr5hkew1IZvYrl1
GsQOrHKeh9uy3Khi4qTxDEwJADYpFy9SczGWNxPQZLsT2EH3MWvQA8POrN7tQQk1vbFvlJrt6dc5
o3YWJ4kXCQ01seut+HTfHyoYiCqYe+ybjWAP84Bp4RwKhmmyUVvqoBXF+2oj38tBUjIowOjysi9h
O72aNOE5J2rthRzyTYCKZWgrhimSOTp+iBd+V8EnwyvzlxSjLlp1/dfPKOXxZfYde6QCM2p/rKso
jAt5ilEmTdEUrVuz2oT9Eeft1UjQp6h0wQjmmdp6qbCyzcMnR7j5yU/HFel2HYHU45f4AXKVRwaN
yFZveVMliffAaZ2FXlq7zmLOhrewtVx35M32fzTnXMrJv82hggWHBeDShUBqQ0c2LZaX3xaDxV+k
UfS0aXo+b39LokR6R4fy2PnsbVyp5+ugjEU792Jsd6DE1EToo0f+7W5ub1+Z8vCIVAlvFb+MtVyg
UqRrerynIiiyxpsVyVOO7hEIrAuQxTvGPRAkhPEyuHGa7q1vUf/5ealEUt6vD5Bx294/3TWu9wtt
kj963Y9vwZ+AdOxKSDiBFxMK9V5ChGeLp+Dv/1pcL9Di4a2tuz0KsogDa3zSP5JYZlcypt9dAjys
TXg7KgF6aL0n00X945B1o9IGuHG7djUWB2P5AxOr9cUVQ1b1Rphvs19r+r9yfqZOGBY/lfzkM0ck
DS2LWQ5o8vp31fAL8kYiRBDm7OHVPmcrgmwdmNTzSzDqFO2QGdecjfXqtqnHe0Xl3N+AdFdrZ6iw
2UFLrMDFVBi30hZ6v2/gd1Efr/Et2LvG1GhAKOteprX5h7o4DoyggaV+QlilQUUxE8AQq3wfC4rY
kINo55ZKmDXCRbok9LgPX6FSae5r9HcYTld7mYwhafEV8KqRuOdrJ70NzXBAz12M7X2OTIsYfrsJ
wO9pVmxnuZSzOoiBPYM6wGrdPvFAsYF1nBIHhrJ9ocKGhZMDXSOloxpDundYIK3ciie5E32RG445
KLlvvJ9Ex1sfx0scVvBhGHRI+lfobMxyQQ1n7IRPUB4c9pv8uw3tIfdedbc2aOJJse1ADilgKTiE
ra7dvjephRcT+dSlpo33w9GZiSCsAwdnfOUycQsrKpqfcvVVaUz8eyayeW2S8cfrRrvWniPTycoC
AwzrGHbBV1oV8dF1ZmrD8BaQhdT7Sx5hTaeb0yDRXUL2d3aafLZSEt61Ery9Pr7056Lm1fRDwlBB
2eRwyIAZ/lM1yQ3KXRl/TX/rSVT7BygcJMzdbbqJAuDMaQokpM2puTL34uhPkGFTs1j2cXlX1xh6
4uxOdwIL1GHxj4R6eOBkYaZ4ZF3sOgWA7I7O2HMnU8mjgUXkil5442On8t893zUJhhBl0J79AOeL
zhCb1H4Xdn15zHK263fjU54W+fuMgsI80LGk/ahw//wRzhytPjorY619Io48EV2kAeguC7lC78sL
uf8Pk42eyrKkYJ+53OjNUm2hyuaosGw5MxO+BIRiUZrnl8R3y6m6OmvxEGSFetvzW1p+2pKWCFZ6
qUdbolmz34s5NGfIM6CSrSz+gRP7q4xJDlUFE/r399I0ma5vmIOb8AV2sAUgOwlAkAlHX3eEs99i
Duo1f5lqt8zDX24cnDw3Nh5x6rw5m00/Gl44W5C4Z3gQjhqDZ+v5zXNSNuwSAxYqIQcrQSC7Jfuk
JAFtM1aMmeumh2x0nma9zotW2qz/vjmviF/HDFatQ16RCu87Yu7KYSe4P+dipFPhJeUl/F/uQMhy
x0FGz+Sql2z4jthppH9lTRaQpLMYzn3Epvm613CLBz3YTdnI8pYviHu8SkgR8x96uPQPUyiQ2HcS
PJrNJhhQJciIbP0F46vYhsWvaxEAhwCsri99PlhWuQkqc6tTR0ombVMF/RJy/FI12+lssRavRJQ/
/tMwOsHIDn4qAi04EP8sH30HZuTLPbRnhYQHt/nCN4CWi4JK/mJN2ikNYfS9c461DoOT1faMUnlN
bgoIn+DUrS5RIrsVnHhWfaQAHSP5WyOSQMFR15X0o7Kx87grD+eTwH+Kga7NgxQX2D1u15V60x8/
aAbA2cnucmxtUH+v3xL7RaAGTi7RlFG5RmAKIkELXlYF+z4hZf6s2brFwpSfBhDEASSiCYtv9bKU
tiTlDhREMDn/VxIVODsuKdInWPwnXjhHwBTS/BdAmBb3t+PINqo+arvUDKFYJt3kqCodho7oQa2o
MJIK1lgYNLFuTt9CtQZ8K1t4wB9twwCQ0l6/szvxEcAwv/7U4sIgaVubTovV8iP82ckfkDB6xR1I
YJm6lzAwH7ZjC289LRpIinJQHYBhd9H4kxosQJAAB+9LgrYQ3gzX99ySmbLzMcc5D1JGQZsyJF1M
niQBtqghvU3fkKN4kIW34wKXR7YFXNTb0tzrDQQPqNcBbO1zHvHpRmkuHdrdP9IH1YNM6iz0xVDn
t6gzPV91XPAQjsxpgHvuhXVW1+Awky03GdvZ6Xdf/3Qqzm+nSkBZbvQJukNL8DbgLTMRxfGxN9fa
/oVS0s1LTRPFuXhenvK4rY4Eh/1lZfXI+WA81TCSRb6NW25tYtVo7q2Q284yQvqeMqGFeM6f/yDm
eBBtjzteN5f284/bccsOXDk3mXnhL77wl/22PfuCrFlSswq6yOQWV/s49OoOGqIy+MMbSGjlxvhL
+dvQaHTJ13f0Q36/InS2kGCE5JEtXtWqKXzuiyBP74Il/J8EMERwUT6HAjpEMZrhxTkHMV63vN0G
KmvHxB3mte47yK2W8XyP4Yt3l407bEvVkAJvPrp+I4zZ/18VgkIThSA/Sa8Q75QBYakEDci2wSKX
qtp2lsgUEhxcL9eAxHwuWKbPgi+aan8Mp1R1rPdc1k/hf9wKaLwYa1fPJGnLVfcihpJwE6GwksQ3
5wWtUuMejQzP8d/sKzYmnK/BQvioemxGnY/BC0LpF2vC24qJLOaXi4WUfHR88F4HYuAtGA+WyiFd
Bc1ijNItu2Cm8PkWNodxEXN75bBlpA+Tqx/zYWc+D8US6YGsRkOpt1eSwnt2VlI8BD7LE8RmdHjF
iDKPk97fSQyRYW6uv4O7f0i3Q3xnQWcNGbyXWzlwNck/DNCRWNKHMGiCbci/zxGfBMxXP18/9o9A
q9cHhryZTQvF8MLBkTPUn7HDBH2fDMt4MJCXAsbHQ/akcAPVKyRcgPX+H4VTyJc1Nn83oyxsULr7
DCAKnmqBe8E9hSAlV1jwrmZUCt/GXF1ix0Udl5feXl/Dvr6DGF0fJoausX1GMu/xlJR1X90t/5CF
dgxnjULO7bDEB6gxDWuCdjZonpeb+YglCh8wulcPEI0o62h0q83W2eRcxDiZfL2m+YxZBcJFD2R3
/31FbD9aHlo+rSObMAnHhnc0JiaMVWmjfIWaEppWsJPocv6IyZjrdfzLOlpKZj2KY2BuJEUZret1
i+51GuaVTlKF6jHtmgosEh7crfCDwb4i4s3uyC862zur+bTpYtAtEPYdxXSH/0uXYBRRyw/aJ32Y
RRwRlYI1ezE8nXbKpeYYjMzDp9GGeZcZ9XsWTlQwrgGfoKsDlbYBg3DdsBXB1kWfvUoFa5t4hH2G
yze3Kl0WEXI9Sa6nM81WHqFMkkMenSsBHG/HkorFx6FYA3MbJEI3ArjrNrtgIlseBiVULxLA53kP
HQBWEGZGeY6CA3C6t4tNO9pGhEGfV6X0flKT7Q9t8lFwmwhu/gLIdFqy9FyeE15hmeDz3fuuubTY
DHwGHo36eJrCG4Djd5vjY9hd2OX2Z3Wt7jO2Hgr0lA6kEEiVQJ+gdkaxyXeTgdrgTWTTrzAyvhDx
xzppD9FHbDRbiPMY8+BiwQIY8UaPaC209mLeX8VAfSD767EG8lGLEPsj0mlOYAHGWaH7btoCgGw+
B2+mu5tv8wKXUXTLZkvCeX4YukNF1OSy5+WpjzibKcTWWE6hKceN7pSbx0nY1TujI+r2eaFhvAZF
7wkLmJC2AksEhPm/VZKTKmjQ5loEezU3fCchjxz48axOkFK2M7WAdnrzCYR+D/yvmnVgvBYvHvxX
h9aOIydgf4BIAKV/pH64/4VYTEMm3eO1WhjSf0SkOVUiMLriW3gMsKPuZkam82Q/qp1Gv74guefh
3OckPDFtgtcseaf9PxoEQ/SltrkNw29R1+qmSaiYEtGVuq0NHzTZVqCJxrXY4ykzUoJtHEJx5fJk
L6BuNUlnfR/0wxIdVZwNhxXhJdp6ffK1bOulHtOJtyDomaRAUUWgAg521Mh4lB9C0wCLYG4zrCKe
cb7DX1tAEW4t+xasz9Bl2ZDUwzgPPCEk6++76jIsYB72zGt2wtVLWx/DdOiVbt/CYDC5AHFFyaOW
EUaoe38MzSY4Cr6h57nrtKtZtNOoSo/jHflM9nGHU50iPSGZIfVi2LQBN66cgFTDdWXS69aDCGgb
p20LjPvLfi4185f5hibtKQFg8x2CEYflJlrXuflHrpNzsjpuNJhtGSQaySXfDbRWv4jUXXL0uojn
0SwCyV+dndhYkCx36boTtFa2PcGu1Aud673alERyRr7rpGTs5w1Dqi3hpqCofWxs+DdeBo3XZajF
5tSNBATRKqks+6RqcutzNe/g+ByWZts8WdQpQCwhwIaM5WnzkQAFT5CG5fQmm4U5q3IUkbiczoaW
Afoa7YAR8Zmt86qlnkfErFVGCVITASH/J3I1vu/P8M5T0qmf9ab/gW3afcpPECecVa6PFR161a5N
AraY2C2kqmhXhiguQi7oycI5X0Chb32vQnvXEWg/xs1OjceIwj+LrkTVqicVSvdLmAFFpJW2iLEr
xP2oF5do53+r9t37pTM5IUvvbIifIgMfDqF/27Pa2dYXiSLr9Le/daVyqvjPiTHBf9NXNEasbEp7
39F4ltrzoMPmHSwESK5Eyg0gDgKS8PON/MzE7iUusHCJwdhM5kgQcR0/bfweTjvpVerYQKPvd1ko
M2M7GM9ZdvwNzmhaUVNP+nvCpni7kVqd8jsyvLImarMFEfHAf00YH+ViWheucYb5oO5yPczeUv/4
AD6h5AL2AjlCVoi4vFoFHnkOKc1v5QW3xWzOp695X21kyUnwZGjl4JuNaN3yZtQGp0aEHsrIt6XH
OIj0exQHiTt0dg55yMXwx6aeovWZg5U1hfqXPwecYyCcAakgZkzKkxqPvJlSkR+lfQuu6wnGHpo9
X72tbZandPTXTN+bDwiiimyETLQLnBopRrlzvI8I5ZxZWxWLO02NfpxfxIKZlstqr0BJ6cH9m0rM
jGd90OijRh96tejxH8ob8HbyGrKJ6yWlqJv0oKGLrRmczxJRxebeDr8jlDne/X9g5SsfgQ2zNMQm
12TG8R/MfdzfwJ+nowjOEp7IosYsLDTQsIB71N0fujS+OQhL4VlHqNOoai3YHepdJLb1DSMCud6l
P6tvNJQL8G5vXQs5XWH3KFqTE8NBy+Ja/XxEGVojF3ZKEudDs9n5BvEs9Mijzq2R/h5S8tTQG4IO
3fBDVEYtEhqDvNGFiia/u/mgZnPBp0kwUF8UTD8fF6wU7ZysA5i5G1du4jinllh9BUpYr1yhoK6t
sg+IDCsknN7G0qwNWjcuBcTFzjZ+bbr0YsIWeBk7MuM3iyvEeM7HFEqqN0IINVCvKKBDd/y0fI73
PgtdqGG7KTax9OyT52OQmNVcYahmSk7NW+gjjTt1mpLsIPoc/AiGHK2J6DcqkPDB3/vVYOPdbAjA
Hm6EOXGAl00B+222x/mDIExAala9w/RiybcCcVgB6CEOp7Ju/iVHx6UtTebum2SSaqoJvYN+T+C+
WjHh3JgjayhX6c/bxsmu/CFAdRGGlPP/rxwtkj0TRcb8+tqL0sc/iHUzvjpAj/Lb0ZQ5ii9DrXMr
cnMehtuGTGDcyuNyfuksLp+8cKITwBHsC+EL+CclMsugaNuaYyGJhzVA8+CwuG0jZ+vjMfwLve37
v8LyNiKT4MHmxghVpAJ62FdbokCOukcNrBCAhrhviNeH/KitLmcvmYgcxjurUtLRkQXlnc8ggflI
qSj4MGF1sZfgSa+pE77cun8ieHGGS8Ix4SzKixHTGIwiCqvRMycm5k/UoMonvNFLus9JGqUnEx7z
3VORbE0mqDbz3HEmABYbzJNUva0N0Cw1gGlzsMdZe7SolKuH7iZFHPrZessDQrpkZnJuzwBCUKzh
icYpTL2sr2SGOXz1zlnzSMi1rFtQvSn5kbAU1vT7fNogYJ1pCG0Law3hkA0ABsX4P2PPt6bscskI
N1og3aheogVWvPB4Q7D5tyieEcf9p+UOx+vKq/2bPzpXRNsvBFxNOMPf/qeSC27JF4i45FglRxWc
shOzNREV7+wBZqLuJCngySrLj84fN8xgIuxW72X6WdkunsTxrroKeS5Q7975mRaPVAu7Dp5mCHxp
n2dUbk5FL9Ecl+fhCcFrdNVuAozXjgGxXHDmy6zWP22zS6tM6vhQobEy6fR7AbA7afWEkBH8Ifco
FaKKA2YCTpmHpWZwn9QKtRPJZVPXOTu+6vTzNBn0flH2JXhizOwWKefBvJpJXCmMc7R3cE/s57gV
09en7I4Tc1uwqnb39CxrkNnHUlVehEqxInvJMlaul9IKrUPZIRvvbw3E83B1AVilW9eaLXDrBpeV
hp64bJstVllQ5OcCRe9meClHgzwZTy/jsMe2vdeddtHWvxpMvbU+gfbGkamunZSbN24cZz9l3sRy
qUD4pMKqhE/wU0XDfm5GGSiMJEp2bhNITGRoE2YvmrDjLQ9oFd0WTl5pPfM7Wb6nbMdvB/14wk2T
a7QBix/PTtvc4h9LAK8auJhJmQUTd9QwDNRK3RrEGGRr+3LMJL31L9/lyAZFpm+uqvyZy7bDlad/
0QY3LPHnDLGA/hsc1pxZEpGirA4PKVuE0C2uO3h4Uw1mM+U4gEboYiXOhPGBhxJ3BPXIpr7aNxC2
lfbjQ5G1yhvr9EmzgJgOoyaR9H6xs++qAaZxNYRtwHlvh2OsYnbUeFPJPOwf5bsNt94b6jCZlfTl
Y0Sgop4J2aUx5I8EPAmylw9KRAQVy5lqpcj4yz20liOLg/kAVkSM4Jvomg9W/PlRg7nhtisaSRrq
vhd2WhfrtNOQA6xpw3v9WPlIraGt6nZxSzrh4nD6G6OJOvpePISA9wo1ttAp+p9amfNAnn1wc4ar
dG0LagVE2cTcoU517GlaHgDixaRB18hwW3DVqgfPrERowZ3R6+uPxyT0UxG/ZNydalLQf567f6HL
rUUkGkmmGIdj1S5MWE9EMyXPGl9JHO4jYZNQz/EtUiVuT4KYySTmVIK1rZzln+2D1T80fP93z8cw
wVrEPZItTSrZxWj95c8RnyJ7xMpoBHAcedyDUpSJYD4PewTWDEr6hBVlLwtkvd6g+V0iB6v//T7j
NpyvpV3v+0HRGhn6vK3HPl24/U10dVVg7zsD4Tg43NChF42JpAh/DIozvSZzyM8PvTLtUkxAXtAo
gViUVqObVuVM8IR9yLHpJdWJMjb0Jk5Hsa3BtAyXKZe8oPEs9f1Evzdsnt45tJUgeaFWgSzBGKbL
Q91iox386nqVeIPnDxOBuE7KHp838kT2fGX1rvqz42A/8fFyINJd1PPW4CF40ockhMTMs9le9mD1
T/UVZj25KpIt1ucT8lfc0sNSfdeXysdpGQCTpAxm+GZpgWtWP/yczvz2GrLYLh4tkLnt5GQRbWzQ
zD3FGQXOs5tzwuVsM8fgH55H93NWRaK6J4ofShFck5jC1TBDPOyKk2SQ3WD/iO3Y9SXv4mou1AOX
VFvY/xBUgBr550GL2CQtj72WCnu8F9c0lmeTRlyu8huh7hYkVpGgUHUyIavZAvE3CrixXBGACiZw
D36w8dkH143JhItAFNmDS6qijMlt5IytFRjU/QxU16267kfIyUpGeTba5CnamggHZNlnDa6TZl/i
eK5/jlX+fa53Mnk5kaHxKOywnfwjqnFnDxI8fuYJAv0zeFortbbZ+F1ecX7utXB7fgTV7pDwQKcQ
XjKjJO9DRTB8HHB68yoHfoph8O66Svez+fGpQ9+s5lKY85GwwmaGhHI/mn9maf99GFWvw2z7Jm5c
3JXI00CxeuufUtVBGwRMWkOMwIU7S476bdlKho/w+DcY/5rcXggrN17MaSE1ATVOIXJGG/vo58KC
O5C93zfJvbUwD99HiqtrrWDGwM4HIB/8MzTomhlq9dtC0LXNZ/h35ZsjUCaAR/c7+UT3NKTjBWoE
3tZOd65y6qo5WdxbomHG7ZTi2rvBi7AUD+hVMn72vPXPQUFYtt8eWqxZkXqcMMBtOx5BltR1pWnV
4e+U6hBlEcQuWoSFFONo77p69UFj6suVUA1QA1/x8nIRTtBAiX3sXQ/7t8tLABV8A9P5Y0QsrNYP
nW+JUTTqLzkB8J9i878CdLO11jtcznu6rH0eRfCp/EFeU6uB4TH45mh6lFpGoX6sppPkyVN4oEpy
ke+Fn2RApTOEWMpAdPo1EzNNvWLqNTDgleLU1VvfLqm8xv4J42FYeTC+xbtR2hngXHL9tUnLtwS1
6LVDQJZYQCB9M6RgVTrc//3otOR5g79QBvKDoo5g1kojTSzQmwLWCc+t44ePiofXyNJGoJvOic4i
GfvljUzyqWcg7ykFxGTBgCjge1p5Sy2WU6JVCQFrjA4J5gxh9fx/PB0TKMh6RayxKuzWwe2/yCIN
CHTmXb/uep9DjhNDG1MYL+HxSlhhugTSHvIqyioeNUnbz+o7GE6/QJNE8/giOm2uPo0S7QDwO3fx
OFugJinOdTuiGlSiG4CAInrK26JANxAIVcW9hnG8YSx2RNUtaQZDPM7i3w3LyQsddk+moc64k4Fv
aV/UV40ettMcjUeBGI5nr3mYetQ7Cf9OPFc6tdqwbne4RaOieVgs4KNfRsQtxKhQpNyRp3mWi8fz
j8H5E+6ZIi0gkHEmQQyHoyYQon++ERwO/EuFAOX/Xb9mr+5EUddkri8pfZNRy0LNxEvZ3zWgqWcG
zo1JccnkOZGwjHhWcXwpqKNuNhylppqeQ5tIPpizniH2nGRDzG9juvFoB51r7+yfd0G6f/ZEGfKK
35pReXO2FiN+ncRbfqQFgBzSoQVinT4DJHtJA5GTRJN3PSOMYyQZB2PJFd8ZD8KG5ohtx8Xd69vR
EZgdLTjHO1CEGghEqZ8ci4QvRw4VMK6+LTN9sB05r5fj/l473hB9TBPehtBR/QY83zdjhC5H7bGE
ertjh21HknfAnNAv8JRp/MPkxlCxSC3UA8lYrRjcv6Je28f8ZtJ4M4QFVyxHjsZfmG/OejVnM7b9
uMIFfpvLOYljAbYebECqfEEPu2YoOVO8u51EuYzx+zZZvAV38wtPBx+1W6HW2OuVsFyZOLKMWSnu
FjFq+UwMQRIS3HVcOgbbbqj0BMqsZrqgpS7If3T93SzX/5fTUIUcI1pZXBxPclvYpTC5sQw4mW7r
80KuX3BQAgZQOWpnBq0JaoWZzRgIJUuziuRYChD7wNljpdQNE68tqfxNc0LbQcws7uIG7HPWaodb
yB6tvP0DFjLNjIscRY+Idi+iHwti5HBpFJzmgoEeBt4gVR2GSweNMM2N0YIjwBcGny+INsZ0bS/R
2t+UK/GawnJ0pKJMWmlEd6Q4MvM5MTUjZl4EGeS2/zWOGzA48cUYSwMkSi0g2E2BF3NVUuoaUcYJ
2r64IMP1e18zRHw+eu7msLR3lZm25rIYLJ1id8V8YZpiECvvqO87COShDxjp+89eE3CDqZocUmik
RKKSsu45geZj7xIKMvChtDlRMb0JD1MgFtNJ3KfzyeW63VdCkpV0eQwylGEZTUVLscdu+3EyIFuz
T5y5rApIvVEOW7ucfbvjScdrkT93RLgDoHgO5TIN1dqzrDhGb9PnNL130rbV6snZAJ2Hq6eTwlMf
3RaFgAU9UQ5y4c/EB/UedXX9S/O4Fdwl1dNIYuGTsC3GPm6o4WY/pi36kzGcQqpNnDOm4iAwsHlN
qLq5A3e2Pc+P5yBHSbgn4PE8WOSPBZt+d/gF7nsyH15CykYHJLoXqiLQQuwi40omERxhsDAHZvNP
n4Cq3OyGbcEGVwW9EDk64U/F/WdfzXDftBoXfhYAMPN5x4PkBamnFbCCSkxgJOjE5fr0ddvmbdhZ
/API97M/Sgf1emVGEgIjt07ZvNfyn2btnFk7MJUetOAU8NE0kFnacK/QsrcwA06N/6u0rdLdYvfq
QaZjnwli5Wxa+lC6PrfEEy1UtJC0vODalPYGlONn04/z0dS+u5Vs3imgMvtLcdRN67yLFDIhUW9h
QKfJymPY2o6XgWN9irYyx0e1+Cs7VBITnXX49Yhn9c4L21PnmeVyGnEjp3Hg7LZ5oZX722nQj/0w
6/y67oWOH5ovLdHj+q0YTAKD8uqjtlU/VZkXV46miIASw9nYTnCDDk5BCjw5n9RY/80Nf2QznrcL
EmVdC8fLC6PuewnTOKiLB1wu9nE3KybUXTA/eqNxfZPvubjsW41bWmhT/81EO8pXKWOcH8dXHzGF
GYTV1YEAalzypDSUJfGHvDZqBd3jMi5Bz1fARgTtszSnNtl1F9Mri6B9pti3BC3bWFD08RaA0uiT
hW3qbV3v7kGNKf0n69VLfWqx3bH22mfTqVf/gWgo96AlkR7ubz8Kp0BVmR3lGrJjzl375zrBjXuz
nqx70VDKct48BXvtk2F0qwCMOlJx7k/kecLnXrkeMTKgv9fVap+WQwEHfyEN7VX6WRm8A8SNx9Cd
kn+UqZWeI8PEe2/mamI3UwzvYYF6XUaSLU8ZpEJKc/SrYr/ploq2WrPQdUfBf9j/HNRC89sP8br8
uv0c4eZZlv+WfsOcTJIVKRVeADqIJG/FaB/F94E0lTPOEBL0k2i46UvEOeQXoTH2bDsnzBh7Fb06
AAO/7cBRe4GQeh62Lmcsebj1XaSFA1EJzX/49SB/NpiEXm0aiFgxB9vZYHY9mVxdM4V3wUAvic4u
DKeqWdCRRfLUXmOMIpShz6dMiFquFnMP7LZzM+Z9AyDfKUh7Vl/6+5FsnCaZBeqHnwhL+iht1R/0
NS16vRwR2TLjjzL+XVyAZs1cU6jlHFQr+laJg/y0V1Ibmajqc1GQWdt/P7sTcWXVLGg+/zKrAYnq
SHmfYlbdOUkMIcvpNFMqVA/Jq55gIqe7bLTcmig/fhxzhHFEfFW0KAiAQyDBMTQpwyQfNfk2GI94
mvJoX6Xr56nfuVy55X2IWABA8RBG2qOR0snI/Hr02gGGG3lgi2E/ZIrm8yImEVnSTfHpqVbeF6V9
R25cd0JOpPksl+R77EjlCZsJwQzpMNAYqZQh5YfgpxqsFVAaNjDk1Ff1Ralov921vF9Su741zuzh
Y8qVPZt9BjlVP0oOyUKOkOTcA+Dp6XMmtBK7vTRBF6ioFY9SnsKq7XKqsJkA/k4R/JlZYwN5gWEZ
g961uvPa399upejyXWpTzcWFQ7myh+TX3MfiRW1wBjyldvVenyQp/1LOh6KkPFlRKA+q3Ef2jg8y
orSXyYuy7GKsgOElELmQOpYqqAQ6RrdVJ93dmo9DGSYRB6Rv0npzLKq/d2da0iIXYmepeRhLy8TM
+DW7W2eXd6qRRaoy7x58X+UQ0z5FXA5TMyAOesV45m7JVPahii5dLvHU7z5ltQZyq+JvXkZ7fg67
zE3PWtJdBp6eHaT0iXyPezUePQ0VnilBsYtmxS1R/mFKe6jaG6wrjR55/OOAr3lHiFzTU+dZASD/
adrfnP4wk4Wm/uNmFcjlP7Q/pJJjiGYMvHfYgjQa0RkyHrvlhzamisfMR9d6ZxFsHKTc4kPzKzMB
Yiq0LHrVyCyRbuWpkhylzmFbqRZPmiAYxWNd/c/oL/2G6HAz5yO7NCtk2qjKys10sfIEp565Ig6b
CZIslSwV5J12tNi78Wvax7ErxmsEJfMh4WbDxuKolsnxHLa9u8nuJGsxV/3r+qpcgDxH1+HSglje
Md+jLa8YHW9/X8R4IqQyV+Ro+xTUCwHyG7kEW8XLK7Rs7LFqRglC6KYj/OFmCLFqNgf42nPnsMfQ
mbx5PMTOK1FNNir9raEkZIGbzShWqxssYkJ52tqeQlFAPDM5gkK9LWUOCxhcJgfNm6HfU8NK8SVx
B3b8sl0rGST9x6U4MEacP3AULhi5aMEmn6b9EhQOOmSHh7Ba0S5kWPviQpFZNrLcjwLaVMb4YHLy
PKyxslAXM//WIVB0/bhRtcdBBUrlqwERy2gNZzjiAiO0zP7hvkfxf/uMF7SMZfGK2sVyeqvQdFVO
aAPXX7cBI7jveyW768YhD3k6Nfh8MGcwbtSsJi2ou84h6MoPUScKYKz3A0v72jXm7ThYG12B7NaI
YlpNPudq7tzGRs749cF6eqAOoB3HktKZQC0CNB1jfNLR/LoPoitv7OH+BwIMlxHPnXNdn+/gW8cM
hPOo4jQmiTGL9DL6zUTPKSJIILh+YZ+uEBl7AigQRSWpjxADyZxaB/MnqdtF8cOFevOsKQ+zpEML
GxiUJftC9HzLeux92fsX7I8M78isPiWJNq/W71QoDmrQwjDRyJz6X25ZdpcB4tDewa9pEFY++P/3
QPqTN7V8QhAI6Gs2nC0hCpoARQpK/6AQPJSSulLpA3vzUGKeo1hqGlM4WT8W3e7SVpN6UxWgZTPT
rpjafYKxNUhNnFRVV7RVFAgsXjTfMhFsDmRgdOfyAKrkySBJjUPfohO0utByWKc865apXDoed0gM
895oudP+VLa0RxgcMGITsNiOcrmldr+ek9jssIoPy2B9qZcqsWB3zUIUH5QoMYpHPm5fbIEo0NDM
yzIPWgsDWZXCCJqwn7iG9eX8I93BCZbXX3OxzYDmVJ+9XQz+353VRaa16wROUkiXoLq47we+sq3E
PwuHbqB5mpbqE4oeh2QawGBKBt0dU9Ct49oBMbqtsExffLICupdQ4+ZqPbJToVPhikeJSu+zLroe
9Glrx11vzn37haI31vnAHZ3Sk47Hoy6mfpmb2NWyGwMbqSxv83VRWLGRZpLaXTxiXRUYk/4C5q73
ciNAdPJ307N6s2qdjQNxQk6Ny8Sc/dJpEzIe3AmJjP4gPNiWyQv8t9O1Vp7PlmX8T5h7bVZqx4pQ
JFZqXN1iChQtELnbR4HnF7vEGLADOT2RVW0tHWUzPAaBvtQp+OZ9KEhi7u//727Hr6eTzRUmu6cR
V4Vn2CTIywvRMAI+QcVfxhyucEdocHIX0WwkEEHBJeH11ZrNv3q8jqR5u+7iaaG6KmkFh2zOCD2a
tsfl/OTBPzmOLKP6TWGJkr+YZjBEXzvFeZl0iAzpGtILxle+YexAQ89M7+yim5Y7HqZdp6gjbPOK
FK2h91GVZCLKrWKU9BzMU1NFg7IYigucXHQL1fwKcwSfKR63emlr/mdMGSU8952mNlPBPujx/2pf
GN7SFNJisBHqBXQe2ZfJZHDR1/SymvBevYoEXLNwwAWDnevofclr/+DoYnYManRvPm3/FEMey0fT
3ahO0vZaNtTrNzXSgVSYlQ4+Y8NMzohxHseSIn+x64dkvlEHm9qBedTKb70HFDKXQ6YRNw4dCr+L
R7el4ZnoxyD5/1XXA5fNl3xSiSNzvU+QSX+4xEuHFk4Uo6vnC06ikoo61bGS5OX2tovYdA6GKK7a
Z3CbkNRqY5ucX2tHesSN+G3W9EsMzuh2MaToURL+ecbhPmB+zKu/xm1rNkGLvSecmYYuxGXSVErR
e87AB9wfeF//UMycgRQd05nQcJoXTa/nIWcelqYjuPK8oVYWPcuOrw2oJveDWTfC6Sqfx0QLDdG3
qg7GWO/E9vSUygpCJUYhAleHgc5zEV7qIG59fKsJeMgffA8/GaZUhPVPn/RgPS47RKeatL48YlBl
u6plr2sID4L0gYEQRPz7ippp0LaiCyX4f6yGNCLr21JPZ8knmpb1Iqx5Y/nCxLMAPL0tie2DEH+m
zfUwdZvzBkULQBw5Ui7mxEX8echqlE4er72s+ve/YCxaA/9QQCx2UpKSafZ7YR3Ubh75HY4b5Vjd
ulNQU9gRifMOi/3kQfU687HjYnoIWSgla0pJftwL5FG7bEhQNXsUzq4vwJmRNpFXzooeDZ4ofUlP
1ghQYKU9Pvlvn8O/M9bxpr4exzcIsUAuaDqlVqpEhecon/qH5mdrnDrUIPHp/fo02FoYZKEwo0ss
ujK6z58h/Ww9IJShlB7xTwrHwM7DLvBi2omHdVxznhQ/ufaJr2w8/q+Yngfok8FOgnbLLnHMj594
Cwo4qxf1eiPDc/y7NmIxnoDF+Kx5XoGfq+Iyf5NXTyojYPjZnvCrfcpTSdUfSdC8atRDnGB0c8Pi
lLFI3YauVUu00dgpxKWklrCiaj30EgXjToFIgyAfXabU6QmxwLipCS3KgoB9sAyPsVYsx0yNrxPr
MHbcQ7xbnJtpdOAB7NeFnAJFlxb03AK2Sbh3T7uofFSd9ItnvzAUUAnLTJ/A5vHRAM3ydKrDgp5+
+0cU1yxesiSJd1IlOE0GR4dq8rp6w+4hcsVUiVGMBB4xDfFkVZf12mlJlTS8WYQ2gNMeZbJqQCp4
ScqPY+i+rr5UefgO9vTvIr6+D7rzY2knUlDDzB0xHQcwx2Igu/5tiL4gKyvsVQMxfqkr5SwoAZJj
fZunAvsFjVg3wc2oU/yp14DTL1JVoeSbczFZr5cLLVsdjE+X6k1lui4RTF7g4ocHnjVa9Lj6yZ2Z
Rz+caQq8bsdPA8NeqzPhN8Zbt2pLm/A66kq7m99uzl5CKCr829mHqZmuV06tE4VX3oPRzZLFMQ1m
firvEpfqG3wlhkYLGbYqP9GMdy4xGPzdjFpT+LnoE0RDdISXgrrxUkpPGIzOF7X05LD+s6jCxjHG
RDBstL6RcdmRDwpWUcoYCV6Mtg88LWyzExD/czA/VJlqSQJo4/lSd5HD7oe5Jq0RPUnFEfZ57tfh
9GeyYn4hjkO9w2p6+4JtmcTQ59ASIHQAU05SA3Lx4yoxz+fFQsxU2xtJiabJ4DpZYNAwFBc5/xpZ
dTyNRyPD7mjAjYptNdBsSpes6ZdgMuvJ9MyFxItiot/fEnjUdDAIsT/0HvCmJr4dz5a9pZKPhEw8
0xW+w/xC+kDV0dPK/sS3pc4Zv5ct2EpbCICVXywPbs10jNlkLUHhOM7L2quIeQynwvEWkeb7lFsm
T5mGn/LV7aDRRB3HfhVRrxjED0bp8EvRnGKDuNRVIhpPoc1ViKmQ2xiJWszps0iUu8PF123B3H+1
bF2Kw/33NjX73lRCNjuolY7l0K65lWOnDB13WLD+L4i19Dcd8uQw1ihP1y8xtTR/dsxtkm7Rm1eJ
5myUx9MLKEgE9ZOmyn0V8YJKcnX1IpQzsMV3KSAsqDRoO6bdy80r+5fDJTuu+4nlV6nyhaR3tGy2
x4eXzuA5qzzqk3hk6Nydp/6pujTpyM10ySiqXXuC/9qXQyBZEfMSRWnWhbdBuMFFkTNvFm4YpZcj
nC6XEn66OxEr/66+8Wqm6un8mkKqSwiqj2M26ODDE+HkdlANLtDQ6hQqoLleum/j5DHtc71LZHgy
sy09RKZk32x+1KHAqzbNRZj7+ARA0lVRapYNORAcO7T98RkLWCXghg8bXsFqdOpun07KhdYqMtru
9iwPUjNLFELpfxz/LhywdszwhaAIhXdwiz/vFaZzD8nd+gyZpN+ssafbY83dRfnWYJoWFrHCdvPU
mLNGCEdRaWicH0+9CGDOo+l3L2+Vpj0X4XUgqHKJ9KcFMyNRjSdR41r0YNX5DeWdhn/9yUBo2okJ
LeQ3V14lBA1cTntIAXYHBfcR8OXMVYS6bGUXG+PjXUgEbMWW2TUXhEqaUx7UEoHZrsi4X0PkFwnH
Bmu5EwZ5Sb2i00yZv3MNGrtkk/Q6LJFsmUeL8sMThAlZfdugUkU/+aQW023d1rTMRIzcFqT8CCne
Cy8+q8WwGAE1Z7VCFHqvco9IzOSjvRQMLodvFL/Yw7HkQSnlBUGQGrvXp/XuvF+wfWDoZKQqZE0B
gZWyDRk6XzJPbueHgNCtrr6ILzBrfHS1Oj65yCj5wfcikX5mhOQkoY5NAgntHzp+4YSiwiFjbxvs
4ODekt8f/OpLpqvCIRS+SyUnDyM9TpanOr+wVgtf5pgHyjrQgojaRWDH7ZUVecAZKj2wCGRJ2YXE
H4W3a9f09UUbMs61numarlokIZGi0HbFCgqSeIKzJrgGcUEyvGVfHthbU6hwccBfn26exRodYUtP
PpouBh4lNjmtzvmCxcSDigwLST6En4r1xO9wK2ag8JJbAhITT6gKUnyZxLKam323RFRgTugc5REU
cKJDCNbtm3eG30+3f4TNSnIH0mXAU73RoVyfcM679z1sFM6ZMI+PGgYy+/BNQEoNtC20YTK/nIHz
caz96SsApFyKN72Kq3SO9SMGjgeGPr+O+FFO7G2DzeA0XEXCz/uqeGzG0e7rt1gazex3YdCXrgAu
Jfp4JQHt72di8coP7joDQwlZsE+d1JsPi4qNCfqjMnGx+MbkSdt/fp8nDvN9alo3vHgSlhAJqyGj
A/7XONkpL/scGjePcn6TQ4bao7Iess5K5JWsqoxqIDtqW//pxLE72n7B0QMnnvU6bJCZlEf2YzYl
YHcDNOGy5tCc/fO3dcSTS7NwTRJ4t3jOOLhxiOXltzok2j4w8Y8vjQyHI4R7lP+Cgr47EpdwKlJr
+tVyaF/42QEY1PZpCnndqIbFQlz3fpE14CT9e2I4Nl6Dnn1rYobtZgYzt9NopD61fYVbKs4kwRNV
Rct9vIEFMub5t9hwsrEUML1w49iDSwZDn3gRK9u81ooBKZ1OqyoqrfXc+k4kMlmkQ8dfVIEUqnlI
goTeuSeQ+Y3LqPqNjr606cz0X/GiM1hBSYrvixA/Q8V6zbmTkk/H+kKR5zjdthbcWAKJIaKtsS5T
UkNewllbtiBjsBN6clxd3B2YUzpm5BSFuSvNjlumsjY1TFyPcLZxfonJ8KDoTQeOiXIX0fFFf57/
50mWHrowm1bW7wOnxzo2u+2k+hwPS8A+lb6BXEQl/q+KBqv1tYthl22nUrLZpk0T/O8Zr9iNhzVa
1yNjzwTVKPvzJCs3z0mWsBMBO4CMguAUdLdnY6QNjpmM7g+1tX5KFGDivKFTMW45RnR6/YYr2mtR
HzQuw0XELCzmJF3x8XFe8Dfqk1xn9UUrVFTtmTQFQbG/RIRc2Vy+ds3MIklOiEMnz/+DvhP4TmQv
NxyeaHOa4VOe33yMl1DAzUtPL1DT+1sKTsZM7IOx3w9lG6VVcG4EOeKY6sqcuixHjKZrai5MZ4aw
oO2UMKaCLSdw2svc0vnqy4vpjvz3FktHquBkBIL7h+7CqEnhlV6t4ucc9i3NEaXGZHHf6TOwcYeZ
sRbpTEK/9A06Nt8941y1BjiVMAQ3V8mJQeHR2r3lGwyKs0UAyCIZJ9fi+bv/+YQi/UFZcEggW+dQ
9HE9ehj68mLyWtMXiG00gUEDvfBCcUIgGoGo3lHMMh/QACSzi31MWHfvHheNDlLggFJF79qUPhyQ
T9FNYc1YC4wh0lmDk2hPGTxJxpWwp3ulYK3mWxq5tJqpv0UYQ8hELq4E5NhFMgwScMu+fO/MRt/o
4SOuTsnS1cc2ogFKw3Cf1ahMYH1qz+93T165HqpiE8aHhqDAkldww5KK0bog/aZX2jZXbIF6QiZ8
ZFs0uz2atBAy3hY/wohVHXkxlsP1+0t4WicrCZE5TEFd68Bw9uN+eGOTrGsbmSSLwNdkJR/MxB88
fZkJAjjJGNGxFVH3D7EijqgStG5r/iAHffSr3ZzgdkIkTXPedn8tJq3b0K9ZzSvVzglSzWMdLyej
Lr6x8SQRVVWXZf4nTwIkTaC/PE2iZHSETOZLVpFLj9yGQnDwjofJiew2qXTJD9epShF/Y7PrPNIb
9tpzvaq3GUV3av5pciaZoYpGb3SyJe4BgUn3spHEQwbwxZinb6sdeAmlNyL8bEquYweGHp55BeM6
Cni1OdFSuRXsYd23iBZ9Ur161UYE5X9QPJ77Sr+TnB55WR60GIzaFtvNCHVELuX16MZHG285XvjA
fRtVVt2oqX1OGw8lHX/+uOGa1q5V/mUeUwehh6wobN3KqykkfVQqvJhJBTCTIqvCvP4MkSckGA6P
brcZzw2U5XpkyFNSP7MAC+J+cI0lgN/qxlbQiOTcKsz1L2+CdhJPGV32HU8d2qFMiWMa8GPMYLKI
pbJX8vuC5t4b5hu2B6EjMox1OTT0BwPqI/d/hanr8eDP3C++Pt+GIPsu1lL61Q24uB7ittzVNxr/
JDucf/Xey/WjQVOu5y6/O2Zyfq3Jg7LcyW4aO9DolHyeY0nKWqj8lJWQL9yyJkPe54DJ2C4Pat/w
v23z5QvU2BXamKIW66ZfbKCzcbUfh7GpWtKLJ5rnMBQXfnygeqIgwWx1Q7hrSxL2XqtCN9qiAszY
ndT2CyeIve5zf/FZ7Zmn7I/cziiQquMkoT2s0yi8W6EDZ6EbJoBbg196I7/CE9XmgRub+9uj1CaZ
v2N46p4BTx2X3t3lrfYAHwX5k/f7cRaMhGoyMzufcNfi9BgPzv9kpQTFQhO6f2TJxNon2FNL53EM
R6mWeGHGwJiyXUy3WbjcLYED6WqwhmfJ3JXemQIEa8KWgtOrkxhg9Hri9ctcTpzmuBy+EkHt9r5S
2WavX7EL38rqkF5vGF8sTqH0EQcyAkUDdZO2wX+dEB6riOC7MsDDq4jtHFXkV8yBw8zBQHLnac0O
VEFo4PXi7EWAAmycTmYxiJXYZuzkAt/186n25/4IXz2BEfWekaY+49osNZat1rCheYlPMt0BJD7F
wLaUelDh//FFxWBwYZZBkQi0C4WkL2nOZdzQ4uwMzSVEjxy+pXy6ZLEnaYL1YvdJO1AQTzSQR84O
yCoeLLvjov0G5NJbU7X7PEV1Ka1xDtC4pHpQLIa13S0wc5R5CS4hXaCRPAFRk8+iFHoKASsfx976
9eLyiWh5DegW0ZUQmsO04fQfyyCqkhuPfXct5Tzc2XUZA0WTM02PGkxyjLUCnA5ptNgzb+pHOChf
Vq4+z3biGVhOzQyBRCGhi7dY9YlojjzoDZ/RY+mE06CKHOM2R3/9DmKmKpsYqjW41dAfNfdTJsYp
N3aejwJV2eMDVbYFVYis//02pPI/U9bhfUoRMBMILeA/emmQ0w0gbKzVJE1AEzQnwkJOShy9QaUp
rMXhvnv8PHK+Q0YjLueL5JV8eM8HvvQpadaw0vYb/nggKSXMyeNqh5fIGdqlORswQfKqlzGyPX69
oBaA0dnLySmc/7g7YLNyA1NMG3F+4H3Dhfe9/rCe/TkFKvmBFfddqwy5uqT5HrqHu9r2IJX1xvat
e8wZXjudnz3Q9ebpJCXj9F8n/6l+aWC7oQllfDDPszxmrkEHgczI0UHeGbt12FLWgBetey7/YXlq
ng9aJf+FFzLM9KOFCw1YP/AbjqfDwRwrigHs5VyqnuC6MfXIiU/kzuBvAm411DFygQhHHgG5rini
C+ktT/olTzj5n+QugGJqQ6BWckMGW/6L6qKeq0ptkFJNZOdqSWua68DeJMfo0Vk72MGu8iel//LP
yZR9d36LdBTlg1mXV7ShPMXQn9O13z1l4iDrW0AZxXVtSpRusF6pSUrPlDXyxpROrXk8H2Niyn4z
hRwL2UfXCRnM9eJh1KtSl61hvqgWobE+qAdbH0rLX6Ady+sCp/FU7l8aN1TPY7B32A+ySRSWN9wU
dU5ZnOdbAowa8QiOOeCZf4JDBLNV3jf8C1XiCGHWKNuI+HECEWgJoS2SydY59Wh2j+pZfF11enZJ
9tUA6YmsG8p/2MctpXJAdDcNpq9ecfOSV/tZsLr1TRoYOnRETk3xPix39K/ykE/bnjKfrFHs3xXD
l80NX31uZJkL9PaVtA2U6/1M0WhdKjrzts/Pk1+sB8HESUmOPEoaC0znsPyP3YxrtSktEDBFzUvI
AJauprgZpAEu4wZFfEJ0TXzUaasBF9/KyZU2tb/8HWgRBcCks+qPQOTVWlUt3klFzbQVvLMy4w8F
lFS4BPF+18S/fqLLKhytlNAaVnNMEP//p6hrlHzqc4ysOBeV2JHLBhe+7iLEY6yHCxILSQT6z5CV
XU7zDnBKlzWQ/VWE0x/ANFLOpKPqzx6vNm8+kIHpCEmB7ZtGph9BvKPIrbjDecURVUPnykluAoLe
sIUQ82jc0VPPG3Ng6dhiI8/bV4F8PnDQJCSKu6Xjx1musDpG7Xf+BRad3cdXVdhTRkOwRuHhC740
MNNRg7lZtXb1F2N1j+reMYu6LrVK/ZOjpc1HNq9Pi4abiFkcQIaN9o19yERW44Vz81R5J/Od336B
/Tsfgsev1Abzayjr4lck14VyTsmMee7UzPLjmnhr878lBBIWvfg7mcUXNpMxU4/+QPDQ49y3ObMg
KtAxoqXO/OZ6onfAro1wo8D8+Khr19zOnBbyzZ0ZU6nhUu4RCdgWWOtkmyV8QPfyZabdCKqnH16a
ZBuZdogd1LvJ3y2yf4++DwNXq/qEMDiQU6b1sp93u7jYoCulX7F6ghkbyccoh0fj93zw717B9A/M
oKuIrf8/AvS4Df6z6fqI7Yp5myxUYRNdy+V5adCxYAK1C0yWnbBAZrVJwqtKNq8FwtfVhrdyvQeC
wIAs9N24V7y0vzqznZIWVJyx64BsxNFCRm9Yg6xHAgJfE9gVSkqk7ddQV4Gd59xsm+VSe2xfPvNA
B1+KoKsXXsF6oBm3hQQLo2Z6jigaHVVHFat7Yx96whCE/nAe2wU9iTTALiRHLjSFTcZzRUGlP929
uaZP22GHAmz3pmX9iTZ4Dod9tA0P4rkRb9RWGbHup414vAqN+yZago5WMVhreGSQlVvqEzJXcbnN
9ZWKIBgqqtHZ7FslWP6pZH8CgHa+TAhq0aJnHn1cyjhX9KAMqa6tiLCG/WwMCjnxowbDYsXPc4+5
7hIosU5xUVM7f5xitQBVQmJ8HRZGKas5j1RQSyjBAaqsFnLxUoerN7r1u5Kljkl6/ff3AKWpctgY
0zR+tNpuqsuylzKQyYObPCnzeciczH1LFShbkZZLcV/xvDIhOfoIZy2YuXcatkNQpSUttOYbwXkW
Faw95mIE8LuOX7J0+PlgL8ltj05BLh2/3mYcDT1OBu1oSVMHuY44ZQOaH3Hj6rcMI3sxaz6DSJ7v
ekA1QNGQ1DALFueV4824IGGDf6WST6z01pUjIH1hDyPREUKo3TYRh5cBQ4JreyQ36VCD2q/7vfsv
dxbG5nHEFyVl2LDoMiFAqc4j4Ne1uaWYkG3hfQ2ZdMvPpsAY3XgEMUrHuVMiLGM7xJpGnIUzmSjN
MixKAafRSzuHWAcZpY7HcavSVuJOxOxPueJEhmk5LtRDZp0zPmls50vxZfJC5YZkHZiEnequKhVs
DuOEDoHkPYAjzA+Rzo/7BINKdzkKcDRJiHSB/LfocrpTqeCgRyZSb+u4nVlyNoDbL8rCrWH3KFNX
myOxmLWCuweabgO/b5z6bS8x+tm7vNfOQqHkQlsgUlU5LbuN3AMPm0sOW/3PlGD0tIXcLloXISDY
WomKc2lrQ7lfP/J9a5/+QQ+m7oD9SbnPBszjq7ZXl9MqXfyeX+iI7gANFzbu/8m1/o7V6NOKQfUG
Rokq+rec7tsCtOu/1ewqRfy6hau1IlChH2MfLGzPRIjTdPVVPaWCM9pI/+k7jQj5mwKik7n0ruyQ
ZNstOy41MbOdg1T157l3ZWYkWNvecAZLfc2wFQUji+TA5qaZ6YkL5zLTxo3BVCkwdoE97FvR5K7/
FjTIGJ6pbcoWBiR7Xas3Yqv7n3Dtoo2B33hEygMofy7Qvt46U3MT6N2UQkOBRQNkaCPLX08h1koP
RFyIIougOt/QE21CmgpRj3eOLcsGYt3iM4v8CJyBlFsly03JaHqTI1n5EPJUepT05i7I+ASJ2wmW
fcWiNJi98Pw2fQtI0ZnPW1HgqIgH8ZPfUvuls/hbmPhaZVJjK34P0IPy0aI2GR5J6N1Fy4guAfGm
pqEBPsb6wXnQzIcFGCNEY858qN/yiCKA864vzYw+xYuUfl8POV4rX+EZaJvJTpbSAxzc6oeL72fF
jVXULexVqlqQDMuZQhDE90OV9WtOdrMsCg46Z8ZP3zY7R8Gp3jqc2kxxqblfT9nUZHHsgkyUnzZF
eQmOM+tNcEd3CM4RLn6gqfFh3ADJ93Fj45QZV9coBnV+UjLevo3AgwjeNyuxh9WDYCTNSlTrSSWs
80TSr/hyHRnjNPxDGCsa+wQgdtrdk44SGzHttCIUMbCftTqNER0aaLkRJ5c7WLRKVeyBxPynVMEY
u5MCIEbUZlM1E+PPrSq4awJ1CTLMaWgfQg9p+ewYUKiuy9kqJjGCeyIxOsClwMBE0j+BwNRuBe7P
SyzuUDf+EK60KyGFY50zXvwpG9uMcMw0EscvgflJ7Y5U1ogEX/ylRGDvPRfWysYEwtX2AJ26ucij
oMbfmIdDf5P3vca1hAu6xRYifQRTx8Ad11aqXGF6dK5LWr3OotcNjOZS+St4mgLdsUbNuxxkt/qf
49fVvGIio6zyDf8yvRfU4iCTlEgkqMMDF1vcXL3pqs1Uz81tP3y7ua//4NyZIE7nZdCDn0AqhI1Q
SmweicWZA6j9yDRBAIB+aRY8bgde2kXOIxs1u/lXSi8d9HX+iQfonsJ83pp6HBN6QzO4DbRflFWN
lnR/5OkBqIa7BareaK4m+rfQsdjeQHfQFmruAyf33Z1bpexS3bjQpfrTATxpmLegdDfLwwUfQmNh
oaxLFUxPCslqhilBxNhGhB7rYM3cc0IhjVrOezo4SoX8C/G0zqq4oKpSWjHfKyygIEDDKPMpjjAn
IkhM0z93UeF7ZUU+zgW0MsmRtWLSdcVCGe3ahK0MIDg7q+mpCsUyHMRBW+dqDNiqAEV/vu0/DZw9
D45gvc6eqs0UEbEdcxGTWv/fbnWlhU1FN7BoP9m1LUl11tLPV2vfBknxUJ4FmIl0Df8G1SEIEO/k
86muFjLscQ7iLeZuGJi7RHI9HARuLghKGPVXanKWzYYHHgh6sXGuplPcf0XnNvrkr05EfaZxuY4q
CtVYs4w1UsyY+Pp1LINQavLkJKwmMzJCUz04G2WLx2kliMGpHttvh01PvN15I15taBMoF/l4TDpr
kJQoyU3BG68B+hr2rtqJhzYK6TQNuObWy5R14PxL+liFL0GGM75Wy5leYpYSiYtHeJTt2oGnxLHS
MrQb4AEYl3Jf4uFXKr+N8c47rQwxyW9l4zYmjsRSywm4ZZVaIvr/zgZX+/ZCLY57DrjphENqBqbr
64B3ZpjAYHYQom4hc7zILAkJaOQT8AkpmMCnKseB02fd37gYpN8/gT8gFsqxvZSlM6i72LZeY1oo
uc+axLv5q2729u8Ot5JluTAdn4pRrhFFBHuoQCDc6bfL3MsZjDW8qJ6CKir1+hNykeBFZm1FLp8l
dRBmzTctPssKtORMoQXHFtUkwQGS9DggRR1OVMGU7WN/HNm5ZpX/By3J1Y8fchJ9xGPdy/lJ06St
SEEuSA/4FYGfu3yiVurP2a5Nidrv+pELse9cfMOI2xMP8ybncq+fIY+QTuM1klPemrt8/Wn0kYTS
QrqyujI5eQQ8c9pWyowZR+w0mRH02yG4YxC9XOeNhRwqWwGjtR8+ZwRTHJUYAGWp9DFiXJPLS/ym
702iuZjmUjuQphkGuru4nU/P8yF8fTg+iWXilc4BDiFKk+Mpnsputmc5CUsz7kRY4idAfHj/nD+L
VoZxUH/KHYWLkmpjcVnHe3M+tZEmJOimMr2w+pGU1p9upJ47mluq3mwcCV4TpPgRP66fikLzgEFJ
vwfrwLhGSP/Xna2Al0PTFoYTsNdgicCSpME1UCU527rZpyKD8Ib15pSvxYrImCSnVuvJvuHyTDOk
OzmW8uLpwzDM0CEMOVUm38kVTN1czFwgTq6E6cr23a25QZwwLfXentC5Xb65IJAoIvlokkhNfylt
De8JkNdgjKwkJyE06AACJ5MN8gckeGcvO0Ul++AFjInQK2rSL82atSf5V1x22aQZXkHcA7m9lF+D
+TGxnZ4WnpsZCYWuLPjyGO9qebITvju7MJ1bWjoLMOkbMgBAgflTl8Llqt8RnaJMX8Q6WC6B0AMI
5Uwoj3bnkvCZ2VgaQFwTKMpUPPKW+vyV5LxsMjsdwyJkqEgf2IOKlnDn6v3h/kdOaUUdY1E3IDMr
q3l152GxAYqhpquPX9jcwUa1r5bFMLSTC9m6P29tKHylo7CAliovknzvy8ITQJfr5VoOm+a5pzb1
jwKV5+r4n7K1XD/1W0ai6XXiTx25ovADmrC5zhCc2wg+MSrdu2WoS6BI5JYOyEAMKTjrlZA3/vo6
Bx5x+FAOdgSG6nYvpe8Hb+xe4z0S7kcXuiEpMmItnFw3T7MiI8BxMCCYMij8QF+3OevqSE/BaROX
E6RhGX5rT3dzCCBnyd1HjFc3t9x2n2fBxwqKdeVBt9rdSbUxirJEu94YAbIqjCAkpnu+MFV3WJN3
+GKj2rKeQje8GHdyWvER42epc6H2R9n5FFLzBWbKslAFnO4O9hNpxjKYPOXErNUSoMAhBUMA/xMf
QgtKsp3Y+jKfiZp0xZS5gVVKh5tT1mkwW0x5lcf8Twdls2Tp+RzWuCf4X4lSRs6UnUF/8heaYzpD
kBW7OrTHXQFpWcgT59MNlUx/5X84Im+nW94AC6TEAeecxQBXE/UkdyGLWF527wnbZ5n4Ghj/Sg4p
9clBlWcFT6ypI43n0OoqpNDJfbgafONxQhhu1Dr/MTH8sjhlQyhq9jOZDHJa7x1nbn43Mm8KGFSa
70/9NV1sBNvGSdMUn3CD8LQjXQjL4gEK8Ku9DObcifkjmU4ef/T8qF7Vh1gALQSnGxKo7K+gUPjy
wby5sNshPVtMpe7Ju4LNCSOMwpWLvZ+fAjg/vndlinDiQJ32SLBuxslRpVd7IM7LNKvflXgLTOWT
ULPXaju2cNjZOzKahYBfQ4FQJRnZ3JYZ61RVrAHtO4SzNMswTEBgui7iLp8M9DXqZMxvroyS3BxE
nQeLFPUXJYvgDSUmkH8ZopuXhLAq/5uYhHKJ+uKsNE8ph8hfoNOwzoE8d/Q/AgileHgBvKL7UpfQ
513cTRW7Im75XGMbdvQM5+Z+jhD9AEX1VCHhAa1eUIO0R6taQ3dWYRfwLo/M3ad11kDil5f9Wq+R
jCHJNQI4W9/U9wGAyJXYAMdWISOvmIv+KP7IhlKYmFeo3P3/OyDPu6SqtHZbj4kqUny2PHNMWk48
jV7AZxoyCfjR70B9EVNWIAvZF1r8JEIeZ3Wm6Hu50feaSu7R72MOyXWs8smie9Lr0g6mq7jVBNta
qmPQbR3RLWGmotzQsJQWVvzlgext+1rTYbskNS5VlTF5bAds/7uJveqoZI5WVQaswol07T0zSfbM
uYu7UVk56/MMOPUbBERlghYbibn0nNg+IqMWUtd0TK9L+RMRKJl1zVOkp1Jq7KUTc+BWyyan5NmU
r1q3g1FmyfgHlqPCabT1WTJsly6rX5WqkndG2ZOIOBrq1hEyIT5wI6Wh82Mk8rPIsicj1bqX1kUm
+n83gTBu0Pz2xw59L33oEr1Ok4GA7QCHcyx8+kzPkoIBQHRn6uxLdAzbnnj1u9w7lY/P+8dX/9g4
29T5+2/0wTyGTpf21KQwC2HUoDLDgrpDXRkGA7/WAlFFR1+SuxotbAlX9PWQMKa2UuQNwNDqZ0Ss
AaHLvhWrcErAdEGMxDgCCSik6J0JG6KWq0c3/+lPJnvzkl4TWiJj7fulnuybZiZaNs50xGZxbiGI
UwkpNlwW2uR6khXGU8kJ3KWBiYKdT7lvZZNvZ3+cNptj6dITYjcevEGvad/Y06XJejhZlaUTMDUS
C3IcnF6Cx2/upmKDpOmaCDASWFjw62tENGhDLGlPs9H9t3Cb3+INF3Z0KYoLCGH+jicTBF1EwIGX
C1yPdLn6NK51ndnVdXBdDpoFgDE64BFx5GO+vvVmB9ZYTWdl4VBA6AbmbPQSiW9zb55EbyQcmBER
MkHZeeEXjSzEgA4kYj6XbV/jVzkNg5EftEc4hD2R3k0NRmr4xNg268HyFNljYAUybYA91Ps82jYA
QnSEQ1gwEUKL7rrPNRhCHhnnhVMzI+kw/S07WEivFWU9Jn5fwl7rhd64xb+SojocjPRUL4bLExnd
6tGYIPmON7qKO26+i2zcS8ndywNvIKHHs2Wv6Hs7GThJrjxhBbvf4c2rQ+inmMVVB+oVXd2/7vS3
zH8o2Y0lnqIfOZHifcBOODHEspQY9Ne8a+6HgBIDkKMrpqj1YkUIAVfQHz7YYR3taNhMcMHGlnyT
r1KTyZUDHjy4XBAewEh5hTtkfzPsOKGrlgDCwiCHBI6EUWMMS47bMWniVsFQX3/q2Q5nNtUxcs3b
x2kg7fuJpkOnndEc0JrLAMLFhBr9g0KQJzYLSb9CH/S1H7HEGSlAH8x4suo2J2jTlGQwS1cIaU8S
ylwsxf5iT5vkUMRrUeNjdUZYYX4fD08dHQVV86YS1imAT3FJVS9iZBFhVc1APhHp4/dVvm+VvAvW
BXOdkq4hT2Q0TqQE5bheghJCyLyHKSNu/wSGUdsazWorePsejClDzgfQ7YgwUF1yDXhmYAN8PFGt
Npd2EML3A+1XyX7nhUBTXGUy1uKDbcwdfQFUsZbYBNGk0lAExyRMvEEnmjd8X2mD//AgxldxrIzJ
GNLSbzErYxd5F4c7ye+gJFy+ZJU6kIbvNTQ33RfVu9GvSclDRp50KeZ802ivYU+AXDDVFsoHkCHS
w+H0SLcT2EvjUPrU0YzQ55LtjSGjKRTjJJnxp89RDtDdh4PsFSDMzgka3jMrtQMwKbdxVsJIZy4w
v1p/AMQD+BL6pbxn7HhUEl5Wg0XOrJt9QaW4PxekawTyLE2IeX9JrD33Z9M5zCdeNJ7Y440s50dy
HMJBUZgqe88mTrVxrv9AqYFlwFX0qVjYoPABGjgCHMZWeJfUtw1PHxhuE6LTq9ke6fK2s/GRsvsJ
uS/4HxVFLApFeBeY5s2JN0Eh03nEJkV00LZwxxJ8YsXPWh4AILKGdQrAQbZTleBHUCx7M3zSczHy
Nax8WtZ1klQTGy7xHcWi4S7mFHzKaGtLKDqNcImzv/foF6Nd3zZ/hknMvlDp0uHOySqFK5fZyEgc
w2VWSu8+r6pdPYhwILlsuB9ARfy7Dn9BcMMiJXSO+3wOmHtYPk1J9qySvorHOJdlQNLyZDeC2Z4x
Wigxp22kWm87J1LPfhn35xYv8/pMMOLXbI4gCcLR2/La8BxkmfZkyqW05yqEeAelUHHl9C8dl+eB
8vcHF1U96SAe7gnzbvWrLNCSEjJnRrdef2v2JRXh1xA1fXTJx30o5FTKT00vp1zSrSRwM1O2wZNe
4l13b6K8OW0mKNf3M/fOrN8cUVetLD4Sw+n5Cl/cipKccIKCHA35zNO/2RQ9581rug5N7DLMXo8d
ERL/3e9ZRWNa8RuzWTDwJZkmJuhtKTUgBMkQM0EZfKrVELMFi1YIZp8LSxJ8i4kgmAGl5O+YvLu3
GGVdjpnR//plz4Zk3wv8S6LAHTdLSIWecEg1aM3xJdbmQdpeL6tKN1KUHXTEvRoAv17ahzmqKgNX
HJcHWTDulyJcBuRyzDmaRVM6g7esqzfhyJaGVFqEZFY7KWSp7DUDLDgF3H2yUSQzUI/ZkJJAKeI2
lTNQ+wu+e6EPRFC1g1GJWcWRfZoYopymNAlwm1dUk+296OrYCfsvq3jd/PLbEK07+9+6O9RE0AcJ
VJW0OpWJKdj4OlnNMNbzRmDdzDUQIcVYVM0+ex9tUr441a9KiiEBQXwipAMJ6xfq5xlECqXay/BY
FSMCrZV97Ed5mU0VEgllXoClYInDqVhhPyIHWKrl2VtVWT/wzGScF0v6iUCnpEBfSvEIXdh3VfDJ
V2P8tqN8S5TdUerqvvYSBWgNTjWlUgxk9kEQ4Fg4oeq3sEwWsNvd3m1pP4YwvXV8UBASEN8uH0XC
A0xvxWK47cRQtVaDzEyEoCwNPnC+NLlSLk9hUFs6pwBSag7g0JmW7Eqv25yc1KqvOo3ZvKzZdXcR
8hfocm9Mhnp/P7gtK/Bk+6aHXOYPJxbu1x9cJM0kmNnsqyESPGSbNl4mM3X3EbUA9IeLqbJr4TXL
ekqS/+F17o+zVU/8+yNtqloK4RmRMYI6qM2oRcl6Nz6MziGp6TBsEG8zVvwTaRqQsgRGm1+gDSMc
X1d7ymks9hB+JGqefEXE02Il7OVkfufQrFGpR/YIIW3byOKVld+xUe030nV8bd53Qm4xg+FJxi3Q
cuSBrw3SVWbkdON9jrqWnApeG9CZFSf1ljXiju4w6m1hMFFRA6pmPrk0FaHbAOxxhHmrvh19eEo3
QQleM3vKEa2ML5FzzFKT73DUS4HM/klJmqu8/oAYdjAfbQtsXbEXC+5uJxcIDpL888s7d6iDP/Lk
wH/cQaFEO0Ll0cgB9aWRXEo8BwctDyQsQKRFz/WfCjq0MpYgHToS2SKBBn7y1bPPs9wjzhv9mfGq
nG5LNAsNWEAwEqnye//PGK+OomPkT1/bs3aYadHnmVo+htttV3TxDmt3gLCOdV6odqaVHwjw/cI+
IFdfs65vygyj0PiWTi/dwrjDACjlZLON2S7tOquF5aooFcEtb8WsBoXumIfvRbFiTAV1ypK5FFC9
j0NXyWahYDYAi2uZvUn2y/m+/2yU1OmHJI+Cg/vm6hWgiPK1u68Pp0DBDH80Ru2sSG4bGrsyKDMo
yoE9s6n45jIZNDthBus/tU/zz5j8IRjDLSfH2FlZQJOx7/+vcdimwrF6cj0YslJwMS49TuG6cz+J
OAHypdkFHY8SK8yDoOovqretmHoIRZ/MdP5nEifg/3XCnt/4HgLpYYddYwdgX8mNDvEv5QSJtfKx
roq91X/K30FPUOOw4ybP9PSKD+/D+60XgP2Wu7EF0WyZ9oNhhJu3bw5UTmC3h1+xXAyerulx557N
yU42KO8E3UCU1FWf2i2W+xj1DkRVhY7LV/FRc/SnXLq8N6ndbk0F9zyOhxvR8bAHORW6sr/nQDRf
oGZgN2v6Hj2xeoekIullJxYJf8AL3uA8JBSxpZIfDdMh0y5VRfKF4FlAMuxhh8elHuf+GqMPEjLT
PrT+VCzDY9fmUG4Q7/JFxm/WrFmbzwslVyOmOi7/hLoUzgKQH2ARRPqz7n5jhvffTaPtciAqRDCl
LDULvhOeWQDXL8h8/n1ib/DYqwuOU7MrwnxSriHkDbI0/6xpmXHWVEgXgF2XzssyF0aV2YNhep3p
uDa0kq5pcvKiMT2Jho60hM/1M0CNBarS3QEHJobyGBorWo0mSvsRYvcqbTK4YoqtdmnDdy/Tgrkp
cyjD4qqNJt65xj7hk9qnj4MGbwiJAsADgNBa/8EQAJZ+ZMvKOejBxy3Jpq+nXx6UuiZ/DuTNHWIZ
U3psdGjPnGnUeC7JuAtfOHr/r26UiFGHyAaXlUkmsJjYGOji95u3xO2ii29Gom3LVrEh6xz1aefA
sR2FfNwfJ4lA6dXZnCFlRUMrY1EKrCP9RRTs5BSQBj3yJ5Wkn1hhotzY9JHMrw/webAjZTIVUvNW
JaoXR4QwWx8lnkOa4xzvnSDL8h7t+9kXVBZDtoZ3wsf34+WYfAQotYzPyUM17ZB77iFqC52qc9uo
2oz99SJlBUBiYACSiwbktVDZ+FLg3c6/uw0iMVXWTz31kKaAeqXaUs+ltkAnZqsJE5dumHDl7eoW
R5K2LZ/mBE+MZnC+AvIaHw6vUUFUFVVhN6gQC7STsFDXor09ZV8jzwwv13tlBK6CCdL63DtltACt
wFF0DhhSsL5Ifb7FWe/1cKmDAkAClrBfbNOija5px24VV+wC7kwHJJvoGgw575FCVUXpOeqol+rv
Svf4Q5v+2SNgAu0/dV4UMhPcmJspx8LFkGYXCJPCHCJDqy9KBFtEoqzFWP97NM0syrs4+tI2rtUj
5VUvWhSapT989exARcrhiFxXQZW/wokSgvCc7FghnYGLjZmVxUcSfaFpM+CUlkLES6+/CfvjOGYo
VKGaVcungJCgvga4SEGDijrguA76/V6NBuHJF20QB+qAZWdMAKV/VjBzmY8lDRX1bVaYmrSwv46K
IB8H0p5EBZmq5lhTH8T2KLgFZ6ZjShDYiK+UhxVktjhSPCtpIeLu2zvXwXKPoXAZEtwlvdv3LkVS
kizYmH5AoTKNYFsNgVEQEtIbu0Yof4jbzYY9HKQ25J1nCXzT7sr91AGn6ZNV1kLyXlSmZEczirFs
WNJopHdPO6ynx0JQ8QDlmw/jEA+PF3xs0G0afyNvVhVv9wrFPeRvUlQmisy1BsIpzBXgB6D6Ka0p
g7s5hY6nUy0GC+J+ZkKg1QcfNuobEUDTynRlb7qYAV8bVTarSsKejtRHHWhts18m4hCfzNK/vWeX
hWVzpwbL96tbxVnVqTBnyC0/42Okmv6UO3NByFoSOGppdJKhcCxXnX4IzEtNvAbnSsgM1+rD37zH
pb2zellLwTR/Fhem+v1UHCv6Kykv4p5Hu05GWy/KFGEQ/zEpIqy0HtbCUxODLiBa1GZpQOzkUi7/
hWh6FmWIraMf/lClWdfFkM9YT874IJ9UYVWHSm/ynSA2U4Y9Irb0IviLz86P6lh4aer1GsFFf0XN
d5MjhTYlsBOKCFe3TE7FkxZqzXAE3GDm4jQtWeZTTtfu/CvZMrr1xCXRISleWp8nMl3TnwiyYXeF
90fYg0qUSGsKpQU5TOd1wQJF/BIR6uwJRNyBmz0VLbapPhu9M9o/KLIKr9LqIvLaipfPkQ1KCFte
HQB/TaZbHUogG7i16JlCoTyEf10W7UIgdshVOKWOvDuzeqgnMKb09QeD5i6ckHWyD2ImkbopaHxD
z0Tb2PYnJ3d2T1cW4FpV9c28C6puhp2Q0G7+/Tk0bCYqUW5QW5ldXDn8TGARjTFXR7mHa60JZlLE
7+neV4fP5xUKoorWDExFXsKplNpRzwVL2Jn3JeRV1Y9E9EKLNVKk7ubs4ZckyInPmPLHC1SLhF7R
8KzQEKdXHlj80T90nF8eBB/qEPDOKHJQnJG5bm608wyYoKnaf7ASH+7PYgBKYRUA8fV1BR8WLrQ5
DwQGT+nYtZF1acKsiMWT7id3XyGwVJEu4sWuhCgggrJApR1luvCNqBwx5NUtK5s0W6YCw6IqNTZk
IiDo3ArQJ5q/ecNNWRYxOMbHDj+v4GpYY+ttSwXL3biOZRbZNPxoVN+Tqnh6SLap6rCejWYUQLMv
Oc7uxeZ8HhCVdQ4pGGSMpJ6C7JHJ5+ppYSr12Jzi7iNXoYfJi/JEBfvTcDnK2vbCMzsjpIR5KbpV
dQwPU1vwKSJgju6Eu8HCrvFQyG/SOSct9IKpaxr3VyjJMKfMAi5q+FISIORqWkmio1gic3CDh9nS
jr9jwkIhBXzRlV8LOzHHw3NVfX6GlRsiFSWX/SpBBdU+pvcGvhuJersdg75pBRC4eKvSwJXu+2qJ
SgyOYU9eNoVyJFcDm2IualHXog8wS6H42myakda7TpVVPQ0Uso/+dpHydcvV+V/H0VCC6h9PVaqa
6TbkSncGq37g4ZI8RckYW/w2+6rA4qyzceISUCH3i+Ag5RDETYSwU69GPJUBRKtESDfo9D/2i6+Z
34pKwgdoqYa/3pzax4L7uLA8qWbVL6SrIRUpuOyyfINtVUjwM+9gXBDd3kXtSnBJwMoMiV1U9Gab
KMNXarYbegW2VBHnZuQpMBi720l8eESyKIn7ksAVjfRoL1FfgHEYG7qP/AcgkkYrUmeDGXmSnpLk
W/ijTGvpA12xfqIwkIoLOjybnh72XpkHibN6lWvbFYsIQxUGvoI9YmEY3NoenrhagHrlI5bqHcyg
oLx01zt2neie3F6gLlacihJiWoOkuCPdX6Ta/hbmyQDVJGXwmXmUVtRkCcRr9jXRc5Sxz3GzoHXa
1W0Dfob5JxswWCF0ZrdfSDRvwKEJKXPzlp3Dgz6a4oC/axH6S+zs1CUKov4xpySaYC+8SciquTKP
Bw3qvcScd6wigGbZgzbbUuHxq5jrA61+2ksdxZsGBY7Adr2ztGFYrhvXiDAkQEhWujLAPFH/Adrf
SHplEAleuUZCfxSAoRF2+xRRAWhmK+7ajFtL8niCh/WkuzCWO5GgXaIRld9VeP9JYX5F3y9TS+Sq
RTE5EynlP4pbX/topfELeu9McPxhWFDTckqkU2leafW3z9PY2yMc5xEJK1J2ZVmzdEcpinDJfCoV
vx/3rs1GC3VtnxB1XeMlonOdwH6CuNVHmkeRjSh0Z1h0cUutwErI2d9o+oViPtkkiyH3Pw9+g0f4
ierPSc0Jq7QTVBOUIjvVJko/0JpcefbsoCCWnqZtk9pPUB5m+bZecRIcqbee3Z3o/DSSsCEoAqTy
kYEIlFzXq6vYykZixj1bolYaP2XO/dctDL3WzY+iuJAsweJHz9u+KW2M6JNCd7QUzGgZakpwBaKs
x40QrviIOKfq0vXfdAN9LSyeKO6jx21jvWXLJKm3Wc/v6ge6+l13B+qA3pec2W03CDZslwpAf0CA
xKSsV/DRJLPTY/uqYl5bmWbB9/n0DL/Pv8Q/FVwen3XQ/Aq2Ki2coAJkMnkPIoGeP6qUp7n+jbKw
h0QV7NJg7N+pExwGVulZ1n3GjaRmZy45xfyqgHlKDRLvK3W1a/9HCA54d/InD81YqivawbZCDIWO
RjfOV05tF3Fy+xAl/O8GapJ+MqB4X1jmy4Bk8I5zDkHuQbY4VjDLNoeZC3IaXi9efxiWYXv8M6xr
LxoUPHJNjI4H1ulSc2YLi5UPaHVUnVhQCt4vBrAS0Bv992BiPPjbA7UF48zD/gWtBQaGMinfkdRF
1MXTI2nx47kq0IzxKtnZpTIsp041meSA09KMmFyPjXsbw6r3e4qcWZgrjdL9gW1YiUTUcvevyR2G
dG0HW75Dub33sLNspgDkDBTKr8lI+2KRmft/V7JFp6O1ObH6YsPdGltF0iVEsUldarz1JNeSGB83
Y3uQ+/3JXHxwnlz15I7Bhm3y92XGNZYJD1MzkgIcSzVGQrcNQ1v+vyahG55F3LB3Aa8odSjfxQHg
efrMc8y5FccC3o97KZHsTuC+QMtk2ofUlR2qOP56W5SWrarbfACG2N68S+s7cxuNSbKdYUaU+FvZ
xqb/ZyPsNfThQmEjqj+jXee9FjD4/8HNQFUvlKbzKhIV5ry+TcLvZ+gwiAtBdYcnJ5NlwZqnUdBl
w+WxK1+xyyj9tCK0Jg9vQ9s+5MXKsl6pzzJb4JVk2uQ226xjmF9YnCEXv1180+W6vWkd8FDoD0Vv
TWdgvq/oSQm27gGJSKCKF6YTFj/tzuem7eON430MNt7T7c+8FjvbXFDHRnJg8PcqCiMHnjeY5t3Z
T0PSqluEM4tS1s969IpRlY5NlIQTVAPktJWFbT2aL3ORWaA4Du5ioQeWFjrei/PnG+nK6jDC22xU
AbZQvMNtdgzs9MKqXD8cJ4k6wBFrR52tHxM2Y15BvHB+Oq0feVkEGKUzBMrOp8U3ga3PQbR4AMRv
fLY/t6p8KF0KANydNdJiNx6ne5pswze0V8yt7EcyiwZRrocFO49kUq64G8GV4m1RuZ0EDwfh9A6B
ygHD7FdTwxaa7CMFPDDtiqnL+wlMpSyRfgfAdqOakH++h+DqheGZmw4NeaIZabQLZUTThqCCq6NF
qzikL9kojUBGzXFbz1mdu3EXPWhfyJniLqAHAzDXRSMHB6EszFucBtu5EMfo133XFP3OA7SyrNKj
lMrqmduHtqaD7RQUyNMq0BzjGg8UmRdXi5Swf0zRANZYs+7bGFKTbB4ivukzGekpOvcmNZcIVf1S
6xW8VSgKL/lhJBBflvuJmW+rZ8XlHJGEigBaaoUZR79126XAaezRUdOkmfJBpAFeViVanbPzhUFI
R4uKCr3hDyewi3nt4GvM3KhNxqTesyfJ27xRZuQYNIAY04aMz9qjEBlx6gNHmhRzAncMugdArgHi
Jtfq3UVoYyuwW57P+ljRakAkqqOpvf//4I+7V87ExzEgG6Av8Y6rTs5uX5gUrFTu+4CfwH9v6exd
tHKXekrhnRN7pOafoFBDkxT6digH91ofxuqC48qgMNzuef0AU6kB3OURwTW7qkUvjy9jXDfwdgtN
wSJl5QU9Olkntq+1fiuyo+S7xJYhu/JaEIlo2igu6uwIQuJ+beHxMbdv6nFUHImaIOUDwylD90NR
epeG7rSC76FPIborbxEh7JiecT4Ha3NXuDtTfrBzY4tSssh4dbKChw9TWkDlQc4WMPajs3USps/j
voeCbC0/JebLWd5V2r9JDropdZ/f3SHJ6pKq+EEQGPB4PHvp4OWu+3mk8TYljpyjXHktVLoFo5cU
qXznqNSkRwPSCJvooxU+rvYFdowyXydiB32CCccXK9aUfZMt+1sB7Q0gVJpg/fI1PmRksz4aD/1V
WzpzLcUONV0nAVkgXfZZdnN/29FsEsFYMoR3MltvXExCZUHb5k6GIwB66u8sZ7glaC9G2eTHXu/w
LKIYPVodlFT20nmgSzzahTjAvd4Zby++bl0oWzqzgvnp7SMFh2B2KdCGjgl9DBVs91k0AgXOL6nL
yRJgZkUjuWhGD9h31DOi8f5amPtsYDqncn8QQv44Fp0hlw6/7sXgbdCZ64ifxA4g3p9Vdxir3tEf
vsxUr2SaF477L4hZsFCJivmB9rBMuSfMjwGQroVZ38lLH2OSktJjTvgv6Vrt7czvc1ePr/l66Zic
qkOu593IbgnqclqOBrBHweusAmv083XCs3FANRwUJ05WIZ9/b9HRqMjvX11M8oe9VhGBFiODBgbt
o6E+IReGXQidZ7lZ8+LWonfo5xblYlpZUBct2U0Ms6rniFzyvC68iFs8koloPgLKsPaM8l2tX+/O
KcQxt2Lk11J4K6hY/OwxlldluWSIcmB8cVuT2wsgV6optVn1foWScpbUh+Mzf1w7uXc0SzxOY5Ej
dRWzHTp0ZWGe0vIPfaysSKk0JeDZdI8J4723Tutx3eFVLioGdmVldMXC/arl+a1cxyFwDbxCTKs/
fl2SpzPOjntctlFyvpkpeY8UQ80WVfPVzyfLJziTOZPVggsw9rQXEoy4Pic9CHi/eJIt7yOgRhQo
MvhdIeei9Kb0MfQXmJs23TK8SKo6j9KRYCVG8cMETuWnZyFJyCJrnnKKsdJB/oyK+ajC2NKR4IAy
eRb3imLjD6cHBJ/czmDvfb/7o71ecwLRGpNXrNvru6qxDe+w7D6AMZKjfdK8/4uEfUGV7r3fYhth
+RsqnRr750lnHF306vyEvquWq7QX9htReyd4HAcldlRB0qO2xtYUe7XNTMforUK+n+oaJuDnJkMH
w5lJCASE2UVPRlfx4ajijxpsQ9B13EaEzoQugYxK5JqI/Rtm/h3gtaa8hF9xe8GIZY5GFDlHYjfv
sXaKHVF8HhXHTgbUoZHoklqDM9+5Wi08IMwGEfraXqPA+2Mzh2ubgddwicYd5tsjsfP+vAdRR5EP
9GwgymwQHfaSa1XbwCi0v6YU0bezPRfDny6ql9xZ7zmVcdT5/OJsGD0bBn0K5Qq25FMQkw4r/98q
V3eRDkYn+Zgs9f2gV9o13gouJ5V7Ztm9eqAkgn23N6bb7DCeqmwZxNd9WEAwS7ia3Q49fqxsOG8n
sdBFuZvtXkU6DfxrZ8EOcHRLMDOKK2hoGsKrWQ5KPEfxLI82JK5amTJX+udnqB81/Byco5FLBy3H
U4/BYZBS8BfFGT1fBs1l69oNdiS7C2jv2MWO+t8m6pfIhoBYOwfz48m206y130Aau9G4otoFY0Qn
3SQKvFHoMQfT7FEik9rgNSxfB0BmKeLxymYaCRhhdGvpaCtOhGz1K4/iYZOXwIV7WKmpug8Sp0fs
itVEBoS2MylftsLMq94Raoz1gvjVUp79Yg2e/EBJdpKbxNzP9nkOhX0eKvSyOJ6Q9iBO1bF1uMs/
I7JXTCnlbmLQSKpO398kIoIRoYjehomyQAvPJgMTss5En8i3ZNvx69jWCFMaZ2IoJY03r9e+086Q
6xieBMPK0WVam7+cKjd/cQYENS5jjWVCSid1v9I4j43+OgggruuHEm/ocgaJwiXIJvfExbZ04MOy
Ns+IvFzv8o1yXUfX3RWQ9NiacyErcolvjjYE9XyQesg2Cvvb+5wt6nda4nbdDN+eD83CQfJxRG7e
ow9+rfmxjHwtkXlh4iHdwfhZ+ED2NK+y7LA4UgeedsB2F/8ZWSKqtcgp3Pe+Emq29fBkCnNfKPr/
4tN0nwlJd1+tWErYtuzIufKSBVS/qfG1WYQRb6O5n50vxqA5r9PoY1/ZiNLiCm6KUF/au8LtD+kd
pj3eCBRWliUp9a+8SH8tzFa96bRUg+8V/QAzw2v+yT/ebfAKZAwwbS2rER0OS6JR0GBRg6Gkmfye
8LyXzq1iLd4E4iqERWwV8ebn2F/6TH7g3TyLo6fd/8Lc6Hc3+6prQcxkHhGQ0U7IZZRJhtkWk45b
3X9UI/1MDsU2im08mDvd9K5dG+xQS02kL7aCnV3GXsQlyT33bf8QP7Xeq4rDLcIPmpKcYOtE9mjr
y0/EzPMPDxxNSkzd5IZaFXERQvfXW074/vIy+rktu9IwrcwkfdtDmUlEeT2VR2esKy9wz8Fy7vtI
il0DZx8y6sLS0cYPLJTXobT3oYeidVnrrK+C8ZctLgowSomoXVVJHR3Tz6dZGfy+k2fAnfwJWDk/
RyHd5Jo7W4H49VCE5kbhw6LY4xbZQak4xTiAQzitt8t06fOWM8mX3vKQ4J9N1OTAoGdWOQw+NsfL
gYoa9x+T8xUSw0dPP/1vZYgJEG9ZnBS5XVQeolrK9YjvIdUrg8GcSu7tRrGg7fW0i1BmfUY7cj4B
HaoyYn0p9DEvbcls9Qs20xEr22qc9icPQW1eqOcalNPfy6HBYYAY0t0QTFBEcfVvyKmjyenc47em
aQLEabRkv/6OlY+hVON4G44OVM/lz0RO8ZBBkzxg3tAvudGhBInHHjnLjWOUq730Rn6eYV0DWlIk
8fagxJC+qp8UUBeFVg6KGwZkPEVKFCx60K6rmfciGZTkQE+PpPHrXEKYPXDHHoZG/V1brvznjG2o
lxzHAM4v1R4AVI5E5BMeConFxvgPp0ajMLlEdJJ0mweN0AZbGmHqsyCm/L5dqwamyDKFS+jybe3l
0r54B/xECL+s6XNRTzg0U1hminrLshQMPPATwWr+APLqE9QNBuGp1cLmtoHwlHFLzNQG+ZP+85Ru
jrvbhKSIuHBmE+uOwHGztCF9BI3r4UW6KlPzChU6SGoVO9TPPXLGlZLZEY117+sxz469HoKY52I/
nSPFX94Li+t9IJKxtqhd5g8iXLJAY6wIcrqyUBswJNFFRHbxNr/1ht1YvL+3QvTgfPra6j+EDIEA
Zxl/g2rXpJwdA9atQ77ZzV2jRqgu29k9Fs+QxOjMjClSW6eYjCIBkRaf3heQGFqQAInjXgjeyEc+
YyapGaNWcuvcwglRGP2dM/XiBznbreIjDzW5k08/V4LuJRRwuNOFZs3YMDMIr8y/q6izkzp9/IXV
ut2ptGVsY06Z4t8iRnuigtansovLmgqx+watrmLOF1q7CwxWZ84wcgI4aiJDbwLNbPuSOAWM0w9C
T9qt+AI6FsfIVv2LvCrOstQl3khE5AEbUhlPhzws0lDWdKyu2xR36FE+WRyeZFnT2L8rxaP9883m
kDueS44AJuZxSVNZr8y9gn4fbLuKMMiuW9E8tsEyUq5d0ZsX1j/SlLYPsy8QHn8AXxwLFEs0uHoQ
/fDg8rg4yz+IVP/9ManpSRlMnTExtMUsr05SUi4STiAeqdhNqbBXGtIpqSDrwNxCDiJmXDtwlwk4
VHd76IReBFdMEq8m0oYLYxawJAoDnvXl5ETuGsiFI4mDzcCkqCRnp5370jP9WYU7z9W8vHMOWOt0
PIJOVGNI9ovvrXILr2w/NIeAK04GVAFrDA1Cb8+mpd69Qkj98QdJExOsgprqBtdHD7Ic+yE8QaDy
a8caJOWcCd0UYrS2rSGyCA9cle6UDWHHomCNmNgQZxCH8nN2xPduAqnu+pqfNv066Tbz1siraP4N
6fC91TPTTmFFvdFLCCrwVDOnZ8vWbA7732hTARd7n5w1dle9aZNhFaDxdMWNIwGWw89xp8Jc3ugx
PPNnL9r7mfL6J7neIxX33AOTgInXPVEy4zCHnzZbF1Y6oY5tGeuqO1lZMZqijtFCEXiQP27lnkOg
DTDisgsefvlYPXeMh1Wn3NO7UA9NwNAxiT8YRFEAJbWDJqYGu5XXdoJpwBNKgkhRh5fDDyp6NcFu
2DkkvvPntsKRlNNcWj9ra79e27oYJ6OFhUsfnOgCCH0XMrtYlUKDWITeVEemtT8qOgDis8UWH2VG
pZEYraM8Ll/UnD+wu0pLLW8B0FvejH+wYNQ81KAxKmZiGHxFTtHB7SENO2iUrrEHcZ3PW+r6KNvQ
m/w3xHcpQ01qYwrKNeuBbCGXGlTjGTi8pr3fqTsDRAhgB4O1XjnIMZJ4ozHqdH2GjAxc+l5iNMru
M2sf7zJR2DL9IxTC2e0sDo9aN634Ainpb8lE46kLtUedp497uiik5XTkKJjFoFGR/eVGCLP0B6iV
RIBMFhlRS/LeboVT26CLXsiUrfjm5gYIiCvXNNFeejb5G6lItX+8qGj1b9V9FLVdCCdXmOe0ttHJ
J3w0WIfnn7LV7Ig3AgpO+HwmNeh1+/79LKR3df5i5mXcGYK1LIxATBSmbAbiUxOOIxXNO+FyKMls
s4ZZQbAwvzx1vISMO2STkNn5F+VmbejHn4yaQRIe0l6CSTjNN1BbJga8eC8rpluV2njGhXJlos8y
Nj0QNVe1GH4SWiA/qVoCRXA3/CzdrqvAcR0bQHHrh+Dy5OfbH0fnPgpEvppkmPfCetUbKI+tV/++
3y4v5mVlXXxxU68xhS31ItLp7cKVl2mjON+gTTokbNNSZJkxfjA6N3ZEuwadMY7AHLB6+EWRtoFw
Pwcf6yb5n+Srq7G7kmRIzn0H6EKP7XYcq6RRIHiAfnUbxOAVJHw78UxCh6vRkOLo354lH7IjOrOH
NJOx0T2TSz7/+1bPk7l0mW7/4YxCK2alWplr2d1b20Mhigugaxk1vm5ZHkK8ZxI6mL+iFzY+98IS
aVPKAQxuhc8NvwoIBc6nrCyx/mpgzPTpWckcgvVwW5soXWlnvBf41/OuQBOsYR5wcYUsFHgpWSsh
AiYt48zNtAwdXoJQI84/rAJcfeYtBylOpfZvenGpnq7rQ1YwrdYmvkS1UOPaNYK558vRHr4u7KZh
ZMrpS0nCc2EfbOyGLjuk37rTj1jbN7lFtMwePZhApLmWABcRY7qyU8tdQem2JaCawxtf59w7T2um
wLUYzYQ19YXgTYqP3bcvhH2RQCScTCso5OHQm2i7fK43UQpIUpBNcX+Ut6E8Xny9Crtt4NSQtYKQ
vuxwyaqSkJuq09TBdfUWIl6TVCIV1XbRYkHV10LK7urQKYTKZSvIr3rZ8Ps+beApQgK0fhw9WySk
c3lBAfLT93CCJq+3tmZfHO65DaONjynQJFu7CDJQj/UwAA5s4AJgHLGmywbr0Bj9RXHfXnHtHD3X
MNhWIDgmtmO1D8HEsn9C9HBNXIArHqvJ3r2rWUCCfsO5Cu1aeDH/0cP/7qMoMMiLpYv26RXF6AAr
MlwHKGOCPK2v0WH6Mh57phERBUk6UQlgMiyfZ9sgUpJ+KzUaEhKn9TgyL8txUAoXAIRdj9/iaplL
UrmnROAH+1NdhOX6zD+aUdE4yOAsSlccdUVQfpDjE5insimJlLcMOPcVfXc6GoCOrJfMZ/YQUui8
jPQUrRk+hJp+1g+vNbMXx+tZSY7UeDc1F2JF14msxYMPN0mPh7k4PJVHOhVfsth4MLuHM2Mpabq/
80/pIpMN+Ny3humB5834xszY8TmZ9/r7MK3kzMr8pKJAwzAliVm1cFMpMBXLax9VXtOOwpfdl9OQ
8+TBBMLiOtfPF6Z+lBuErPmUFPv1omdttz4ig6iBqHZdZ4g5d1TSEFH1zwiCCCllm3R4qlTdB2zo
Vb+oSq5uMhIhTwIVaCrNTwuWG246R4n9xBRois1TTPMoGn5/DjHt4426ndYRY8YtRm3uPoctpVSw
S2rL2goW0NYAEKOEMo6EY2iObL/86g4etF9Zsl7JhAOF7iVHiPkA+2KrmBpm3zAnO6AB9Aokmwei
X+E2tbQ6YBwrLRVPRVR/PhNKPzcxPdHPu9yDhnlSxxgN3Z5go1hn5kv6uLbvpbPOrOB7GZT4tR++
XxveKXmPawXxDGZqwczmbFimu4CsMrGUHIwKt4EMwp4teM/GdxrfGZkdLYCjhU/ie3pLe/gBuDJZ
O/cqsOYcS8aNH0k+P+0f1BXK5Y768RygpYfHjkmiFswmca+oZ77Qgf6x0yoo6vazP5+6IIqNdu/u
8QpgqS55KPppheftoBkI95eCy+OZYVPmJ9Py0r2h0z5upZu1dotBiCtjPLr3T2k5l2q+fhGk1LPM
dJ09+rqkE9AXPDw185Tdo16dNgMar7ctAmuNNuuunwV5gz3Vo6BzEzKLeaxj0b1UQSr6lMfmZZo0
g7Pky1PrNIoaMDeVt1sFHdNx2OyBxSmQkH9rS5Wz5o+/pAVvABtp0+FdjI5DEZM7+ikW3TbPhrh/
P/2hBxFvTNmFUHy4nwO46AazROrP8eLY8wt6D+Rwg3LQLJhApstrB0c/IIUsdKIiLySdjVhMuBqp
9J2ECgs2mPEbczxgTRmuWv8zFZJrWmgDSWqZxBVAlVmhsF7ujj2+xRoF74HCcJyr3WXE7aWJwNmA
MdoxsLPf37wYh87tLS53jQ2x6lpizT+UGWudGGYhbSGm+Zr8WvgG0a1jSM4buj9VlFBPgYI2OIJ3
dQ8BvWU9BRAv4dyUCgxMfXx0F9NUSGK4/xJtdnoQWuY5MzZ0dz8dGgAe3sXhxk/RnkdSq4H6Y+ZJ
s5SsAw6QW39FbbeXb6vlQJeFcK+ZpTxwRNfXfcEkcpLB9rft7wycNJBFL4volJTTPeW2GCIcIzBm
zT4rKXwZ5GuohdVxKMvcgS1Y0D8fGxbdCMRzfusuGWk1PBncGniI8l9/KbIoDbjDtN6Q0/AnEIF7
dNflFbLtVeRtzG6sj+wvuXmUV3OmiJa4Uv8tr17Youio8zZkNZroAbbA2OlpK6VilbV+5dDD7Uxg
cTecHvGYugVIhCha8TFc7hL0P5XGeiPZWjIa9/218tnozj/K15paUmkcaxgPk4gi0u2x8EFZWInc
9OqHX3GaD5uwuiewganCB7OC3OJGgZXZSpWkOSP63rFExWCRaW4DHLaEtA4s4WcuAAik/DWdMTJA
6OqYGIrQHLKzKvtQccgqfl+0uEhZ3uNK+TL0PJNksjzWCyO3MZUv9bE2Go5uUzVdeVkHoEmSgOvw
9/I7yXOvEOK5BnF6WsYuf8PCK8IxU+rB5LUMmqRRLhUxOIxXtess0YrXPKRJ4Gv1PBuxM8bl7dOD
UIZkkgEdxg+F12/cvl+2jZUzZfFV6vBfIWurzfogK+vHkcApzKWiyg2tLc+hfrMyf39ocdg1AFvs
ElYsP0oeUfhsY8maNdlilIgsuI5SttceQrMxDIxsXN3Bp4uifeJDMlGHGlyBDpqCwjP9YlcvK+bP
L2JPiXGer1fO3I3aWShZM8Aw9IhaNcxi1jQ1IuiJWlrhXl1zxbwA16l5DzJcLVzWtCxRo+/YKUQR
zWZLPrIl3VN2DeLTZnBeOKJ9YyB3ojwZ0+zC53knQhtxTjiyYtRWOkZEqWIjP7G7AbopfulUH8u0
AN2xAXfWjsQMfJvvBmMfDbajktt6PuANv6bCBzQ/wAFWkruGY6Mp45pyDX8dk29v4vNvKtnOt/lN
PZ0MV1T/N5YboRGfxOXu0BY18tgdMMysIh1o2vd/GPQoU5MjiDZ/XWydKDNGV/hoUy+xXI5rpiee
oyzUpjOXogVz5MjXfzY2IgAUJ4FVH8ssmk+XaUTAGRhXy2o1NqzyP4RLQyiVlz/15bjmK+B6syo6
z4DOiruBWcnC02kc6Wpw/1qf4RRZUP/mrtybCw5nMlEZvf8mmZpwzWNJMOaAHkIHH12vPDirXJgO
q6O5NN9Yi1SnKjzyAXuWlv9uSsiXdovEnYjJNxylgFg9Y9v1/tP2xf/gHjIswVhb1dpYyN8ylC+w
yvzmeqp7PHRLkks6MFHC412wxh40Oc1Tz81QnOTZQTRbjBJ7/Uf1Xrn3EjbIxogH3tQ3uRgOITxA
2MNNywep5mJm7uvoSCpLMoxUDzMFGxNl7GD7jcCW8TvF37YiiaiyufUiz1G6aWAAQOC/W1vlPNZn
u4tNHcXS+7saeLIQY1W6ENAXEtzhQi15wWPqfQS/IhdSj2xacN90QhHLRV2lfUtQI90JUSOCZwAf
tkjwx3/9hh2o9z1HXMC7KBg9p1X7OCZkEwLEuCIQZo0wZ2IZHFGp6zp4dOcQq/x1GrAPShm5QqI0
K8FlAA8OWnTU8ucHSS98/FQIbozPOX1NdzmqDzILribE/aU5uNhvXWl9N85fqztQY+kvJnBG6BAo
n8FxbLuq6JsrPDxPnjLQYGXyFIMU+Ar6cjyQWCKD7omg2GkqiZ9rpi0NfGREPd9KtXdkIIZ5ceZ7
DS1Dw7iGRUFIfZ6DdafIK87L3zsNX3Dd7/EEopY7Fe9VFMZ6xOdXo0p7qh+gWR0hU/jVxinJy1mR
z96ETwZFhFxaBVYuiyxzZTtkxLpyznWc57v7xTqv9F7QxwXGAuAEk+vmzGWH9u7UVQGlSi5IvsFJ
OgJZzla0U43lQTiGBuu1DqNC1vaTBnxqqYS6b9xdtmF/6fW6GLPDLyZlhguTMNKx2u2myQWNj4uq
6s/W8/N1A7QT038t+vaJLJ+DJKcZsV6UOWkT8rI2+Jv90IsMOqsjn+AGch8UMYAFlRA03ZTKSJ28
m+2vQMDtr01b+GB+4zqOwbs2EUWvuOb+xnEWYQXXfQycixQBvtaZNku2XTY5/fWQZZbRM2cXpfwV
Mq+4G/kD8oFuFmXTAO5vzMdMmWDgBNek5mgnP33bhY0F8cR8DwgtXS0yCJ2N78xOUbmmw6h654IM
xdNtMOJXaR6VkqCltq9oNIgHoCVnLKgVm6K/TTBZnm5u77OIX1FkboSskpnsHD2sIc6EC/Oc5vDq
f6gXVGFh40piAlYRzFeraUUjakiq3jjrtgzS59qfftTm72Yk4KkiaHtIG+GJkJUeYkVwbx2sYrXQ
PXCss0VHfaWhioIMvhKlcWwR8Qi5Q7lWTBQe8w2k4Q1c+urmqjpSLaMB5Q4HrMFuquQMR4XOBXnE
mcL3B0GZ+34VgW8GnvsAaab8WAkwUW8T8pPkciP3rYGKjkuriIYNwYgklUWTAaUiMDe6VCObx+XO
rrPPQagBZwBVH3QSypTUIF12w7KJZfA0YnaU8mqz3bALy1Xuyu3DCBcabtzWlNQd/JgBQS/u+kd7
Aox0LzkVXhTAHahE8Q9CERWEEANjeYZdntxat6GlqCWTwis1ioDuphteIyCTF0uUgkYiaMFgFgpt
bG31+vxHRFlwDGDBn/k/QRKLAWl0XeTTR3aHF7dncU6n1Y2ZJrVJk7IRiVB6UYQMts5hgMOmXFrZ
Pyueb30d+PmilLA7wHrJw8sVW4sE/cKVOkK+r7qOaCZedQ8X3lIi2E0IWcUn0R76NtfwDuMZJ9Ey
HDHnD0lp000z+bdbwR0SL8VOql3cQgjmCUL8WbGOHEP0/M+NgJU6d9j61tiMXtt9kDH9YyazqL3y
Esjwy/gdvpU3iGuJDnIiiFR0v9+gvyhVWrI8EutozXpnWf8LTRkYVFx09p0XQPzkYLAc1P1SucMb
2L+DazjD/cf/HHvCkzqu4wv3/ZyV6+lfDGe5D8aWpeSF4RD+nwvGGZRI94KQq4x1whf4u/pq/Z8B
SiLSP1+hxYrlQiHOXjQUTaAKRjmLbHyrAejAHJ7jG8sZ7fEfyGIgiMKZU/tXm3cWGz0AKq0eZb/I
FxQMSGOQzccQsKxcnDIOi6U4knq8NpOKopEAIwQ2HHVrQK5rmcdDr27Uip6KWNWoBEL2k3AaAZKg
eQS4GxBNoY/dhN5bhi4zRhtnLeyi6gc+g+a4fVqSmTIxAHXLpsB2QJOceff1qar+zheTZCrOcxzg
WhYkyfFWd0+j1EQoFSyiy8ha+/q1oQg/rQMFcGiVZXcj/o+UKHM0G2t6BnZRhbNyHUJECSGuqn0t
SdmcXqPmbcssd6tvR9MmTvkGcqURCm/yydz6BDm/ANHHyEPAQ0lc/NWWwoBSxcCSTEWmiHbC/PAQ
xCXiarfMrduT/PaP4m/Je3Q2QnnPIqI7BNIkTlEq76hVFOwO9KfbVI3TSm2ZazeKBaTmsO5I03sc
QpVMiONB87LAwBeMINphoUDfXrtcqRuSedJsarWcjvwoySyV6UKRao82+lniqaT0Wnj54gVi0KKj
WsUjOwKmp2a8xq4Twfyq/YD6Wys8oaFV0FqFD1/qQUUM9zrzR6Wd/O4c5eSmz+k7Ap+j2nDfyzhk
9tOW2zhLB+JYSJdDSrNWHWaap+b3b0ePsT7CjUKQtzSw56fBqUEjgGdtfHhi1FO5fJs9PQ7q5/mE
T0+dN70WdNNX0xqUeIqma+XLg9ut2EjyNm4xqBDO6vLgjKVPXcWYX6dtZ1GaBtxhPUxA6rL3Iw4i
v3umaxG6oWeGKYw3RF4ww0hXj6wPeP0KMtPFcg+xEtsxPXscqf7dqonCXlN4o5d6VI7IsqeKlYoQ
S3Hjr8/7194OroWik1h9ERqhokRsownc1nNDd+OjHmaLPl2OXDu2NmJdM6O9bCTSNbQohCnZ3rEo
h71P5SCnLaofFEVtteVdCd0QG7aCzmqBwOjNd1/+Ua/xoOw+CODuoM9ASU4ndWS47rWv4lXmhlE+
a4XEIHAYjScJxXs3d/7A+NfsIdZtqkJUa10rcwQ2lVALulJk3iLzC8EkwlH33tpWYue1CLNEz0jk
kc9jjmDJjFDpbeQ67Oc3ywKu4HkGL+7RTLtaojUa7LmC4UDDayu9fkoxXp3BBpeCaBqUvz9l47rd
aYLKfTtUENJkJ/uEI5f/7lluEEeeF95xQyE0NbPgKeNk68zCiG7xsUehRjkUGzMpouoJ1/j1DqHh
u+jtsUGPr3oz7/cdTtj18v9VpDnwIktIfRbKsXpmSTITiRC6oWOiTiCr23VqM6QH73Gqf4gvIkGZ
5u3WxLVBY0jUH53KnGE9lVX2S5giw9ogUYNNXp1ZeRfzTSMPKYZJpLZ7cloq95slmMYOo+QQOaHD
hOruAHXpmGU0H5frVfJ7JYOJFJ0Inhw3S9GVlBo3rTTVxZq/hlCdGpGEFhAYhBVFxMn7LSCanVp5
a/GDr8dxZ/ZEkdoVl8G8oV34t5WlvvXLIuPN7tkNnNnY7OilScB74yV5SgKWZpxCsnS+saLTyVyw
nux94MwXounVSHNBdw8kMNew8C0P9BGpZMq2RKisPzGatrWDGFMGpAF5bOmxeYjAWnC5PqFQ7Pnj
oFQ4egCCO3d342mt3BCv1NqT3nBu2nYCa/sgJ22lC1PykZwXnOePc2P9l+XKG3IK9ZdnSXsxM2lA
Fu7CtpPy9umed/vDaWd8+iy8Q4QTAsOa954+OR5mAhUso/OMT241I/If25sFfIMNjFuJo/uLTbZ6
jNZB+JubR8z8N844kTPWu5vqbVdudVEaDoWYhwcm5xPv/kviTzA/EbfsVtc7rw6T2bPmlnAY9Hzj
TvI+FAUHIU1AXtQTKUBaXuTGx2aUMEViHO5rSkiS6GNU/0xF6l+mO00ZbPvuMwn/QLcMn+xiIriQ
ige6ZCx6pVGh423IYSNs5ghXIRBV27LkBA+Z2CZiRs7h9ktBRd7IejRJSEV+lZF9aMIF96nEZktd
y1fVWfqVRZb+4lSPZVme9/+zdA+oSP2DMNACj89mnfak7EvfuMJJDms63+XiyXoU4hCnyCUZLfS3
TxA3jyQA7KHAHaVCX0iOLRAuddm1xDOAV9PmSd7C8nas/HEraJqiXQYm71Y/2bcU/qdX9oHietMQ
/DUHx2oLLIg+TFoxFBpFrDTGbQxqjraWie2ebJ7V6/9e3iNgye0Im64tDUG8zAcGeXzWKb1w+eL8
7dSQSaj7mrBn3JbrfWEVYFxVnIM327p4yJf0GDb6Rj7Uvr7IpU74zUvTrdD4xfRv8ImMXOlFY/mt
cMV8qMRQp0NRU82GP1xMOpVE2bZCWxmCmwCF8hsZ2FuzpzSsVAlQOQHrcJVxpHOEaRjUQpDZvyWZ
W7o1Fc6Rg8O3tpivLXoWX5wQ0gXWb2z3j3zpSMKmpl5si3cC/c+loBWXwszYEkJNxSrsu4BMQmDq
fw+FRUtMeWqSXRIZOh4UNO1fkjQCl2CSEZCUeLRQuyWB1RNU+gxI0e6NPukSNeWmUrsgL2HIc2NY
b6iiQEPmFX3XSTv4R15jQw6GAjcjvbDdpQBbmXiGJCBWbhafq4XaSUc/cQbS6reJtSHB4hAh944p
0g1roshm7cVcr7Owh3F+1MsYVTtzdhcCWggNK2tj6D54RpqmvPaxE0JdY1+/emBAFGO7qGmGnYz2
FC4OZD0A9LlYnYj1c0lHhqcViL5+Srga2Yn2nzNsaf7ATBtVBfX44FS34ocSwQ57Mfa0IXPH6HRW
G5MVed+MW42S8Uqdrbb3CzLrgDmgmkYNsKM+mjKSTcs4sL4ffCg0Jd8Letw9vpo3ApLs0c/jaVZI
mJonY3ZuAvA3GfAUcVx/jx3JB8pVv3St8G5gOPIFNgaVV0giiT9RL1o1xlOXevDgtVdF4r6dOgpL
EwPg2P6TZLoCncSvNs0UM96OlvLAwJU498PLTGRvoCiPLOkvjPdNrDJlF0yRw6+yE+XOPrje9apG
plPtbvOJqRrF8jwMXKgATbIyY+9wFZ/bkz28UJAE3StvaNaVqe6Tq3iKvmKtPK0Z7+4QCr7Mh80U
q5+QNyxkiZ9sy1z148iZtnY8ELdSwJXd4SwLCYU549lpoqdBeLSkAr8KGlAR2eirqr0VHoSs0LV8
Lq7rMbG95EXkSgkrdPOyHe3S2jz8jukmGq5OY/u29/OdR9XKom9J83copWew5rUELOfxZh0SsJqv
9BKKNZ6Yb7MHTdwEM1+8/YvER1mGhjzjgxUFkalcOlcuBlsPN6ww87CovIA2KchIq+TseBzg1LrJ
x9Q7n8IilB/vT0QaFHJ6J2PspTaCXoK+evnstgGj5I+sMyWFslqvrnCWrD3Q8S5sVrui/6Zeu9pb
iMasRDkyCnv/gEp+qe7AivgMFy33dBiiPMpBaR7shKjHu8eCNSC2aqLOiwrYh4KfD/qcjqtV6/fb
riVkj+Q7WTjUAG1wmzyUhXEOt9tDRwTrXbd7dtUZiRWboME2DbLkD/V4WJGa6+Eu3HND8eLhYaVX
CDgKwio9wU9gUoQCYoHzSa+2oe/mHRZXV8A8jmf70+WP9NBVUfD03ofNqBYKrRCqC4rI7TbZ51o9
+7KXoMxoZ7X0E6pvz0BgPYYwj6IznecpcvVepcsISJjt/gI7Bg2mbqyyRsNDfS54f9YWNHxyl/Ou
7yRAY1Nz0aaNlYxMhINV9pMDguyq7oLlW4RSg3MZ23rWHaqcHm3RpnoZIp777NlwabuAhW3XnI5+
zTrdv3NjS4cCPUqLPfS/IXj1x9XJkRvsuGZuAlIvoC94DCVNRUjvxPrGLOQ8J/wdN7Yv5cmx6Lb0
TFe1xLzS5g2cXI1c0A6+qBomtpgwsJYGzx97Dmh6qjVlI/KySr5EOf8LK2Ah9xHI3DToGT9n8lLA
4zaqgTwfxP2+bSR5XJIOL335M+sDGbZ+x2oa4iM+y4QDl0Ml3oenCiV2kBk//Uzyvn5vOcn3uwmo
FGbB8wYi8q0I+YqZO/wnd3RWdBiOcU5XLNuzBc8OUdP+JfRW1JIlGmFhgmqcjGU2ssUulKJ2+Xc5
jtUy/hThg2NbynJuNANWlh4orFM9DAdnucUqdgjYZmG/7ED1NpsyZ3mp0fQKO5oFCBz8rjDRQnp6
3IoKu9ieOTkSuW0uo2DCZT5cteon2g5wp9kdAgxlHcNL8p6dPTltyRtTWZg6NFC+neKLIbTFPU1b
Dqh9UyxoybnpEv9L/X0Qf/1dNUVG1Xljb5t7MJAGco/9XV9fl8DmNUnIRXrQ4ktwbbOHLHIfTV4G
pyLUwbjtnfeBLifDP27IpLsIhLHAYu4guYbIqoRwGo9NBjpn0sVQOEpDGzc8jaYpxOzR+L2gukaN
M64JJFhDpaCaXArcW6rhR9x9FU80icDX0CGILdQqAg3bhpXIMGZslGlaosgjZl+adATs++aIyth/
nZNdP/uSiYeTkm3HVE+881KZbEBlMw4mS0LNEQwKTykinXOPPuOwRLJit/YT/PS/PZPqHDFwZ3yh
9ZnS3SWLmhzGjWkctEzf9poRZbi5Q9y17PL+QIPHYXqiNGSEHCjT2dX0MjQFEQSzTA55RJq0ghM0
eC+khTaoIw5E4EnDpqmoKuitOdSD93ahBcEtWXpa5dBaxfewBiygtAyXIOxpdTg8+GbFNtck0wx6
Bj39mZA5dheCPZOtZuB5Hfi0VfwJsLmxGklxn2sviiuaoGPQ1EVcfUWhVWmgf0GmHwdSzpk5ayRP
rauhOElmagVQwolhGu+8YfiyW536jE4LXsI8bd7/PS6qnhDnVZQ6l2LaGa3tXw2AWa7ww0ml9tO/
LRNeiyGIXb7aGKvtyI9VahxOSNuilTkzvdefTMZ+kffYXx7NADDwVq0LBI/VLXINb6DAON+lDyPe
OcEPOUeLM83ttGmueAqevT6doxt019Ckg+OeThrKjIWOWpPAOp/SS8ZUdQggOYdN2gdIPoDTNCF+
Bjn315tVZAikdxbS3ZOovDhmCUU5SiNIXfxyqmuTnr+B7RxtbYqQOetntNbE2UvQUCl9qew/OweT
gwCe8CUL6U+Li7qCcUsVt64vzN5dMjker328cK55yoXDJNB67BQHzlvbyqukmNOA9dMjsNF++tKo
2QgrwQJObQQcV4JlGoMYgI+I7jfchphhRr9nrovynBOEKTSkiI7pSlP9M7sBOxI+FcUebsFscRTV
+pU5g0YPTtf6SIl7RgZPKxMUQ98krCFBpgxv8cg2aYxxNF2OrZYaEqnj2+hUGCNR6h1ZZ9fcw15k
tOyegTeahnJnEEBy29gG9x+35OBJaWSjc+VuonPZR6QuC+po0u7+kq+Jz1rSDO9P5lhdPxi/qD9p
j6etUtUQemGlNsEZaJQ75HOTckiN1BCeSekV+xpbeLBfXMLXgntTvY3GMAX2DDHEtTYdYA6Evj1T
XKjLqP3pL6ibntnBglyRNTutPkAYvsJOIX4ePQVTecMHiDYkxDrtpPdCYZON5hatoZOShMTrpXnW
jZRCz87SEf39We2ow425lZZD4sAAIMlA4SSERBc00nnUBKjwW/88cREJ92SBDMZAP6AfHltTyLde
XQaIjcyKBMx3DlPOP4rN1N/4ZBN2oRwig1YoSWZOBZpsZk/ibJdEYye/jP2WyovOg7dwMkB8KmkL
M4N57Gx2lUpKSOz3m08XdIhbESyMnYKr3OrnFHUs5hrfJc8W7rcixOFc9AH1EciyNMwi2TgjxY9y
f+0bCEt8TlVT/dSZs+VBnkDIB2FtMP+nEMcj/VBH5JpuL+YEDPGcjv05/hKTAjh016EVep/w9jjQ
AheB3CyIlNVx3HppDr6XLPDjtachaKLNkE7+4FEUucs5e+k/ZaiIFPHK7ORKkLhGOvqtZyEKaMbI
SocqOf78ALDhpWI4cVx0g8WULKmWK29R0nL73Bs4NwcAGtZWWJNE97bOMYUZyBRVvt0OzONMnh8J
MCQVknocry7JnmBGyTLkDeE8TCJs6CIr3VvQC9DLfxOWSEgo2zgW6pYdoARM0twBXbrbLYG5hoC7
RSk+k0rWMCbpS7Vzqz+19gbnYXpJES3B8s1AaIts/kq9wB1ccF6q+QkurUCLn2e5efRihDKrfafr
FWvHJCCa6eqsONCXf7gZrxYF8VX6CdnODt06a2zVYFS2NJCF3w+iZlTONizrrCQE9G0iBJRTJFFI
zF3Z+iZcr2AhYg7RNTjKPj6wg4H11N6WuvrmPjtHAAgVnR8jzm9mBxu0b9RSG/u1DWcf71+lTmwp
3hm8Ea4EGbmRXNkvyjXCkD+3Icna9x947cK7eQgjsZZIbJadhkvvO34Wgd1U2Dq9RaQD7Z2S7dr0
XK3wvJcgFGIFd8+yxHr0tIzJEs6YFDE7+gUXCqqBaP/XT4GpR2vwDMrdX8j3H0eqcQGSR/JKotZN
WMlG94/XFbFHj51hOqSMBL5TiWtj17351zligS5bT0/hANx0U2887ZmblG9a9aK9pKQZiP3H+vjC
mqGz2gWsNsU5cg2hntnhyYGC20bvG9prayfN/DeaEkD7vwP9OqVUJ7wRrGEz5FpNYfcZft++Do+M
y70F0+U7jxLy+a6uHLVOGpVD1lBamZlUfNS01FCmnP4HlbEzekVdIHNYmqJ244pV45ivVw1LrVDk
/zdgqyy4crBslCSUJAbIMRcT10eQ8Zv5FozEtsEwWQVy5ECASZBYt9a3WKOZ5pl1wZrfKeuF7EMk
YwthC1I9hnGJ4+0R4jc3wc8V4BDJLgH4WAQzITB23oyvg2YAI7UjIJn8teka42HirRBsQlw/3MEY
R91tqNh94xp6Ay0VtGSFaaC8o7KXCrR2ejd+15w+R9eIQQ4zBrPWuckJ9/X1U9Eiyg+9YjoeAHjr
5OHPkKsWzaKjw6F77Pmgfj5OR/Nyn7FHGNTTAtE7k0YS3jUgjUz2nMSgurO9MZu/3MgihR2AjyBK
ocPcixS9yLRURf2+6EqmPfmUFwO7gggmhte3NRNtEajvJHS2I4WK2F7Zke0eOFElX0HGVx5Va9oo
FYQDSeoLKPOLbSGf8Wx67J55ZtmlhVzFEz9m0hxfOWU523P0b6gX+Un4lCiIWS/VtK7qXVYKTlCa
JtDnHo910+82OteCaIx/bQFUu7rH5hFZKwBpUpTp0+m7rMUWsXh0yw9KlsfKRj14J9w3jb/x6rq9
I9K/g14HR7/e8kw+6jGI7avjh1s1AU27SAhc/V4UM5awmm2zyPUc8icqLLKznyp4yUmlRWNOZrIM
1xq8OHqN9IXemvYNhuZTBGoSEyHC/uJAqerN8JbLBWaHFQItfF2GdHFFQh7nNZsz5ZFFzUj517hH
pX+v6rFs6shAF9y+LtWra3GieVJgFBG1f15cQ7k49DsR07yYiwYaGilQQVPk3MbbehOowiwTl2vL
hI2Uy9hvMuC3um2tVwTCSeXKbg5LCM47JL4FLq97dU0QqUquw+HaaXtWg4uyNtOisSLrQ6kAPwck
IIRHS0uQe8OCe4Loz7IEXngFCQBzfauuQDps7/O9KHTVq/sxC9rB/SbTpPVJ+JKyHXcjonvUA13X
X+pzxZo/5wUomNdlqu8iWbrMsrmaFuHQGSzVfDVT3sEbMU64dUe5LwCdlUTqCUaAgjdT+WZrdVnT
4l8nFd9UE8giOusRtoeeBJw/yUTTRIztSVJRm+cpQXw4EXMud3/kGluBiTx85lGFLdSZ4e4hi+uP
tRmtN1ulK8t5daKhwcxjpOchQPdV4t3nUU/DMCDpln4NhcK2IaPOCSzEBfnes5CGZNUGR/itfNuL
oocgEdcP7aNoYfusXQr8oYao7xhoe3EC8Vmq7TA56iN4t36lZ+b70wzb3EY3ZeQ0Tlc0TwsXzR7k
YV9rBoajR/xuoISitPiHSr5TVd2lQxFygi3FYURDjRnPoXB8AA0PhV8t7xR7o6hoe1aSkrH5aDef
MCmvUq77ZH0WGo53wQEqk8vn0eFDWdnzRS3lQ7FwGp1oXSB/G15Rh0PKgQPukRO3amc7LP4+g/+f
TaGt/DQ5gJvSgjw+DTp7kzwphvnT9OXiMYmL93FZuewYZGegrXC7t+4YtYjGmyBQKsBVz0HI4mDP
58NJ/omrgYHldyhcjx2tqUzQQvy1dzWF/qQNUqOcLVLmvwA3gFHuIyZnqUTD4KKV4XtRYnPff1G+
VjXnizQ2NxvQm0GPK/FcKoClCbw9dnMKF/0RVc/1y8NuViRDSPjFUnRL/I1elcSqsZUuu6FU0kX1
MK4014oEkhZAQmut6omg0UI6H7nABzymI47MHUe4qxqrBOG6IUYS5wh9VKggLMSg0EYavd3cMxLK
xniZlOK86LpdUKlULFDqZJ/VUBtCll7ODIH6hqI5KkJRwt4Es8+uTJOk8z9f2SdUrZBBBkh+SGEW
yWffyMtl1yBq6rUA/ovrgHIEV5khnLk3QeDvkivMVZseDi2YY4RtpvBHJiNTNfUe5E4+gN6yENqn
cpODbuWQ1Lv7wCKux/0YGTVixyZgv5tfFhvtXgNyoyxVoafj98iqX5LGUgvDFIU7jelIp8E1lZ2D
DGwvWIR5xgYsQZV1AaZSUQh0E1S5DPdHfRyn9RsibjQkcjJABXpQrNfDnqiPPE9ZFzGiDEMYPiRR
xiCcdqyF+tp/9kj/uoDaH5wFmIKDbPvozrv/HMjhWl9SCT6rIDYO96l81GBc/gUipdxP3GbmvPKC
FRwOCw8kABMWa9ku8/UxkNTecmCFn1P1K9nmuBZEpuLMMC5TXlEDtGq8NZ+3qa1Dp472z644gRn9
eFG+w91PlSIisj+ffEXDT9P44PKQmr/iI0Rwhlh6GXRY1zx3nXj0t/t7puwnn2VfP89a38v8hQpQ
yZ0GM691IZwQ+Ph15i1t3fL/oMG6ocKD8cEZt+LcM1Nb5yTpT8jO/RWjLtgw/KgEWcfUALs4SN6E
pHJFewHJdOflNfAopWO57ffseaVzDtIyARizGn8wVhkIi5s0bj5vck1/Z9SAsRHrXetCAHS8onQB
BOI7MPSefZ8gEnjg2fE1N1bCqKdL0PJy73zKPihufe6aLW6cfxBOOI4ZGVymVZ6UYS8T+tahhVzB
DXyajch1Az2A1Z4KV/Qff+BJSMaxAJs3AF0/t1gYamTZ3VBQBqUeIcC7bxB7k1M/HWnyQ5/7JPdf
GeFQkJXjRGzdsDN7xZfs2FpLIwQci+05qUJELoHiSllvwPA0piXHl3n5U13SUTHttDQtpREfHfVv
p+/DK7yy9iLkK3uvM2yqFB6MOViKIICJ9SF6ZHEsnPPM5OPKWsw3tECuqDhhmTDGGYe1y8+pbYGW
Qou+bzh1Sr6rvlrrJMtpny62niumAOcI16ArZFk5L3r6IgbpYJluuwkP/o/veTbU0TIJyO2OAO3p
hkTvKCPnvSV+u4oD3YREoMV7pOyyhr+OEaVPGG7bfyXk98+HaiPRfJ/9vyW72pmcdnd8VVk7I5FW
xpbIllmXbLigwVKnmN9D2Dd0fZlzZkjrZPV6wzmBWfu9nOmbvqrbBza5yvSOYBDDbXvsC/T/WpuS
SpYnyFbC5V/zpL4fSuOjoGhvjYBggMoQXLfCo8e4naFx6NITHhiT/MHRco58GZ3Pk+KvwKjPHTVl
KGNXWZUryEyRKfgihZmwjH6RYhpENddN0XQpyUq5DLFuillD3Ba78HpqDwTZuvwD5c7gxtOU66WW
XHI4rpA0YYb44WmoVNTFeUvJvaECugf/IJ9DNQw6TbH9AH0Iwc7B/k3idOknMSF6txvMG/IhY+gJ
6XhCymT48dWpGfvanvukyx31A7Ba8mhshNV9HToa7cmzmEqwL5aSVLVqdZy+TgalCaWZvTxbVNAq
jrTGS2/dfrWMTy4hauIHygciXXLD3nfvBeVRAiZU5nfN5vQJNXRdWOxnJni+95Bv/8f7iJhgXDvF
CcSB6z4i1/UXfhzfy/2geNH54XeyaPj0OBvMWTUTQJnx6cN0vlUN5u7ZgGThKvYdGWNkKiC4wNmS
LD0t5pTtKgExxtVTguqmM5s5dVX2QTr6TQ+cxQG6YtANi/wcouMMsu6P6aF8vnEwBJ/yHtKyageG
SVqfdu8UCDgXj1o/aXkFWZIO2BtUDW6rWnv9VjEitHi/besJTmBSg86IbjbFyOkhgL1lUO2IoSAt
oUdSW3NHWMXR+dMo2upLb7bPG87n7bxmK1l70AW6k3K2n9uh2t7lNv5YjMnKxmymz6mA90N7iYIM
YMe2wSo+M90GBJ1osmv0O0UOW+0Nzr9vil7iooopeQy/7NRvSfT9nUFrOd8vJ1L6xjkatElm0kmP
9IeQN/mOtzaEOcd3dJT2EGX0RN2ZwHsQC7VG9pCGUTD+u4n2muCphszIXatgh4/5jIfTP1KrkRKG
+uIybUZziGKJue2kKHIzXjS8dsm/rRPLtQAO/Rr+XmuRzt/g8MAZaNwMnZGfyKJ5wMWCvUDu74qO
HFvpvJWugOyQqA5Hla+I4RSuhzRn/zq917IR2XrE07Jr3qrjp1M1nrjEsdT9JHf0LHe11hS/P4fy
Cnq8rTSycm/2Lbb5XPwbKjToUAygZai5PTuKIk56CEQgMYVgarydij1/L0k/4eNJqMGnna/pAaWx
CkfUbe74dg/fjbbZxehoT+CuEwQE/1xucgrn/B2IK/rIeR1++qbh8u8gg9PMbyT5hmMcmLVGx8DE
HyU5NOXdecwTc20McKeqamFrXyozOPIaH0eCJIhPUf0m4WwL5/lslUWzZ4afpH9PReBuGaaDeSV4
5qwzcCivg1BdU+S0wXR8VsXpuFUzvf6SdRZQHSaAAVO1DV4jOL+kOZKnZf1z1QksN9W+FortDwT7
uBJsPiUpn/L+51VZmwLNLwfLxhYDZaOOMq5x+2laTSgylTxlmzU0lCLiLixY5y9wRf7UUPhs4ewy
pUA/f27DFav7EqvroE5jsITqDqmdL70BhmJUQRcVHoLVf9/IijhlZdTi91PzlWpUuUR8vMz7MiNY
gShejEyxm4MPBEqavHrdqHusU5sukuF/5oE5vF7ZYyeSS/3gbdFwtbqKwfS1eBHgonW01e8/aIe+
JVsC7sfFWKDWl92ERtpq/YfzwlT1lZsGntwCYybh0alQ9YMmV6of00iOclBfj31rFnDCVQg0T7wR
IC2DnCb3BNGCuKHjgfUSwbFCroZ+UewCEO8z/iuc/iLzhFPtiApK6uLkmqSOvnnrQ5n4O5cocTbu
YDp30IGptwvhTdCp97gga4Z6QA9eYiRYYNmqOpbC8yQrOv7SK9YV1Hs850dL5BQ8aahNe8/wfX2J
m4iqRB+FQ3ilK641sDTSxIlCxljDAlxURCKt2AaWTigZ3gRNuKO7VREIJOjn9HdFjpH2PKTsK9GN
DnE32BSQDk5woh/BDFoueqLsNwNRTZqwgtvvYW8oda8X4WFkuvjlD6h6bs05yfcvEiDrUG3K/+bS
pUyODuF/MUW5eKaXoP5io3Oy4TlHXbdulBL7a7NMCsK8bUoEDQkje0my1vOAQznxw/WGlnNp/H8k
9VzYM5RvRXl+0+acKIjMI3xKxdwWtzncsIG8TXQe7GkGT7oDd0nzmtZSPc2amTCGukRxOEYbKQ4i
fRzRAChtxAhNzotedmWVVw9ti74oUcAMdYgYmkTCqeJOEHD4OhSu53S/NTgKv/eLmTCyX/yLsD5U
2mZHrRc5GoyuTWsPb6AXudBVz+pzBjwjKdfL/Gy++KgTf21vfOe+c+NURvFCJrETP/P+30wDLI2A
1jn9MtResVCKqH21OJV5YJIehTM+fTIaARi6Drl/40vaTaws49Z/E5GkwK2AJbod713NkoTrZHnV
U9IBNTF97Gk++HXqNlhffYD2joerGkT4mQQuLz39HBeBbanxJAEUZ0GOgUOXW0yzUFtnvEKSE/ts
J84dhb1x0YsO3jHgfrzvynr3wQ166zOgU1AGMHnrcBy+iroxbm2PPzDe1V1wuUBo3/UQalZgDdyK
pzgjfr/gpwNOmbhQx9QZGHO8Pj/s9x7mgAuj0qjljVERZVEeFmAwiwwgYtpc/CPKD9YFcqvZisW0
TvvCwxYvDXVJ8vEH0pF9i2Eq4HbPqyxxmnTRKluPN92Tkru3RT6JIpUWTZm+s3J9roShEvggRgsZ
YuSZ4amiTohzFCu4sAYAo1SdctFzu8l7B9/bEn5rP0apeWqap8nM2TrrmfE5SLCjof+4NO3bWG/q
U69izXxj3GXkHKMQK+gdxk/n0dJHp5aICKG26WRaI26PBdnZBSeUvoaNNsheVfhqHVCp9ipYUZa2
zG+CCf6HJR35Q3fYx2qGY6SvJW+o9CtkQmTSW5LzAjVOQMjElMWXK52OusKEUQcKBItYhxHlK2C5
CrwBEMgoD9VXPsN1tZ3YVtRWGfb+Rj4LWLA09r1IMAjY02WW5aYhJtXUKo2ULSsdMkOvsCNBZtOl
NRlLfPFOJI0jbyqG9x/Oh2Dp8j6eR/aSdIA83ZrKNaslAMprRXiwqtggzzqp5cII/vuftW/cPm7K
P2LekPXMVMT+Y+8NqyqIrEHulzxrhBrYuysQY9LtQG/EV3QOlnY0quz54C8JDVEAJYQT65dk2zyS
Xg8AB1PJBSUbM/6Gp6UzGFN18YwBQdHzZp4bUGySGBKZXsgG0CLR/E9Fx2Tllptkz6mnXYYZ/8Za
TrgPA0QYe5celj1UpPZuIDX977wfMe10MujsKk74NRGwsjiuMLDW7S9iW3uhrN+OeB0V4Lq70IIl
BZBfWOwmp2RN+462VjW+XYl3ErmaH20e0r5iMgXRb6HcPao1qc/dAUTm4fNLlORt2lcdJQ/tBoVT
v13cEa/nkta7JlrjzZFwRZWTU3kMDeDID0JpsaYsjnz5rYS4vtYPDl0W6CfEoBPybys1j06Bt7C6
8O/V29WSXgA1CqzBYGqOxRoBP4HA9dnVJCmMZ9k/lwXHebtr+bvCgLn/nD93n+95nlpCuEL0ouEF
t+L9U4RbzEoar4v31UwVd4cbjutVfjao7RCK9esFKLM7EkOTKGUfQWGABI+U3wPROi5uOWoMdiyZ
O1YmRHZmlPJtVh/qYqRcrJSwBzTx1MJq8T5xF534c/Di31KVSJJePaqQFMhHnjEKWpSCjM6V7laV
aCI0KvZxfe5MPoj81vxK5BCy+jg+tHP7rBBIYEl+d6iWQra74KJZG2jB3dNVV7w0Knhfolv83ui7
Mw0Pl7pgrQXqzPPpcrzo0MEfmVEJTILQpKiv1gO2Fl0AipZ+K5R14w5pDxshmWpKZDS7ubx2T8Ct
04boMdFcgFu9xD0dum2aJHMk+mTkKbL4QWtLzkl5NoFyTg8Lr0MwzA8BgXhIK04Mo24xPX646vIq
J0cF79sYDfCAanOevKkHcuFg5OSkLmjw3ZkvnLvPYOnmg80f9vK7fHvcsUZ5zaWB/x0TMIRjZRwd
V7UGQVIXRVqOJ6Azq64puSKiTdLsCLjIZp1kgejFdZc0zM6gMp7PpkmQozBNkTaC96khdShfkFWV
JJpj7NbTrR+z0bTBcRzCsTT8vSQ7a/yYII2fZbV9XlKwHyci+7Y+wyXqYqFUr6PdhTcG3oxo3FVs
5VN+6oXaw/KvepLXyFmgEMKENWaUY8sIKK5Qoe+e4lsMRqA1fC1EcT1iBS3lB9jmrYASa2uhb1jg
4jKTptGmXBe2B2hfSjPkYzMLAfqYIchVtr5G4hpUC3Ls/2YuI9/rLGDNElMUctUNF+lCyDOusOZB
Jif4yy02fnpScMNCjkH3O8U14FrPtP3me/tRpZvpMp/CpPzMbAo8BLk6CNlXhDPfDCHRElCTI10V
l0ac7iSVnpuder8q+aeDxEBp75d/vXVGw3tfaS+szaxdwehby5B1MK4EgxIA1tF/Mqsi28e4Ncj7
6j64kJRI12VBEGXO0BL4OgENkvotyoHm3NYPqdwdqfUMuLC+Rdr3dSOiU00Pnr6J/NcVWJUuhl8i
VaNc/KtTebu7KXNOVqeSr33ZTuAPhGjPZAWbBbuHNdnOuqzEvaj85OH5l92hbtsjpjvPSPMCQ7ZI
qenl6M11d4vsRSIosn6TPfurN6VdRE7gYuDXCk54QaSIYM/q+Zz5AclRsc2DiyJMRU+hhY9llo5G
+Rh0gRzBQHNgftKqLQquVlDklXyTaiqQmNHQKKKxgL2ygC7GfMENV+xMsuDTg7JtKv+IK6/f20F6
LQ5a252rgH5AcnxAhY1iDlg7IaT++4YEHvTNEYMJDn3KbdvC60m/wGDlJxHHyLut0JlaK/6WrSrv
E8cqB5z79Lzau6+rlZNv6Jn+ttIWNnpB4b8FnBpiIMN9ahVxRyghc09AfA8fjscgbBg8AzU7Rgko
wUpCyRAsJhTzHaU1aiAHoCtC6ALSH6y7TPYPaDXXgij1QDJC9ez0PYUfl/QcSLFhyldrobIPS2fg
b+X+fJ/nl3GRrCN/W5Ff03raXpysGlTPAUBydtk/BbwR1JoyuJM+sLSEiIKZPrzM4e3mivRm8E+d
M+eoKZbtMZoPcau9jVzFzrwPzGazdPaxbmFQHeLn+LJTu0o2sgK4BOMFpJR1JWBbMtiGMF+Pkvqq
zY2bvEdx0E2BxioBmA/ag734PPLX3SX8brn1guKvsad8xov8qDrIKxW97v1gOvrs+SsEjhj+wiWK
Ysasnehqi57lVK46DkriFXPPqSh0CofuUyN3qWBRclnwzoNdllytZn9IhImcMb7NUPKKnfMN9M8o
QNAuO6Atx3WvvTGLcWIgwuusrBxSDT5HYLHTzoRuXV5417YJSwEUdVQTix13JiK6uGOXBWOSRwIi
5+zw89w3tgQGlVF7doFPvC11uOfxQIjN0Y1EUbXdE0lryh+e1PqDzM1Q9U4EgUnKsnuVClnm2DAD
leCWlhyP3jqOC+Dp9riudqrny1LFzs9mW0C5Y9gZmB6990HVAGTTBovwN0n07QjGKc/yaNNNf+8k
ZWPafGn5ZhAxL5Dp6Zz5qQbqnNDwFQUn3pgh/xhG5blXvDuwlXqFb/P4BpHDFKET/lwYBPUhIsIS
1+xXHin3XyLLOOrUPPQNxdsE2uuW16j3JxjRqFlW7EbVMvSq8J+Fm6elEnmpdu9OS2Qfbo7/sQSN
fzWOCNIhUNGrLIC51uRuV3YTKo1b9nmZRnlM6Nfs4JH0ZlhzeWI6QmneajGfqWrTG31kUa4SDaQ8
7nY+8Ov+aOb8yprZqWdf480XLS5aMYSs7wHoVtr1Ege0LmSi8Q5aKhxasJCYK7ghU9EDrnoi8wz5
G9Kuv83gzYnXEcf7NywSz6MH8LAeyzTXbM9c2A9ekxM6wUM3mdcEX6I2PoAjDizYDLSVia9p5ixS
XfgvmwVVdDOeJvPQRBt6QqZ10nd34BAWUGRIW6CYDnMpBuU+SVRBQhsKE22fk7meUOFLl5ce0Hlx
w077DxX8TlvVJU8VFqTrOxm+JisJo4YeFVnIyeWXRDtgZtrkPaskw1r/Et6LwqfO8XQMj0OTmRMf
uoIVvsYl015kK8N+NyyTbn3yRXZ6f2i26tS/xqMhkTGYS7szSkq8fbSrqnEI7EfOQxfqG195vZcD
kOpX7DKrszUOiwNmz96GUy/ogi5uTrYoVgKNTjdtoZJOZkZF1owtaSeqYzDnu6sQ0+tFUnYgHvGp
AiPauI+X4fzWayDONBH3rY2LLPyeyRO3l3CvqpzdfXQa+BeIsTNffBRSQYVahoaZwNOW5cx1pU3d
c5nf6s/A8p+6qP8ONDPuI1Uk7/h5bBDUh6qSBiZXskzkLgp3i+9QTxme27mZ8qYjbiRb+/dWx4CB
NcdSCMD8bpIeyXE3FIWDbQtGmw8TVA4ca5X5JY95s9/6ocbd42IXlAECeAPEnZDfiCX3Znwj5RtX
zN/IVzlsGt/4efK2TwiiH1FxP+vlt7Ec72TkZ4V4lvf0gzhvqv8QI86DKCJGzUk4QWQUlZvkToY7
LZu+nGsMdGBTwQ7e9HAjXjJTdVKuoL5rsRBpexqDdzeHMGS7G+77wuo5SqRM8yL3ZgdD5YHmrGIx
DKJg/mgKm6uHlqEefUKdKT85Ief4MwsIjFVQfJxhqgvnNBthYPDIG38fSa5HgY/qBMs1uM0CJSou
eXJv8N0dIVgZna3Y3+pwNlqgbHOvQEians26uB2EXl4g/xno6vkBmWp3fG1ZbchSZt0ZIe2YkMZ9
h1bugkftk2AX7Y75H4pofLD+pyCnx5EvhvL9RvHq2GTzNBvIvmIm6J0qzVmoGKvBQ4HFOsJSZYek
/gT4h/8hvV5HbnubyfK9pJ6vm205BSvsF0oQVtWnnp+y9l/uj6g2Bu9S+Wqw2P1FZgda6Iae2Swu
8VYj8HZEdWVGZ5RnPTnd9H9etmNFqu1iyiAktfzWHyXbriNf07MB4o5+A+l4AfY0EW+1spm9RAyO
98fR76dneD2tuWUI2afpsVJr8AmUIGnxgDlyh1ecB8/b+PtFyLFvSSVYfe5hEc5kI2oTwRQ2Slq5
KSIW6xC7s6NW2eP+X3iSpkwDW5Xtuy1tnVoemwjXjIZUzHKcZiYHTQx3PgZmsM8Yo1IZ85WNZT7v
UUAHuYCBkkAfjf739HL6JaI0VdK8SK22MH1FbPApHKRq6w1usl5GotfXOdMjt28uzwysNk9uH6PA
ghw3EhoMA5sKSMzZZ6i9ND7EZOWCJIcBmOIk2wwuRTXaBzXSuv/4XL0bvFzEyok/rGK/2Rm7s/4n
gMhQ4BEFI6KLwYHSG5Hv9wORuLBgN4wb7lTb745IQndkcjNJANEXqhxeNE3/ufcFsO6NdWONubdc
X4r+QnDxmcccehWLbSZrt25VrtBA+Ixfp49/aOw3J3z8gAsJE444w8gsPIhJl1RM/BhJtUuo89sO
WxIR2XMoAziSxUpJXzBHlYr1EL+BVSh+OFnVjOJ0axtTx11TMTaGYJK2VnE3iY7fUX0eYHAMo2jb
xYkUMfFEF2Jn4qXL/QZh9AEOoJvKq+G+j0z72GvTr3162yAtvRMGG1azHi6KaqqTqwRB+wApacIy
x1slHVYmiap7EB+oPWaFKWxPdU76hiOPityrifSrN/vGDU5vBFBZCRlkMOfLDTY1oDYL+MG2AFcN
McXLGF2gmXwJpvQSblELg9yBPaY3xdxOLc6DhrXLjuybk7Ma2j6kaExcvBgK/cBGcI4zAJjDVsO/
TI4tjU2jCp5QEliKMg+RkdIoy/h7nVviE1pRsl0QStrUB72A2nthWP/BKVlNP8QIYyA6mxhZIr1c
yKgaoyzXd0zwKpcObR0esK2/i4ErwRSGhBCwgUKHMxlRoa9KidNAplBVzPHctGu2sUhYt0LwU6mg
iI/9uBoojVyEDpMvUr0MsZkMuWM49YrMR5yezjIEYexXfSngXtr++zrLpxq8oyZZj0KhqNOjo3aT
kXWCxLrgdsphV8s1lPCVv0tg020FwxLT/U9qKJh4K9nxaFYAjNHs7CV50o0u7TyIyy1FSMZjIqKu
qTztBs0G4HuIBKOD0qZVGCBhjJPHT+ZIIs+RNe4ylRoJEQDvdKRbLZB5U+lN6XsqhBv+wRTZxoop
FwmHrBVZaiPmw481XsdPllyqv+GGqnXdA/4DCAuacujzMO64s/S4XZpevZx/sMqvs+59J393OrY9
OxuQZ9u7AeZT8V06L7QMQ/pOX2T0qIKUUYZhvdtsi1kTWB+h07O5LW6LVpgwhE7xVsXGG6YEvUKZ
guYNSa7Vo31dOHlNsBTnLdtwQrC/lerBAWQLqVBXWglDkzRqXfy9SH+foTeKP/fp/tOawyVCFfdX
3Z9my+sHZiWs6PT6WbJzrDlcxmrtcn/+bwg4J9pJJe2lM+UpXWh0eHhYpjop3Vlr/QUNJrvAW3gX
sUiR/vg4Sn5bh4KTbwOhQ+B4+xDozSb6bxuK/4qiwtnOCxPFXhFDsXGXTLJujak3xrVej7hGcn2p
3irILgFuWzdtTSVYxEIM0thoCMMGthNWPbdf4qNnVohPSHJ1bxMApI1n1RebrLba9Mnhw0gGTUU4
B7JXjf9Xc6537lIC2sFUHLuBZSThXy85F/n94Y2pskLj+8SSfQjbiHlpnv1Y2mSrhVg/mi4ka5CL
AoijGT9PSVfErXhfukyLF0nW9WgYMGr+mRRqPJ0kEPOCZtnoTDVzB8xCqsgAxjfTWdvz5IJdMdPW
wbXbM/jjOQp8j3cpc6DqHqhb93AeIFJNDyvyj0FHhb15kXQRuVyRUxNOYmAk1EcPo+moQNYAJHHg
VNMRl/t1Ewqv5f/UXKtD6SBRz0d4fDp5g4DTVCjGfDeSoxml2rPnApN6fVob1s+WoVh5isIi9oQR
NA3F7l91vgGg4E2k4BccPmbalozZV2nnAZYtyPMSiQ3cNcSC0l1wKb8nDw1czcG3Mj0iKjYShNQQ
LXJLASvgePwTKJQ5+TW5BjnLCax9xDUAuanplIoPXiwAdNU5h9Ea87P4RkKM3K3hd9cxW6hhar1D
i0YeIcKXgpnloDfk46MtdTNv4YbsXU6Fs560p0DTcpfhL9SfWU5AEdbztsfsoYKpPKjmqoaEzV58
H9P6o8FLoQ/l+dkDlhLcoB5JHSKvzgVuvnSu3cnrBy+HLkGhAO+HiZlIkYRUf+qvEpD7gkFq1NJt
BSXXZ7nsBAn91v5cVJRLcsC4FpUp5uDu+RpbIUNawpOAMELqxVxIX07Bq9+Pdm/FNrXKILP5+XxZ
kFIvKgXpyiG9W5csxzG/1zAO6tQmqNdz1APu+qVQJjQBaCw97GhQ9OVGNKXnaa8m5nb9UuhQmfop
lUB+VAm5Z66QuJMycRDmppi/9KJct3SsY2jYE6vsKQZaxz1+2qPDpQaS9kNyWTdxqF/nXl3id+44
8CAH/7/FEqEfixJW72qpUuyiLun/Kj9xZhGfglqkzH+7/JBKyPpb+AWPfkbrarCyZrC0VDNLUn//
jUbGzwV98pBs9kkEEPCyazAUvHSHyM5yphpCL7ilhTyM8Hajzok4u2tJtc3FXbw6KWYzVO8v0pKM
VeQIuBuTRM3qYCs8MhD7riVwVqGtvE2DpTsXyKBAlfttJVLMzanu8sDvgWEDfJGjacjMT5OcmTtg
XpcSVeq3KqxEH3GRWBzzzHUpG/kKhqE7gk8xJBPZ0NYAMhvoAG5rdU9DsZIclmO2/bynq0zPTBmE
IxTC2zEboadsDKUEzCwB0doeKmQu3txRf2jBwpVZ1F1bSla8TkAEW7DW6AsEIOuzIAqNWr7YZFZG
sMN70f6HiI2D8Y8RR5dqA3Jwqw3CUblAIusZnrAoY/Y9Xt1yxQJMD15EoQPKw5GKzatv0YKDK1ou
edhYT8aBZWIADBczMCABBIMo6rJXU1sgmHNlNecMXMv9F+1SFHtprpjJKQoC6ItOLT6XKKmTjwC6
Z5GoQImR3ZGmuAyIAb3QkJiYuhqk6XvVwuIDqXqnfteW8Ym9rF77EY/1lZf5Nw5CUcz39fluIhuC
tE11NruE26BCx2RaFlV3PMzmOFjAYqyK1VP+Jag3oDTR7Ca+vaKKk61MZs+AxqN5f0WThW8Av87w
WRuG/gIgmTUnxg3EhbSAWuODpTrOKgvarg6ZW7xk7XBANxwpETC4ohx+JgygiJkkFC14caCq+zT3
/1NBzJY+tSGn3dIZJJ9beJAvpr/Y7Tk4Ag7foSVyDEAhttItLOpT4SXsTp1j8LeSXZqcee+mzJsB
BB+Wyim4vrzPbq1r2NRcrKa/MRa4pwIx53Nl9C91GcrCIaIne8kdbEqx/7WKJDvaAANaSg/wX2ee
32tcPNl9Py7tifcTd9Klg1CiSzL+0KjRa/VUtnt2QWN7pWDHyuGBq/wcRI62z3B86JSjw+bOvkNe
b/xrwPf7gm5GW4oS0gNWbsQCEjT1NBDjwRXfZaF5l1cMwCusNxQMKlwN5PQJQbyLkJyRDOPBWo/Q
C1eScahg1jU55j0YmRT9zhnH4TZmeIDwErPT8C7H0B2fH4AkwEKR09Ca/c8HFQfb9hLpg0fTnDjL
E7/TuxvNhdqzOLOLN6DRy7oUakeAntIMDy+BwuGQ4E58UIcuDBaxAcF9AnH7H9IK2vgf9b/daABh
IY4vaXSCMFMPZtsRrB4S6PkKYAIK6IfBlDvJxW5jx4EupL0lXSI635VKby7NmpDx4+eSE4V00JZz
H/DMm9TtF2oKdC1ya7ZQmS2I2QS+Om3I1d/10dK8JEgffOWEsCDegNkwtZJDI07V8MtNrckyqrVV
9m34DW6qFTd0Qozu4jseYqFhKARnazuVeTmYfBQGZgKHGeqeTXfpGrPpIeSwd9pMy9PMAuQCiCpC
i23PKJmYk3hv8vBEmUZ+cBW3S15qab01EPNaU23yX1u/LVqkilVbT7M+ORWeN94/jkx/wrbDrccd
DCBMyP+OeFQHc8dLvdDFKabGqTh3JkJ93tJc3IpdGNgArZpMEFK8SJI8xsWQmixW/AZSlKMynWRv
RQqpUgNIq3TKDTyxJ73s/cpgjv2htWeGy+k6xkoRrzROYGrKdyq6QcJSD8Dx+pVrNL4Y4hV9Vryw
NP+5Za6BQqbAgUjHQKZDW3bsx3RSiNajC9rrLhPpauuYwdTWodamlgPaAfWKMnPXuJyTeaAPzU09
pmmqjf/zKU4vM+TDySEKMm4F33fPKAxpmNFQv2s0yUAELyiMF+NS6x/lfSGGOxq7dSqCYi4NbiuN
jkJpdDuaWKs6Xnvh3r5XocZ5sHzGA2Gj+Sx0JWuB+CeQaCEKxt4iF48SENcL9BUu1NPgzYOqhXWF
btmWvdm/d/wfW+KDZkzWxpGN9sQpnd6KRG1EhHMH27ETMgKBIOVwJeVG85FyonPypZDaEC0NT9vG
ercfZhIEnq2E/jICwtWCk9j+V6zYp2xZGbRRsADh602tcJ1/3WVqhlTV3FTWZHhmr3kaYGNjkfss
MdbqjVlUDyynLY1pPSWOLg6wxPkWSD8ZCA2yXUOgv31Jp8v9S1Z6CQlUWp0Bte4ryKI/kU5lUFYF
SH7QcIkKpI7bzw1MLHWK5FlFMi7SvLE/MdagSg/vJ/sCJ9JbmR5D8qUEyBeIdSVesGBR5XMeam6F
dZdMlkLb/5uZcFn+EWDuWJPINkjIVURxKdJRNImTUEOAu2s2a3re5CDexDUXhPFVs7HnnCCrozOB
F8d+wmSmBUCR46DQehonod57RH75kc+famP5/W9dyCRxOnkw5YhziHoLKYB+5Zvj7seRX9whoWJZ
gAYb9NKsA5DWBYWL2RuQVmtAVG3eZDxgZg+7byQT3tN1ZLhXfGvuXsAZlLQ/9KaFbh9HOHSXodr3
kU2vQ64myW5mgxKP/DBv5kI37m7KqytXkwbbAMS4XZWFHeYDAFfa5IKZaEXEVnQQ1nDp/oMQaqje
ioR0CMu7Jj486fdPWLLQXfVzxFVqg7SgVehyTCkM6aIIAUx+hEaEdk4RRWQyRbHr5ZQlS+zS+Axv
dziSdx8TNCxvQL54efqLAWhKb0vOZkleD173349G+KCBhQ/qr5T3UrZ2z8oFWHNdf4Y4Iln1vKm7
ZWqXv7X9myrL9qob3xhwMoH+B93NQqrjERtlViDKLMIegjfFMHOTY3Qzs/GugNHOIepInYm/uxyD
a0BYjDTNH1NMByR+Zm1pQyhkN3bYuGh8RLAVtCEr4nzgPr60254KycibzkIpU7A4tNrFi4yJH7YF
RvSXuVjH55XermKzjDsfXpUw5ndQcgwVeeCAdGtAsvZSyuA2uxv9siwnAYmLFha14QgBwQ20ydAP
7qWJiizaZnjFO8h4NGgIOs+zKtZq+IKvMRyAF0TX4jxBPFbRRiv6ME3Dv/3BTZK0BqODMs25B58S
M7J6O8aW1qlRDZQNaZEJcR+fOMKyUNwLQVWLz22OQyC5qYL7EyI7TAU+P9abBa8s+fEywiE2vTCi
TMUf63BR1rM3XwHDYToLmYmcTqOLkAZGuj0VPCKKJqX3fL6AyVIswTfkaDMfhOlVyLhjXtjNiLEl
ALooFGO4MwRr7q9AXI9zH4PU+lD7XlfqZG+9P9VrW5G0+Bmt3oYUv+0p4XyWAY/AxrDp97ItYbmj
c1La9f+LHA8BMd0WbEkTXVk48lS7uGDleNmOGxBonoulKHLU4T2JjtypU2fjXBjDCd19Bi9djT6Z
XI7i/2x9qGDlHvuYLxOrzi2vNw1te6GrCnCWt3fsN/+HKZ/wSwwUNBuFWxXqXloWNdrR4Z1z/d52
5Tey6X6y2sddR3vLGQD+2xQYnMJEt9Pt+L0eq81bULnqE6uZM40jsV1O0EqWEEAUvsTeCfWoLttY
xzf02ALdUXfk3bE++lc0sdqaRXBUiNiTyzDPaEYixp/BAi/uPuY2cwwxp9dmlQyW9vQc6TFdFhjc
83CfV/XC2VnrD01rhmQXHoxsqb8jdhZ0Bsnbwc8ChfCf7rn8KozW3Fe9eMzJ9dE6syEH1tiqjr4f
+0K8CsHFDirrAkENTxmX7RzD8Q1dhr56Dgz2mTx0mCP19EM+inObqjN3NLMaUq20ZIe8Xf8KMEGo
AHHPEUSec7VrordpJDNXvQ3C09DMePVXteIm2yc5mbo+s9CUY8CI6G+48eKFiX5M+E1XSMGvHuAR
7XkXF2/3zMLOajU4ZzaDQozz+z6fdH/kxJSp/9FtHAa731OwGPudDHzje/82Lq/OoHdvptogh8za
K1rUBBVb6pPaTxjqZFXo5gblcYX6KOY9ZQ5Ej0b9lRBkui8pO9CYFTjEsB9BOAivp6mqxqQ+w8lR
0EYrF9zUzrVV3YZWRrq/HK3cTlgYksWNXAgisUJky+/mH/eXqaKrqtLbapqpQUmX5vBSqN/E0OIT
yMzu/oc3eVu4oS/iJSaYUiFQp8+DdmP6TGbJF7mjLr93b2Y6m1gKKJKRSr4fPaKqkEH+VWyOwc2x
sdpEVK9do4LksmbBd2SkxrFNOkbvRr2WaeyT8/GDq0Ia0OdmoLOQvhI3MAeh2cMo1y5U5cBB0jfX
kpfWWV2/m0OH0j+4+aCUwZJYaLmEdENejS0pIWCYCH1buz3EeTuTGgBjK9u99/mmzEuEJ7C9bg9z
q5oXsXzyLkuicgmVEGLfnMrSRwjocS7Ss+lV7AgI3H/M/CSwBW5LQv05ashY2JppvNdXRiFdnIf2
su+kpGuuGUEjMIExMoxEEAiXex/0fKAYaV/qGbxPHlXAUQ/zXk+Ffu1810Fsn22r33VQtg27HVlB
P/4TdeLqlV43x2dZexVl2dH1GeAG+3sL6l4mF3R50bhkcR8Lwjm9mdSFbQjJ/IkKxlqEkkd59EhT
MqnNKTAyZne4uQ/SSEoDlQOg3jrJNyyWjFFMU7mdjkk5OsAK+tG1JRi2EzZ44fjuVCPESA0XYRE3
tW4kYhBSamTXvJVRtqHWsEmuS8H9GFiEC0T6kGfnUGNXqD81zl6HILcR5jpKte33JdOl0rkOz5Ev
ukZFSM8mlIKzNzq1mwWHqmPrnqmxpQ5FEsUdIJHVK9O15nmtuxe4ASCsw+FtXAe09zJncir1JUSu
iqlVjpCK978Qi4x6wr4bSVFIMM+a6acRHHkU95KkqsYKZWnBD9kFPjL/sAmtB4T3j0C8s/jZB3vS
+eNcfUXgafud2OLioOsiwFmLh9fJN4UJ2zJjZ7xcKKbLhMy0+Olhu5khbQoD54FFhn4rCi6PllLD
RrJhMCWEJFqTniKCASrQNDNT3/zXWPUHI/4UEQZGW9OoQfwL2iTZVajvm20IL7Y8/WN7/pcK9SPc
42yFMAJLoGOwtm+KtK/gBB/T5CtSjFXUGZtABvcZm8OSD5t60KfhFSKiEeXqnKu6erLLX3wpSDh2
5gXZjY+TYTyjIby8tGU6zCjrrA7alngqVBL3ef1UgMcepal2EmDI7JXjXZKf+dqjTcMsFrfPfXA5
snnYRgDE6nOiPvO8ARj6rWf6OA/USNRxn1h7v9vpVbsrWv3EaziX3X/YoLsysWt/ep5QDJniJisV
lmOrPHnEOlyqrfCf3LV0kMQWXMNriid0VWeP1/akR/CpS9CrTdjuNj2Ua6jC7xmI6PoILPuKUONQ
cISZ7IFIKTz2OzlEuuMX3qC4GNrKzrmbCtUuuCjgZD+oFozkVVAzPs16dAFljyFUck3/xYGJrPd7
HQhDB9XSLm8vx6ZuOq9jCIWa49p6Ybp+4Aren0BGlUZHfZqNMlgZb3XGRsjaxrkTZorZngbU8bnR
FdiVF8lBeNXEuLTnMRRFEKsarVqzEuKBT4xE3SwwtHMMpCXBk04DyugNQq02WK0CObIdYcqplmMD
9WxiyO31hN9/eIIrCOgAZY4LORf69Q0VJve8Zy/yMbE1J8tZgNxA7uEfwBBBOXDR6tEcQ5vwQ7Rg
Nm62dEFTvCCA9890AqJr+FbqVU5WbyYezQ9cKL19t/rxBAVNaGa1w9xpnnweKwQKsqwnQmGZvTNx
YOEjTsANQvhA+VlzWSjVGcBPhIkeSRrpuJ403XU7Q9svyzE3qv11scTICiHdvF5zFNCW1qzE7Ruc
ugDJQ9Szthn7I9vcgNcUHs+rPTobvCR59dvW8QDhgcia1aSj89DhoMpUj/n0kgZMt4AptPP7gTcH
bUrS45JGri+f8jb4K9VRlo2hSaNKETEx4pcWx76Wpu0kicX2LZPbrwLC2eyX6OWrQRyI29p0NE33
wxK5tO8VZkNmAg3k3X8U5yepKA9Z4sBbSg3LtqRoKB6hCwkUVE6iqueGMmDJYrx7Zv+pYbzHeXeY
kFwzvjgjVMVJQyE4D0AX9RXPKlcQUzU661hzdaHfMZF6teveliPsCW86QDmrsOp8y4Ox9UMYu5jU
qW6DGQdSoogQfKyr935RMEHzqwNd9CzES3kABxmeikfK0ngiU3giWebajhmoS48nNzX3s6U/ZHpq
vCr/m3rYDZSK09xNApTk8fp0IBZuhPTh2nlJk58yzaE8sxnq7iSRp4MMBmDTYFGcNFiCusyEMjVd
EMlBXxX2ZK5OBHaJ14HE1mBYSaKyR6fGRDKJVhv/ezYhQ6InLVqq2hSLyke1ekkoadoPVBWG6FVB
edVcT89dQt7niW27e4qii55qrxLqjhMjnMBl8OQ1DDArsulmbdBB282ECf0EIKfd9fR8wH0FIJYa
ikAv74cowgs38l62CPvlTB1qLfx5597lQyHQcC0NY1F8EsmbvYMowDfCIBPVzeyPKDTxSxpeh+sI
gkDVaUD7YlayQA3ojiBXR8AWbOgogAR1wC5I34evqrI9sIC2oOmMKt/jM708C2u4UxQwO3m5IsOl
+N5523lXH4NOMGEk3iI7VS64NrMtuHBE6bvUL1P2hyqZy+hZKxpq4nXrZ3zeqMm2ABuxHDiqqC0T
LnjCvJtvBRv5BucUl2NFZP82zDAAuHeM53hrQb+XY08yHQFcD0q+iEDtr0rjEkSE6y3aQdwcPsP7
GKpeDvv2dfEIDNktHPxYjyS5eSghdfNa9rUV3jnXSGtaVH5BvXqSKyNQU7VdhM1bSnzxkrPo3Z1d
t1I4+pXKXq6MMslse2cM0XhrmES+ZBdRHsxeYU45UblkgtWLLVzah8OJjRJHURdsRGFMsS0vy02a
5d4PsDgwwKTXGqxCejygbCGOGOEPQnbEy0iciogRmG06enZjqxA4NPdwU8ZQTRLtb0qzn+3v2oSz
b9VsOH8nWNig60Lm1qntnIL8OkZp3PSC4TS7tom4MkAKBUTpaXUVxwlrDmvyXoeb7IjkeurlHAB3
5RDoAGGbFPGce6abrW5Hu/5F5hBDcYMgwXHUavro31frL/mijisneMLg717XrTwv+amfgHuj5EEW
dLw/w2z1CuMGYe7dflhXXKFBOJVjFZEr2ed1ZgQq+irrmMdrFBYhQB9S2qLcCPYo6KZ/JNkQySMs
fv//uPZ3sHXlJzbrUgHHujnaAaWMAaXXIIwcJNwPA8BDZIIOG4cX7EkOYgTE9itSN2gGQItgDKRm
hmFVsDtX5vwiLrl1DB3kEs3iQzKlxZhstzTSlftCI4atlLHsDjGMPa38VWBoqMIjoZ+b3/mjAC7N
2kP9PoviYAXy+knzsIo9H8wDe30fXbRkUbSWsgk5RJBOTzNiV/pUdhRmEdqx+AV75JnlEkxQsobd
21uH2g1wj4HL70jhi7qGLJzK7e7sTj7lxxY1j7qrO3I5Yu9F0gfkSPc8QLRMES4igvRMZ2Z60Q1n
SCRBDKdv6irW0HOP3Z8Yj1sdit/K6WOOCtrqgnlbSeOlzqoqmP/QKhyHd2DpzU2yuGjuU2BaJVxZ
P0w/iQGD7JavydzH/hivsS/J0tmHIfQcFSWemJEttlZ92IHnMu/bLChNG1b8RVmBxH5xJynqCGP3
Rt6KSy6nhumk6FGwaGArhv3h/z/q/tzbgG3w+y6AYQs0J6+w2hnyKWYpoJOm7XNk7hPm6egoDZIl
QVovZK+18eZ2nDsUwLBT5dnebUQ2I4VbjOrTlnWwAxLvEu51YL7lW7nJe6SsjhgKM/QdvZvcsc8Z
hwMtunr0IdzYbynFZMci4yspjKAfHtaIhxFMppTzBazFD2+Tp4Owic+yaJKwES0AaJE8LWJ6f1SX
hCkr2nshLtl20adsBLzB5IyDh9xc0BaDkmThsWcFr71Ay+l4dYar2qf6OnAX63/qkvbI9hWOCMyK
P4iYAP0GVozsoIBhFKakqYHrWwBkmIH3cyam3a0qSzd4dlGsfUAew2I9EkvCm8n5stBRIwwlzlwY
MwJX++yJ7UClcF2cVQ1OI4Uh/SKcbVM99gkhsnp/T+NN73hYyAbdlKAUuH7PiwVT6k2XpnevqkZu
Pc0B6SYuz5X9MQQb9JVh/a1Sbo1LRFK5SXBfYvMJOpnF29lQugnNXXlPEbLoeGbl2pDOCy2fqaoG
1OWiinBGrvWXc0JIl4mHrs5v4MmSBo/PxX4G39WkVb0igh/j/aPjC6PtzXIa8ESNKIEZcS/Uny9O
YRS6bLP3gOLiW7vq5X/ErgECndnOtpX3sITeUMotMMTzqWa3vKotK5e6AQQvfdobPeS15G0mgXrG
NYqXrYI2v1JfQ39fcoO57ijWQycWIU9kcbk2YgyYyh6E5aYcgDa+HpZms5ypZNOYey3aeJbJR2lC
nFOdpNqwllOdPfcLkPKoB9gCln/3fTY1bLnBcmE5vL3x7lVp7G7uN+1fEWI8Ao3dT2YKgVgmyIvs
EzTuJ3NGm1vrLk73zfb7USj+oUQUA0xEl5296tRCJu4r2FzSF+gCjiZFj6F4AKJ8fyXuNnnYyLkH
HLChZuEJHzzT6bJ+uWYjh1vipjBu8J9kIJXjjvxxwFo/InuCku7uKZwooTY4VxF2WZt0Y8uP3wLr
fNPOs0gwMG1X7T60J6kPdPYKSLDXFR+/vEpN4Z2U59FZTnnmXlOrg3ijrUu7FL8dpGXvwVCe2nPJ
LVUQ40TIis123KXRl08eKFe4woWmICM13lqlLquYCHGl2Qcaz/VvitJTFiTUeLlpfdAxcy1mx/lP
AQgRFW/MPrDzdo6KQNXoGTQjrr77LHRIgG6PWIdEzF+P4jXaUbkR/3dbAlFGsGIejotwRlEx+inF
ZE01xU/bx8Zvj1s0FAD73sF83mMAeR8ZNQ50thOGHtTFpnUUN8N0EkhaS7A/b4EPoV7CTk9T9fEm
cPuwfufiioXgm48MUZeyW8+uTz8tzvpktBkbbYoccBTxAEaf6KHn+vfiEMJk2YrzqOviGDGsYFUn
rMFJNeh5t84Od7yN4DVtLVlOTueYSUEFkhbR0BX4K3e85lXp20WyDUmukQYZj0IhfSAYznuVp+v+
Ue0OjFnvvixqy/+B6TBQ/9VuRTCREpGSwhjfVZtH/1BQsk2WBFoATLpcnuurG0i2g1xiDhwUDSDA
sdjvp9jAiCVaqALAEATaCQnstHcIZzJvfzPvlvY+1JoNQb7PtIx0oGeDLTRaTEeXogm8yvsT+0Kx
gttkSg5vrQi0i4sCDOdJrPUiK952iihZntfaX+M+lDQhzeG6weX+Ax98o7t6kMFYJlj5fMmXqtAf
l13p/Z9fsAqkFanFfDHZoLA6t1kWqq4UgBytG1zHBqjqKn0fzL/jNP1blct3KDdYuvhwiMvQlTbD
w46zkh0QO1lLHbh4YvLD/XwLRhPEJgFckfOOruy93+wymQml5u9vtjWNOQz6XUUNeWX/dra0KTnt
YdeuHZYrYcuDCeUgL384yjTX8Rpd9NlTlDfAcZGo2YqnYDVvBdSo4aGMzGlFPHq4xHpdzbBzWShI
sctc70XFrhBG1dptc+nakXaoVCxaP80vzQlY/d0cf8eJDLMl4cy7HXxQzg1J0pF6ZH2LdAUP6fUo
hCVWAMhALmU3yQ1ETG6qcPE1g46t3IkYP4etLZTnMKWIzOjAkiwt4aAXIiANR1K4WWQAYNvLdjfI
0mKlBeUFY8tfABl1mnTkogwmAgBAQhz05Ye+u35wWzsh4gCOmWhDPoBBa0qwHHG+aRvt5uA5BwYy
isZlRpsBzVaY52RX/Dj7ZhJDtuQyQDs4wMVgIP85Np0YdXTOijSWniMJVY5/MqROgX9HDR8hVeiz
fUxMwczdYvBR4tHDXLRF4E3zuio9Ms+cBVU56mBom4ZlZqBn4O7caMZEzOxtuhOnpja7WS7tKAJM
0DGzc17E5g7hg7IDCaB5Gykgu4M4INwosoqAE+3W9BxFsNCHfl2XGXnm4JwO4nAIK2xuEyBMgAZn
ZWCetcieZnFTrTgG51RSiYmCAZs41Xy4RyrsQLqOUjlhMThvDjo5ZRCFwiDpz/QxTBejCDJ1A2u5
uueNS555jhbTd5Wb2q8DgOuxkiuhGA4JEVOcSQQEODSHhBYsfZ7I6VuRog4TcyiCVuODduQqe+Qo
F+kmRIwfp8LovJGpEaJT1ygGi/sujQdXyd6d8TsZddLUIzFe7rYe6SEbaCDKAQGHa//uz7z1743y
WZ5BSO5vkm1lS2Fy2M4najpPcurzVfO8CZtGAtVeO79ShSb4bJphl4PxTulc/SI0dCv5g2hJu8CB
5fPJzan08jklup8xoVCIzT+rukFA26aCEfO2LKxMo7EqZObbkRl5B9RVv9YRBNQ78vAWHBDUUzb5
jciB3v9Y3phpGjZnkjKzuYRe40odbCM7YttlLtBYAOpaVYhx0vLFirgAf4xOSQF99OlF0Y/sQn+H
+oEi2qYCpID3wojRP59YtAncZLZSBibACuW3mg2/O20TYeR2ied4eSZVjSrPixnme16uL0PEG97W
KGCB+mintq+RTBB97c2aECiFKbJm/RuFLp2HJ+F1EcG+3WqZPoewsdDh4Fi79ilcAbBNBtHDOz7l
9EGQW9LEv2tgKarVEqZJjG5JHI/e1rSUhv3FuieOIsSwziQ8MGYLhu9rbr1ZqUmEXYdGvyiAk5CR
nWN/PP6TumM7vBN/2Bgc9ie425YW4M9B1sQq7XH0mffjCJgv3OyrdLiTDi2mKqt1PWVAqsdtHd4Z
NQWpCSGcoVjz28vGrek/WE/YNIKYQw+ihiRWxc9NBx2JXZN38+BDHeeCai2gmJkirmF8/strsqmq
maaCrUDzSmsbjv17fKfwqBv/YM+2WH93pRqSzjKHURdAC8BxaVXnfX3Td9n9yEbXK70qpjYzLeuw
YknPGGCg7nQ47L883zuFGJ1kbPJAzyQPMUnsGdCRUSmjzvITbw7dNwlve8TSYcsRknQzsIDwb4EH
fZEB97OvvhxHIU/qP/N49nG1jfAymae2fCerrqL9bbovXpLGF8whwUxv/cmNnt2HEqG95jqCbht6
S+Txg9QJf1EpA+K8EGMblt8BlhjNY9eK8OUKhOjO6xHLtp3Khfj/0H/oW6hC9L5p45OMgGs84npr
7R5HXYGiRSJ77XVGrlUAr1Vr5Ab6WPBMfPui2zBxCwBN69PevZiI7dgXlDAoDlw7fOPmS5rAUbxU
QEUOghDSZ3NqKxhC4A/T0gxFKBvNxjKy5QVsbsoug+xC3KJIfOFOoG3pRMpyFVs9GEVJa/enGF0D
S/jxQrxPqq0TusbGmI+5+NSVeJmAvZFCB+dGRmYEWnmrOoCQptX6pYxxWUlq+kj1vvuwneKfCCS+
sIWKWgTAfccJYw1lhKoVfcgJhgk58PGfpsdws1zJBEB9tKF+q4/gGYwlzlmlg724jTI+H68V5kB+
QSa6hvxH5iSlarM4vwwRDaCz2E22W0+SlAw9GYYZtEJkecjW1nZVKqsFZMxT9+4NnWWx6Ptwl+UG
phhUPUgatktmIZzSU+DlfNvIc9QJmJ57LQVcMc6yhAn7thdtHs71BtPcby4UkaJKE0reQOvrJHbl
Za9D0d7F7AR0IGkXyEgHK90ewP273wjYwwegLm3Y+8/R/457ilgGCuXf6UA7L5XMWSHobtiNYRh7
raqFsMbRRnC/amQSmcwqRCiIF20bOYfl54dLIaJUc3QaMFMLDN8i56IX8AUmMlLJ7Wh1o3N34C7R
fjIC5/8YezIkxhA5Jl6G6A+v/kdL5tnYSPKh05offaier57svNIdtSoys1PcP8Y5WGepK4C+jwiO
iQL9yMoGtpT+e6G1Ka484pNV9S6YtTxfIaSRG+rV6Hx8erHVHLmO6bUvSBODzujOGB3yyrhrDZHP
M74LLSGlrk1bJTlFj1/AwhtYbdOEVi6f4zt6WrFsC1ST1LkA5HsQPv/5dcZVU5ADvwy9aKuaWIOv
toa1gWCiYGBMg3HaEId/95pa5E7Cpj3L4TaxdktdFK2Ky3m0rjMDffzK6HwFC9pqM4s4Fj/XzkpY
5D/VNZ/VKfSVgZaUNYqvnoiuF6yzSjOci/tzZ5y/0n4PC/yqBng2YYoKx/BGbNNxvMJn2djThFnd
aS62iriOkvqVHKMKn7was9n4Om88VBpB3wORMREJe7ITN6ArYwRcZLBlCCzE9TkhcmoK+oYhsrCI
zbdsTzf0J3xoVBLVj99rywJnpxF4+hQ3gFLQEUTx9ST51om9DRCaVKTFSmaIc8VcUhZvUvZhUKvJ
8dlzggRwTU577VXUi+WWJtoGYZuaUVD/+awYg98JlHx5POBTLcISoKLdcVAOJzi+7Lp1U3XD1nZl
SOEv0vAnIyxRTUmzQlym9qNForITqj/dNHJ2KXyjq8NoFH1uLkGJ4k3K+zdGspieZYj97bh8lfDz
g34LD36j6RGKJO07Ey8iR+bB17B3Fn0kQbvVJ8UpVcXH8G4L365af9U3JJObNQU/4P3PT/ExVCq4
4ygL5NHz2QG33ubY3Joc0zmTd+t9MquqeJw3WAtwtw1NEAFh0FXmFhAzIe5MjnYDzVabqP2knPyN
ZNhbdQ6TLqMI+zr5v/cw9LZdtGtZCX7d5RgoaymLrnnguU8Y+va4avyNM6W0vp6OsxFHtK/nW/l4
W1pzb77NRj8pCrVkvLqZBdGoWYgpUY9lZWeeS3stl5FEp5RWnW4lQoqxEW0jm+t+BHvMob6HULa6
fnFtj+vAsqaaZL52kSqxNVI/VDWtQRgFvrVihXOmM90Kg9HuxHZ73dpsrg+xG1Jspxh1qaQ958jx
yuI1r7m0hi/aYt+RvRFutMJU3rvCmGwm4KXOXmtYaNVWnm+SYBxeic0qR5P+TXXAN1Gwo/aU+pJL
n1ANx4OySTZaaTUHCsAghVkyLsDYpe33sTV8KRyRoEsp6Hgq7S9wm0IYqX3/Hf4wkn26xS88BQ0R
3An/CUio0R3Jbc2EI7HIBK/0HYaUhoPTdyF42dJG/k//XQ5tSlwZ32ftEEmqQLoKagGCyyHymHGB
s4XoZcGsQ+5xbPnPsyC0N6OggsvmpbGt3lWc/B+fWjIOpcCa4uGlEdfwJQwwJSgDdFubdCJc+InC
bK4c4OCDxWTVL+J9eTITOqz0PH6E4rV/vaSdXVosKEzT+YG8M9IsTPyBPJp8UaPBHiiE0LYzap3R
Nr2hWIdBkakj2ZKvf+qyu4G80+mEn+U6UqbRBAaiUWp7zNLl3XfKYKPbZN2bSUEz2pNpwH/e25H7
bkQpz/hwyPpbzydCNWZ22v1fEN+1S2OCFRc+MmQtkhm+pg9um0/mvozgelYvSyDkM3Antd1cWk7K
G4kftcQ2V4b9bPie3TY2s1H9YejUYad53bw463XY9SQkzVnLsRdWbtHtXAxeeoEucQgvTQkd7WoA
TyyLCR7p+v9bSvrv55akxzmN3GYr1yMpV0ZXyR+EOQFAuAOqVEWq5Eqp943OVmTv5aZgFetRMn6y
AY0Fi3WS1yQ9pCqhGQzdefqs0tLIDkojc2vmDijwItkmiZ7X5e5RYE3wskpoCg+DY0NwWURhK60Z
LT/Gs/CIdeYxADUSNE8RLgh1+bi2A3rCiRKCC82o34Gy8o3bygLoQ9yrqtm9tnQ41GuRPw/4uiF9
ooawdkydjWcs573PnKyAbDxyOJeZ4h2+b66useLx7VMIx94Ap/Qi4XMCzS7MymL0fuYr8Mfy+OB6
ZQWYJ3M1p7NEBV+sTCul0zrMBcJm8/sKlWl5zuRIdez9+yEVy/7r0i7ROBjDqi3quihH1KAzVe1X
d6YZt1K0MLeBThSTclqlOPXfXdqf99oA7pollXsitLyQdq6f9clSRUhmiA3zAKKntG3876AyNXlw
XtQj4cPhCL55wMB44z/kXSo+a5oD5VftyCtHycye6scWIAC1Dd2ZKFmwoUogFDNI5IQUgGJoyhv3
dfkcmosBlKKO9+WYhmqA9QgClCafXtCxHFItTnXqHaiuLioUqLgiaIbnKqOZoS/gwsyFnzAjTvLt
CuM2mAmnYaF7x0/SbF8LsdXOm2d9ikQV14cyyM+AHrEdjHYla8GnQn+MReaDa0cCPEnUo3yZteQm
P6la84Noie/+yGckJoj6RE3+6VbD6P63pJ7rVZX5/WCNKxd8/4c2TigZ4r869FKprLwUALGGhMDK
GxotDFg5bf4WIX0slEJL04Y7FSFXAeEPPRs0fDxkGBr01LSM6V6/ykPrUW7PCYictlBqwhtbvX0G
glISBgs82mxyzlpQg5IuRl5kDD6ZMGwYE1sBDbeDsX5N6GudH1vp+qRSeYZUfnySzGB6zVOlOmfv
x4C5prMMqkZlYp2WPIIKQsnC+3KNYTyJ7jeES4LYgygRUuaXcdc+6pIBG0pzjkFOEdfG7uaiOTyL
JUEL4de7ZGL6fYRva1sXB+feO5KhhdTqHLEEMMH+opqDeki7omV6/LzgpYnCiTgn9rppYxjofACR
zHUnaVTRKFUz5u0Rdiy1z+3KW1UK32P8XC3R589bNbUyFAoKej6bcNcmJ2CT1LpupUq+8aMm0BwJ
T1OyDHPuS0FVA/Mg8lB+UVXd9Rh/SuEc2/ceTU3TmY849NVPidWk6S3yqmfWukHQOuUBbkZq5d+g
Vr0RgOqAF+Lw4aPyzndrbi+SBvuDGTeVS6nWimT1F91+ELSrH7tPKzHcaAcEzx+hoQaE7J1v990O
Ejw8+JRdnh6fBRFbsOP9MgBRxB/BeFsx3kDulHeUl5e9OPvPBCLoBsyJ4ti3t+0GJo+jI5+W7Ydj
D4rVToJcMsAl1veRWdlj1ruqyDS08fYCCQ/kQqGJHqtjQVXt8vsdMvtK6doE/8BW4Es6pV22EMx/
/xgn/YFz4/o+vCRkR4fxefgxAceLyW4WVxR1AmcpN4yyTTFGX5PvCu78Lsjoxejzgi4tTxHhAy1b
Zh1eivGFmarKwJ2jKzdailxypL7eRrINpaWsFYcL6DojUAHm8SsqkNYfpD7yW2hu2xlIQ87j4I9b
RXVorFFJn07VJU/PvL27DmjRES7ozQUrCvza0Ef81cHizoyZb+x8K6lqgTn+KYeVwJw0EanWhfQF
38B0zYO06zVuEcOfdhBkYTQXabP36rhoe/4GOC1N09RPx00fQtpvAVMgHsGkG+Kh0Y8Wa96sdKF2
2JtovBfjr3U/UKghN1nVLA8rDW70POKRTC5DxnKDdQlGngLLitnlmAZ2qN4Z9uXJuZDzjr/Xn0Qe
f71EChC4Xv4uaFzcktalSQVQoM5Lo3BKgOiAB1t3PzVFTbUza/bultrspP4KQ9tjjFYJHUK6BVrN
zNXlTXtffJ1EPnxokIiZAaaYB/LAft6BpiL7s2ZGPwyqLbhQJ5EDBya/RP6M9kazT1DOXCjgtuWG
UD0/AE+cWsJvM8JHobzRar4Nzi/2hEuywJvEOAq2KLMjGkeKbFkzxikBSStNOpYZHj6pFQ2f94HI
MxSNAitgdZiJZHfU2gY0J5qLt86FmGng70Nh6MaTpZN0FlsA3CA8oJhsuwxK17LnthqxLIWsS9c4
m26jzEiARObwXGku6Ay96YTtZxErZ/4koEoIF2L+VU2cL4w/pr65mHqrrA+0VtdYwN0H+Do6Vc2U
+mHzlxK3H/UKqUUOg55UHpVrLOLDawGHJT3Uvi48HLpYBYj7Gnlh2kSoqcbbpKtVyZednDSZ+iFy
zgHcIwzTgQh+xqGR/+nDmmMy7r7DnR+tu923Kn2utO8Q+VAfnrPEGAwkx2JDjZyB8srKqqYFnyDL
P26c6wt2uskTR+6ywS5uzvFj5gt18ulUW69/SkE4wjdZUc7J0KklzQIxgQ1eg1AFzS6XQaSG8x0v
oDdofU8RimBHiIwKwYuUwP+40sOmBLRpKrsscEN2P1W+ZFNz2ymcc9LMfxiXeh5iBft843EjcY2X
Y6lySmzNftdvCE1+6cUvG8ma9zvhCV3TXjke/z/O8dhIWGHSEm0NOzCf0UfI2vpUXA2ZjLq+BhiM
EmC8ORQwCklwofcvf2y633vyxiKgqe9CPAoffpDT1xjaOYenSfwVVfed1HZ+XgkCYDyqm9kVFIZc
Sow3nCM+8KXeCcqvaz1yhy/EkW9MN2vzSDq6jjeBGeYMiRpLGPFQaF8T2BEbQCdY6LWzbzOf6ns9
PM0q2bLWdfOWIF1DxNuLqyVTVvwsPNGUQ5/19VJlxkMI/UshgFR3Ng8mJ2QKv8zlLSsM7S6O96Tm
K2koykofQrPzy9cnWUUk2Szxta8qtgj3KTmSpZ8Pf5vHZQ1hmWXW1/5pfh5yQ5JfObICIxQwAY3T
BUdSm8HJfJuPc7ZFhlMVQIqhScBDc0IWqRtHnGVRNxC0lATXzVzFwTI9swVU22R65THeF7GfkxKn
VlOQ9GhCYM1rrjYHTMKrlldJV9XIZZdHgBw6WSFHlHjn4gyF3ziLrwB94wEVd9wWy1YsgaxEVhua
ZxGfuTaf8CimbfGLkc4uosbn4MlteQfHT2ADw6DwMr3xrkJPseRh0aL0AC/S1hVYE5ndVqvcyWPe
aOVT5AdTbOTXU6UQKZgRPedXw7hAlP5Jv7A2NTlRvVgODwSlRUCGtXakgl0fUthwXtMd1XUPZPa5
7oAtD8KEXoBIbRWwAQSU3jP2ObyIr8ubpeWb8yeQWbChJVouEt+SwDk0XEaiS5nO5ojVI5J/T1Uo
qZP/L1TBxkRg0Yh6bdCYfTfcy4Sym03A58ILZUG7y3od7EnDILmaa/xIC4g2loQxC1Hv1Le+EePl
lRYb7C9GOBp3OceSQH6Uixt6NVxUuLe03YY4ibyopw4nJ79NuukFPU/44WBa/p+CchceBdUZQGrJ
5j/1DlT845pwH3xuxtnIbwASM+LlQm+aQnRESNlFAd4mzuUlWl202EVkKFXUtmEDk5YgpB+uvxiu
FQ/gp2/T5+gnxYnVp8XZJ/7GfLloxEf5BAIukBmgRjKWoOntOb3amiSpnURMHawuMPnWzjyDLU6A
JUCA3wmloHeDas6ijJFBbIyu4/T/+DSEAhHXCLF4CqHs2AUHT+INrAnulC1bI6mTpBO8JknO7YLv
BmUrZCr+VyBxpqA/+5Ol0Ra52vHGpPZBcdiJyD4QR4Y3/uEiY9ufEEBL3PvY+TdGw29LrcWJ1WKh
zOcDVCnPaEn5znS3uqt5lE/2uNdNKnhu1R2WwyvksQId4rrqn00AtihA3JrpRZrhVLIO1LsALamM
cbrXMxfz/cfwzUsvaPHZ0iTeTCgcC/E6NSTBCruJK59leaMyZSmb5cXC7A9DlIIcT3cD1uKCsFe5
iYDRgDT/y7z2tt1DH3/lG4xCYH0i91nRCHudzdVrb4FHH/nJ3bHMk2wA8XU6NwfmHfitCFaNkEQd
Gp3+trp+Hs1wu15kKrIq715Kh5jMYKz6sTSAz4/HKpdowZzBDT18R22ayPZ3tt1sbl0X51vJJ9wX
g8sMAuiQYzvdOqZZw2WRh14uzsT/YRVSyfPN7/8dx9at8DKe4i7QoW08YMJTXpMoKtQWUCxK8KNZ
CI42PatTWK+zqHdUJTSvyPJFkZZqTWSmqjMhUNoukoSarS+0KaHDllNZItjPwCTkY672ZMU373m4
ZQTgBtcCNJm3J9VgSW6ndZ1K3wh5FU+XGm1pD6Y4JjrXb81YpdWXqqNhdlHFEFys6BZwgSU0vrr8
IUEjncs3XpJzxK3mIH/DFsmmtLgfgHdAaaMN1fMV480w3aSCHdSguAafu2QMawziy+SGGqx5sryZ
K2tHuSpR3JzOxXEfo4WDfGftLKipVeNvh7Gt1V4heEzZJzDBJAGUM1NWZdaZTiqxarXY2nuBcMJ5
wcJjgu5PFr0c4Kv/Ym0b5hRtpZA/R0Vx24edgnLJY0IMubB6j1KJOeODcvdVvPpP8hV5HmQ0cZ7Y
Wdia5Z7IjgdXMD8pusBL8TfUU/UEJ/BTE+hS1ys5WhHtFP7k8fG2vStkSMnG46pssy3we4/bKRS9
4y816NH3/18/d1g98xRuZRDrMRR1cGHTdh8SHZMcGHWdsnoMHIgoUMja5m50MSnXZ3tjq5I/aqFT
p73AQWrIh8FJPFgrsYeyXo4Kwp/iuwODuTPQe9wHoV/J4dh+kEnmHPg2o1DHPy/Uh8Q0MayBTg/F
ftyFd4XYGdt7w2TQGbv8mqakJJnh+fyaFzqUybUmQbWopMKgUGV89tpbN8x67dWL3j2ldo7fHE9+
MxYKYDXMUAMaf8jI/uTSLbE++gVLN/AFuI/b2bV8lp2l+JmL1OxLKuNHO4owjgj8duQ+BiLWbt+W
/0nMaNiSjYyBBT+aBYysbXJEJJ2mVVCCFo0zC9TsCRmV2WeiBRR8aFsLPnS73m3sLoc5QH5zwYmE
9T5c5l3CKTjAIQGi8frUgaHhRmrpMEgzc10r0p61Kg9c3RT9VY8UCVHSP3eP5cZ7SczT9b++Igrc
PMpbQ+fp2KGUZAHAKUW0B333c2dT6qqI9N+WOciTv64XJVVfrkYRzvhJsSdLp9DLSOzzKY8BWqcY
E2rIV52pUwjucmsiprm6ME/IveCJEX3ItfPKx3oI1qlBHd0elGnelF+0ExVzKiCsqLLGcCzT3z/5
CMSIFMstPyMdcbl/51MJx9reM388lhRZp/N/C9Jjej2PiVsWoskjUGk5ZCyYbn5meGKBMlN6UJqY
oR92oia4zvOKPfelp+xxH05G8UgW6hNXe5NXp1bqNE01hHxAxgpW3ZeZvxW0mBrMznz91CGQYHx/
KqRKw2W2Ie/84Tb1jXtuaHMKjE5OWJLqL4S7rRMx5/qjrOD0IMhFs44oqAWLMJkksuEJOLRpzUR6
n6xXIBdi8g+M6/gwo7hzxvInX6l4bkdrWB7Bz93FRg2Vr8pALtwhB70mnMKvPeFKUc8de2NYEWxV
KlYrhYzn05I1ewLWBbESzspXilO6l0FIdPEEo7uChyfG4+jsbWNOsjjnsLJn2i1SdmcSbC9SXkI/
CH9r4AWIy5DgS57R5KhK+TbCbC1cuedhODbnKdavcmnZKrn7Lg5HFl3gl3+NWJ0xE14SRUx7QmX6
t8+TdDoLyg/MqeGVoRT5gMjnDwoHhz8lByrXhbhmrbDNXCdVPTwnR1SNRFk4Pik9nWWum3HZwhvG
RHq8W8iQQn5ekkasY18YNaOGQ7kygvNd0TCh+zFzO0RGOy8zze8FoJm5Oal89sWh1LF4jnQqFdHK
sFbQIoE2wCWqOngytFK3PLadufCMOdFr+wd7WGy8nvzDFV0ek+motDdpijaEeqm6F/i1iBUD1Vz5
5P1S+FfWbz6flKhcXKgSImEKAg6bb8ZorDjZvcuNEN7w0G7GNj5ka3mj3xhsI0u9jF9ubzJlAof5
vIuSEDzoE97jCDwNy56T5YMNFHSDBfdS4MwLQ+CCXSdZlb0UoQlixxkCKQWPmUs485CqsqzsI+bY
WoidamK9jCwXB7IuyRdS09Mf81C+wfLrvzx/8DTvqNzkaqIZxONgiNaq5534pvmGsjsKrzj/ZXeG
a/oimVm2BUYjloAMC/QspnNf1p/ve6CBkI8aeCe/snathKldcAPpu8nwww3m3QTv2eWyOB20uS0r
3B8B9EoKr0w8OQ1ao7UyzntRuLOkAx8ajRAXQreW414zc7XnUHqLeJx/+pBoZTkq4B6JCO5iuFtd
O+M42YHBziU9QX5WUlgKv7hszb603j9EW6+yIhk0Fbgnn7wbksV9t3Gs2vbL4tLAiL4HEd0IYLWJ
KaOlHFDz6zr5Qc0rTBH7X8NaFTn2bAacHkVfL+l3eZYPS4gR7xv1ndYTd/ugl3xikRjDuBc6Xzya
4GydsPGe00N67HRkJrlgLdN34GpalovRvFTHmdAQi/zTCgQwCMafl8j4UaH1aaMNSXC9/99+0IAJ
RD3Mp67UETs3b3n/eC70PkEH/7zkKqFRpz2FXzJljJHZ5UXoyN9gA4dqbLcHtBa+tcOo0Cm0HcaW
FhRJIE4PCLjaB9poQxa7oHCqffxVKwSJ6CkLU9vAYyUN3RNN1+1rqzoZqSwrAqi5invWJqxjPCUI
jkLgsRwWnYsz0O475ySv5GKnHB+xCKTzkwf511WF+zccXdDHWfNQ8Qvc1niZxwvggsdv+KRYoqvA
ZyCrW/CpT+JUmcQc5DBD/ZnuE8ppGA4oGSvAwuou3ZP4XIsnujbTgVPrcCYtWfZv2B0tS6yN3Z6j
D8DJ/sqG7ZDglgAiJ8d5ZkmDYWiF2Pe3nx74dm3saDZCWk49yzEFtj4Nx7xRmuDs2xv44B6GMAvF
0i71/l77lgAcJsKrNZk+rS+zQ3loYkhGsrIxRV72EzDvaTtSYYbYb/xT1CXLPhfB6o0uvjkzyKb3
vpo2iIuZVve5gCV4OQF/irjGag4GQqpbw2ll7ZcktcwxIML0tdMUSDEt3kYvL5Q7ZKQ8nJOZA4pD
hqcSyoskH/FLBAQpe/a0FoUG39zK84MHrZSEgxwP+LksiTZaHqw5sIcE3YoXWcVBAxR9cLK+Sry8
ENiTF2T53Nzjl2xefinz5zCL8IQdu7LXEZ7IjdwFP0We204prk+8xzVAC9R0PCfaeu0/PmZC6nyW
gHp3Fji6arrQhQlCrsTwPpe4z08sKYq/xSNsb772rwTsVtODTXel8HkQ7bklQQznAd3lzlvyyiul
HOVozkM2d1Yklp+IQAeNrcpYOUM9z8o70FOe1LDtw4ZzgeYzDJG6NINktckuTZYYoijMPiIwGHBJ
Ou4PSDn3UoWXdJcXCVOHkShTRDcKV3MxQbn4soTnLALOlsvI7O2XzE/gYcGBnd5mdY04iFKn89Cn
WNRH/FlrdWDvHUUW2jsW3jstVCDdia6LF9GGlMT11I27ql40cjLHV9B5QezXlQ6FXimv30CZYG4I
15azTWCpjMr8ABs8pUctHGXlDPZDVAG+Qz7+NUtt5AO7k62gPhcSj7h+Fj61TP7ovqvkpIShQPlW
C1j6prQClr+UBy8eU/EA4AD/6j8gZXYbmECwDmzhLmt6iWFBm+2A4wadhfIbTfv2B2JkwSKNY8he
COma95cXOCsibkEAD3mnhEbzZE9YDciUVC5WC6pcBJV2c/tyGO8ibtY/Fm7+SA9hbROg1kb0LvsC
xbqStLHdV81DLJuiqiuEZ5LsQ6vzBuk395oGtpDl2MX15U42XVfnIPnmgmwpXJ2W0Ef9tG4QkSd3
bkqYTe0No5XkcHTKs3HdWorLhfHUKyXvPEieySbX8Ofkh9gPxIXHqSXIPR413J0qhxDsZooQ3kU6
t6Pgqu8Q7mBYlAUjZTa4xnnpu2opJUHA9ZhgvSKIy6W3xjLg/efbpwxe8p9NVIwIlmo+5KJ+7Xy4
cfYMMb3r8Xvm0AV89Zzt2grSB2k/x/NCguGg3OyDRRjGHHxsPDmk6dEvVDiZPvycr8UADTaRofC7
835Wim9XYuVR4Ur5/UnVtj+oqz1CWSBi87XS0U5E9weNWdIQVRN3iKLlzQ6o5VFecgtHpFIirTr7
4VMx8FD+YF6xmdmvUCekGCFwiUd4ZHi6IVveQjwU/9wQiE+jVsxRxSp42rhamIVpKu13uL/vZQ9R
lucgk5A4RCLr+wY2pF7MVbKEykmu8O/ZBsH7HlrZvA7gbcEHwX8DeOcWarn3NM8O+Wsd3shG+YRx
fFjQPytr0oR+UpFV0PEA1kc+9iHY+6fawbRZ51hky1Ugc8GGGcvuM51SR5gwVN4RQcSAYvz9Towy
YZjgBrc63fRpBx5wBoBXW4L/PqewooMRqe3uK+lulZybL8b5AOOvP1gmBvDAuo5J3ZQEAjgYYHvt
MSJ96IQN9pI/dBMZZIAtNS2UarX492qWGWALOsjR7aNr0GHZdqHL+6vNNyHElnwjoDCrJLKQlvsK
/nIUGVxG2Xz/J2yQgFNrRnwAkN+npXcWA03zU9xJ++IBRVrlevlqzFkWRmK9T5mMUstwiDkEpsGY
qVtwQDSeBU9DgBaUAR6I6t2ySsTSVxNgLHTTkdlLrV24oYcSSeWqeel3hRF1baMJmyFKN99geNZT
tHF89l8Fxwt6C0YJfVLECmNoO12sCnn/ADUXAJdogWu6uurKdQdjEzWt1EmkmE+0WdOiiLHRk0+Z
fBCFJP4e417BGmJFyZmeSkb8NBQ/yv9Fv38h0kG4TEjThXR75nQXSeCnq4rjNYS5tZIeNSWdmaQT
KDEr1a6Uu3+PGNLMD2ED+E6ZDHBYE0YxuLjMI2DUDpq424EQ7yjEmohh6Yr0df0zSnxFEf3nJnhg
EBN711NOz7e7UXZgBNxw04lzXpSwtPj99hAiqAh18E3YU0656zljVNbmQLle2PmHJWkbTStzBdSx
Ga9Cy2eLgMCIcD00BfX7CY8emRF0cpMBXUi9qXjVbNrqkPC777wBnZE4NTHP99ei8tJ+wunCaHAA
mR1rvRqxl6KmYBmUj0HlSh/Sf8nQNdk7wko7CJJ0MCWHrg6HVXe+wbP13HfF8GSYysbHLKwYU9rv
6taQn/hSs+CroW2tVVmDvLaswWaxOy4o46tfWW0kY5ydB/QPzzmE2vu9SYYUYHyI1E3KUgXbqN2y
t4nTBukMLjD742E8qrFG3BE5R37ljY9eLPpmfay+/E8xHHsIcBs+9kPPztNM52mXQVJjUWVFUKnA
KKTsGcDQFv31uTQQdFwAXGmVQAD/7qoiw+HvogfKZKk2jiD9dDwfGy2pDPCM5SFjy0ttggnLJnBz
WmuVkPfwsCLjPwa300abcnPp2zqObUSx0th0crYXWRZbnj8I0Sjaqv8PWxFmpFYWm2AW4wwsMCkE
tZ20WcQ/OUSHhEwAjlBRm65CCZDmd1Lfl4ka34DbOu0CB15QfGQw5MpDE2O4LRAmTN1hHDzGvZ0L
dptb+l2kOHi1IvC/96x+rc/Tqes361ALneOn9YIC+kNWbCYhRrgs6AuPzP+gGVM90PXKUmz4NUMo
cVDcQgbfqcA/EW0s6YQ3tk0/pjuHKFngug2YMF4rClkjGYa0HZgXrD59fQz8axaxxgj61/2c1URO
mRd4noXFdxtXipYk++vUQrPPOp2yp1qrLE0AXRpVW4ooN59JYXWBj5jLJAsDhw1aniDd8mW9dPyp
GWe3Oelvl1obFw0YrHnVrivb+HyHSiFonl9sSQlGfsmAsH40OM1QdcTBZ3UC2yA7b/D1yhqW+7G7
VIwRi2JcxaQHBq9JS2hWus9Sq1y60Vls1nOoun7s+IJiV3Wr1cVnzpHRx/wKJZCsNKe3LwtP+My0
vxAtpfWYK0MPlZGF0ED9cI8hYzKD73f4fci5KFfLoqeoj5aImdpRzeWVVKxOEHJpEzFxaoE92vBA
gGzNHEpx5PibxaeftcVogL7JeK4T/XEU/h71wnANb7/UdK9M6ZFDarhIliWte15TbRsyezOPWTyT
wLuAtjmF6jnBeptCwM7OnTrcqlZfp28qcJalyU1yyyVh5dkeDunYyeNLfy4ktHucAUwmRuU0Q2sT
4+L84vGeqSpcGDbydqmocR1BwYLsQTy38Gk9I8EBSyuQj/bkmX29y1JUu/wFUwppjhXYZm+GphZp
DMzgR7zKREOugSWA0ympHlJUNvgD4rAeGrsFqXv3KxJy4iP1c07dKE5NYn0eVAuqMIKp3SYICWtl
G2IQ8pPMajdzA8u4a/tVKFgRpqyQ78CPXFVqSMXU178Ew9vHOzakveSq8kvjLiLTtVbuxA++lDYR
OL/blYs6okuJag0CrVAD40QekcfEwY8oAv4SPWw0pGnXo2FmZeHCI5bMTxPb/MWeiytXNmAPToz0
TYiLKemg8593GDNy9CZMq7TAXCvK4yS5gfuRJSAVjmiWbO6/HPv57YWATwtEMnqGhnAbTHj5GZqW
eKnXQdC3Jeo6pR0hzjshR9gK6Jxmfl9SVn7PjbrqhK615nAtnF2Owzvq7KwMlY5zagbxpojCU2UG
pE5s0c+33W90oQJfju7pdvzBrHL0pTQERWhjg/1UgvqKuttavw0y4i+RbtHmqc0nXtx6N/XVxR4y
gtZbQIsBiuQemt11HugTPhFhyblUN1HLI9Hy/kJLckB9eEYfj+b7We1M4fQBQcmHOGLRAi9Z2Yqw
wpPP6jtGscdmALKgMj17LTCpmoxq0topWmuSlOD2cI4a28Rda3KtFz7NiTQpjj13v5HiKyKdXATK
tHQz7x7u4AzaYhcVBX9YokXj0aztn+ZFHvi/oCwf4LbMPwxlPX20CXK1clmL1LF5LRU5LcyD7IzS
rN2Tna3W3olpaM57yakTkKM46ed9bT42eOARVjeGvWcV+kxEhhZKROF+d3J8U6M2Wp1osiFsbi7h
P/JLcNvWuZzhFcEt50kLltjr5/AnFAgNiU/4uJq8SQle6FkjaO5/txPord5T5oTXsxvbWMQDVTrv
fWeVLYC+qfhOlN5f0epM5BFC/KLUq3CAFVUkhQhfyDBN1NIeTqz1+djJCfpzhI6Kgh8RcpvDmGqp
oYwDkhEM9Fzjm//s2D685v28w61BJLVfc8NBehe40fIMcf3exPG2Kaceh2tjWbYO898oUXlb3Tuz
MUCAXBs7tbY50fwvynXBQrna+JBG3TELWTVP7ciPm6Abc+YfaDDL/JyYsMW6O+uxTED6/9U5c4Fw
F2H3S+mBkl14fOUozEnhqXY6vIYA3tirJVCAAhLnWru7hCyEU0jDU7grLOQI7ViN/TY0EiRpxK3T
VFbEW+bLYdHGn0avse1++Is5xQrC0wpVEKrr9LaTjGLdZOmd+eQ5yKbydhHzCxxT0X0NNqL+URtj
3q25zoV5Xzf9cVv/cpwzIsi0DonZT17It5Mn8rFAT0F3B0oxParbnoavqxtLk60KDBSHJlfuNzyG
pp+h779Y0c+Gmhwx+1OVuqtvFdtgjU5mcJSk7EZp4c9pqcQIhHMlALE72VK0Afj0vVkJ0EmSZxq/
WOtzBP50Gn0o4fUm0px7WLu4dL16x9BJRs9w8SVA2Ju7p+kiI76DaEs13uLQovfzlUGHCUTrAem2
tI0qAUcGM1NQJAgTuHimR/aBe/hc/TMRHtq5Tgs6K2+cU/Yr23PIQqAeMm2Irl80Oh0Ngnq496+o
iP2hBgi8zNhyVtz9oJOQuYa6fzL3siRKLaw1E9cr9d+wC9v2tA1Rrki7E6k6K/LhlAMYyiqCOkX5
ObQnDkNkYPwG4Duz8p3l9Zczp17qWb1tOQTt9dR+tS9v8Wi9bCtEv9p4vIVhB56F4LfqAZOXVxwa
TApYQ4gkGpzD+ZDQtnGYfmXsXuu6ZnIvhAp5e7okLOEhW38mB6k7prHrk51cCIU0D2WZi2tqGVEi
S/gT22lNN6GBZXx0el2pFr/4KzIKR06+lnzlJXkeTfnDKNnuFz78etYZaU9EwuX6tHPTXb4KrF5I
spJ65TDMaa2x7moNNMkieGiGbA/cQLTRiqGcNdzkb/0FU/PhOWteHMIHWiqHZKaxlZ5NezAiBVvN
OAEhH/PH3kh7dxwCHoxPvtYnXT1VoHY5fKu1BMBvhYVO3g/myR2sQL7Va+CWXUothyQk2IuhIqF0
4qeq6YfeHtpkTVa0+orQBIgH2kkkgNUOnbwOr1izWXcxeLDyTkSK3TmBD9tlS/6qes8fmR++Qboc
eBY79bXqvpU+JnOLhnWDABwfC761SQk+I1KpycWlvjNXtj30ANbtbpEy4BH6d6bFLwyH8Zp0zIx7
xLJANqp9GwJAgayBJ+DvGaC58SgrMjMUJv8RyGdt+e/m+yuuq2HVnY/7ZZ6Gmu10aEOWna7mHPFq
j2UWsEGNNvSOtcNQiEqbyO2WNSivRyrbbogVTTbQOmsmMjM44qrlVFRIKBXj2l7XgRHWGkLVMU1r
poVjrH8jh+OGUqVD4p6oAAkxXqUiSA/zkyu9EjcBx3BgNAlZy5G3E6I9NB+FxAO328cywdo64q41
TQSenJQcQizC8XpNfG77y+LV1u6o9IS4AMdXTCiYrfsXusDQzVArZw6WPfZVllHV1KvOjja2/sGt
2G1swG3B4p7IZRmyOrvw+aOANbOiZUQzb72Hg/XMWK3Z7DSl7QdPGpnHFJNCFKnUyDmjq7yUctcB
kgEw7d9NsfaBoGIBxkeD0XoTYJGPjTVJEXyfJVdoX+CQpA1bxETRaIIVl/uWQy/PSBCIZKQoXRLE
a+V3DJaXGYUvVoApTKvknKAsFtAGxgtQG9tZ6OaZ5WNVD6Ff/TW6RS5n0u7ZeyBVvJei4O0r9wl6
UFiDWdk2jb4QKLp9MIqy4OSIH197N/i/jZBZBFK26o5qXS0wf++K0Kwh8zncraKlk6Oiify8gryM
MVBs+MT+PRx+dC4pwtjYFGW6jk+3jB4unP8mzANgs7M2fNZo7geTO1CiWTnbKkFpaZ3P89zST8YS
JOr5cb6bviRnLdnwcPOhC9ElNq4hEMX/tVnocVprkVHUD4J/Drx4I4dLbDPXND7pc+xE+QM54co3
WNeSdWmtrkQ3UmA8p0946ifkKcdHOZXqdNkv+nrIrA1nJZ0QSMVtoB7IgGQkN+oa1gn+jW2co2Pl
Q7U/CubESlqYbVYymyhF6pr/HK2Kbf9mJWWd5+gbmLKbIi5yYk4GRnCxLFgyVvAGPS1LjoYQFYst
tf543fABTZKuWBIVqKerF++3K0TIJ+dsIefZPsVTTGS5zVTLQPC16zK37UoZe6RbBFHNNG09Yq4c
BBdgzBiJc4i4NwcEMPhwqMJNlTGPoo2o0gkUkkI3/nOzdCIhH0r8eT5wSgcFYMTnlcR+6hsSM/5w
antEQHY3Rs3LMUbxgYBXYyA3xZh+fy0N9RnT5ZkGxrmRRLG7LTYh3uhC+n2mWE3Kknp51vZ3zAxU
MpjeLEuDEF6ebbbII7jfRbXnd/f/gG3by4ezrHy4zWvAVfyKM5ZKay+SKHmaixPZW1uRqv9ekolp
b6jGn7b1T2E9CZpcnjmrHt6zLBkQSbQpaB5ux6dzkvyW+pr2tbP3k7RXVbvpcHiL/uFdp5NUMNJN
U+nRA4eiIHwp61wJ0s8FZ3BMa8Gq6UamFRVrsNLvLzcUXbw9iIcBcBkbk//GlbtLbk+OC13li+AU
wTrg++hBxTzv54CudYBMEWa/XqkqstOYOgOv37n6rd46MzfQGg83/An2l0nhDANo56VPazBxQwQ1
IVn9b1Cx0is11mkMiegr/29nznAqOXPNul9c1kvOAAG86Gyv3YedwJXrunN6VOZkb1f/WIlS58Ac
2WGXLX7J6ULJZgRZfBOk3oC2ZMOmC1Q/qjLc5JIWTUmCe5bS594txzhR+nLFgnDM4yejJd11Hr3b
E9c1cQUSp9j9kw0VZkB0QEokXpk0BykZGkxI0NkczSA2y28LEtrog9cen++9+5umwNGq9zBGquF3
tX2CuzDZDA8ndD/O60puiKId0o7HILNQr5k6H5otai+Hs8VY0Fq8RnDFtwH8c9ikgc+Pi/E8p3er
46LxLOZ4W6vHYqYhubLh+bL8IzgWTHGBmP1hqC8A3rJad02+sfFAuS09gHMm/D/afuR376A65Ni3
pZ6ByoUKueYKUxAHoNouVfbzM5Uy1JBkH7ETXVfRqjrSDSExmtCr1DdJwO4uNylWuz5iDeiTnHQ9
MJqixZa4gbsUEYGpuMT7n7aGVsoevCKQyFqdLEdARf8eTJsZPKUE828VnPqBXZPUmlHKZnysXOLs
q6h/AcGAtIHw1aMO01qWM8mHTTn4yPIA+SwZ2HL090jqurLvBR7mvW9+Fm8VQUEgzAa29tD5l5Fb
lW9HT/Dr9UJO1/ffzXHNETP225HLiPSjqyboFQozQqMvnorYBgQqmsRGdmCD/5/S3iGEcf6ZB4+y
sZP0vc26zl5gIhnG1FA+nkA+xmDTG2ScsLemV5j91Nys07eFpvErb0COjAoZpNae0TAbTD0MtSRI
P75Jk1IGKrvbXJaGX9q2VRTHtQX3KoUpu7xxuPIjthVbkGG1YwAAx0EoEjeYSDciYr9J1eJm9RtB
Qu4AtFvwsyU4pUlzGrDhKS1JN1d6A3QvMxKUviUkXW4rBQGOjS6pX/xnWixPQVBPjEEKkbjEt4yr
u1aygozOMlV77mJ0Nc0XUpcbVInYrrDeOWY5mn2Yf8Xky0CK/l5u3bOGrRt5Gq9vS43JtEuuI5+T
KglpKbebpGCTMrE6xUOfjsO2z0OF+pC8DXrhXI3E6aeChXuO3EGThAe7T7YUQ8F9K8qPL0k0Ta0n
BErcsHP1+KT8g63bcx8WYoT4a3OhciUoP01/hXtLLr6hv1djf2jECo9z+whWARw0eXKoGhnypWQt
3t+OcnTOnxSDt3mcX1BSuk6RtMinyysOaz8k4GwN702AGsMM1aeEOYPStuXdIlCEwxHHU55jj3z3
KGDyJ1hpTP+O9aoyYqwDhVuEP4E45C9PLA/lr5BnDYYwTtKV1Re7uC9kK9bdIx+U7cBvme37+LS9
kI3Tx2hRqOEa0f54MkU4I46QbLZOeHb2nFfzpTnv+yE4lOTJkmxxVWyNMu5nba9QAc199CjAZe8+
/PGzcRYCcZ2JZJvlusUj82mEblDHfm7DerQZgyR4BXVQWsmA/+MzL3E0U3875braE8DampXroldC
HsV7JyaX8d0m1m6lrA6GmvLBq4wioLpzgDmC+EVRzLaMztJLcX8WqpbA0IjZeVjxsZzqx+dX+yiv
MD6z/T3/owXd/5omU/gfuaX63x+a4LY1Wab82tq5eLAJNBIlkcQDdN5AJDfxoFKPSimdOUAoDiZ1
miRfir2Z6+2Y2FyYgmIEBT0MG/apHXfYoWTvC4MaB33XwbaDHfmthbxC3qff8wX51mmxp6lPPQLV
BmMbhPu2Slekdk0YvoG7Hh17uN7OW0dPek8GC/L+LRjZlPEZTV5wyOzFWALinuH3wFL9f6Uo4bVz
skovXKGlonYQap90DT5ThgCklg2MmmSTGBsIgndWW3tCft76KgCfb6YK2TVnaMb4gl+N7heiTNKC
JUBl5y8iwwea8mwwTxLCB0mUIpsuMmUhjl2vQholMsBpmfyfAa6bWwEgNYhsU1HqOmpXMZhw4McQ
/CODP0uZmCHEb11LImvjt3i0h7WRHwtdSm4y3NKUGOEwqZeLbXfg1J4N1405h3Renk2TLqv3xKol
FcdykwEV/QQxqdBOwFbqpYBgHBF5RzRklvrn62znDcE6yRrGo2rVjcqsUyoSho0g3gfmy3k7Bmt9
67Ef6tCmFx8RjYF78kBKh6Ieh2FsPBIzE7K/RxiPb85UzJA5Feq65hKzYKLok6ZkkPBOVhtc5yqb
vPO6fBhpN3P4xUlhXkZJZbcKj33QbGLeyAOMLMxufoPRoqkraF8BsiabP/1l7Y2KEnytVBZFaYO6
H3Bgv624LX1UOu+GF15QA6IBAdqMSqEnbxC0doXD0JbHrb96ZB9lyXzIDzB+9OH9Kb6zPsMHpScw
87yyJAZShY3uJDvJGW4SkcZTMVAkDAuKIeyeppMFo2S7rDCFWW3+WhgbwNJbpqC1/nRnvCwC9Il+
3zJdR+YuJZdl9BRIlMYFAiL1DBBSllDtijKVebJnRO2FMagdiep6IZlozQyTKMtRalkmy+57wfej
MN1gTpv8rK7FbgdzyWm42VmTFBPzVoEN/hJZWUbsKkxgS02DZpPpi3a5tdPke7cRbOSSiNaVk3dp
8TdrQb8eZNNkKpeRX2ZGpuv3vWkceuGbFP0Vvmcms/y+fLlejCyp/tNojA4Oi8RsxVXNXBDpLw92
z90A7Ng8AHCqHtsDaoK9Myqt2RZGXacCJp2IaQMJ550Q4r6lwdKSHWN/VHwo89AaWI39lSimZT9N
fCJNzGPEj8P9Nrt6W+jApwSIUu6gEOXO0Q0lJm7tBwRP8L9bpyMFmdYh2R7sKH1qBSLvQilcPLS7
l6aOz2PE9BOcf40w4hc1V9wsiGo/qldQpPBgGD3bQgxNeTglQ6r+5RMCYS4ccf0JOEUeuMtXG81q
KHfjg7upV1oSfxMTAM8Anma7Q8tQMQbk9bflMVgxHlB6AXn83P06QX+70q9JQ40SVuGYkx+iVZf2
ssmo8LoYaqwpMDdkgNiQqsdvX7mvIQnHKA3E0yFffvVgW+X0rGcU+RizkY58XnXAHupHwbt6CubQ
OfVKSyvUIc7++MJCkSxYI0vA0MTWkviBgNe64pbbl736lxfmZ0gex+KVJaO+u/VaoyFPUMIwAkp5
BV+grMfLQpVaFhOj6SP4PGU4fM5j7Y4w0Lse5sSY36RNxlBlNFDQQuyFS8s2+FpBB8hFwVnyMKGA
00UooBEvAW97HEEdN79oVilv8OSYak7z69vR2C+t3aSu8f8VoYb1kil+LylbDFkXKDHrgkXAgify
p7CvXph4cu2+zWn/0MdRPYVhdDZZi5Hm1VoXc5nV6W7waURUiYzz/U2CilluCy7Aqc+ChdnnsU1V
/oDCDL/5Wfip5kGdwXVeMcxvHx5msghtBBQy/S1VhOJRFDqx2z4JvPGuO3uuj+kI5RuRKNS5mW8s
yTfoDSXZdMZnOKkwjMdmeFtU8PgVcbDEYd6M+7kZHByU7+0SIYnm9UP3JY+zo72YUGbbSzNsxGLE
m2k+2s7Mzs4lFLoR0YeosPfolwl6HWehIJSch+1etAf8XqvdwYLudv+OHnk9x+jaj4L6iRbM5aW7
GBt4HAdSCmARPkY8szRB6qPhOsHSt1NXpPiIBFF7XRpi0EPp9wE5BvKJvlsZcBAsjqgqRuWR9+hp
zYw/v1AzKzpWnfScAJaiEOV/BHkQheWRx21e/avs1GzNoqyNxUmmfioIjm51UmfCD84uSjEncuJp
uQuQ0mw1/1VnO/LHWle5iP90cXw/nGkglamZDn1Z7GedlgJ0SqjFrR7Ifu/5XQ8Jdh+KS5Zw6XcQ
7i5t+XNI7ksfuqLQEvTHKVvl0h92SJ1H7V9XnzRR5UoIUog2p9EMBpvU+xicAOCVEmggehb/18n8
LtWP2PZlGkXwZrXBgHupdYguni77U56P+GGKrqmP6CTcSrpE8tpDvfH6Yn31zmxi3ykHs+7OOKCi
lGBTCoNxocwZAE6sDa47I0dih8O9xHQDOW/5IlJX4dXACVu+Z7gcbRf7xNCGEr0IUu+6nCY6ZnYL
sZ6YHVga67YESJie8gQYbuDQCFA6Q0+bqoiXHHbz3fmSWvNfjLbXX44X3fcQyPZaVWLz7aeWpwfe
sBIIt5/t8tSCPc7rFWHxB389rhUH5/A2cxnQAwdBx1nkMfKWruHfWaIcLcPThtbNNfmaoGuJjc9K
/kMWb1k2NiXnBJuta5rhfGtcrmJqexQDW9ppl2qN9Nij2pwFYhiN8tEQNKS6llO9cF6mzLDXOK2e
weIMlS9oQ8tMHdvCLUZVCHBE6g5RiZhwbpj4UbwfhF2kNax9SwutNN3wM2ECF753OzJ2Xdegq4eF
DMotlWwcE+xadY6FE6kQNwOKCZj6tRiJlraAmj0atdHcVWS4NC+aeWhf+H/IWrwnVNuMueJxkg/L
0FZykXrhyVWBASx3TlHfNDtybQsCzo5ccnXqldV9lC6kOZd8ufwKq05Ukf5o13i5j3ypSyvvu/HF
jFYKM0/OBT9epNK/8BXhEnYEJEfYPezEHc1fKQ9mXPJUgKwBi4E9kIOfFta20GrViUGHia8+anvr
aXMLB0uif645k28wLzNAvFknlrsrkZVuTOk2csn6hFQrkz+FAF+fP/QTfhyMBfJJfcMYLoBIlyCy
PCaqJQIRMRANGAxV4BvnOxm7oWBXKTZ2JIKeZV9Y8F+3XbQFwhrr3M/cExgvLc9zRQD7/E1AqYb9
JRYjAUJj+QV07quyI/UliO+N9b88RjmOjfIP3JC7K9Y7mOodrdxveTP10yxS3i1bhvrUeX5YAl8U
LAjPwbNQrs2a9F88JSZ4LVxo5SPx1Lmkk8xTycuKOtjoaN8Dh49lSa9OXWCd6bpus8jFL0Pnsc0x
MIbLxLzw0rEygy9io6m0bU/sJQrc4OnbzeyVagox04o3Bn5bJhxWy67p0rOcTiNmNEcT6hbIhiHc
75axleTtA/u3kqOx/P+SJo4ef6TtrN7BbvvMiNSVbRDpMlhiahRklJWytL/L0KDzl0i5V1utlr9e
FCcdxz1R78YhZEwjPDWY/6WtYNg5rmsb8K8Qm7vrM/dxCGoiulUKVhQuKwerW2o6vxXq5EBxQ1ar
BA1BuaRQahIg2dPKr6PjjhRIKto5Zmhs7RzZICwigZd9+caVBVnYYe1OTmyO0CZLZgJnwvH/CcV3
K5/3qdxqGrsTogq/s1Hb4hxzxDr+OmrgzNZS4TAD2eFSMczLyygYBDJn0+eBOuTXBW2nh/3phFLF
Wqi7e9pMGkFWpyVDc++1ICdsg6xWi5feok5Tms6quaEqMdl3k56tbDbgP6CxPfrk87ih0Y6VVs8V
/NRbYKk+UNgBk5wmgk2o/IoxCY7eaCdrUyZXKD6FozMDyeo3a3+RriTniehUa28HkhPqUsaZiSEG
LTVRz00ZcQHDKEuxhXYTbGWm05msGAUvr4lm/a/GDWuJj3jWBJrxgiO8yJYJ5aYPRci3+LhX99CK
4Cco6/lPzeHrd8ZTGIh9oiXLQR1Cgp0cBLvk43UB0AoMFScSJRUcu82fDTCC+ri9o8uEbQmRCDJO
eAWOUxhZh3ce4goeQQc2vX00FUjveeZAdrhaa+cIZqCIjEpP2ELFqnP2oSbKq0UPv2WDfEs1fzSW
7gpy5rcPISbxh7V8aif2v44s52diKIsCJBOjZNAcSj/ZrRPUBAqa0suRpRejqY5h51gF4npVRvRL
4DXWUfYVMCFXGSplA3WT+E8QpbNFlBOx+CxXZNE+IrYPs2PZGZ/iDMrx31Z5cCXeQ2TOI3knymZm
Lrg7ztpmrs0tp+/nZs+hvBTKqlA7H8LRDS+qCAaxiesIx7a9zZC8bYOAMckWJWFlVzhUf//1zJxf
oRDm6SJbEvU05crjSeW86GqiQAYGIRl4QO+/cMnTRU4olHp06LaMPUhb9QW2Bu1z9nGxfzNXtMOS
FberNDoprEoUg5M77PQrMdlS8b2LC0X3AS0NDi8fVtI0Br3PWACAJbFEX9U/b5yFHZb4LF2t+bx8
REZvV9hHZUnhzyak7JSyIDdtM5CufggTP918uRsKhVc1Md5FjA/+yJrvjj57b9R73UF4WGIwYXXX
T9aZMihLX1YutTKctnan9Ll7P/eg9jFIUxbgj5x6DawI0/NGUKaXoSOMBKmSPUC1OZAbWWhAqE/h
edt7WwEeSMQjOQd9httQFZyGrXugDqVCyYR7HUI8+jDN21WaOMmk/vt+NYNiER4qmVljEfrBuCcY
pMgdokrJ9ob2fUU6C7wgH4c8QEiA4OpBKoj0ssKnGvwgJY3QuVZyFUDGi0DQj5L1DdoQ28ecKnP+
ZfSpTInw3058FNUA3XvOInuEEKeSau1/hrTgx9XvAhE6fp7Jc338k2dd4Qr2Hdcm867uCGlPAw4D
mV6G35HwO2vs/xgPLk40HCycOOPFkZseQIt7gqM8GPM5UQYGu/+e3rF2CZ5UpuovyK5tO625Ublm
MMQYtZTZlbU9mbiKLN697Nq9h3ugWmQSz2rhsUxoI2Avvs37NQCoiHf+jSwBCSVoetAzHfnOxR0U
aaMJwo6bj/65zmLV2KEMaNoRmwJaqvd76Q2dBSxdDkrIRMQR1I8rWmaqK2FfDXTfv+3MiPBM5tI/
Q7numFEMG7lfjJjKlFFE4FvkRfsu82mFmZIaUBWDcaurLYJrlM5yjDnRSZTR8VhNKmjyz5BHvt83
DGFDbLpCk5AJaJCkS5bJk/MAQKFgxsc1Ov9OioYtpRDV6ty/wLoqjcMTrntVfqaRuhpZUScPNoJL
whgamPHzA2j0AD02tmMcw2v41pihk2rLDqQkgRDDQWJ1iPp0Ortjsw4CFqyDuE3NFdeoZrw5nD8t
gNmZhcg+4cH7KrEJdyrRfV1Eury27rDQRd4Se/AV55WJm22ZzUJns7IFArFhRmQVHaPQeHbS5vMX
sHkCAJGzOcOxwpzsZqI2/jq9dPuQjSrqi/yBvU7ybCjnBQUOezmzZMLgTyHjfzgni8BsKXhXnuQ3
hZ9inEmXp9+i8CIJsbLaMTRJJYCSKkgB4HuLxrmGVffn25pIEesBP1plqq3IiJ7lx281taAhWO+R
yc5DJYctlxaLE9M6dxWKKgPcjCgPTzory6k+i/Y4B312sZjWoCUO1wP7nrWckJbl4hCP73EQ4Axf
oKIruHBDzfgy4f89X7Bbrb3S3OMDlUckPJvxSPVFjaRXcUGTqDlW1JtykpvCC54IK6E3WTj/JEz7
yvZ0I10VDYyrz2WnO2qstZRBA8NV8vw+uUxZoRpESpCJk7Jq9WfrFRZExJWUBNfiLcSYdljEoI0M
mytSq+TsszkmriAUdlLEe/yHo1FA0YiPsS3xjusP0pwmVIVRteZsM8d4Ljlpwd8tIvIFC1/x2KBO
LazFtbMlrvTL1SuRtalJeXGh+DvoTxueiQzK7bxdR+H2rRGyy0jGjek07lhU8dwxoLxvP80q2TZJ
07L8XntD6peKzcbAuunm5pxmJ9+RwQakgwD3JNgEltUPZ/7ldjR5W5S61l7MnQWlvB3Mc+JeQE+u
f/DHGAQ7xXJJQ6OyV5bVX4D2Rxy5fOT/cMZO+VU1tDTaktCD7ngPfKEJkR9TBKdShbuecr/736qN
U/ZGTK3ibfN3Dfx/FW1mAnLWeriTda9jW3TqIZa9in6PHgLLFVWjKqbuD/4Bdn7bH8nX+JO92EeV
9U1F/e8N2HHforOLC22ulEWqvden2gbmDIxjLWzcvJOc318i8O/ZjvTdUXqVdv5MtdHOmyC5dYaz
oe0BlI/Zb3h0BHqbqxuRI7OB61dfCpG1DJcTDjx9OWsOr3NvN1G9lFNK3fwGUrVX+T2peAPI9b1G
+RIauj81zIv6uQ8fYaY/HcaQsUMXVphA2ypSnrRpgtfpudoiLijNq+ZuAgAlwsyqmfy529lq+uww
6g/tJirW/NnEOrf/I5ZKCI2M9sn4mfwzTFnZGUe0hkilzBmO1rAxvGRcjMwyLT4853/6bA3ad+5h
FfGoQEdJo/ytSdCcGfUQfbMU10inOouia/LxUpOLY2ZzQ1ncqKp6cl9y7/45dCr3hP9tXryx5sIu
DlgazfYjX+pZM3KtX5Y4ZTYzDKt/wfGFCAtEJ59XRzp43kdG9dHTbXXEJn3uVicdK7CQGszgA4GN
LYhIgZZMiSfqLSdRZJLQ1Lgoy4qL75hRIEHex2rdxX5ljorQ+ue3fc9yrYUraESxMZ3qulNr2hRk
gmFoENLvGTbsIejrGLJpQ0rhZ7oUWOoDlilLlapGoGAv4BHcFPDaxjQNMWqu7yM5b6ykSwFLp9Wv
cDd+46JsvaJUlqPsYNIL1mm3sKm6uzdx5nmVr1slu4fG8wV1rK8DxQq1LbDVhXwk5N47TjhDHdlL
nsdJcFdlDturopzFWt2HEpdVIXuwg2BTwnK9aPrQc8HM29XyF+YZt9CQuBwIjrtg+dU+pho+POnt
oH+7obrjae9e0GKcawn8VpP25KuearIGLy/uoOYSMgeIAodNzOoz2PQtAVA/ULmsTX/fZ+Ra+H4N
2Ma2769ZGacoDJJ8xYiq9+Q5S6bghwO1mK+oPagMxVf89R+LieMHZDxpF5RkSWqA45wE0IGJunlh
9HqLJ+z/2do4Nys6O/AyaqlGg9Igpf3eobaJVx5z5OtAgyVEy22igcouP7h1rN8RPc4QFrt1uQ4A
WycZshu25Sm1cGu+iT0XREuoppIFyLb/eFABHWbfaq9CvN3HNmBs8V7xCIiRLgD+r6AYgDT+gF5Q
W/sKYgLx+Ggml2I0d55iAs3BVzDdg/k63Cc9Hyd8oj9B+2xaAAAdTCJMj99oMfcK0WSRcRm79PXU
TvoFqF3EF+6spQfLJN2bD5o6Gh1lDct8k0r2ljypm9PyUqK7yZrxjBsXt+iLEeoJTLA2ON0CarIt
WN6Bxnc/XT4JTg4gAD/idOi235oeG/3ZAHPCn4QS8dPZWGXn4Pbk4QurwQLQpo/5B3GV1eti7B81
Wc9ujtqA96KvHWEKg6rBoN32d0xHZIAoEGMU7GhAwWaU56HV9rodnKBHOR0Zgz/jEhME44GJ+Yxn
ZFtRbceYqR/PTfNtRNJedcTI7sLbdeaGTJbT1305oCJHVXf5BkPe6lylQtD0QrF9qSK3jKI7MSik
DVRNuAp6Wcmh/Ocgi5Ku+c33fATdS3dtKK9KrvrOKmaBByFcTtGB/7yB/nRi0R1qHhsDXBtler5x
6Zhxckga7iuaqnCREcGH0jQIkaeaUPyjPezAx3mknGREvakM+R1sZY9uZzcfumMuCWymJM1islcF
I0FMxFZvyKIN9WSyzHYVL2QCO8sDs2OYpLrdSp76bJGAhRrDoAO5Dzkz1uaGqUIiwL5XPzi6lMJQ
pP/69l5EE8kgayMw/e5/134DGlBawOxpnjdMBwchc3oNP7TqzeSa3WK7a7gTLZNOMg3jr0WWxFCH
pSLgj5H+qIclHy8q69lK32lj+nB6otKdnLBZOlcj48eO79AxeSY0e/rUPRULmwnYVzZFjO3FcNLi
qpsWNNvL9Fa+QuS8yw+dhf7+sPbIp29QeuGdgDdGIXs6J4yZp9cc6zRcLtlYWRQlZmonLrzx3lcI
bw8SRBBqWmo4k64ZjA/0jY4I1cc3T3ICU2BsDcU6bkbLsZq9ETZh1t3Jwu5Lop0r/q8YgOOFKHPM
oZ+Dkej+UA4uG8rDsN3N09Wkrqr7TA/co5rIW7DQMBYPAsPGnAQcjJL4AFu75x/8pFAYsFmyKX3W
KiZ9HKJYhl5FrYKZ1SIcGNKm1YkQjzs7BgEcZKo+fj6lbHC8gloVRO8ypQ2krSITKYVIS/BCuZOi
txkraQJgiUZpMJ2oWPcSA0QgPlRZO8PvVmt3NAPOkHWPGCgJdqzzugdEYjiNuh2UyC4F9ZqbU9jF
jB6oLtjh53qT4yyJENOi0gy3TTl+x/eeHTDFjE+Cg//qjZFU9kuDjYtpoyNcSnEuKL2G38xsWpJQ
2Wwu6fbjBbmDX4gKXjhxIyMqffPzsIe/xnHZ2adno/AH2zhHu+g4nNMlL/4/FZOSe0cHCtEwKzxu
HKprhuZNB6cc6pHIqm/fMmRG4ifACXdF2AOiAH3GdPWIA+k+yAZFfBjcCrNbxBrcCI9ZIAMeLoUc
R+X4xpCY6r/njdWhmNFByNVutrjNhr7uREYjDHziK9/ig6CB86djwJVVl0vspPqZ8uXHzqDv7Cim
6TQeRDCksLJnIfnN45sQPBEDwWQ3bLvZ7TD2iDsRPKzJrCEbo34zXP5VSGC6PHCPhr/zcvjRQYgu
2CMvdkllrFfLK5gtHu3/jaJq2DDzEqV+T+qCwvCyrwbR9my8W6gukOHwErfxlPKd3uqbL0SYf02X
hr4GD+9AGSpnyLzbPE41Lv/Cy3jPNbz/jiFrQApmPAYblWgzj0vITdvnD3xUQGW4UBilTMeuJibc
8GGN0SCfS904EOzLdPRlG1TOlqffaKmhZeCSPJodM6WDLJs5qczJ1rN1YYdpj9/kmAfWV3Hd8x9n
U5CtTCG8G+fZQ6MTy2EzCc9ZYqR98FZ0WInDIf72wUhBtVlB8BRFGFpcr14McMbYd4P/FjH+zpuV
OmmdybfJQ4yZjBiDkHyJwYTUTNVnIqX3wQsqDBbPm/iLlflMnNiXNt0BESGJ6GGGH2AGIU/8++J+
R9lFNhHt56eKMmc4UhgQzOZPWMYZjTYZv3N5xrNZbn58U2MXNk2n71iMtd6ee2lWSJlVJMmJps98
PHlgjvHDM6Z45HV6i4yn414eRW+acNdu8pIAGStPRatipbjFKVaojzTYFM2odCsCTF/+OxUnvlRu
MQilPEcUdjM2mnsI9a7S90fEDMByTSg/8EzG6Zj75x/lFT/NkLpyFVdJZfVII0rrnxdVKOetXB0n
E5Aa9tJoLVuacziLVqhjr/BO6QmBQ0LpnP0sYHHr7Vk1m964+ySNXXyInBFN41kIVVAoIWdugixe
5u5n7O7wEA1nyP3U1oNcAZAQMve8K71XAzetXv/HSIqbLULtLEuNlX6wyftkrRrjKL5Bebjxfkiz
/UwoNh3mUPBffeda48WzQHUZatpeWrSy69Z9YcKfGB+PZWAw6feMDYazwTxeuOEF/E0q9ft94iW8
pXa1ViHV8wniXixh0GHAXPPBdGNwK5OXlDGV3d/lmdl1RdoIe/6a3tPnN9mvEyPF0XPWrq/4uf5D
AXtEyNlLQti59jKQyu86w69cz3fYF6xrGnWS44pxvhK9ySnvQ3M8/0mYiGdDR5pR/EQCctnQrkvG
HWBWksDJnYZHfE9yHtOo4dXt3N5il2Q/QjBS5kNZRWn5PqXBy9Ch+me5pmw1za8Kw1pPLkIzszEA
zMXNigpewWmBO/8Kso4HTWbv9nOym55bu4xrYIsC9uJrzjuQAkrl43cnUWkOpaShU7Q+CHvD0WaQ
06DbFCmJP1Yh8VDTNIJOAcTfyRnReVPTPJjVGft0z60ZNrl3m9coboICm6FrnWY647J9BTfvLzsJ
k6eTOFGaqrhXChoUIDi71e9Ydjo8L2H+hZnmpQIlqzH/7/bkqElUpUBxFVexouUGbJ6NRm4pBg1C
udgBZg6YQ5uecSDu+cOHuNhKFdTjx+FL6uqroaKdNy4gGY6ueuDVCweDDRAa/+ZdOZFTejBP4Q4T
SmBrMmqVbQHKKbcZT5S7mrO2+BWHCnj86RNOYTovCld1PC2Dcb5JfuIDB07NX4iQjBpCL04NZvoS
fI5nk04Vq/uGW3VMPYkLe48f1d5qm1guo7HCajamUPHPyJ1KqgMibwXTUWKjYFlNcFior3NLp2EQ
5GMTLDxrTlQx4ES8bqObxpu2cLWL4onVn91hvetv+VUwtciDUMhrOtyEV0DKowNtdD25jqkgsRkb
2AHGSY+Fyxz/8qcLtqo3TRNodmbhtyMWqT2GHd5I0cqYGclnJbfMyZfjSlsxkEM23O/7miLIeyet
OwJkNaOAtg2k0m/IK+Rb7Z2GUrJaa5BVM3e02hIpHsiqfl6p1ZcEtCMEp4iaFxRZWs3pIR+lbtor
pt+SYsItVX9LEL/Kso8BDvjU2ivuXy/wixuqlvhha89sxCtu2PAmHkY25/Fzk61hcqLWQEd+Qosu
Jrx8yzwSq0VzikvlpnVllTviVwJkqesz+tM1ek5GKeXJHC0eVt7A5C1ef5LRg7szzaAIBQ8Rjt3X
wTnTAl4X7I4gBngoUiI6JnCOsQOCk7NVw8PXGQlBqEms63j9A3jRbtlBaEq3CB9BYfhE8ARgKdqf
+mMsQb8MeYwYCRxW6sLIDEAMUtviuxqnHLMpT4hj5kkHjE+aalOnBw+IIMqQYGtlYDXW+PMslfJw
xHUZMII1DGzBpl3H08+OO9UMjqPNOfvjtRnnTtdIhsPgp/td6hcmam4wqZ8r3KppVxGRyHvkYuIa
QSvsvOcVu6+i/4dTDOt12Ynt53HmcExU/tEYFmKoilxHFh1U5obnlYF8psI+V/bXdxkqWa1P8WCB
Z5d71vTxu4v2AmTptae55UhyBb36Fy8jEe+aiUT6QzhrLEC2KimRhpyj7IUSge36KkqkzvPbEbQW
zlyqRx0qvgKdRq1izZu49nxD8qCFx0kRaPehXhuI0lFaAQTPWv3pmDMWSBQtW4bYZxEH5diPNHzL
fIYDrdsvcshTAL7QvPmePlWxqPm73V39FMNBncFrgl6bspFqBR33dPnEPuccNfqwtQicaNyUNW3n
u/FROchBCyqDA6fJADqvgr/kGjeNJjGKRFFTnj1FbosKvsC74vmOersSag21o+ZcjP0Fcuhzla9U
hfLMeSkt21Hx2pPaKzcoxZamc/mlWXmQ+I1yYfV7n8VI5aBobmHieKcoNuWP+65PK8ImUVqGfk/1
qYkmJUPF8HPPAulvunhXhT7SSEQT+pviXhwhV1bhMfxF86b7k3kkwHDJi8n1WA5d0gG3N2pZgBBc
KOkW49SJCkmsQYYdGcFWmVADjjinwRIxHEBAkYfcqGrtLkSbogUSqixLuckxLs2MA/B3JE8C899K
93zrOGW62Fgc/KXPCz7ru0v3OFWWW7+vcQky6hpFz1p+LBhAYdCVmeJIEtjSoMMkyt2/+jGHzTu6
ByMfs2icE4AK0LdbZyVv5x9V0ADjGHJFhXgnPbbQ+BrTtpLY04AFdUiB/ZSr+S/m8Y54VLeiGWxZ
SH6ZFM811hSWe6liPE/xUMIQQ+PYBJQvvcTX9mFp9py+oqIxILhBBUBbCyWDzza7WD+Hi9Ck3ay0
xDVHjBvfec2WUlGKMkj6LXY2GFhGaQuWfxUJEujbbq9a7IFTN4ACpDUfmkfcEiYYEwJ7ifWc8SBQ
hNfMF89B2XwgYAtXT3QnzCM6Jh/Oj2g9cq72QA6Cxq/d17bY6clnCZqPzbRvsDgvZhSL+Bu0MpEQ
CdZn/O4v8ne/1MeOlHB+IreXoxu9tSgwMfZZ4b8yE67/PZSxmTfkGzT0npmE8Q+AC/PPCF8taFJt
wpP4uQBH2PqhQ+kHFBVC3eNkmEybCUOXEFKLd8G5WUl16f+SiUbsHsfaIY/WpTTNu5RwM/t4A+8Y
hyKyiOLw4OPb1YX4Cz60d4931uLkNhFcn3ZnAppil7LGgmwUS3drQBGC1AgAVyOt91rrDnxBabld
MuD2btDwU5Mnh0pkxOj2j165F7Hve0a1Q8w4IxNDGYZYzAEZhN+mJOwmcqfNOWxmU+MOsjQt5zOt
iCJY75SLJi2BB7VSm1jOKW8Yv5cXGtrLUd7xWNvJP/5+aCB/swuWfWdAfzV7qvAVIDrjEv0jpSXn
v0a20Rpw3mF8zFGAkEdtBqa2O/GatWzOmaUidwwsg07aRkF4YDr/jhBdCoe+UBaXaNNXkWA0J0at
E9KS6kFLsnEEU9Fu5VKvbKt0mcHsFymW5QOD+H6BVRbSHYjPTLzoh1Vhs0V2LVLcpvYFFf8CB551
eHWMKnKdRB7RrsKCd8+vXr4czQQt+MuedTbEnD1YnzYqgtTa+Q48S729zbkLSfpdUh6hnywaCg43
tmvM2wbaJoo1HZmEu8G/EFUwghqG02CjybGN5yPyINGQj+eDIsMhgA0sjigMtztxo8QxEDUCc/7d
z/jcep/jkI0rE/pWIbX1UZO9ptwzVaUVRUoFbPJ74PZc/ZA2T2Oo7ZvL5lYK6LwCsg3GOyKujBrR
Ra+TchuPueat/ZrMPAqbAoM2yd9Vp8LEG1agLVN2BNh3LxPD7KXU7jPlgewXmkxhpUiq14A6cev7
Yv/Nr/Fy8brA5DWb5UzhGpSqYaKZ1hMT5qnpJ8YrK1a3DT1Bv3fqSJoKJFlnrZAySEvRiEAmAOmL
LqU0ytl4VTcwx1jrubXFKtOXXYWT4dUhyAn4AG+puYiDx2/DlTvfAQdy/PHXoJPAuDjLQRAUNTcy
jkGA8NrvmhW8m2TR3n/tEmymRgeGggnkSzOFh7NljOVk7hP2ftYRqK9RQoBZcmMu0JL5VZ9LyOwd
qdpns7T0Ak/AoDtcK9U6zFT5m3xjF/tXuMUZESKf7pewOPMecwaEihcaaOV26tGG1Gw4D2rEMBm/
45AINmt1E6AybN13vsUrRNbyz+WrpKkGdg15nKcfjs2IweOibFwdPFMGg/yyMr9vaz54XtSBe1JS
7wzUfpJs87NEcerYZJLsWSgQXbSlKtOr9DX5k7BASJSoOc66Un7N3CYW5igWEMHqGMGLin2AstWq
pERDWWi0JXxhanNsQJUcBAsucpRUfv9A3nqPBa3CY+894Y5di6pZBWkO+1W9BirHAQ+r8aDSChMx
TKE8QH41zTaGHHFam+/ZvCogZwKVi10qOS1DdIdBYr0F8JKc9+DvMS3emjLA6rqnfziZaBnKTu2E
/SUtn9yjXqoKckn45+SyWC0932Bjj9m2Q7sc48GZ2iNGwwLbl8P2KjELRPDn1Ao2agLVRwl+6GoK
EuzaVUY8TlBYa75THzwnQD4oRFuIcjwzLde6clbAVr0UrQM6fBMTOWXs912NKY9dhsvcS5Kr7PZT
wFqYlrLUzPP6A69ucniuqGLCyPWEPLUQmkPiwXl1LXWPfKrtweOmzCpepEWy3EGwYZr/ftJAIw+G
U/X8OYsy/VuRtteHJegfP5/PQb9l3iHLEvklTPxNNl4FFPEs9kRJIAdQ0x1ELIR2XFscJ++kZVww
c6wPxlQM7Y4Ohb5ezR/it1l7rxnG4Vw8wjBZpGMR4UDsZ2/2Whz0snKOFfK1OQwuKT6UQgxH++nf
Qf8sTiIJeILQeqkJgZKfrT50iJfFGuf5TBh8iLpdhWF+cbOJr8NQkyEfDNdVb/UtUt2CYRDNHiLj
l5lOx18I2tRBdvkmvrbMqrRugv+S8e7XeLoIJ1UnGf62a7sL6VSCQZKIR0bYMBzxsfiCsYqjrwGI
FGl+Q9blnHXqIQIBXfsU+zUZPmsqW5+HjLPlBDkrOFE8M9OkNaNAQroM3Ggp0JJE+hMu9raH2RDx
nxTTn5YYaXfkM1fZC+6MM3g92iufBurf005uRSMFoKZuLLjc2gZciLaZa6yUCxpOGJ5lgwMj3xfi
av8x29vr3Q5Ixah5gmJwrUJo1VMmUj97An/RIrlPoOJ3gs/uQONJs4dXYHXEEAkbRF6QygCt+a7u
tAUX5nXV+zsWQ9vJoL4NA4AJrBMGsf0mjlJme9v0Lf5WyJg2eb4OEejHQkq34LuYRWaOrhrLFVoK
aHNKLC3/exNXMtMqpuKGlaBPFI2U9Eru3g2QnnukiDpaLNN6L5jZde7xH+n6KreznsWFaVGsr7dT
Zh/KSUkshp0cL1c37+eZUKAWOieUysi0SACQWT7U1wZrfF2yuVnk1WGBFenSWOjhPTfYmrYCW9oa
INywanaBXTcLn+CZdVn8uq7oelPiFikb9VDZ9rngaz3J4SlhWqp0EeTCkWyF1waNJf2bD7E5Z27M
a5IYzDVwLkzNWhEfPkLvk672fKDA5wlKh+k8i/f+7fVtZ0E6Ze6fsx8zImk/bshnQpE2sp2tAuvi
5RRzfIpHUqcSxh7Ar+kzyg3YTCHB4bH9cylH1HVwhQoigpLxX35k/2h6uuNABAQ5c3r4kpbKIpL3
1rAh5JgwGcDBk4CuCs4KyMFxnHTPh2lware4hB+4yM7cQLwAblWXDTZls4eL+psWdEybpFbGxr6W
qtA9ovwd6Qz9usCoFzD94aBf0LAncFxhJb43aTHQ1qKjar+JbhpJnTGJqP9i1Iru5GohLEE2tnVi
zCoqbpUnWEKWQs9YsHDiO4AGUbeFDs3/FBQh/5imk6PAOzg3otahEERULgLQMvj6pWvfNGRuSJ6D
DzTVMMR0lTfVHU5I89DyPGOGbqpVJHsm3ErdGwPNKXMbZ6J3zGdnYwj5wEqEzrRCrj1ApKnUHMgE
S+RGAbXcNgblqRQMAAKLXf669VqpMmbVpi45cwukDZ18r8BbJnhqqgk17L3HEObD1IkNFJs4PqtZ
y3fY+irgS+Ov7AFSEcuIXyb73lMFrzne79istu/YV6u2ZTLSS5MiwRdMPDcyYJ3j9Y+TvTnqsIxU
2kfdx2W/HGIDHHNcuMHGwmdV4gXefIikynW7fID85OEKVXmcYI22MdYx96336mWTQrS5jI/wnk3v
3VQ0ROWdF79EvatxKBPlqB1JVdo6zmqsWSo3MIftVVsixMryVSuY4fyEVe/1yy380Buz1OApprES
91/4bc7Jvf6Wo4XXaHb1XMe6Ms9jHdFvh7pfiiKkR5TT84Pg2MYVrhowk+93vQvYAOnfTZ8WRYVW
XdNW5Uiw6yUEHeXVrZ3M9n+YHUIJmL9k0e0J0mRcHoYanhQun/8QqOJTW9PEl7Q+lcUr1v7pPQfk
vKW6teeK1KyFBsRdduEfOg/WrOY9aT5mAhcCHXv4oLiTa7z0hOnB116pEoR+0oTOe54kROuR+FU8
dy47sqrfc9dhj17biZTAE1n4Rc8fZV6JmldBsEncsLcOwGfz5gcaXI7GQEGPkb9Z2FXwZ7/DZ3Z/
mPEwrGM7FdVnMoGhpD5awWDp5ysJwgZ3aky1G+8EyEkDog8LuW3aFHOQtlfZSKxubLqZAlIlSFtA
S52jSn3SbiM80J7dqVtYQ4zQlOyxaJyaNRFAXwAEa6w54NccE18T7rj5QSgcuLDSdVMYgYTZGjFp
V9xVucKPUUNsnzeh4tQaG3iyAlczEinzPU/d+wnzCDgnH2a9dnMGn6+ZJN26rr+6py+aAAIaZLlX
N1/JypLr46ryoHMlji3rnnWw5BGUYgBiiCrFtLH3uNWaMJlYoAWETEaI9C9N92xEIULALMPw33Gg
I41rLhqJcwVzdLf0d9mn06vCWw8VjqULOGlOXfYBeaA/vY2VuBu+C+dw5AEWgMS9jGrQAIgUCz7s
aYkO4JuKtxAj3tcgZxvq1+1uDaC+fFlszP3q4xioymnF2jz5xAoTQg18k05U1xg0LFpiUGv5oUHZ
LPBgCP9mLyPUW7QjCVV4wbGo65wddtsJr0cLo1rRyNJyH8F7+Y2VacIhEBtnpnFzWQ7sAMdEQ0sV
vkSYeh6jrbgkI4Wlj0NSxi2XMZDOlmIqEU+4tYaOfX1J40sKxqp3MQ59DyhswYW9C3hlla9T6n7M
YvCnTnCHC+tYTsB4zpRpe6k+ad8SHRfy9S22qv1qUKGHsWOhOYDOH8j7rLb3t7w3W6eSoGbHGzut
r1j+IQ8bA3oUpMl3ZMPyUeCFYzI0mu2F0E8sUyai8/MyQBZic52br6lBgTEr+m/5RrelrpM8RqdT
8PJ6UCJeGtpUJFkQKLywz+JNlHjZWnlHxGqLzM8wiie45200nySMnXKt5otUDQSe8MPNWQ0rl6Dj
w+UDPeJVSDEVhEDgpEDYd6HU2nn6f8HwvTKZdsASJ8+eFvhoi1YTfcY0ACjzVfpDuXRrddgpAVuV
n6liyc4EiKzXuh6OTd76FfQnU9Lea0yyeWY5d5TADUPcSSy90XkAT6z8SLW7X4sl6GFc6TRHnFfW
DUlcLGfwriw5u3hzURo/DvqNBoKsrS0FtVP/3tV8cKos420dfjrRNJOlRU8HIJN90ETiFp5HxFSP
1gRR+tjSYk+mXvcFey2QOUpq5ptbG5aFqhLu9REJSuJ+QOIojS9UIpHdsERX8FXEKZjPLCKygTGO
RFTnkSX5ynbMimCqkiz+cMn49BRR6XdQiOT5aGn/ndecvnJOq/j0k9evAQISUS6KP70U+CcOdAhB
1aChM1fLyOeKSH8Pc542lilWW1hsoi0juLo/yM0iMSDr11qI8KqSGhuPaK32HGvzSWtouuAZ6NWv
TZRT6iPd5oIV5+OASzABDQUbwGIiWvMchJvM89yTATj3MIQ1keKXQ/wTUBdp3WUcvH8t5J4len+/
7isap5Gjr4Sp8iVEhpWgYLoy7+mr33eUx+iil2zCT5PPgzWLOZiX+9BWw8W7tsOia1ZVZBhxuLXs
GVPnhEmsdOMr2eCxrG+Z72EAhmwdnIL/KoujuG4cmnkOB+/b6BuFRCoc4fc1XgM4Ly8n/JtDDGKl
GG26CycWUVW+WOy9rfB9p1WfZ7cC/SRlo6l/PWYa9f9yo7AYWU8XQOMUIzH+4GaTQxVMs0AEkT2s
zJ90TlQfREqqQr9cgcGmBpWvCVF3w2LWxVUACZjO3GrU4Sq4rU4XYxQqjpd9lfe1qL1Ie478wzf7
4kB2OaSqaml3xvFcgRNqdNGTobwQgMpOmYgj8H45dwiA5TeA45u/HbqbmyGSAcBliHCdooasScge
rLxPusWFmQXDzTv1x61qmUwA1PM3QBJf2v98uN+5yQGgnqUSrJ5Cmtm1Ssx16fMekTLo12YMgwq5
E5miGf1hTE5rkdtM8aOeKajGCS9yGnUTVJ+GsAy/Ru3ZNWP/BVilDOv/b26pu1lLbK8E6XNlzph7
Rn9WAQViWwiWNHYX1R3B6ieMU7wnr3dHgl3dzdDG1nBY3UgSbfE+HZyfSo3Rx2MGnauyyJX+yjkE
Ft+5vOlxnGQc6Iup3aXO7/DVg00AMhpwLVFi/MNpT8A4JrHIGNlD2xbeXgHn3huGK1dQwt6UhAt6
VX2GFKnbG8GusuZnzb5bkz9SIwNrg5NNVBwxJlSwH/XudTFF8SekuQ8R0vwo67UCbMmY5vBJleuK
wE5WdiPtiN9PgtKGC4kV+XHcIj+CTX8YV8gS2XIXx+KMxhFSril325BPr1h+bUT79638cVym7nYw
rE1EeqbIVkeO2DqX98WvsJL4T7AAWR2dJbMokCwn/iuzV3RhFMeDHhx6ufYs5/K+cEceUpZcG02o
HDliD2kSgOiObzJrv9N1NCK86TaKoH/LCwHBiGCByucjaOsiwKzc7AozY3otBZBR6TDpG3ZI6l71
Q1plu1+toWH/jrnUVm0u3D2kH/YtS9rpYDMnSrxIehfVENaH1jfKC8vSxqMCFCj9sS6F/Cd0+xfK
b4PYizqD/jKQnlVJace/riHVLNQ4Y3odqSuSSRyiQ3ShNXzgCSBsgqVj8smnweBJ6cFzL13qd0Vm
vGVY3gga5BlH/ndm09PF2DUTYPOGCj590UPPlMoewAoGIxjapozRjgoKRIMUpRNkNkYJZSum8c8D
FFG/rEyTsre9NdMgbjPzWteF/yCL3I82uSgwgGOB8SjSazWx/ukwJIVoO/c+9to5FBbgDOuwDmKr
XlQwVBUq9eUPOlBsWbXznS41GY5e4zOiapwUGKFcSBpiDNjhn6fEjeOg+2lXfTeCB6ovG8+CtlOj
CygtyZSxnKCzbVekkAfWVJoGhXyeLQQmgjM55p7SU79+kWXSNq3utjYR1zXJbeknxpaUDbzEXIXW
tzqjNz5GCAUPvY5ZyBr5EA+k4bJ1CPC7GaXMrlZzI0z/C3THi8vBHLT26hsPKU4vz8ZYM6HtzuUP
VKTzPvs8FpdVVu0/LxSQ4yTfvbfLqlfH81eDQd0iedrFTQRGrxr9qb+mfOHmaI3GRHgVRh1SY07B
gErh+1pRmGyYeY+LO2DqIfXS+iiYcg/hOyWY1DGqqCtmi7yeyCJQo1nIoN+Wa8v7V46GwExttWNI
LoKYivAuZCkOUS/d80iYiPrFWf2Q/y3ZS+MSZC8FbJHTQebaiR30y4ql4cFPZVDP5a7z5X+RoVyr
4nQhJHAgVzg8/6kckIlD1xuZNwhxmfYojDwR1wKH6pad2oDMhsxz9g2N+Fcjw/VYPTznbOR/2ghE
BaR2fe1nh01xhVi2UlGuIwiYVYEPa9OxxVmNEoxb9yO8542laYpia2GX+hC21cFByKvtRJDzLFnb
AcCZgVhXu0PHMh2Y+fE4xDk8GK/bXGyn7OtkG+CieGIyseoCHY/KWFuLKKjAewx4/Nb6N6WuAYXw
05fZG+eYHbAC/iTn/S5qzTtO10A3Zw6B9J7sT8gOkghlcl+jwWZh0EIpQigubN9B4tyMHMPnhQF2
qjGWF6f9MUumxW0mNVTbPhZlYl2yD0FY5T2hNEL0NVf0A1x5IvjFyDBZcKSQRp1z1JaqgA6Rsu+U
ikT2pL8+xf3bFC6nWVeVG8qNNP+6c5iLE8oJ9wN0B/TO6uj4zJGZVzg0a+iQ5BABTw2M4Wkik6Hz
6DlO8ooQSef1jQzlfoGFRpRlcHIrKCpuIrcQdoJd1FZIbhkOXpIkN1+y/IjWd7Kb6O63pSeySYNd
IniBxTNxS/mDlpcd+x4LDybVbv6oKix/AffVN1O9wTcGEW6etY/gSw93Evi4BQd+PiEXQvsuRRtJ
A6n9EZ6dR/E46G02FheDBNV5N3isnC0YNEJFhXHXZpCE+p8svXiKg4tNSHKbtrXQ2A2WNsh7Uun3
gifnaT7peAwSUck6u02R4DkWyKXctKcPDsD1VElCdBKa4M8XQ75KbDspcUzTvtRglz8PBshhcOW4
Z7nkIR8YXeAiLGOccXQpfJtijdDtqgGGG4wjJfVSq+CUlY/wcJJKzeN/PDBm8cXizyfPZpYr/BQd
mzfZ4uSHBn7skELdkywmavlvv9KJkNR6bWXnOApC1RGP0XeXXjkfa7xAgiaHc37Ttu85SYbf+pg2
3CaTQWHbncdGozQshtzbzkJCvxWSUXzWBLjOHxkmDNaQCumJ1eYt2lTyBJqrIBd7OvkI0hz2zMSl
q8kNNb3650cxqNvVZfITANjea/wAAS/z3Dflmnzj1yhMM4tP9n2A237OTdg9Uhp9a9rBOgt0fjCb
PvjZ8L/lJ1zQr5Yz11XFrJETXpNS1joX3PXqyQZY3DdH5R6XK68SLth2k5etyoX7nk4yB8h8LWQm
E4ZW0XAX92r23JrfFtfv1LDB8tTvV7oDJBikHXtfqrcizuxNAYRoLV6+ULtFYwSCz1cuwGW46+RP
+mMACHCFYDS7zLSkD4CEv+vZ1717uq2tvWDLE4b7VW/WuRN5e7cNeXzaveKfANEIrLXwHzTgkCUR
UK71SPzeVWjTMaXnrrzLErNSbuWiE17olivxytFwTSpQVJNYYc5UbCDmxcFT4DmLh10njI+y+wNw
VVcvGBDQLlkn5Wo7ZC3yL2ABpBzilhWn3+s7AvWZoDMGJjT4OmHGiGSAyrVNVzvxttRJ7kOnnK1g
cRXAQB/7BRiI8qGfcUiv1sxujtO6xX4Jd0t3a4Xg/U/4TFISoq2h1nFWBvRH+q4iRunBOapRtqd7
+0PBceLuDrAcvpqXIs4cEQJf8taJ4ZdNArMTbjQ/wbii8KCSEFhqsToSB9+c4/3RDD3S7PMPYWaV
D5tCzp6KQY+38aztml/HSXjPFuA/XEV71xH6ZWZheRdPMmxPrIELBju5W3ahg0E/WgVYFvpq3FNk
UHPzkQlydcWIn2mWzwzHWnQ89hE7T1nd+A1Li/12pBreafiYZR5mle45Mnwpy/D0aZAo5ixIDX9f
83AFtTZbYHdWL61AkV8BV6YyijYtEV0H44OU3Qm9IVFQ1s/SnlGgtkuiuxiVaujTW7Ffp660Fp/w
Z0xJRPFZNvZ5s1SWqKoRrj5/DqxIO9xyi0mt14cN5WsSXgkYz2Cd1/+jsAnxe4xY4QbFMSw6RVl/
cyRDk1JPOK07O585dmPeRKOCqFZAQ6okENXxh2J8MU1f02w1FCG2dUkMu6j5u/QxLNrMl1qUxQ46
E7nQFtEirk2odUylj4zs0P15MJCIBFTDkLfJFREuLrVemw0QKX0gEErv7EtiOwxZOVKp5BXbfDpk
THIJRlYeWFTJylh7Ws2EtE32uhGy4qhqZmyp1HM1L2NDOB737/v5QfusEHSZrwY9HWlhLJCdBk+C
4BPmpdWMI+UpQmSpBB43JQmOCk1wntPeDzx1PVhH1k/6Zj0V/PLqn88JkP5/JWCaNVS0IXqW7b+R
ViLPZJ1FxvvThCj8sMa2ISnvqyxF2Nw2inKwACaMTQbwexUgV703GDxqababCuxXRE4+Z1QFb7UE
Z37kj9QWMLg/owzxRIoRNwwwn9S4CQbH6oNjtVhDsqZ7+nZDRQfL3vihZtHCJI+tSYlZOswPEom/
N3fykm9KwxsOttnHcOdumrXow1l8/rSO14zcDRVx/VCQIn58B7cRTBjjYYc2Vqy67tnQqiopVL7d
WKM7hFKzD3LhPtdLJlV5jzTYbX8GUTlGIOc9giHIU5OfuxkV4USnLTQiU0NmDiIN5ZzYaTGZ6x8I
RndVbIRJ+uwfCBEiZSr+PkaZG9wvATygG3x5cOmkQV2cDZsXtu+OdbfWkTgbNlUSajVI4d1TTGMh
Wmx4GFM4mCAq+rmMre8TN7q6yTV14lmcCvBYvOsCUYzOET/ZQyUSY9bPPwLdaGmGMuuCBfAwtzYC
7xsvW6vExp7LnDludV5pE3sR9LrTeJ7b+13nvX70gtAn/BDzZAYc7upAfQZahgeUI0HVjqNjalse
NNhd26Lj9K5KZ9QL54Prm180dLj/YpjBN0Y3vM0UtQR5qPD4sfNdQ+fIS8B0znfsIGM/Ief9etMJ
WMW2vS29bMslULxcobOrk5xZWf3IXneM3YvN6B287BoUD3Q9gqvPGwWut4VlrfAngcSsl3BSNI4l
0sv9av8qsaHDVcoNSU9UFTMeq2AywsUzUUfKC5Bq2bVvQR0xyiYI039F/fnKIZ2lh+0676glFSsI
hOMOzgu5KwXCq6LKkqzmdYNvWSgchaqsGqcA9WaOJ5CNx3IpisVbZTCZSByC7uYCvMk/nqXZfvJF
nVldldYeTUNpMJdHL9XDvazHW2tsVUroATs6AeD7/S5lrLnyaDdO1YxFJ5pGDYidHstt4WD8v3Tg
h+b7CD9FFtfpHtaOupzWBoHS8yyQ5t6Hq8RAHPk8xBDg/3EPdELC1t5huBXsrQYc/0JiwR+6yV7w
c729RbYq+nwYZRfYK/ANENtKuMxTnILLeJeFCqM70vWxtBjYtLZ0x7tTdV8T/lb48X5NUfASB49N
ZlBnZS/J7pvnTuqLpVKmOVTGudue+cqo5qvI36m6jfWic6R2cF3UXktWzhxEIe4FF6haTLUQt61/
jGR3Db0CAW+QF0Llghh+32Lsl0LOCiFYWgvPoeJ1Z5i+oCBE49keLD2bM2rwriXHnT4vekiNjrv7
E1VcOHuhH0KSsEwz+d2vRUs5LuIeO54TfAbTlvsX0envYsJuIfIoBCUq8g7bXKAl5pZZtXdfiKWj
cg6jQBdBWCkE8mi2FDCXMVmfNtD7bXVHDtcXSLV0V4qOrn5f0HtC4r9b8qQ2xk00MFWYePa1jN7U
4VUOEJBhr8pCIE2oI8FyT8sIZ7dpqPUY5KNQXde6hCIqBa7PbpbmpqO82o1TKzbj7pD1kfyMrErq
5kv/3mBY27i7qZhPxlna0KjMOj9Wc60RaWHEIhblkxEM/yoTbpDxIQSqPv4vVhSS77SlSdNHRpFI
cNE7DEAPsgnxFJbyzneBcegshSQbNHKAQoDoeV+oT3nPwfYkput2PP7QXzhMNPKhwZa2kYUGkErb
eCvz82GfO7e+/A90OX0YkfgoHwhXR2ZYxUzCjMLsk5cjXKSqQ3cpU9nIbNVDbOyLOjJLjgk6kG/G
OEb+8A5ADrSZ/+Rjf5+wDlH5tydQXvHYf8CrhhGv+X88YucRjLS4Y0yNv6T68OZT9XbSgss1iif+
xCR2nRYO+ZjytKj61ay9zTyYAtw6MA8kz9TTjzUxKaEGJRuwk6YCccQE+rZgZQWaSOwUreUDdvCy
6G3qX5+natRbR22VazyvXdHtNWjjewMzeAht3LO3WDeHDQDTruqDtDOKWJL6gIe1NWVMziN+Xk0y
3JpFiANCcneFMAqXNsI50oSo7nTMrsJ88r0fO5qIF3S7+qxdJ1PH3D+5KZhfgsTNfuJgtL2fEOuD
78LY1Fb+ImwpgIODN4K/tScouoHKmaJKqeB8pifMuhp1LosBQonP4NOi0+8WoSYgLbfWtdDtRNmO
HjOByC6ymc2TfDlwyAlc/nz343vW5UEeRZj2k7oB+XcOcKInQWwOyqyAJvChpdi4gtXWzikrUzRg
QOtNKdb6QXX0mJN4CFGkrCPcGR1d9KwWMVgwWbG4oJUTPWxS9W85iXmn7bwz2i3B/vyMZEdeUJDQ
hScEki99tSvjwb1uBZw4N3eou6/zGwPI+IM8+WTOVKwuib5unOlGH6aPdUFAjHdIqWw1lcY8khMO
7opXy4Je8oiWEpxx7IlB/4dNIY6JAYNoTxfR2yoseE7w9PHdZjjfXIb0whZ0eabTzVBFMjTHFgYC
o2iF0DZ+4I/onZZNIWda1u0f4okJCC9h+GATVxvy8owpBlQ9OaRv9ZFOQtKvpSUx1oqlGU7cZKfp
v6A/yihIhJSOYcDvhQVFuQuglPPg5zyJNl3gvGKGCXbuLLkhjpm/sqV+GC7vvx73pDRSEC+yXuR+
SxjiHI3qlShKFQ56XSmWVVCVa6wF6qRatotK2BDDPmg9yH+k+wbJCxinf1/XWavAjpSMG/4F+a76
nO3aHl4piX4U1/RqIoqTOk9ufOnMZ9dd8sFF6FcTAlmRWMMLvCkAnCZEfQHPaDw9IRqQvPsXQDeU
ZZCp2BafuAEdtC2SQJ5dNS7M6kSsxOV2nwFWYRi3MASxAKpVt1kDYkHbuujgXbAmPcTyALZuQbWp
Aa6Yu4TnQXut08lTsCjj4imQqIgCq8f1XMH03uHRq88XF7R6PWs+tfl6LEk7rsrHtzzEpgiO5hXG
ufuOJ5abxYdD9GWYxEMRxd61ue24ZzK/USopb0XWglhJu++/2KS4Vs4Vs553XZeTyIys1SCI1Wkd
2WK4/GjGeZI8f1h8A92dKk918+r+kOLgcR57edUfcO42+YIwdsA9H+w42zCL6eUsgR1zTk055PDn
1ao5/WN29smos2YIyLKecf6THt3VPE1gczHeKbg/yvWGQkHS2mB2jzAmBzO/xDv5C4i/6LaBDO0E
LJdW6bKuItjYalkpzrIdUgXRc3DZ42zmqa+29om5bKL5PZWTQ3qzl3ZV6o4k0gTFPaNjxy18+oiB
DFbyi32mInUwpGktzwl38g1m5AQfnyu/cPcfIiwYTTDHqeg2lU9nHpIT4RJHFPLo30PMd+OWgsNl
c3Wv7dnbJ5gmArktc2OF5AnL3YRApqxvl5TSFP3luHnepOE5neCz7BdtCJeNkA1OJdTZDG5XTWCc
c3ybXpqx+oRJpse5CL21/aksYAYGAPH/CwhRgPGau6XoQZVOUfukliVKEnmIu6iCsEOY8xIMyzoS
eQegX2bKB7vJ7L0B5KAu/XoTtPrXKDkjMuyhnUE9BJRPois96xHP8nVsLEwJmIL0uhPKhab8qIip
4q1Igcmq/dRvKZIvc/bx90Rmby3hscOb3f3xxkKT4lF2qico7mNBg5Kz09jzYnSRSmXD8Slja+eN
0TyWAhakJnkHtZVLJVoIwhK7Yz+BibZASxiTQ0VjneXN8YelJjX/By2bdkcisgHyZy6bAP+6QZa8
prhCbFhqEUJt8hkJ9fBVfYLa5tdRwk2/H6Xdcm5EH4nIhM7K7HpYKiYmqnAXNtUeDHOSeoLxQehD
ZOf4EAlhGCgLeY4EQG8uZI1ApO5KPH7/floVtF7YGvZDGbaFQoObevy81MyQUMz6/Srew7AGbg4u
Nu+kBl5ChjyNKgNyUNIZicowhjHgmIID0fDf+aEtV4CuMBz0RwaouJmAkDhBvEkp7XAaqa9wmLGk
QsJuXZrIVo/RklF535M/YLTWn9XTyydWynAUa6OIRTbOVfL8Ix+IGs8KhTg6LZ/twK47+ZLvwby3
LOwR7Lbbh60DjDWz9w4LnJcx4DKgA/bD45qoTAo9h/8sCqvztv5lkg3bZBZmM9LGQ9HN63ADnUTS
uPZ20F5RttVa/LlpbfrVt6wcWZ7gFbq8s7bBhEH/vZqXZl+8BHMbo4wF+8gdW4qCgBZqiHrImo/T
LoklrQaRug2livHx6gKMPQ2Ath11K1BqtWRyAh1sI8ps4Aj2CemxtFiGE3OISm9ELEbii5kwAwnY
eqgi9SGn0jC81vLTlwHEqLrJQQ43zmrqtEQ4YGdFwugVuE2VUjqLXZJGx7wM9Hs6XiNe2FOVwfeo
m/3S1rtT0exunwx3Dpm/jH0Vdhd96Ul0NSNf4xF9DqBJ7PiZ5dflkSP/bq8gjhMWdnu85HUNG7/7
3nXsWuLmIY4RY7MROwQCDK5Pyld4jX/K1pRVZQDI0cFqSenW99vk6shzZSt44+HNq0ivXN0NFg54
LIVcW+XFNTyMnAEeugKZFkHZi0lFHLfn2HnjYz79FeFSq2ZlUmgFDCSxNaJD7SlQpQpEhJhxsbT2
xSHBm/sd4vJqauZFRSvtPQI2iY3Sftr7NaRpBc96myXH7rqLz+0myPV3beK/4rV1VkoWe/5KEZe1
PaetgQvzq9HbMnm8YiIuM9JT01O9feu6mZuf+bpsVb0hckxhRLgABLvHFddmuGer4CTj2qGmWDW6
IyV+I7fZm05pNllGXUpqSVYN0f8leh9sj4IJwENBn1+3w8paoZIHj+uIrocw6tDDT4G3uoglx+Km
+upQHwfP95yd0EB0le6P2jwgsIA4jZnQQyMvjEFta92r61hNa45SLdbjZNvP6Wmcy7TWAfYOtS64
/nNPWL9HdffjzRB1+dXjgUadXwYUYLeKGH6r/TpQ1SMA9wGgfUMK+DILsOnwWzNSXmgPe5h3GgCM
l6PBpN+XsubiiU3y+ir++1ePFgl7VRFtH5YXDLrEziKnBC4Plq5hBQkk8GE3E7EgBhpYrmv8bAOx
+i37r25+M7hGl2idDxyqQ2fidKc2f/y0FsTt9WaeKAq71pyoXyU74sOJkBJu+TFM9PdmKDlD4nQ3
aCd9iWGgEn495Ny6u2gQ+XaUbLryXyAhCJ0PXjj2T8ykL9lo8SZyFGNs7g5hq1CEzHWZWNzHolR7
RHdkUjbYhtMVDNCdG/A2uLlWyJGHuiEIwRZjL+B5uwZvAeOZLbm6N9F1LfMtIS7K27nFDAowuWw0
5joY8Cn5SsUdyXgU2ywmKWp2y9VdN0F4IVwzJjW4ZpoqsoKc410j5VxXiYzyRsuzOykFyYAErM+c
g8NPbeQqeyPk79Rtzw1G6B0tePndAW19HExuX7GIq/sb3d0jtAKNYpmP+HOpAcWHsQoGIlmcqzTt
DPjvTuqtEJ7WLjgBp1s8dZkbWyNabp3z5mxf8FLJh3BLzZKrNX/mGMlSPUZxvoAr48aN3XoRc6v4
QcFVZAFuk8BqL9SG0yl0QTdmYHIg6SN1EFoXfrRMqjqS+s0An0NjcA9EraQKtJffs2ZYO9VtgNrR
G0xbv96V+YZoWaBcuOffGJINurdnDazT1R4PDgG8Ofia86T3HtaPxcVNEk7xdn9wc5NTyP+4hfOV
MpLMXNXtsG3y77b9quveHTmlaJy7pKF/1c6PIurEi5lvYmsg3kGeZmwr8u129cEsWm0P1zoELrZG
wueWzFINaECjGLhq9DDgN12jwY+d2F5uSsYjQHPdnMsjvGwNbg/2u37AYjhxaD0nnBYoIli5U8c2
NXPXODTqzwKg2xqsDeyVT/C1FPVw+rl72LSf+ard827iFhGnSsgSOUqF5VgYDxn40vZD0iVnrffz
qaOW4Sux6R/5WG96wn6j0AZI53PmcbL9bh2NEjb41/uYAEGbQs+pLOon2eaNXFZZG1agJrT1HncQ
LRBwUB4doLnHH+0tK4HeRLdrGQgNhLukBszE2w2fV/CUquFHZSm5yBHWXEhAAoT4bZI0P5fKjRVf
L90u5E4R6pxQ/dAfPbDx+rZpVwuzLYyUF4N5Tld+33hmcNv2hfNw2dltIWDjTn5iZgLxv2rGr5V3
w1iNKXKB4BmQ73EcNavn2fMBX/ok+U1kYuIRNy2rCzvy+1aV9wP/3mN3XX6rTi0YAlnQ9qFEIYPz
vKILYJJJnV42gttygPyo5FJgYWIN71IEOTmnylYeNw3WG6UikLIPJNZh71KP/sRqIiefoAcrDXV0
K10f+4otfxirLBL1fbPX9c5e2agmFkC7jb1MW/AHwGW4nY9IL7vdqXI8xGBpMmmsXg0b6zC/wGa8
VXFCdbO8qf8LfDwFsQf5G4cV4RVU3YMMtd1B6GMJEwtmvB53fzYTXkwHWTWYWx3jL8CPwPAGhp2F
IuajRfokdNWLecz+abqcFcI0WJF5NP3Kgj2ZwQszoFbd+BQBUl40dSaCAYBzm7YJarsQwA+kZ/Rp
NYz2EBvgQb6quhUytenhEU74NHdrpwzXp/w9O6SFyDDwRS9gOYmrFpPjiP8lH/3Fd5J//BWv6kBN
y8/GPpYP5G6/E4Q23Nfr1g+1Ff6CNWI4OV4y6BOK99G6XGQutp4mU05d8mPLL2l7hTK2PM60oQ/b
CEppBIjcHm/mlAIG6iyDZS7lUgZft9kLvGfGJJRXmHnWFkicHGZqOThz3MuTy+uMt80Vx8+9kKpI
W6F7Y+42lkZY9YHZOF0sY+9Vi8O3Zy72GIqlqbZhrjrlZXSM1s+xpYv4JTSPLdRY1h9YaANFJs2i
KLRGR919ByBryFejmwv4Bi0OeJJm5LR7s30WKkkBOIZVqK4uoJjmPq+Q9yuI+2tFhBsuO3h9MvpF
5Skt4VxTUF3IePfaLaE2mCX+i6F76GK2LkhK2QWGp0J9GNu/eLAOyRln30o1wyRbiEJ15ZcAF94z
nBc2aPP9xOBMoFiM0xEnogZElZmPnoRUzMCMJSxcnOIizVYqmJ06JtQkOxEcDjbR9EFpwHT+7sl6
KuD0/uFk2aCxm+1bGZh6+7QxzvJikQfEjPphXb+04I18AW8140rJ4eN+YtYYGWwiJrth1AdZ7SpW
MiuYPsKeJ2fH+YpStAFZsw89me6Z8FO8+K8bsN6f4YlJsQzM/zrgYaTc2jDvPiszRXd3FdsnFvsB
E2wuGyG35wnWprWG/1WYTulsSOm8wXv3XSpGPRC0RGoHVpATGFIzDN2S8URSdsj+TBAWqANNRYwW
mE6ZgZAOq27JUaAu4MiYdrIBhU7GII4WyNFJQdkhV8sz9HSMngmOqVUSJ8UycNEGS8lw8ZF/mcOj
hLRlDWUB9RuOwBS9DN/PhnXSCeaDJ3Tb33zefXFHGF8OuxbN8XiIr4fgx5qRry3FUIYiZprnvKvm
9QZ+K5tkeu2AViLIYAHBWGUxjnK/8jT5XZwAS3sOhmnFoB+7oK02phJQj66eY2RM7GDJAlysG7Nx
onFIP881bCri5yZySDPRee0ZGg6CIJZCdyO5oGvv9K7+CAaHbtZVBM1/Ryrj6eXXx8xnyVax1z/N
K1kJ3XIA6SIf/gkwraXiWT59HeDNUmvbDKpm5PNjX9+xGI/WCHQ2lTlCBUWkSJ1knlLM7dqmhImt
rYOIXERaksdlKt7lNyRCVXMTldz9c8h6FqRE1+AX56ZL/wdnlASO0VGXv95EYuLzEamOtcC6aR7p
0Z5oMQjgG/h3x1OJ5uwfXweZ0+cPOpIA5bjPglIMVBq0wqW0AKkFMpy/FI7wNYkBxO6LVTDm7hwZ
N0TdJq9i0oevlb2Z8ausNHc83OxQmLNbZiLpQrKKoyXh7TEVry+DMjh2UkOjWCgv7WfoIZ2BQJdJ
BpWIYOlX2AMQsH3jjKQIzZHRw65hDS4WkZFlAYYXncQvW6uCxHMZnhlNxTWzseWWOa0LFWkkcmAp
wJTb6QXW1+13+Z1QCVsVwJP2ywOn6c3IVNZI1z8fqusIq5sZmDWnzxnXNhhIzb9xgvqSkNrmih2O
J3qBDmKt5FIjSQOPnAJX8s3XvJgYCbjfM+IX0Bf0McAlovlQ8VIpBFJIHPfiqDtIWD57FlP6ZTKP
n0vaUOlVyAp7ZWHDb7yDFDTkYwEL/L2Ii9em8TTqx4xn6wSL6O4kbl8ctdl9+ED0aNpeZr6rN73l
uqg+HOZFT/3cihW2Y/uPDbamKUbb0uDI98sv6DBSy4gZuattkk3nAEqMkJ4OexJzmcBTOk7S2pNq
L8PyiSqwtBmxV7cwbfNKwTIM2LX82dNWkvseHIaGPRLl1e19/lAzSjKmQVnRQjTXoKkHS9Pe3IVU
jsiv4GT4zIzqLMmaWDBfWFH+8HmYpQBPK3m2A1LBPiSMnHcjdxvT8qFefTZNzyV3f5clFTVhLVxY
0JIykka9NmGCzaE3AHtMM0dw5BafarPUvY9RuQ8uq9a0eJGM6gRWHxRtP+peMHyzUQPQR0L/a3+C
8aQ9QWkCEAsB2LtjYRWX6hzBqStpFwvFqeJ1pcH/B9xPTY1pGkRpu9rIy6Ir4cCGlKCQpTGQ63Md
nxVXlsMDCmMBhSwIYIW6mQl8aS8SxuNzYB+balceaIyT9iArtNx939+nVmtcWvpjkfWiO7puUM+r
CKWj2wkCdfQ5wefQAMHGQBpSlV82U5fa+EPhL/0dH6Kxk2iB4HZvqBaPThTqM79QjqEk3hEPneMV
D2YcoDwcDGBndLN1OZXb0NPG8EDVkxPQw1TruWfjYmL4YbCkQ6oeKRwEitq60SwdHbdDDl8SeoSR
gYyAWcZuT2buCE3UnrfNDaOx4MHbCm1naToAAJeedYYcrAZw4/SnoSR6oXwwFXaAKSzZe14X7noJ
E6FJWyqympx3wlyc2/iYDoUnJNlG1tF654E3Yww3UnEL7u1yeYWv0nQMZl01LLajXiPQxTzcaZHB
qnSkh0OFZcc9gkVv/yo6/tbJ1JzB2r+DS+JF7HwDMBb5K6TuYCMr4RZsSywHwHaQ6JvIHw44zIvZ
kYRNk58EQQp0aV/3mi2lk5SJihRVJaNV7KrsmRz/l83Pug2xT7MIwDpGlh3UtEIxav0FRtG1Q79i
P4XoyIbsi7mCbfAsYQI/5U3tp7YZPzfHb1cWHXmsmNdNFwZrehyLc4vhYpKal+peHcmPcW8dAH8+
wtTEgI/EBcuPw8yDDzNO8SLZ15x9oVvA6rR4RLN1oXe9niEqY86J/fBTmQlsKglYpFQj0glX98yG
ygOV+cDlGLMNQvswks/PrZ/M+DyK+ZvMI+/ZU87YMgTyjtd2aFP9/DIyASD1yhHqlLgmD4AvC7Cd
+0Mlkljomaz5UWiGDu7QauDHKzWMbm+vZ1kS8Ve09osHZtvQXvD04CFbfTi+k21ZLeco2OSOHTev
mkY7CDYWFnS2NE72bkj1OH8NVFTHNBkzqq4i676Q8fJfK2Tg5vz3i86XZZQTqeMLUvCkNbWT8ONf
VGFR+RirkfFrC6X4zXxBVve+MauZowvjockOMR/0I1mmsiDkIa1vpCjtg9cv91n70GgBB2pVBuzN
C7/YesNAU1hJTgwks293CDH99dahrAvC0TN8OONwSU4yE+h0/jlkuKruC1cg/g+RKFuKam3gfWAI
lqRf5VWZjcq6wlsvTaAzgDPEKFjuNCA+uMuP7DXufl6JRAD/cdQRJGH1cGSlxyOzDrVJi7qZn5rX
VwioU2mzfqMoaHOS1vVWfqrHgEWlSfMpIa4CZAI4t/voKPXHZ8ef3ovaSM54UBlN9J/MX+sf1Emf
9jtLZU1eXT9b0O7eZlzqh5ANNqRu/2hPDFVHvuOfuzge4nGiq9pRkJFjSkp3fkOZ30Y/PMANMNzh
jusFVRUOKYXHOrwKKJlaMYQ2f3CozdTEqEn+TW3F/UuPfcJ9kGoKrrMK7QnDZ+9k+ZMdWt9Ce0eG
h2YwK0jajUXaJNdrOBqBtT1IM4noSp1WtRuaYv+jJuZywImykmwMsJrq7+wIDA2h14C3u65xA8HZ
1ivjhzW5Cu+OrHiKle5xo4NqlQhV6O/50flo9gDJ5zhjB/pR0eDMW9517EbwBWXCLnBSW/PuzBDU
qaYYipHFBamQkQML5gs8E+JozOAeMAwNf0MXkbd7bjDfFZgX5f8DeuDCCX0FA+OhfdlV3BQ7CKHD
jzkmHiyswXDT+SMZQVzu4CYvIe3BvqhMKPo6A4USoLKyZYyKwjid/E/y0SQ4e3vuJa6WjbLWyZ5Q
No9l8NhQMRQDZcq59kY8C5/xMan4dRFJNuajFO0YwErzX0F3r/EBSDDeEXYAcRLfN746pcq3rJPd
ssHBs3CgQ5k8WlgHYqlqDATt752D5bE62r7jTECmJdr30Wsu1hKvPeUa7KgufMCycZ9a7KnFO6co
XaNE7epXoaPMFzCXus6Wr/cBckWv3OzZR8ZI9Wfbc8v7Vy7dO5ictBLTuyYhb5GuSaxt0Gx5hpxq
zqhQ8PmZZpAqaLZ7SSEFrlDRbFdDtjQqPyNWFoD96xAa+AfGGAzHMFa/nanX+VPxpScUbBUpTyix
qe9sOqKetU7FV0lHssSuN8cl0mmeU/ZzztDS7MypWWwmQStrlY3bo0DTxdmV+fx4jHsCDKtV36AS
H3cVT9HaMGg3Do/CMIDOpuJIWYgfJCRsA9ovGd23n8A/sLfZdmS9VBl4OFFuBeuKzCv16sQnIe1a
1ndKaBeDPO3DvJDbzTEUyZ6kj1AKxTFAJvmpJgLzTAeVy28KNchqWPYlBEgamCv/+TzFPsUAvj7t
hj/CfajNde/QqLa4r2Y8wHhTXfq00uqK4hDgNuEYXeNiA9l3tOFYhvu4Ms6lK8w9Bj9VRBxDAHUU
BPkU+wnuzKMgYk1PvmELNLDZOwHK4F2IAKSHJnqLWHL/CDkOthOLqIN5IzGh/QwIPcaeH505XD0n
KJynd87PIWlDjvChThjbrwVQi++k0zVCER4n2Uy0pfbuUdOUbNIVJJmjgMak53OPpxilJclXez36
bP0FOn2ZFthTssmfNrhKZF9ZcqFGEKoRB+5nHBQwkyZfWu5Bsrl+TDQq886Janz0qB28cHHgVXi3
v/DGPyXoYEX2O4BWhohpZHOQBVY0tDVqxjnebwFNPGJ5xHuW8upChv+i/AITn6pr9veSNUr3oR4Y
o1OyJn/MiqkF1gAajBWlMhi/Xbv7+eyL69Xq5b4WjVknRb4gRwbroXM3C4bqTHW2yyx3BQqfFUlT
3b8TCHdPdIh+BlqDv6wO3Nrk7PnFD6o9f3WdL69zuLypLrB5kra3RHJBCg807MGF5ksm6u/r3qAs
6kwxq1ktIfrc+4j5Sh3/qrBB7QoCxUKV2C5lNXms+6+8K1q19LUFwOYkZpBRy8qiMpY8H/zrIeMD
F92H1NDHGfjpCJkLXNFnlOo/StWmoXmgGH3ZUIfH6YP6Hru6IxsqLPXT6JiMmENoOQuFioMoPDOQ
rR7ZS+JgEAlZZUv+3YNzZuXjh/RncjaovBXQNKc1UX5FXx1N5x/He+IqwFVaNsOrUBHMjC+bHNre
iONWk7kObL70xQIPhIqqKsXzOzmDuobQUptYMLhPmJzPjRQ5+CP08agE4kSudyMD03eq6CE2HE9W
OYKdVKzOASiuqKcBo6LWSL/JVRR6hTa+D/HHHorHvmzJHiJ0pjakYLrNzP+tMJkgSlR3BH7Q2ihC
UsCW012N/zTsJEy80v0aadHN/zZ/bz+iCeI3EDbyjaDJxzojpV1VQgOGglSYCEM6uifAIXJkp36n
3oUixtHTKuqXD01/c/7Orf4pZ5b0xPlBFz2MGdf+mOADX5sqDz2RA0KgGleOssTXJkFslo2w773l
sm8uenHpRqF1HptugxdpkLjQjRFq7tx+QqjvYQtJpBZXPpx3lt7i+xbJ8lja+gjsnptKYB/vsUfQ
OaKPIx9vyUgkPoGrnpwLxsPQOVVB96W++2cbmJEaijzHts30VZGROqwa5Nfxw/oZtk4IJ2uiOLWp
MtWSz/2CYus3eC+YJQHtPswPUOCd5DQ97ulKLr5P++JtJxeJWrK7YSGuHKcBGjQXx92b0Br0k7ls
qSeW0JdzptuoJSV0iCnRZY3JoPNS1sFhv8J41WEf4zTtJdqW2EcByAcoY94Aep+M8rkBTzhbMY+y
HEQ5cN8bhm6SsM6hQIhkWSXjJTig/Kson7r+dnIpqOEyoCgzrlPCGa4NA499DnnhnOYLdy1IVv6K
XK9bR0+K3W4mtKtnpg0Au3ep+mIXJYlg2ZQTeZS5EdjtNJEzEooskaMF0omoi1wWAfNwUdCSlzzH
fpLp3HAx9+BJdf/oMRDwIOyoaeCmW1iLT3GSPf/yCsoquQDcaIq3W/ZRux7I6/2h9qo7X3fUnqfs
RWFyQGe02Rm3ti0cFAjxwxRZmc5RF5G2l/Zj1XLG5rsoBvSWYvxaSBb4bocZoP+ta8dW8RTaLU3m
4bXfaURXUJwdjvyLnj/J1Xn4NeaXRf+qhDEDwjCXwHxu4QZpYMBxqp0ZUb7/EAFaVjWxgO9QiRsQ
qGTsATsaizVU0gjtpEx7WAI8sZ/dO91CnaYogL6hoYz3vlMpxQ7i9jM5ao3f/KyA6CExsPuawh+q
E3cZh0TSTfmf1HAhIiCN0p7uT3P0ILEjC9EJsME9lmo5L9pz0mzZ9yyeTLPtyimik9DNBzDld6/3
aVmn8IpD0DKEjiPCmH4o1C3dAJm4RfnDQ1yTfAsC+f1NPJ1crSuc+Wh1rn+CpZtyrTEhvi8VlGAp
95G5m6VDdiR/Clmp4TOzwfNReXU5MhuI/SKlMWAs8caJEoqRq/MsKfn4BZlkqCwmTJRgiyIWVMou
TfMY4XDdUHjMzzv7+nxrNjpYmNFDjkWN/543PSG0w0kAs2ijNc1m0MiHUCTwC84zS1T9Sxbpk0UO
BQj7e1OtqRCL+epCRe8dmTTcNWk52+gJgf+ZdtmxiHmpxDmQbxjuQb4U0I9ImNK5006HrX3QuyTY
gJrJ5HZB2AC5BbqAAUX9inLO2EonLEuDCNVuUSchagb2qqDec1o6qiRQr+VMxIN/4G+r/53vYooZ
6Q0yjqB0nffcDCqWj2D5MPj/n7hHRrvYT3TyUxLOJCecvYYv/qp91X+cuWNSpIAGW76HiJ9v45Kl
DdaHh6PINAbDtKCP7KHW2mFbuN4acGSGRz5PeHZczkLros6AYYa/K2HXJYYz/eiM61h/6EbdQW6Z
dYoP1ec8i1i+20qJaY6xMeS87XK8aB2WVjFKYXIyO9wIAMowFCpue3hVIzC5/UDIPvd8je5l3fat
sVWGBAqSS/YgTAMnEymv4vjE3E2CqDzINlWNn5lde3R4+57DTLn1josVMlpxnIJNUsPDI2oyj0yV
c7HY0bkdlppT6f6p5nSnw5uoCvuURhHGdXuOOSu9XUZSazb5mB4pnT06KQmnD7twWraobCN6Go+k
YL6hTGecOMpaOzzR30NUAlL2JNTeaZ9DxUp0JYUkJVvPyJuTC1irWXvYDWpWWgK+b6RtrjoX69eh
SG5Yd1QbzqwUyU/lwhJ9T6nJ3B9lJd4o3t5ryunYTHuF/Khs+jof9sg7KMw5xWveN4egW7PJZdsB
oVQOCLNNPT5uJd4AMb+aCvhJd/msc4l2hCLc7GbyUS2GfJcLlTEhFITBNvQUtbtLp0le3Qo/T/4J
T5C527Ox32kUejTViAwhQKU7myZEcykMlF3wxaYZli8Y8mQWD8sV2Shy5MQREutbTEgiYORU3K3D
apC/DiCREyvBKxV1oJuxqxloII70xgru3Q6/yd0A5ktDf+/PyiwN8fnjSM47FEmaBSu6UhH3RKqn
Z/fYgiD+8NX/I7DVtgKXIllrxUiJEsepNEndP+eVAedJJZ9Ct7WSceJ+425qbCvLjC0QM7LB5PBF
hkOL0+GFYl/W1fH01Tr3IafHV22fY93GVsxjucMiJ0xPRvEuqdudvcusr8AyuY092pfS1q5AwC3Y
wYv57veF1OWBZlNAqcaGKjAiuwpFyRbArFeMEpeaswOagSEYTs/2KehSYKFMerf4WfXrZLpPRQSm
N5aavTulJbElXqAsIDAFJZCcBB6oRfNqdY1iAHTkkvGXPXFyPkjF28mObKRawShkwiHHlE65ajUk
mfXbCT7au97nf8s17PzNC9/Kr1Xr8TJVsQDWKCuhOv4qaIqMqh3n8mJ6mmmUuYBzNHi5V7xRXJvy
SZkvic3o0trd6qEiXZAz+FaztFlvJ/Xl5/1+ThilndnLCIvCk3UPdCpSYx+i9WbYNn1n0+/fxJbX
PSxzOE3pz6Nzx3gkG520hEDGFPKzQ3UOTDrMdhE96KkCVzeuaIjUeK3aW3xmdE1bSsV1cCAeU5Va
bbtq/OV5WZKPMpl/sf2c0riRr7cdU3qW2EBhyGs77RmDMteO0V4nZ2Mf3RO++/A7682XFVE48R/g
+hby3zbN34xugVAZUDG6AbCeaTcZUdWNsnA2jYK33C6+TcOjNjxPQXBnThcor4oJgx5CeuKSpQub
Rguhaq1vOpktzdg7BvoUrt3LBbHBU5OIU9o5tn30xfEk1DZXdvm83NnQR3mghaooVzOnvKB+VDG4
nFj0QvddulfVcHX+03eLuWGAIg7EMogiM5ToGI8tEZ+D2EOc0Q/c/lsySFEsRwyjAB/cSHHmN5Zc
5k9KE+BjMYg4EHUJSbwyDAnCFFq3HVGYDbWmKdL2G9vn1rAETmZmbCI7CPp4r9VdyRFRd01rOd7o
FDrKu7Xec6ckq5jRtUlQaFnqUD3F2Q2fB1dSC+d08PSxNYYQTVgwSjQsOh09xbhEcLl5C6A21dVz
kIsd+PTkTqttwd1ZBIcPI+Xpkf0kqa43bzRrwtPq1fDrugI1OG2AI1BEkg8wP1jlMuVJ+rRGyz8h
7LJB6aE1gQE/pZP0t5tRFQz8eDw0QUzMBh1sznS8f7JzjuXaLdKv4kYcn79lBiaz7NjBQfzLsWoh
tLkANvIFbHCKuekdTuImJVRfD56gs2PHf6rpt19N2T97QM56YX8Vn/LYEjz6lZ+NM34N3qHpblAv
mnO/uIuKtQjV+Nid19oByFxwexJV8Mnd5nUGvWDngTBYdO64c2aN14TLkAAJvbbcphj0EnIoMC2h
EDxaobKAM7zRsJrju0SZtXfrepG0YIOD6NIazCh7eQCZNsgUiyGeA6HIcuJLmLoPWT4eKDvzJNe2
bWt0Gl1jj+1M5Ya+lVhzXl0di+JqnCIoXAmp4HIirxSYTwRti1WiF9xfugHZz5Cu/6DOsZSrw7Hp
A6fXuU2W4jFoJbbZ4fIfgBJXaJrzgAQawyfBvV0Aqqb+JEDpVBoW/51c+Rha2TvwnrduWzBHsJp7
khnqjYiMq4gSBC76tyOQo+KgoQwQ2rQIQAc0tesllPBI3XExgyvhYGnJCIX9xq9lHR20VzCWas/8
xoMg+vvdXiS8qqjlu0vGyxt9JSHYEGxyAAujR70x1nElEojMcmZUgIGpzxipE17npEKtL0A0ra+P
mz6Z6l+GOiJ3reCK3JXsDy98fH+DZGmJhAWS2HybovQTauEddU1ypn0oPtoZ1BEm07tyHGS8M02D
6IdyUPlMaZBA6ckqrrTLolXWvelHQsGAtA2LXsWFyklvAT8dcLe0BV/RtT9tXlt4KsQ935MpZq+k
iIH5EMmVh9jZ8LFydzjh3fiAwB9VOQmd0Z0aQaoDG2JIU5fheZuu+axWW8I2Cp39n+4/gb5cOjo7
FUcTsU6/gPIpU0T1SyNY9w7675mtM549ijOcEdoU8PtFG8UEdQ0jkCjxx8UMlK8aNYJsXQINZb8O
3GAiD9zWIuzaGqph8hkqjdEJ+F6mZrw/8K1GmYroyc58mPOwbsFk/ofsE7R8FqMMnva1xhDduQT4
VBSGm8VOxLdDaLI3QgSA5DFF+GlDVqKrYGKlUZjF0wY5gNJffsaGKZeQu2UoXoogCOletr4gBEAX
OFsfRjnf35Ln4Zr66rh6ITpgM+Vi0RKhYpe0oUs3+TacAF5edLnm0AVPTSgsRs0JlHVIOrwBya1x
WQb8sGxUQKzcaaksQ0XjZe+l2Q/3Sm0rS1VYzu1lBXKosglDOKCMVBDB7hm8Qkd0W4Y0PmCxCEP+
aXhSh1rn/hgIKnBOPa2Z3o0Wd7jycDfuScBFid0tEitIaNfjQnGXe0S3CDAfHPtolimiTQWxlQZR
fnb12PJYikVu5mvOv0H3B59AlHbZmDOznjfX4ysG1WRGQIEgNyLodyY5iGIUoGm7GqZJ3kGGeL1C
6mpDCGU7EJDWhi6R/6nm4bENmtMRvvTzRnPldt4HdEZPQ3ODzptvBs8yUPC2hY+pJo4ZjCwKqUfg
T9n7zrUbz+/G/i2G35F5pwAYXcugCu0FnZ5iVW4WSrvn0Rh26oHwC8h2TWpLn7Q2SxdXa3TvTyPL
CKdE7KPj0DggoIWsUoHr4g11HGNAIKGI6S8UG4NDagU88qcHmWm/CzTTipy8o9rwPV1P1zUilICE
6Lbcq58eo08m9duPyU5pTEid9KRV+GPSBqHofu+Syxcj88heH41S+HruAfA3VYqSX2davkD8vKMp
DBS5pzRtTp2a3ol8ZXHjE9crhmYnl/yAN7bhDuUtRCbgEIx8nPzuyPPcoRK32YA4Gaf3+xXmqnDj
T9WXb77QIK0BzUbocNrOWO9wxTfEal4dBpyLA3qR4NX2PcQ1sdrRtHEWZRVGRFrS3Iuf2K8etNud
IMOp2mAC5xW61qmv1fL7mDa18b9ixUIdfk7d/DeMjSsOsO1cj+8lWaNp3x35D1W/8x0PWNxT/KWe
ymQWzfJ/2I/btrxMzDHDKsH5Am7EvK4vSQG2I1UyfaRpT+f6cWcFb+pAEaaenqLvIarW16pyKYvw
fcZu8d6/0Bt7qDsYw43oaniJQaiFlwoYi54TQAcxFJLnMstsuLGmZ13/y7BkNC5vgcmJrzvHBica
xUIhDTpeS6E85sQ0Zt0Zgy9DvuEd8eppWodBTs0hdT/UsdvbA1soLhAB8aZzrusruk4lWc+ZTM7g
0trxK7vWSdtuctNmuarIH8Mvv7GEYImA3bhdzQ80omy+cNUww0xooyTMDtt0QM/iV14rp4X1eIep
0CpG3WJJm1+OZdrruD+2cKxeusqedNh6aYvppbX6tldCtylqta87q/mFL9eYsuqwzJyWexgpxHbo
mFwH9xkWOTvo9QhsOnVqe4aLoQ58fnNM3MAhMnWH9BA+0w9taSLyzJWktISO5AUxV6McR2UU40g0
aNNDWW9q/7gg+vk6NnTFLxHnaGnINrLzlYQe1lI3sYreyqujB7h6xNaWGvQlOxli08PSgIYSvUM1
5Zh5krlcrwh7iDUSjNhovC80rDsBdGhTGoIxEFrXuWNAcGM0/4+XJbjGYOwE89ZJJOJxia5/1oGS
w6vjty97iyneMCBqnj548zkaAPX/ZWGRS1LN4whjCgMpqAXOxpY4wnO8GTQESt2/c2g3rz00OWl2
4rzMUtCJXuGFjSBoLdv+XK+NqPFPZiy829JpU3kWS9XtfjK+tMMb06M+IQJuQ1gqFdudwjaAD6s4
ffD+CCJAUPfIdl2Y48KzSA9yoUrgcAUEKocDQpm5TGR4pbz7H9O+n+3OPZ0ZPomvsclaCN0/esyE
GsmkTgARwo954UWoDYqHWU0jdUDOsuuwTJcoCAdJcMTBrKtJFO4HTAhpvlmWXTpMiBov40i55dRa
kJJ8F2PZ8lMvQptv+m8LItOcGop/9riAKkg15b7WjKyCjY5wv463dUFWtIhj7bHdt2PmMb7ll5Ki
ox2dBk1+l+vxwzZmqjs8JDPO+G1XNJdx4900EX/K9NYdb/cNzRLu7X8/i5wCqIW7LdqW9ODjlwpy
fFAmzvvVDTTKC7EuxcUw6VXRj8BXkh3MsoH+duQZbRQ4e6lF9gsaeGbAFOeUmSDCrE1HNZM/aiBw
0WoLd2bbdPk3AGHpHyBGdCxSA3AYV9AAGSrgf14MpQvkNfqAdH7yYCzbEYTQUXpP8Z+E9aaBJJ2y
SkeXAcp3lYTz/q2V8dJXtREUaX9R5OKjbCN3u1oFwvDX7visYFmCqEvUPBxEkCdBsSf3cWz2ivk9
xgRlbUL+Rs/HSnn09LfhsdUx1yyDMADVmMP03mFkk51rXZbZbrzNiWdudS1z7EYZlntJFzpU4sEc
iOromvnLqQHCqM4NkRszN3nQHj8Er9sZivetTugCZteyGFMhIT7VGNu0HvzwNM0YMUxev1dX7GbZ
NcAZjr8TScaPfSVp1V89rvB9XqJ9E35+bArOeQDmw66v1MyQEb6p0lu/M1f886FUZukuRRUA3+ZJ
Ce3BxLFEeHC1+yXqnWdhn8b3qrW3covqcOmd2TJjJQXQ0zmmEOvZarC9YSL8pIcBm31Wmso5uA7g
y01UUlvU5Q09inXrgV597zdRZl42JpXM47rQ3lOGvWPJN53txi33tTGkQzQxBLeEp5to6Rhy0yhK
mzCT9LIfa0OVzxDq4HoDRiAO/+f1WWOkjajYe/6ysO3ZjkhLARZdHquNT04Y9Ql+/UuUHPobC4MG
3GXd93/BNeD1Yn4EijjP+3oD1ADQoeNv6UOOpg33chKcp58TBIK/vI/8EJqWFD2tTLNocZraQBP0
9YEEbvh8iNAn1zQJDIr/uEiSieWNGXRapgSo1X+1OTIQrYCZcKW6EB9G89WXxVdUBB6lqIPnjCsG
pJtK07WgjYs/6wWE7sSzO7GFXLo8IRWDDJTYc1mSGyIovjtDP5fjoj+prLAjREerduZqpMK9W+Vj
asCRWUY+a4DwOK9X2nDZ3W8FVP9nCMhW0nLjjI+Nq3z5c4+Z+o3eyDbHz0S5Aq9QwSW2vG2hwRv4
8RL8Egz9S6emsXkyNvJxYyOBLemykm9F4yqi71KVj4Y0U8e+33Sdi2z7FyRwge8j/gDrxZu0TMil
6/xUCkumjPtnUI7mw2AGflE1YIjwCoEQJi9y0uaVpiwhox+VdYwkTJeyuYDvNc+Nmhrq5HGiAC16
AJHuKzQ/7MM8+yRcfkjARqaJeE1FF7ImrxpbSVNT8ljGwzuruXd3UEHDq9yTlAgPpq+tE91PcdMx
4xYXnwO+LhRjDaKP8EkfhGWrnd7qPD4S9GZAwilnnHKQ0ObaRh+jEq9rmacJAL3cDIsAcYWsjdYS
VPJZ5wqxvgTgKAkrMCyfHm0gnpP5JXGpw2xR7YCtrKZIk6hRcu2FiFcHVpDFkM6YtM7GLujZLz0e
ArviQKemMYmRwa1+ri0fVHYvz+IK+hi8Gcz8BXy7fSCYpSU3rFEDUvXlaIi2mO6JJsKedxy5LE8L
4Pui4NS5/UKAGzFcHoLXv/pANly9iJUBJvnuvlnyLJ8wgO50/LNxbLpdRekw/J1/VLS9RnGpmy98
z8EHAVwJVvDQTVddUonswiuOmyz+EEKlqkPYb62+kUqc5OQFWZI3OSCsThVCLu61XcdiT9/13jxE
QbQ0Hdekg9/qrUzU7Lzzp/9fEs4bpOS4LjGNtCRewZ0n1oP5Rw1S+L2V3AupAFb5FxCanC9oIHSl
LQT6yhhu/4LJHQC9Tp5gn1Y60RQrm8ogsxO2DIUZQvTWArmNJf7HDTHCohwOn1kuS4xmhqX2eMxU
hpk3Rth7wZGzTsSeOVR3ELDFLb8kQ+5P1Puapo8I14KZNYZNRql7CO8ROE4tL24EO1hH9O5RJZWj
aWlOiZ3i1EWufQwmhoQF1DgNw/gYhQ610bGmhW/gzTyapTZ4tfebyiFHysKaO6LR5LaZSUFrdo1a
KzHQkg5QwMfLWnRJZ2XJ/N/pDfl7wDAywf/oQIT94lDJrUq28G2dy3l6Tli6dIcIZbjH3bjtqR2b
d6wlLc/ylMrW2SlBnnNxRj6BcwIzLZL0zNxhgsVrp/iZ/redskcRYvhjbhfwKmWFdDRUiATwytup
FdZKJnrvGxhQpTcOn4o9VkK1FcQ9DW4RDImDm6/FJwZEyFPLIOySRkT7bl8ywG8D7fZ+Jg59/6ZS
fTsr9lRZpkHIbArp2J3ylNuukkZiXTyXoKzmeoSQ17j7DKHgEVUCb7Ng0kx27USkoj26zAAtWL4Y
+kgWSi5NODe4tx9pAUM9CFvywLhq1JnqT4uiSDfGvXehu3Hc2t1UbQR8RcTK0B8qSGURVEkQPMdB
xkEmvwkyifZLaNJSN0ss9fWALYHwNPHi4CljBg9BKwI6Im/be6LaVJGjDeQJ5UNu+Eyc+G1yfwUC
dykzYLC+X77Uq7t0X5A7rkczVyHZEqOVnmMlloiJmPoPENyEKa5+MZ4zhcIy/77TOD6UhYVym8/v
1veTTzvIKA+OXJFUEk0PM/oUv8uB7pq98l5s5JsmIekkii70Bnyo8ix6IhtXCUgIppqnzmilaOem
VsXCULGVC2O+9O1c1dIOBb7R+oxFq9rcFoQEZmLzWAI+zhoKgJjgDd0CRgQBDqAeikhjf3+bOAGH
/xLbWEpUhbFRd1wwC7XU0w4+HPEE/BjcqTMhhIB3cGLTwYO/061oUuJZ7Bj/kF/JSr6kEulUPv3O
1gLgeqn9vQAXDlnB3slx021p9JFaJ44/yNf3s3ioGoLUdo/NCW9+UUUlLx5sJA+8GRHKsiOAXu7N
9Xf9oj9PVopP1rKohDUequHrL6an+A74+aQtn8WOntjL/llzRt8SoIX/c3l+HsS9xyU6xCyiMwzG
WePSP7ctt1C6Podwb39B0qkyBx5BWuYo9YLAro5jlUv4Mjv1n9es3dqIs1ApzVuqzQhsK63GjHhL
ND5ZyzZ5fPJvEUq+r443nbfC9cBYXCAlRl1MZng5DYgZx5e5fvoYWOo++44VAwxIBNvMlLRaMCEM
5oDkMcKFIKdJr8YIDLmzp1+bf2GdOPT+G6REtC0a8GOWzB7/6Cnhq07e5IvWCtv7MMIX623QxFqk
CQ6nhbTgUq1sjmnVVfJzmdHOatTUkdWJBcQzIre8lKsOFwMJarmXPZSJ/c9DWCb2n52qPGG9qzfR
M6kof7Tu6/CFexq9ZCQ+qJkEuQjHY9umLoef4WaK1vPHyp7jrBU3fSYe5Gxt63FAWZExG30pqkKg
xcRpiCkiMqMaGULts7h+Eoo+mKaRBds2dJPuke3VEVJ8+8J/mCwvga2igSqc2h4Xa0seSjATYJne
iTs+lWgAhs5mrXZ0HK6L51fXFqewaTzplSLY8N6GIU0Ml/e6/P8NWjaJ8TaVFYslE5SBMVPnCth7
NYF1PIRZQdnK23iM170tyKax+zY60m0Mz4L4x+CBmUHHXK1ohbDFVz8YxdusWzEWp996ZhNwiO99
EebqF8wNGfaruFQF+glZmrSxrS3gm00umqi9qo7BwIXZL+o/iACAbSsfEidybCPyhyN2DG5oBKOX
DvjQwBeCsvly7O8HeHP0Owqap7ta6OAXTfsLiB25A8xh2pmMHtgTRtoSsW1wkBojZvrbH5BJmRr1
w8FH2yDZN1yFfu+s9dFZRzEGLh5B0nuq23e7suBhGmCGvmALQYQ/Ng6BELNLSEfPmpyOSIKOopID
48gpjTMhz5ctsJaXUWv6arorX9EY3PkRul2qSGbsWGmNU3yxjodB49QqB5g53aUtwA2fhj5smqg9
D8/1HzXVIdIwWpjqDltGn5N2W9uLx9qh10GvbvvU0cbU7ijyfmvOvXh7MFkY1bAO0H/KRqQRmR82
e+weMOuI8DGZ9Iaj7WgGDrZK+PNUXrUHzGiAADwZSS7iPvEgZInntIyVaX/EnvB7/X1wlNjZ2eS/
2o73V/hfhy0NG0TFd2R2bkD2gXDadyQAvEjOQeR3wvm2sEuUKIaR5k4WX4bcVfLcP5rvJwpDI9Zz
rzkr8ecRHc1eBrcXoLY2P8m3pc/rT3TCKj5wuOQVC0WbdrGlgxCjUXmdKFGhFjT+w0hqOBZg/jdb
vChAywidvJSlmBb258rF9OvH9NL0vBEnnxdncqKWDaDgDfyS6+JUEbOoJXuWNh3LQv6oK0NaVWqL
ICU1lR14ZO2EjPx6t8WXCozvAjnNdFhdrFLd4B8W66U5ud8JEdsIO9+/11szLojv1k7ou0OOMsyY
AFn8J4NqILXeuUq/wyIvuCVskCl7IeN4K3XMm1z6Yl1RKemhWPMLzjA3dZIiKlukaxaKR1FC9Ii4
xjCBM0reowv9TcOTDMulYD2Jh1LvPXgjSBBYIyJsAKi4y/vrYZktvo+dxVCzy/e4v9NL2xNfAJnV
fLHNN0QYOzm2vnrytn4hry0V1KAbO5Nr/oZKwSVN5zNffpgEaMwokBF9oLKOv2Q9RnZmtFD1RXUm
2mtAqCoH9DEmbbtb6gBMOnSqoFndsUGsLY0vi1WR+Hbm6Wl+iUcC3q5fB/iU8PcA2du3ftSiW7rA
CAJSm1zJbyxaYGXj2fhn/tzx8soOCyGplAlo5c0FlWAFddOJW6RfATKKNeIAP+Ce/bgSajLSSjG3
cLxdwavVsK/ulljRI57wC03gFUHEJX1ocm5OzmLmPqHExcUk5fqiE1SohSd8UWtjpS7S5UKYFlAH
BWsjRpDL+XyBaOctJUejgY0b9ccN37b7Mn6yOjoJVP+UGcDNT66SfPwOC0ZGBm16PTJIFxjtYTDP
aw7j5xpNGzmQecfkdhIkXG8zbS0pMna67yetn4SgmBTIqFcySDMI0thsg6nGX8K/QOvma5sdgrIS
W3YozaN0Sw9qRvxdq07aQSw1yq5AZujXd7v/y9b6J9TDfhexHQ4vKa1cs3SzdD82G+Bsb8G8MrgV
bTu1N/BGH8BCOGwxRsnmqIU10W+bT5ElK2xKdTvm6NOqVaDaFgix36ww/snzzsceYl6rBP4dASEp
qMibpVvkrQ+/l3HYaaUwK0GdSuDTL0Dwuyna/NOwk8QAd55MQSC/KWpDSociSC8UarPCrO2r7Bw7
ddeo92CA2XTrpsROh1p0jNmtyKav1mlnqcr4Q8ETnHETTw1UztfB8i+sDzqRofdacWlKkJfFRUQ3
fWIPj9SwZMIOyCF1G3eEn9Id+7K+N1bJVBbSnInp61NXlV6fPdab3NzSvAHDWd6fuVUwU4mx2zKY
lX/jVmJe7O00EE84eQs/ABGz35pqWuZO5dzbnHNuaUunIOsChkCSu6KC4wcF3e66c/YXl138ZLHz
ZCpW1QXMU0eNhdh1rjJiJhDR66KWPeCG2/B/WTvHmcHSGjE40V+YIpn3/wmFOt07Oux+1ISItrx1
mrfDEvo0FT2cxQeu+sAFLWQaxYKUQDdObr8BkRpMe7WlS8ytjcUWnHj6LNAwxzn+gvom1U3uV+yB
R9SWZ3BPM+ZCv5Mdre9sdQTOIaTm3amYsJrpRu67hXNCsvjMCIv/OpAVVXH3nG0cl9uLvpdtWwWg
UwnjV2ApNOgl82dUywFwhIsbgNBfyrVUWwn4ShF3u6B8SnclpHFZm/3uwuIFcsEesTnD19WicFrw
NvohpJbzZ7DV+INUwcH+1y7EoWm2WRjnEai8JZnmRiERuiU4ovtnUs+EThaGkipaxA4N4vCM/8Uo
489W3q0NJXsD2RLYB4YlabAEeY5ufFj7gsRjAcSe2UrUfFPp7z8SiIFS19CehheuYntw0Y+CY6eO
90GNYbqhwtzUDDDrbDotuVpwGTMLDRJePmIrbwv7VEDU2JW1rDRUScOTxV8x4tbgOaNlYMEcy8hD
CVtq7CZkFIz8T4VkbH+fuiAf5wrODutFH6E2qTWNvgb730Tcb9+8GlNQkAtBT//yQqAA6Syk7AyS
+UxHO0eAYN8xJHUTGXghv4n3iKe+l9ULEoSTwdaAn8ogO1U2lzUR58JXBCCLJsA9gWgtvbW3ecG3
XJgqm77AMlksPblxeymAOdvAQ91O/WAyRgIthC4hg66rtbQmHl4KWpqU30iF6VYLGEfqs8le0omt
0nX1u+igwPI4Ax/BU5plfoOnjI6IyR6k8cCCqP/m0lrS8CW6ZNAyv7ew4G+DJJ4Do5xPBQRPeUur
RefgrIOUmiaxzt9tTaptzPvu8Tmr5CbGlyYo0WuT/6ypQe/m5lBybZK8Lra3MHd1OshxNZsqPaLU
mq8YcDl18+ESG8pCl2LbjcVhpm8fsxJII/MhjyS6WUfh+1ZSVZxuD6M3ShDP9r8+JFWgzVyy4i84
l2BXqO+GNCeH2T6AotTwGCcJ3jUqmEFgvmdvzbbEt3Gb+xt1k905I+I3AGelQ1UtG5nWKy+SCSzh
07yIasP9Mb3RGy4gMVfprgDQvvRK6ktINMz4wEQvVEWMhWa1XG82CgWtgFqULTojb8cPnbMlRwT9
CLRzVMgO5MDbMjQ/NO5EsEy7clMIUs5jGS7DuhHBo9VAazGHVdvM7cuKfvh88WMDt0zxFgJExzoA
mfmhQI/UPnvvuiH8UprCujvWhjkE7ISye6JicX0epRx90ZjCRsIk8i3Imch3TxVYpx2XlK/WUYJ0
XXJ5rot4NIYzPb8/RVtTnnTYCheOwRVigwXPrFTDSsdejhHK2sxCwTV/a3fyVxETQZWAJkYJwHZQ
wLgLzFgOBRyqizzgsZVs2KItCTbHCzy6FC/tnQG9fbRZ9lGrqR5ZHkYBkILKuoAG+o4xtAhi/bJb
GwdhJVhT1KK1z+5tXwp7w3LDkFEc92WZJHiDUOfGL1/8dxayc1jloJFGwfcA4JYXJxMKF8p0TgCA
xbZBItBmOmFGiX5n5iXo/7pWGeiJOg8T8KOnShJo6hfnSiZtYTaBu5WJxpVYvCKnW26wdQ0GE0pR
mJrJA4pJU9Tkmxqu85wVBZspj/G4wrCgIagAgvoMk2laYqwIoB9eFYMdJXCKllv7jvCWOLBvKXiR
GaGP8ILnS/qQAJoB1TyAO011Kt84zONUwTYFHXE3bStETZbxiz2oEw72dkXSYUyTocWB+sO9PntH
D73sVAnj715bSX2w0f0juOXaZpM1xdfCCYCNF64XpSQ/eROjxc03bRMHYZ/Z2KezIhDXb0MFhMtS
G1dK0zUA897gMEGYR6/W+feqL1oofJhgZj+PnBQmgmslePVeSv9pmgoBUTew8Sog8w6ynVZYuR+y
1YuePpOXiVUapr7OJT1NhWlhOE84DDPlw+oDN99Pe92xt4iB7lgSNkcR0DKlOZG9CoW9NI0jBE+X
PHg98oHrVvfuXBWZNCT2Sw+jayLfYivSG8qAVku1gchqOJufE/ZJ+e0yiO7/NuEd0CWzqXoHqJYF
8uk7ARL8xHvxSdE0MVAoyYeSNKy4lc6hLTL73t9q4dk4MPlnx1y4yzuOA+vYTbtUW7lmYcmFsfyG
ec2gW3pKqAs7umVGEOJiTOm6/q07yK4zFnNaqFeJpStXLtWFB2fLcZm/aN1anl7qHeBKHgMSHQ9R
gCNVxm5z91n1+l+FjcULRuzmS1C3wXkP5quQOXdDT9Yk+8ppbt6aA3tRlMo682CvI9oeUmnPj+FC
W7oZnus7wI1ImgksXIlP9RA9ip0bitXi2+gyVYsab5+dkfDhfCxquOz+6IJ0Et9lNXI7mLhZ6rvR
eJGw7Nsf9yuZvM+OLQOHwTAUCCMSoDJ35ZNQZFBmBcoChDqUvgmUcS/TAx9fJq2tA1FgdYNvGi+e
wNVJNNcEy4Hlvbgs0wvmAfRUVlAQ9I7WH3aovpHDVyM+ujo3jsr3UCFIhgeZV8YmSeMfzcN1/do+
PvbJw8Gk5XH7h7u/eS2J/k7ohxhYBWIk+cCHmTwTrOUVjVFYp5ZFNsbbEd2Q3Tl06MtSKqJ0xMdB
xBs1rxz704tKu4MXUkiQq8KfnDuKKjYHdRY8F4+YwftqTxhvXTM5iz4QQdKSzoymcbmsfSDp32Ow
dllnl/Yybrxe9BuK8X955ccf2t+4yg1EG2kTXGiXtDCWOyzinKiqgldSIlEYF6Rve2RHai/5KMQY
p0EuCDIpDR/oWfXxZBXAWz384ifsAoV5u/zpvSaq0vqW/F8zlfKiL3VJFHdbJX+zv2QtGXYbT8sr
+TX0m+p/RAPNgESi/65urnZdlGIoXDaNWKaiZIt+gOusNPNBMGValvQwhv9YXPtO32YCz/TLXlj0
ZnFBIKtRXkGm/J6R/Q/J/gEm+vsK+nWmKfLaqiWNZX6c1s7SVO7vcr0+4dc4sliyvXDbZk8n47uy
20nxlaSrdobfUCSxnkZLDVVLkevkdbzHkkgb0ZcXRRgM69YkTZNscMRWaQuKUV5/DDYnk9qGdjSl
ly8/WkfFwCdsqMg9bDrUl0Abo0ZvrCcvsYI7skdqeWtx6N2ZeEdg4w2RQuiqHNUlBGiA695tPBls
5OdnnNpGESH8RIVe8Ol7Yr1FMM0B3I+s+6LPjf3sjP6Sm7i8VD6xVd6DBIhN7qDotUiBONZ+FRaz
O5/YNU6+uxTWei63DFKkZFxUxN/VcCzYYfrPe0TeEnI3zMvewaLPqK0yi3gp4ZTQZin68WfsIXLV
Bj7i6qzZyeMnxNCdHw6Fbk+0xj47OgiM6raYTHKlsGvEFEPi/ghqmDa1kAL2f9ldubbOjPFtuPu2
e94USlB3qpxF9la9vrJ7CIdE6ekFVlbRAboPvdF2F5ws2jdLJvvlOOs8mKIYhdEzYIpP6zOSiJgu
R+lNeDfQl0u+bjCvAY4Bc660RFjYYT9xGVKRPStyBgK+I1WI7otNaapRgfXLW2usoRUGEHiUCthj
q87JqTxNxGVo6Ht+JE1u8+8fLaP+fzy0TJXoR7Dem/G+mp76sMRW8LYKOpR3oEP7nW4iiyYeKqBW
NKPggK8upHny2P3MOHFOC8Dg4sblAc8tVOMZfzvwaY3lbbmX31aQBhu3bzr9XaNvhQZF5wz5BeBk
S97v9B9GuNMfpU9iDeBo5OWxArU//UdUGHEHx067f+IzSSr9CgBN1BjjvQ+uEGnLSBPcYYzLJ1ox
TQLpPUvq9228tpbP6KcOJvkTF4vyjpiOMpUDr1KCuXO0fuq4lU8TMJqEhHxPTMAtpG8wb2FDJGKn
oEPLq5czxo8UAqOAFjT28blCMX9VqVb1F1aAY/kXHBMbFSXpH4ILiWvr++0sfDUA9NiKVW8TJJCo
TJ86n0oUdZmy6xD2Mi5XDvjVwPJUHAwYIw6q0rcjPc3stW280n8M0Cp/tdC+M5ayNrXhYgVE7EKU
V2fOKMnmgvLAlU56VufcU+n1HJ2ggbRw1Ak0lSrhNXeqMDc9JV8oXFSz5XCgE5ew0UOupOgT01+D
f5wAvm9qdPiYFfFSwIW+NpSZOJftcRi2UPhSLEYEGBkkBVQoH4HjxMzrInbM0fR4iIFGCN6m0T+W
OObE1xbTBdrM8pE3RebYzsiMU47beQUmllS+CXbCQOAyIMrpO5VedY7U+kEtObNsqruCiYj5RsYk
XbBewOZdn/Eh+OEysJottwfXL14T9scgSgnwHgsMt1gGa9t3lfSRCku7s0NZmsJ34CSqVlKASrPA
tGRgHSX9m5ErLQiLg8YHmGVhovBCB+9H4+ElNryqcKKucv/Vle1T/emgne1dYXWKHQpfnwtkxqfy
StbvqWK8cgvuRFLBDisfPuRxSLyoaq+LyT4zk/aXchfr6Kt0h9jz3CogU3Jid/aahg5M64K43vwM
1aCQ/bxfX7gc7mD/Wsbq9sScdidYpTWymf9NtnWbdf2ZWAQmR/0r9RyGejeLOtehJdwM7uSw/LsT
xb69ujitccsVINCVq0hKAhLAdXIuMW4Z6ytfzjgYbocEfrIq5o7Ua9cstVhuuWgPzQF1h8O8untI
CnWR56uLI08Q4O4IRKxhefDj8+Ska6pb6/vO97jC3Vp9hwyLSBL2n74hD6h46IADRy4e7TqkKHF/
JrZvzln6ukCMVL/qUexK3ikNvw8Dyk9DDE1zbGCzO4O+SkEEIFIT7u6VDUvJkGwWkdd0b+OFoBjp
yQe9Y3n78PzDi4ET312E6RQVTDROvfCXh8coqoXseZmLVp4T4JbY4sz6jS0m7NQ6qlZ0Tg68fT0Z
0Epz98ot5lQl/brXkRIxbpadeYpUNyxnyQ25uniuZUBIoCGUHcHODdPDYKMNTErRul+vZk8da3d1
U0RIgNZAIHjZhOWwELpZyVqeGfTDGH7NacnIgSw+TBwBiUy2xsXnyW8DR6vpEIjIuD/7/IEkmAON
kyPXZ9qEe+ZkjJODzLNxdwU5GjJopmP8Mnfzi29vNegKNaeYXGZ+dP6k9USluyVSe+Eu193y77oP
wrFcXdkm6nwAM5B5SZKlF+sPvdyI66YGfB4qx0nn1muu7ncTC8MEsYo2VLToxMcFW8Xneq07ig/d
dVPrBno/E7mF5s5mVfMqyNgqjulsM658jeNIUgpmJcmNQun53wCrNaye5bjAof664K5TiB8v9u/P
x0u5XplclaY3y0+etHDOpD1cEdQm9T6tCiVV6rC1KVulp39wND6drKhess5ZZtMgijGG40wh3Yqh
p2ebUz7uKwvZX4CDI7Rfcone1VFrtXf2vT152mR6PnB5AOB0rknv/R4zoCVHSsW8ODwzFJbahXA0
RkuYbwErpMgc+kEHyWLOfbtl0P3ODkv22x7qFuL9uNA0ympueWLexKJtvWzv9/fxzhtyN7D214ty
xUxqAn2c5FWbLd+2tJ3BDM2ZNpOorbvISZ69SGZojYzawAk8HKXyTvp14vqb3tkA4S2MUp9vOSuP
Lvs93XuDSUHg3DrYk0F41lCsNRYk+7uiKK3/4AbEzg7hctqKmQ1AnGU0CYtPdlbxwXViDzw6v/Ah
JbwNPX5jLYadNKF17cAS8xn6T7L/uY7r6439zP3wMNuaNKQbZQ/lfLZMJB+PgOoknJb7bCHWvuwY
gk5doHSMryFl32n/xnYx5AQeHGb/D92Yp1ljwzfqyk8nRDp+3ynWJg0A5LbpqTUVCzANGJ/UcyrN
c9kOlTPcKnW8C6Wb8DOJXXtK6Yl/htdGT7kLCOiQ0brj9UR4IUQgctcxybjFz+aBb6tWq03Y7Htm
jKkMaB9L9P+m41tgsLJTtWXh1vXcR1C1OXDqOfIMfPClPGIHMRNV8oqgT+qXLiiKvu+GIX3Bt5GL
ApSXPqK9EujJFLf43oUan5b2KWUDjapijebDAZbhWrLxaI9hzrNs97Rf1sSy2BZ7nd+EB9Pw13OZ
jOHJJHGjcDWBTYUuOUeGXZHPUMMuVMDomPn4XW+7o+Rp9EROHGpTC7KO8ywnktNjfYIFjVhtWQFd
haScRjE31pLyprgWKN4A/n2k0GjYmeyuB/TXE7n66/mVfuYP4J+kTAUrngk+JnvGud5c/LE8X/LU
EZO70+CWWHAyZiZtjgKw+Rch40Qto2nruC4IiUSXyJyuvgJ/PfeMbLl/ZlEs0scw5mLGMEf9frA5
egVm95CYZfBxYQRBW1uJQj5wuLpfvYdf0EGMPR+QFzg8c0LYAxz8LY4KuIHqCkDY8/cgjtNTuxPJ
n9YPJo3ddUgmjGsQS4IFqdr502KgL/h3+oV+oHicaw3musJFJ9+HD7oxInLbUjeL6eulkTGnVuqr
O7aJDlwQRB0MzKU9w3e0g4MHAC6fXLd31xCtvVhTuQ1z0Z/Uctv52E7rTWMqAPdRjscXYHrY52qH
1Ln2GJx/fv+TyiHQHTtL5MS+9fXN3Pt8Xpmt8NvVKo7S4R4BPqDn6HE+3Im1JdRjrl4JAkS9BESr
SNUYZTTk+JHXuZM+zUos2jMq6VzKJhdZsAJFrYSrtlCvC3fhlgY8llrf+Z3g+A5CtGbQ8379Il2R
NnbnaDXzHTR00VMa9g19yAvUvwNUUGbshzcdKJCTP9M+LKMkO2nZJKag1CiSSyUkc6A3ennaYiPc
aXWJGPFozCKAImhuQ3rQ38TJxfdRzwkOjGxS1/EVu0vCb+98gjNuMlzQmOIVAnL0mU+vO2LtJTS9
SKcfNV9+GRwV/cF+z6ALAiZkguTbV+RJBK5hw6eMepHy5RqmbIfmz9v9aQ7Pi1FnUjffl1AuYEFa
SAWkRoPPiwKpA4I/XzzSD36oglJx8kCbeHIyRL3Xpv/WPLk6a4c6Ksfounc8kTzGaMHdC12TenFh
o+fOzzi/ad8ltgVky5R7fpUfE9UyFGG1/PcLA9OLW4Ligcv20wkWA7JDm5xO0FG28kBY6sDMEmtn
Ruz+9JFSKoDhOBF+6mrkazhoZSQrBodsS8n2VWSV0bLVonhCWaV1CFNbiKKotA9h3eLlCZA/MHcf
6e5GWoChXbP82K8R4+WJx1NlBUnGFKHRNEPs/c8VPZNWDdnq2pwru5a56dM4ezDcGzYCH9ZsTHrg
uJDVzZxqT0UcbPFpV+oMlMOUl92LxSwu/MXFLZz1bp0ZUXM4fik1Pb7EH10MDqUkc6gMoI/S4dRZ
BuC/yQb79Y7bBDt1pvg90ljIObPt9zr/bmKYdHyrD6PXlWRHsOEFTlcdHecrHwy2HNedNG8E9KB0
MYR6NjC9gZ+wUbPfdVnhDRIUvilIFBvEEgSog6TTfp+obsz8ztfNSS2c3U/PQjCVZ0BM5p851aZM
WqSnqRYiRPaXbf433/cMgdXFTFIGQc5puijpXP/Rdh1JjpDOBA2AnVm///7JJ6dcmkO3ouwXFldg
xf3GIO6Vk5HuolmjY8RsJSHpScgKaebmGRbBgOowQgsFdHtfKKwLBZVoVzdRXonnXmWFyQ+gXSln
bMbY6mhZ2fplF+YI8scXu0YmIRNA8EMzAKC0wBMPkoZW58WGldnWUy08ha9G9nKl8Wlr8zKn0ELP
o06EtRR8pV+TPeK1/rU/Q4wLR3odKNG7eDgZwbJA61zX/XW11xONGpzFMv6CkCHgO8Cmwz0ri+2D
Eey67LXhkk2r4FJpnTpGWbW90G1eqwZ1r6Ix+U1ZJ4WUcFibWYFI6bSEbTfb/rmQIkQq7x4cwzpb
GhJJk7LSd1HUNg/uzzvqy8xT2cbwHOTKNb8ltI5F64RuB/O1xLLDj9Mk9Hhw8x+2oCuF+E0nsiTP
NCAyIFwAd7N5wAq2rx+M6DSV4lJrtRu620elWeHN7iG/J1+5xZYlGaZyJHp/t++KCqiI9/hsKjOD
nuqJJLzGLWHznONMPJLeEcZ+u4z9b2LsWVlj3m63DmsRPpgJczFb7rjYsp3SNQVJ5Ujcjmv00FbJ
mIOItJXE+ARzI/XT7pgleil+sAm2gGwIZrb28oreqwF2ulPwp7PefGdupGSrWLilboff5XbI46Cj
aaTbpZGPmrhAApx9kr0JT2E4qRXU7cMM27SzMyz0nAKzoDatDuVO+n/0DoFax+snEZTGBgHfMS7w
NEaFqwMCBuaATMu/jFZ7EcDDKRTSKioGDlRYoSRAvHv4XJB3cMkoHmrxlxyVHAOj6GY+No3hzZlk
MPxhkxLoiU279aiwWNyYwDpmaUop70PxYxWwIzwhr5i3sJpSTkx4qWg8d2PWTg+Vt+5MMakOzLf9
E0oqIhDYwEkPrSyTSWYj+Sx6Rg4FFkRi8JeDhx3ja0E/msRj7G0jhinlnnkZ/M6Gcv0rZxBt6yDl
Uj6JoqHKUhd443o6/DzBTvOxnh9a4b7y/ZZLK/ih6nTdLNP0LPMKuLshBjppWPSfmwSrHCCvZr5Z
0HMvMtb99FI+htDqPKUxdATIzdiBOfBXdhOAEvlRH4YIxMfO4zTpmzaw/y6Pd8rTcDpun/veiyNh
44VQnmFa16DAG6HZvYP3VMr2Y5OzQerUJzbN9VP7jJY5cqgOcC+9sbMjmMNLfrWJCxK/177wFAmh
U1FZY/HXan0v8ly2sGo6VrvtF/qfyZSC4WLcn/L4I/ntH45GW5ck53XoE9Mu2gIdQts64m6gV05w
T1d2aPjpoYSkCUvpEIBil7QVKgyjgUq5U/CKOryTPwiW3pnuGCVa1mUThbjKQpRdfcWUhrmJLihZ
JRwMJuEbvscLr8ZkOFCooK+JAFqtWOzPm3+nrpRpiqBjl67MWKScQ9NBouo0o3erQmxLbjlf476K
qJvjNoPOQjXRTJfj3ZPtB9OiLVv+xpqBhasO6vYJn01l//4/dxBmnBDtQ75JSGDLmLIUim/s4MDN
ZC+l35GuC432M3jjRUm3XZe/qDihs5bqRndJNVCIzfUSybTPc2Zsss31X2fR57d8dJ9jCgMGpIRy
XrSFoQccNLFtXApdIibMJRp3ToNB/6ETXW29+GU6KpjnfoH7eI8rX3Wn8q03Zj4sg7iABI93d7nh
q7CwS6WCsmIPSwC5tW4dXbazs7cuj0x13YNdz6U0g3Euv7LBZ807sCyRuTWk4GWVHC8vs9VRdtuP
YP1deKItfDSrMvHHUm3le+Yz/+xPMmvEAeR2XXimaMwGLHxsqBJA4cKuyS/AB94+T5mChhD7ovHn
yyKuzkhXuG5s644HoyeF3+xLFsbFlUoRorj+5BHVdN/eUQxFyeG5bNyXvPTStB8O6PKGKh74p7Ue
stQW1VRwUTkTLvugAStXfPHy3ohoBaFNMInFfcUI8Y3g5qIi960ltYxqGwFl1UXTHMwSPOtBwSxq
iwOTrAHRI1RM2ho4nImJ4tllTspwaGa3n7beFdpT4WWBQRSnW6oVQ63uNBVA/G/M7xi9bo+LZoxr
p1J3RvtkoixCkSuFr+QpM4nDu3P2yMaMJfJCYaEWBY0GHFGYedPyzlKJOk77V4H1OaEpD1XrgBmu
Wr3hXTs4ICdhbNyKbBp0HV2INB3guRIzslX7MJWiL0QfEFdaoxaPh38oVGaf+RMkCPMVnkrQAOQa
i0HWKKY3etEsrF2bMZfazghy0FM7ucOWmr3R4z+hAkt9d+tO/kl/MmraM3z77musEs7cCOGDw+Tg
9kgYxei38O454fX5pN8q6nYUllEhfBGLgUnjQ6IZYWG9A3V9iHOiKMam3QSelppEkhdexAwZ7v/9
zCsxob4Xq7S8yyz38OuSBsgopidn+Nd2ddl2IWgAZ/9tP3SVIBsyJUH046hC1Fq+R673XDYe4sWd
Wtg1NM1p08fuhg+yPlrJJIX6a7DSLOhqmTnbVK4kwyzi3eCF1Qj8OFjF3/iDwXxyNpdvj713dBeJ
fMIpj/2a2N2DagSeSxRbqBdNj59/W1XdEZ6wx5ujocVFNBr5VYvlMaAkpR6D+RlhnFOM475JRHWz
LCuZPxd3RF0Z2NFXCZaUE6mI/YVQi+mYCDmt+I5wXE/TbCRPfo8Tt8lURVmSGavOSLSo/OVALNlp
zITFozk6IMwa67bOQdtEO8O5o+iD6fUjOo1csoZkhdIl/TGBW5TbZLZJJyNrcRNl9AFl1SSylVOZ
1zQ2B5i0IoIxsaSqFK6uz5GAz3U1YqYZLNDrRa6KFAXmPanBBwHFE8E9119veJnrmeYEGDQPrtjB
29rrsD0mpUym7rTr7zJz1n0VAwHwcCEDo1k23TrelduXUJ/GyDYwMUIqhETNAGk/5nRkJUYeMD5Y
qeoYYinSlNaqB0cEicL4fboJYS8wXMCauFGiLzAtcFouHdxMvcdqXI45nymDu/VcR7PhIcfqOqKo
BNfkH+JhUIyyUvRIwfZgrqLBRoTA2lBrxHbnM4/hJ4lT4fHHIKjJYPTR/3iPMrgCCPcybJ+/tFd/
MDlFYA2tIqCHi2Ko8V7fgedTs/CkWRdx26vCMMgLZfjtCPS9zke/rzRIMP+MEGM/xzqawmMjIzVQ
Eh+bfPbkiDC5UFSlEHvaL+8Zub/UPipp8ZTZUhZadc4n4lYdPQUE7Nfu7wCOOUS+RirYn3GQcV3u
ztZSd5IhxeRz0VFcfKXYHhUoJU7XD1qgSM0DlFYHiGWyRNbXa25Ci5t7hBKl3X8hqpEjkf0iM7Kn
IAk47YUYavxJbSwoRt6YP4etuZUz9LR/QfGnMpewvr7PweJqyCApGptC4p6LDMJqpABYDGn+0NiV
2plNKoKL7zmFF4ppc5dO4YLZ8pYDmVBJaq2I4c/NIuZVE0eOjmTB7dIzPCMKjH6vtO9yYieoDkrl
fxlQclpTBiO1iOq98vMi2yGWx6CXOcwwJY7Oq+0CbuSLV9RajDAEEsc5fg2tsAuPYWn9H93pzRr2
xzyn/RweGjyEeW4wiWw2PxUf9Waft4QxfH9JeaOrIRsqxj4C4Zy179Z+POm2UIfwnYNJ1xkK3x9b
LgRUEjiMwkUGVBjF51R5v66keKHD8C83+yOfb8uXg5erLnv2mvva6taRvD8IaiWmeGgZg3QKnt2Z
1ln12Zn+/g0fSMBHIaB0W0jK/ox4IM+cIrf+wZHVZ03iNexttNZ9FwW43ulAm02N9/cyUY13uBaY
Bgw0Xhixq+CDLtD19OXMWyMO1GQE5TJYkz3dv5XfSOchd2JK/irE4Muen9DpwCy2zyo3UJHw38SF
ef4iECzzhz/FmO3EyuzfNSpPnsTwCnfeTWDarD17mfalXpTeCyFHG51nQzBjsGTtR4XckqFPHcEg
2hJrEbkElvJQJyZjdy0wkyz5Er6UCGFg55fj/xEpFksf05JZLdvpyEjNUb/va0BZC6EHmZfgLE5g
M8xPvIJYDh+WufA6LdOY3K//oY/4RmEdcEjoppXigS3f3lkO3qvBqnXytxOOVGMhc7uHThypRg90
kESZCdS5mk2Mm8u8DiZWEzzvBWBpoZcbRCMrGJ8Iv0ywpNnnpP5eUJlAx+7UIz77TbbTw+rcGQ2F
/miFTLI0QwsUbVsVtTuG2myLaKbRywFqtXa7frf2Ylmd+ID+xarOHJI4YtyE4JqGRKKFXCUoINb3
I0xAjCJZ62hKWn+V8+3SNRzwx7+FeSTQiLvGHaJfm1g5ulLNdOhwoRQw2nWp2opJ8qcjtg7o4czD
iWh1959He9pTI5i1Ju6H6W7XAofSVPoTANk1qFnLYR2c4qiFaJni7y8EjRNAHX+uTndeBh5+h0jo
dYpMuSGL9V4SAr/KwS4C4xRMSEelWIsXQgvZaJPZ2dF8EHH8JXSaefnmDY/Qw64k9bdJXNkyzvNh
sM8GRldug+f5UxrJE8i6DIues69QKgIMDkqbtsHaSfvUEeBdZtg+g2K3dmeyeeEO2c2KMNoubps3
T5X/65IZtR3/LnTkscR1go7KMfhZiuq4BTzhYTwDEmfBWUKw3+hUSV7MjHvMTPPiHekZSi6f7RPs
9dU/KG51aPyqYhs4rw5XoqBSvZQd5aJi1w+KdyAx4VfAaens1M+K0+jHVeRRAErtwiwNBC9i+DtJ
5jh8c6YAHJ14/oI4HnTpFypW/qdRtepjE7XGnm4X0yNO+K9QbeWsoaFDrGJZueurtFjZVnzlCx9h
m25HMP3VXKhadg2spgemdJQtzNZtpPppfXGnjxlgNG80YDnp0eoX2271RQSW+fAmLh4vvZ3wGVwl
cMhOisSvvWgLmEShCocP9cOgu6r7mXJHXg5UL+8hCD509+m3C4aQZUEqo1d5Z9ZzRGFI2//Qvsr2
XGlksUNEkgiKld011NZEhT/uUXOsysme8AcelAFCZTs5/ZwGgjY8G8Ow6YO2BVMOFRFHy24T+nb5
K9nT5is6LrSHtK0Abw37KUNSle8Aauhvvv8vmnS+81Eo7DCTx/4kLKKd3Fl+wKDU7ZsyCgZ3nqXJ
g9ThZWpXpdniYVdfJ0sEG2hEOrvuVlrkuTIt1MaefEDPdN82UUq6oJbHeuMzdZ4haiQ+ltGfbw0h
c8Jc/oZrBvL1GACJvLhPjZ/FllHcQfW3CGtlrRNJayifHML9mfYl9LSO9JPtxWdBoOLNoSQRYk/M
+TWK+QcSGQ1cxF+Qk6tKtKLaw7ofOv7QTwi1TsYHEOkPnlrEHDLqBeMWVeALPbyMtlJpiBTgDl8S
yUuLjViKqbe7Km11dit+Tnrd0ubDWEzN3XCPX7iRyc26ruL79dJjr5iTZctQfB9r3Suk/Wqk/yIN
D7fTzY5X4LzcE2DSpNbsCNRxUQhzYG+mdtkOBUsbUzGLSsyH/KQJURMwcc1JATtlKhSD+Bn+QoC4
bo766lQh5Fk6LQPXxHU08+bkwi1DAN8Q9Z4pWmhimvHd4EmPNawNjsocget1VURGhXyN5uaAT78m
IB8HXLZ4c3zrzSQHCu9dXSQuRe45/8hcnaRS1qYUfySCDh9E49nvFmQhgKf7VlSGy4zql8aTeDK7
wCxQqLNDWV792UWi//kJA5/Z56WvJQsdyWAnXMPFFNJ3OeiurZ18BBD512TMzKLMH1jBkQB1LiHY
htCiETDmhVbLyunEHFkBhNLkoish3zarWd1VvsCNNoaWwdv0qDhc/07ohK9+cpUIu9M+Wsxz8TX9
FUTxHuFlV+UGOnDvtIOHl0X3Q1DbbT1DR3eB6csLsin02GJ/U/5NzvozuYVX8QjK5zGkQQCURy0Q
irNs+EiRZCxo9p2Ljkh+Z6bQHTrlGPzAv6dLk1O5jb1IrnYRv2ctbpqr+P6puEWSWS4NlOguyLiv
f0pPJ/fWRvzfm5B0ShqE+86LqqgSLcjCjo60UY32OJpCcNvXQ+BeP+TXMDxMM9NQ2sfCkxQkeZQ0
g38wgwoFJU/sbyVyyPUWDno5JBM+/P+vneVFjKnsck/+hX6KuteqKtaL0bCLBptzH0OAuU4k0cue
VdzDjm4nEPWtH8m/Yt6dGibeIFA2iR4XEAWmqJGS3pM6guW6kz3Z1CiWjV7HR5KOnA1LSC917pvw
kk8BizdDDZb3gb+F3PE9gtuOmR5AOrEXKRwzzsHf9ed0leeSLiIkFyCf84ZzuBuoZJW1VqbVVtKh
sz4+IJcVlXDRi8C2Ujs56KjlIy85gXXuSn2IpEQRa5ARxil3Sn7kbZNetCpa/8dLlmEhTm82w2eT
yePezR8F8/xYhtDE23qCtO290x8MzIkZ28jP65iAH4d2MywRW+vPLgPOMkib6RJkgrHpcWb2Ra7S
nQT9ac10WkZGh1DJ1J/dNURdWC+AmMUpe8F+dm04d6jZSPYNVaFKPqYlXUM6ygM1fTpQZfG3QH0J
UWpqFWu0fqYc+V0i31eZmT1ykcm5gcAUpxHBEkrp1nThD01vHZkoyeiLlqyJEDd3sC0WuJdIIpL2
bvtZHL/Fjzdeq1zu1YxOAdwom4fpQZKL13H2eZN44HmBvj5kURvhlg6jEDXKDunRl8QLRCPQYuqU
M0SLqOAxqCzcHlomhcTFcv13D3zWK61vu4ysMCh5EuNbl2n3SrgpPIjPNGnRKBR0R+LRgrnEtKxy
tiGLuuqo4SVzYaRU4GVbfuQttzhdPVzEDVApbXYV8dCXWaVXdvkXuT4+7VxaCLOno4W2XDab1HPh
ukPejEmJgaY/y92+ljW/HdfQxXnfvwoX4J2f3wb+HHS9SxeMbST5xQuk6LBo9AltYmsFn6ZJI1R4
7BCWtH+Gb61dyf7Jls1U5X3yVxLUoPX4/QHAKR5NYB2br6R5Whr9e/o8BdU4ncYYHUWUMhu+LciM
k+ZpttNOUARBJq2jp5hY5m4o4hzUXJTvV3OGsBaGgLkSienTsiiNAB9Dc8o2VZiVDgsCaPR9+DVR
SugudFkz/A4Sjppb1njhPN9SDsg/8V7BnCclHz3Exr4rZoHFuAMI3AWWq0lbpv7fUTAN63Pk5buQ
9veFySlrH3etvq7oivptOPFQ2gsyK3h9PU+ou2zfMtCt7LH19dRo9/qHzbP9fqVwEn8wwNkjG2Bb
6rGXyLbGobSf45nQZ5QDqyQmONbJulMJRIoPrdyRkZg7345OHSEHPo5b5JD/9NYQv8M4adWBVDZH
TaJwOfR+RwO6Ol1wsL1UUlThZbW8xeKLtt2x+3aVxFk+3/4t1BkI2eC7Yl3QWe5tRj4j0QMoJzra
xQkZlmNMLW21eJxVrGi3eii1jy3eLfkJBeq0CwgUlq4MhiPe68mbO4MvsIwNmgbu07LuzhbO2qMH
GmO087QpUH+Dy50siwj64jAR1adyiBTLSFNGsEz2QH3RRViPbslzDwCQcHBP7nngOO7DvPCi5/om
uLXvo9GwbCzpraJHGhhrxpegmrH68vQ8MdoruYglFxjeg/hrUy6LJnJ0mqOfR/QYsxNXQ4SENEYz
fwEDXqc6WlqUiBZOxSvGaP3mO2E6sQ3Uo7Bv83KAOam9Ho5C1o0gu5RRQYAcoh1TdH2RH5ksLzPW
aDGwGopnan2tM0fwppLBDsrFP+iE4QmbSksSJCrl5lBUQRiE7wzKobtja/wcAW7KWgu6kdtHA/WA
qIj3Mx8Y+EJkNDmwTQKbyI7G9uj35uReD8TsafhnDATowArWPODCJgf8kdsPG+VYyNhoVqYPc9XL
bcyYk/BW3ina7b93Zh/LeBLZJu3ivcOeMrvM88WVWoqqEwDkINgkiK/NYHz7nrvmdBNgau07AXZC
GQgOyiRpw9Q9mpjqUCeg4co6NiUa6AVNC+1jn8lp7oT9k1h2GXNxQksu7hTbMs94+EGmVOmROFQP
y2qjAmC2eDmoadM2X75YjczGtY41hh+YRCriW1v/N99mTXF87nFHSqx73mmb84yn3SqfmwfmbuMi
CB6ROSV5+32QQQqMejDcW7u9LA3A/DLf3ABfuooPOCp07KgrPZYT5ui/co0893rWxSt9J64iv34q
6LKYslUg1yf93iiZZhLxspCixotkP7DSvw7hy7VN4l9ucbShvaPzvo5gwvEB8i6NdBuBa9OvLaLd
frY3h8VaOHzQOHtc7gBBtNUdZKrfa8bGl21B0yNkL9zUPA+QWYIckjcWkzXqd3NlIJkhPb+jx99Q
W9FF3FLtzSHGY4hIfkPlOO0OfldWorHU3qdw9KOhoXRBa+Ea6+qtx1DWjTjB1OtoSz7wSqLFpgk7
J9WlDHET9ZkjHOz+d8q1GlQS3gVTYBmWISra8B9jL3slhHJH/q84mv3LPXLqHBw9zJWcFaMIepx6
QSdOW/tZ5VgcUDE95rOk4YVTpfvkj7XSP6F78yxlC4vcFbNsYysr/5ceezg1J5KskVbji0ROJPJr
ly3ZbIU6T129/9F8XdkVSKNx5WkY9fdek69Wb0Tww8HCB+YObBM7np26MwqgGABoCFNkW5OmFpy+
EAXu+rYFNt+DaUeyQxtmmSw585ktWYdgPB5lzRlpquaeIqvJYFKE4kATrYJmD3nUho3Cv9+lozXA
Q0zWRs7UBjQekY9Gv8qSTsoyzgC0s5CYKZS4R/yaEIahUxmT8s2fPBlOVXae4zuMFfQTFe8/pyTp
6TWwDxp3ZmFTRjEAkPnNqVpTvjley4TURalq1Z9VAzDHKcQRMalIOENiJNnvb33sYGYRuzI1f/zB
8AuTa0Mzx+gXuBruh/2jAzrgZg2Uv+buHCjJxge4AINjsedDuo+4Larj75bMpfw9qI4NyezeKhx9
oRel0yg6AkNaH01EpFm4AIsQVBNt1bgArqbvHMjE1cDp1UP6JmNnyzQi3LAIjZgxkmBzznxopY2R
1lwiDY7wu/xnG5+hyEhho5lFXJgF0yl/t0r8d8nZwtAfPcPXAlIGCIry3ZqMeLy6PyVRblQl72T8
wQfDWwnXu9Ah+O8nDTd1wzDUX2FtsDVwhh/2gNmHIn1eH0CW4UKWyrwu2YuCNSXgljKm3fzHc4L6
dMSRTPqQ9W9zn4Fo3K1P/mCQPSkekvpDKDcuKlcpNbY/jeOqTfzeUjqFHZwc6hDkSfTQCN8IHxpW
kPpi7I+3PoBN0AtRFmE7GSWxN39bhg4RcnyRJKON1wuZPBxvmJe+XAlbwAzIFJ8gOivYGTBFyBEZ
kc3RQnRf8JyuNjXJV6gHMWHr2RV+EBOdZv8GH9KtWNwXLOWhLJMv2V7nUjlKpcQwZGOpUSsErLPo
O+3kr2g4rX++QbeyuYDzGWHYW3oDRLX4r9BQp3CJRkagTt51/QbNOUeJrAAhxuCC64Cnp+kwG33K
dqzO/ShrEB6bWsq667guus2GQQKrfH9P6Puxj4UHCrqlWMbvs1xZ1EjIUdaeNjLd9ipKBa+cV+al
OQufy6weBTZDQqZLMqzQW87Da3eqb3wyNH3BzRj5pO0PyJiO7U3na4UYtFAMYBhEO9tBPJh9meTA
DPIJrQ8tMmBrzrIGbiHNZSY1+//JNwmNdU6lYgnb7min736XTgP6dzRA9E+PPpsJPd+GkwDD91q7
S5scLaLZO3bxGuNYuMGjIdsssSPTdJcELsuIRNKjiWVkAUUrPPhUTph0gK2BVL2IqTmSAD/Wbg1g
FqwE3sIAXv6l87l2KQ2Iy4OYw7sAwxsc3Gc5IoVdg2BJ8r9CzQgCgHk7TMlp3ecU1oRG8ZbYoaIo
cnBD0wAE17tVLWeXEHb5uqVIAfxk2NXzGiImcy+x85YUs3RhuI5R8VhSjSH9ImCvItGb7hhKfDWx
ISIQcooLxifrXEX9lNF8CF03CNfdK642k1/qt9SV1YXPoT5w02xRJ98ozLT1Zv+wVrBfA5Y/oqOp
Y4su6XwLGzCVjfRj57OWoL6wK0KMFFBodNxqJyr3pfyINmT0upGUJt1i8H+xEm7Nkf1EmWQYhJMP
TcNEy+t8ahVuQXWddeqVGoZ9vH+YSEYd19DmY3q9E7chfB8btoVBvx6woEcrmZKvHThTKrQOOTd0
KmQ5YM+J8yr7Czv0YjGGlL28+kcQx/ZfmT2CdygG9tZDJZlUf2PjJTyCW1aAktZGoCq6VqWG4yjd
1XSrKNPWiwxLUGeQZRAowoXtcRubp7I6l3k1KqLsU8lIDKMs7ediI0qzImY8yS2Kwd7ZunNd/dfH
XY0eBADG3btwEAvkfrIA55CCsqyH7ilQIj2IeuKHZgnSuZe31pKweWEE+s4RZcNjxhtiYQ2zR7I4
ocxHbt8uk7+hh6jHPCfXAJ17sfNQnPp25vPrI/m5aOkroCiffiZDqDvLfEzrzPHgqjxXuTshfVZI
KKa2duU1IpGG+dnDaWtqdCaG9IA6ZVjkK1vnXgGQjMicqb2IDF5ljZmfsjWA1TWl6t6dapbasusV
+Gaspq7cBvBKc1Uz/tBl8fwiBhkO5jSGvu53JIqb/fViPsfTJ+V8gfa52A8bfzHnIjiHiyfj6el8
MY43gmMeYKTPy2PdfsQY2msZ0STjStsTRzSG/yvjuqS0dueL5M3zzrwY/D0tlq1RfGZjl79lX860
FJUiqUHGzzngdcd6eue/uxQV/OBrjsHzpUoEQF9K1+QfMIU5uX71FqGnHIJHrQNKffQS+ZixoIox
tHlA0Om5Kp6cbFuzI1LOKpmg87HFCbT4oS/CsjNYLpQ6ga09NT+FllI+uw0IjjoWNRHhD8xUv/gz
XuErtIQn01WfEb7cgVo5jluI7jDQp5TnI4BmKVRrAOF2sMZnTBiJqs1OXo4FaREyQC7WFSsO0fVt
nTkXWtLAwOYDwiGv8kCBLfYKhXzi22NRWiEslEtDDMV2ef2PtypYKrTHUkn4rhlLFqlZ0bGNVsi1
iWsZ5vHHH7TiWcBiQj1VjzSjjaG3hsUBci35ShLpvwE9tG+8apYIZ7dKOUMjG5tyWZ9+4hV9jmTw
JCG+ylncgOo5seIVORxCgjTsb4WOiZI6dw7+DfT1n85qJby30xFdKrj3QdhHpi6MU6qqxdEuTzJj
yOHvvEk4ck/qSdpQk5NYcNTNESq4BDtn8OpIgQfEdJE59rg8Nz2qcTw2U5wGgoo8nj6S5XagFuEK
7CyqtnygyOf86iiCX6fht9f9EBnpA8hG9Ft5Dpu16z1D0rB6p7TgYjnao+N2YqRmleOEPQE5aq2f
nlCPnyxO/EVwqLe++uVUqbi44Bv/S2TKQ6ZFvN2H1ngmh8leLvq1iPICgqoUvFPpWvZx/EoLoqA0
ZVptaQi8azs6KaOb1iDkuIUe7wYDAIj6ockT49Ioh01zmSmNEVKIO7FN8de9Lw+rDAiAa1qNX8OV
OABI5HdonjYVT4u26jGizxvXfw/0zCG5KjOhRfCuZsdwmY/9eTYoxv+2sZ32VjHpoz1rKOx1VHUS
OhtPoEnI5f4t6uYAmll7eWlVzwtJJt6J2ql0vrTCcO0isvIVk98djdd5AbgyQ7i2+oODt/IHhNdh
0N8Lgky6ZP6lCueLuSHQRIN5O8SGRf7uCjCGve2rs2sKca9EpYkwTi3FQxOwhYGgId3H1+8fJJTJ
RfCietxeq4Utg04IBrCA0ms1wfKiL2sYbCr0UghNDvAlhGGoXPZhdIj8rY8zdt57qAa1uKFp2Vh1
nvlJOOJHIB4Mu+rUzjdzyvNZQ+cx5c5E05s+0Cqu2sPrv9wGAHEJAAXCszYsD/xzcMdwSD4N+K8M
y1+nt9z/D02byROIQmCJ67RR2q43q651CuYvR6Z4DZvVc7zSAoLkXVXQ4Jet12zbShiVM32wnKoM
uoRSLJLFTnJAU/T4+M6M6cq6wiy4iIv5UHuD9pBYqVUsnfTiyzUh73u3EOcZSk1ZC3aGEw1P1jG9
Uns5QyNvTpo9HTBWIsJ3JG0RBGuCSMtTA4P2NxV6JaCphmdXKClNdVttEIEEkGgClw73/GbEBO+a
D8boIP/03ChzSxbcs/rr0VqATzve7lNGdmSYO145832MKW4XQ0n6LKks3rj/e+JJomSe4NQSXaQM
BQI7JkHTXA2PkunjIZPnrVNlpD11Kc+8ljT72BToU9QUDR191GekoeqkUU0EP8Q+g9OcxcDLfzGo
YLYfWd5omhgrAMwHz3ApiR+UoIEmKdYfDKYHdaDbfI9C2cDbuT/3NEd+96UJkplAxaLUaMOJ0AbC
UZPTLm5qgwdOYbzzk2AWvVYIiPH1l4eP8qcgpN30vZrOfBYg6oD3BKDq9njXzD8KvQxMYCCOo2+h
8itzV/Mv21NjLx/wmTerO6c4lZVdM90lILB0i05rWTxqlIZOKl2S9/CjzB0rPq077tm38vXN4P5y
5+Tm8B6I9Zpqc6jMoedY0TIlPzo39g1GWTWaJso2DQaPVxxAD++JSRQurZQ3QLbbBpBOQYgyWmRX
QfqToZzpSoNhWvYFvAR8PxSc5ivTgYtZuxdjnlcp6fYYKXMcrRDnUh6yOvJd1dqUhE/TKOwCIk6q
TRX+fczWYyoS2yacUi8724NHjw9bZjBEf/7B6PlOAHFCU6nxI+0Da2ucj8hKHHsF6VuayLMGvL/3
VugIS48rWnZpB65PTzomtsMkPiQjfmozt8JwimX98SdJMlFNEbMv1PoGtchIZoOTrhnj4HlHUOki
Et/3DW6qrnqfaGANRkGg5jzqeDunAdJxd6L6ZNWYDjz027JB9DBh18BB88yF0Vj52sGwHPiDtlJK
fGvlvblxk9hqjmOnMY30PETN5kNRTHxXigjVfBqyGIk9FhFGu2JEOEAptQJ1UtHeLc7/L7qiPI5e
iDA3xcYLb8YwbBHkY5h0SDwWSrohEsFOUE1q7bnHXYXyij3B++61pmXozflL+DX6+n+fQihwbKQ5
t2tcLULo6eeYTe4PkqeRwO24uZo9k2WCH5w5zAbjUhDmPkO8owVPOREYaHR151bxE9fwRoRnma7H
GKCwgCKMm5pC3/N0jtmZ2qX25h0sUQu19sTVCy+da0KCwksMF5OtFBO9oMvgPiRgYw6oQaEmtyYg
krTejxhiRqOYIMphjKcXYoZVRNBzGGBGyGeq0f4RdzxgSYgjRBvNkTDDHzP1mwpx9VQnpMLJrUo/
qGeUeX+NBW06lfuQFs8fiyFjkJRFHOhNhQ/H/Bnpt9xzzP2/5tJyfOq57VFXmnp3/jvcufUZE5q+
88WLthDUwikIMNpQh32hCtwqAwbeZyOHx8z9L/iPcRXJD0atPRdVRcSBU4Eia8F8rg95fzUHwsjE
A8LXnbxUA0d144VFpbix55EawJ4hqNEvJLunLigAoWRSdMsfR9Yi7lU2+NjAhLIqUZGb9KOE35L/
BBiFxZ0r25FyikztlmoiQepehdJ6MkWcvNcYF0FzEyom1HnS/GVnfdzmpEMI5EjO0rAffBh0ShUt
8/AZ899bNnyHo6uiV2FU/UKAzTJnc130TU5pboiBYuZxCdsHIjIe19g6t3XYEwccTpLNnBo3nWDe
hKhTbjW0jDXGbtUS27Sj5jYbdkuMnyG+PERXjm4nsw/vSAF53i8HN8sIRSUd3n2YWVgIVAOalHqH
qkQrha58sUdNWtbirv8GAvc8H8U84yb0wxqeHx0iFXi1HWI7aDTgD9FH+e+CzN9fRtTffp31d+tG
xPpvKSCWd/5nroBHtDP29a8/kG6nd2T2Vglm8ABmX4t85AmC69+2z1QFtErE8MsuclH95MlFZmx8
+UfzO890bZETWB+5phpUhNcU7jwROLklTP7kibehJXi7ipmhHorh7OPMo0XoW4vwgZ+fBDG90oM7
Td5AJ34VnAeP1w3qZ9RGx8HWx6pcSYu5G0sNgjgtcYOfz+ScXWfDaIJW5xvjnPoqslHYvVxyeffW
Zp32q9nqYa172+nPzujAaSfOfQdLyt/KGfvoi5pB6w1pw0KVMZ+Ma3UzTjqmXfqfZm4Xt8O27HvM
xE06KhQjjgJ2hhlne0v9HcbdeNxAYNQvREqarc6bnvc3rklxo2tFSLtBswAr3Zxgd5v8lTY8s2A/
l31kgRNd69cR0Ow2iVEW4l8PIOYOGZ+u/QkGkFiPhFiKQ87m1iBURyz18yTMrwK9jsAxR4Hv9ydg
twR462Zj26Aea7sFKuEINpWQBP3zBJ4rBz8msT7l15ciNi6gdBOLRG4xd2BFDnoweROce6wDTz3K
TBwOdp+wHIg89rw0tVlPk0ro2WEg/zNdj+tww2eLoFsfaYunnqHSAo2c/q54QWop3oMlk1ZRUro1
VoaWFieJOAuF1+Rnmlwm7utlC0hgOaqNeba89Jy5FEVUNh6B+HPsK6m54qTfFVQ9N1EdldvhA1Iz
aR1XiRRygNn2SRuuv1FU7iyMCkV3Gr1ZoYDDtwQdp+SPbaj36qQOE9eLtU2JUW2PCeP8Jn7jpRFN
qqf5hNdNHkYgz4uDsF8RB2qMs1Ikacenoe2LPTw2vSr5PbQs5ab2NXWT4gsD3WVKFCN4X2lRUQZ4
khq5071BOtSW6LtDY3GQGnuKyc4WQO94yeYg3xL3S6EIZdq5Csf1kHcUCBqDlZP3whV+kkWPyRGi
0NeYnhO4TI6B/mzaWUBfJfX5K1d+Yji9AqIJBJEmHTde8FlnKOlkDGrXkVOLcMPXOp7FSYEhSjup
KXBbd6slq9r/xv/J75a4BSN/xRkquUfv9ZGAKvaOaZQR9yD+OWnGl7EigwM8NSFFktGlLO6V6oGf
MWp3Ikk4RYIrdY1Ql5kteVcsG7tfTzzxfLlK/n26DesoabakdBBMddUJBgSjGoTzHBh7e4+7p25L
1WGnpe014KsM+DXLwD31FX2yIwM62UEEXoXyIuqjY+WvHRs4OoS964wtfxHhXvmBtr6+bd4jd9Ed
YIsEjaT4X2LzUeRrGitkmmP4CHGG+CFXkmPgtd98RwhCxCfuaDk/dBHvXxbwuKcUfOd0fNqSHify
R0beOGmYG4piXZJRlVCtQs7GwMfZtI1utvFZihS/a0CEedpBfZ1MfJR7Tg957aol/v5drQr5RtKX
epIG9klOAFNSdYNCa+93efeLMYCQ45QuruE7yfuM3Pu0ylbNGccxhiPrgnl/4srtKA9Y63ibwjCM
jnU3CBHaUCGIX+//LXB/s37duI7oD00w5OqmKp77RUACpvZQCvcHSycOeE3lOCadgp93nT13mV32
Uc4rYu5NwX8xV1ZxfZkdC3PE8atEy10xxuH8RZVRgJIoq4nhKo1m0Ey4sJou0p+iopbTgoSra78X
dVrvfEJbkUU/x1Hsm5F2A+Q+LGJrAWIh0Kr1IAdQFHFZNN9/xVLyolorSoQJEhzntPkvPicHmfYK
JcZvhqqIeFRuAIWofj1tSPmOw9GJTHY8GfrPvjG1E4cOsrb+Qur2pvM4AeW0NEZYPKkWggt85Gya
XcTu0o/InBcgNdG6eEIwWbnM8MqfqBZE7VrLaaua3BzUPjk+Rg6x/fMZkn0DV4cOdCtYROIYcBkD
PcQV/gyh5xZOxlbeFE2Up6JBhi810segi/fIjHlEvAX8+Anfbj0Qw6AAbYNn1KtODteq1fpgEB52
ID1vMq+2qtXIO6PtAWwVku/uvaQsZViFbYqiOcf/d33KZVbRB2y0udMUU9g+xjpD5jXOfDOc9Irn
kAWKl2STwKbt0RZ0AvfvUn0Yj++r62dhBUpdFRp4aGFk2dbc6SvCpW2sz0GgBYcJVaxorbauDUex
g/9ezjFlT5d52rRXZeZvq9wmZ4c+/s2JDCb4p7th8Ayu/tSROREX/QJD8A2deSTwVsdTEWoaYGnA
nDYvsMWQhPE0BNsj0QBO27PQRDr9kephoZuDw+RAo/eQNGE2BJ2RcnvH0mCZd4ru6nufXv5XRZNh
QT+La4w4LturvZx2B4bh3nsgiva1mLH5Os5XF2iFkHY/TtDi4Lo0Ie/h+OIyqmDuqgNRWUw29d7Z
kZtdiInPTDvIR8NXIAdVUNOOeslkNHOwCBdrbffqgwNVFjaGbFnXD2MvbovKkrtfM9VigSuwNMSd
TxoDYhr9QwWuqewt27fs0+OWEwiidkgc9moGKqxiNoDESGPHM+SKCbYil4nNProQ8kCxyeQnJokM
uhB/uw9UL20wJVES8ap7+eahiMVeB0onAPR34co6JT0sc/dqYMILnuBrPr0b/bWhIcNOd8FeIi1t
L99jcrdnXZB/radmkdzOUHMf9Weiu7WUKYvLK0dBisJetjRW51OhqUQuuuXuPeC/7Z4VbW22VcVS
HElBEbS+ni9Ch83qgON1clk+KXLBu9GGJtPwyRxPpPMApSpbYcyZ0DPJmRndPiDf1zpt0Yi5jfL9
ssbD2Jp/BLHo5E2x/ZUpHx9ZJHHJQm60FYhS8ssdfULW8R5TW1TkjXsEwXWv2Z04K1A+8nlpQMm7
fr3LV5B+SLuRA758nTSqnnzV1VI/0ZjbgtX7vgaBEVzjR5RgHHD00AWVMVFWkQc90jtEYHNgHMOS
b9NvYrnqSKeyysn0iiq45XHTMPXocnonxk6yATAxApRcKuQHj0I4YEbRobbJ5dkjmPsFIXBjDAiv
45V7NoU9m9Q3Hdd2dmgSXMefTg98fNaOZBX4JGeY9YJKipdjE+Gd6Rv0bnhyp2Uh3iiXD2FYQaJu
TLurXImoIBAdMnEBjaqc6QGfnVbN5xvQldWXlKt0yQyEwPUltH6dgmYYegFbuou90mvJHre3rTEO
Ww4Nqi9Idbe5uwG6JItSEBd3v0pl4Ai5oM3oiraO5AfMW9v1kGg17mcZ+T07x8jsiKj0u9E36Lc0
USe6SsoMA+kA9fQpZIVGrHtI80Np72SlGkgAa4nWHRr3yK+KsfRaf99f3zi/ftOGFvIMaWgx1jej
9tB0JqifNtyzDAQrHhpsT/JQ0XgTAvnFEJk8vryeBP68dTx78jkk28VLHrjp/oFfimlNrTVPCP6P
djSFzYP9zLUrSZiK6cfsOSIqGL4EY5TdoN9bJJ2bPSXZIX9dMV38X1fPLFqbIcLLssTQayVlvj4n
Mzu0VkwN1e4Emb6StnXBuHpv0yiXx2yN3oL9os4UD+oMH56s6QcJw6r/tUD8NUCuEKurH40p9p2S
ZzQMfQXDGBZtOurPnZmG6HsYVonRLhcfeZl0VDyKQ78h1e/9wsCUsRnYLMDt8v9iJYkbkkV03/cX
lQSlQe8k/2NQhk2QC+tUmqxnrj7/DyN56u8Y++EZxzslqBG7hY/wi5oklB7GvP6aUlYVSO0ppwNe
rfCxvtiMrXdiqJKZ0mwBdcnozP2hNaOKCzOdyiwTsbE/KkFDNXBfGBX/AJx4MSqYc5oHoy+B/P/P
GgTbQ/c59DU46vAbML1rCu/aFUCxXXmTdghyyovbJ9/N3rGmjH/gQJEyJTstFJqLmW9YY37twPaU
gRsTNZUjgPHQHajnYdEHuZDWWmyRxI55CjosBizBWrI8l5e0izPcAscY9rM6yvvSaAcBUS84rWBg
Ls+JcedfCd3ogCn/1kwikiKsa3oRbAQN8a26Hrn7+uGpV0qXXrspRhj/+aVsuU0/N5aVAICB37xN
QPocwBq3Bf0iiaorw2uNf+CIQbNhIqhJIBSA+HVRQivPEaLuTZn6qlK+mEg5Q3HlP3/8NVTm7N3F
3SV5e/qkuEDEhxrmwFbeQykDXe5t0QGKU5BZ7tjp1OK9w+zFaOYd95YyFV3zQKuEanPv4lOD3d3P
auwjxc/PNlLJw0dnvdkhQvKlepY2w6mIEYZmyeNyW+0/F8YcOGzjmNz3AWtS0XV8BCMWCJKx3Lde
hkSrTOKCKp94fODWwweg1pXGMya2/ZC2SR2hJoseqAwkZe8mOxe0a+Ryb4AbE+PfAM+CYVIwmGT+
UaWaheNJCGQ0fNcptNCxqfPhZTWqRJD/Z1Yxc1Cepi1gjmSV7z3FfXodnZdt7xAWRGROEQmXTwGG
aij3/tjNWRBBIusIJWramGLCKjXShZDHLpETQ3qhbzsQrEqSzOhxdmjkbCbgAVTnpssBlnChmu7x
SPE2hmmXdRiCBCTiAAzYj5vJiW0tm2CbRoTnvcVA4/aM9u4eOiWvXBCXb52cuYHOc84B/juG0sWK
YaYFrrSkFjMXNnSzGnaCIhs0R2aJUWXDbfLDUUYJx+X3RH7AIWF6RmEbszxK11MDaUjVrW4Pg7KQ
vG0ynytdIvO5Dfrmd7IZw4HO6v12Cnzp3eyNXL6KbIQ2dDugFnIBPD6KcJvYkH+NnrH1SC6zMM6p
nso5BRCs6pXrW+BP3+2OduDiWxHnpYtWIY2/gZiAM44PoZS+Uc93wDsQQDpMnORW8DONNQKKWz8Y
UXUrNeOq8T+DzxjdUDOdNcO+VH8V8x1/7PZfTDBtglZK7gDbREoDEV+2H2XF/dd8ph6a5miOSqgo
+ibR/hc2B0eeWkAoYUYwsHl2RMSUBbQxPHPMH/Kd6EuQBJ2JaLTipKFmg+W0QM7q36sHJUpJv01M
KPTBaI+RzHkX4AGQlwvZK1amj19frGWwFyKcuRBp6MqvbkH+mN4m+ejjwYerzh6k/jOlVcT+jT+J
gXqJUGhbqjRJHWPMdLONoviViCqoxDIY1MjkfMBbRIdGp9jqY+t4fKwWmwJROzjvtu7M1+WT6rec
agm/SJPuEJ0X70fCsqkznjTuN8nekFUCeohZ8f2zzyzDvwykx4JBPj8s2L6gTe5hzL/EDiilO3zh
ntBBmb1diD2xGG+H7GgE1Im7GewF6+7xdltGID5Xl9onRdBSf/2kjnOgh6sQY7RUNvF86AulMJEA
sn/CakT3QlYXUy9aN0iCXgaPyGONtFIhpbwn1IgU+64wNt/oVKa+YraqSVOc5DNK5JZyrFbsfnUr
uLUYE9kvu4o0LXLCsk+jUMOBZIkOu2vIqHmxED8cQQV1ngBZrXYOClre0hZKkpY2NTmz+Pbp3LUE
5o+oRbbxKdtbUBVl3FT7sKK3VboegIcAxrqFCf4YI19/gTU546UAWPWCAL0xNfIKoT9EzgYqkKpF
6GAtnttwvBY5aYR8deGEVgL383fkBekD8Hm4b8kpzi/D7wamAhO8FR0BZgedz+r30IllJw1kSrNP
YbvIAtBYOKvC5rJGOBjK0BZ7ZK5pYnMlPZHIZqx4FRNBn+gJHD9u66QX7VumZ2Sfi38vfrXD88s0
KxjxL7uRO9YB0NqH8o7tccFkdQ6vjclEi8ejWOaIGS1KP8JK9f1ECyX/wNvj1V2Hx8EW7Bghhuat
uLg9xQu4oiOSj0YxONHctB/9rPS09768owG9/++V6Kq7m/nI5Mc8WkhPU9gYefdh9faNdCCGtjIO
yvO3mnNAtggpM1GnwrP8IUJAezBLy2yhYvB3imYnB7rglyUWk2T874Am3fmR6GkkoDPpxEhPPG8G
KlZ95AFDB9QD3fVyDr3yWdFJ3/46voQpw3bQAOjYqTZZ3GuZ3qDBjD4wShr8KPuT86M/6YjqkB+5
GLR5oF8dXSO64tBYI6DRp2xQYr/LMeN0nnfeiiuJv4n2YPgXaBK77uywlZzI45FLsMKHI9p8CQM7
GKTF3rONSfRaPqIzPzKoXAH51352Ppmb1njxiivx43kUm4W59mGfvmX32za+f/a7Ql6Hy5FR+M9r
GHS0F7qk25X3sRtljc5RP+6kdq018rs0maHee6ssJyQDltstXziVEdLUqatJQ/kAqbjngCrckcpb
KJkKtT2ccvZoZiVj0AnR8WMWssj6wCR0lpLtbT/4NBPatYhO8r4jENeoAHOXbh2xpzgC2vuScQYa
gAOkOKzTG/8u2851TSYGyTwEybiSNbUndTby1VQl38Jdy4StDy5htNZUJD4mx9CpUfexzDLzrMUa
BiiQZGwgIK+ErCnieizA9WyOkwy8W6Z+/K0Zvn9My3JV0T6lOWOi09nMj+6XTSAMN61BJbR1lPLg
/XssQhYpE1LLBMQGugI+URir8vRrOdn2ZFjWZxhor/Wn92i8/XBWjhD+WlvyDDR77yW1QnLCqq7x
FWpK66AvH8XA2qjcK3xPxRTm/unAJK5dx5BJeyv03xiroKWJzPkwvFGKUiKJhVjPvUEbTS8oKV0E
dnTiesc4uIvJgZGM+MCEEfK1eri4FtV61dvD/gId80IMduiQJrDlA70uXfAyusOmL1G3hOivjhqJ
uFG9qRkUAj5RCtD1x4cYHvbdQZhNg9JV4H6Rs7sCbCZZ7UqgbaA7m9neGms8m432Djp+loWskNN3
cVDQYHBhLhoKrdzSADHdsH5HRpgtINesIhDyY1IMtlzG/qfNw0z/ik5/zRYzTyXVrE6twr1ZeWJq
VfDqAnA04DXRDHZYL7IInvPxCogfT+ngy3JBRpw+fCz8xmTjCL6QcxXLTDLmC2x0z8gvxVN2ZpsJ
CT57fkkG28PXbCSgkiTUig7RhS3hvFKata3gGp3ghU89pEnLxL8drIBAMUiO0h+h7UaCzkZWYQsX
jfeQSRxtkdJMiA+9qjspxfVWMHiAOYr4dkyUfm1S64iqFkF+B8hd2HUbbcpoWbrYKlJzQ+DkQU4W
xZmlBaRpsLezCEY7t/mWmbPotKg9iMrfiGR3oN9KrwlYIZC8NLxnYLaUhPiXfAbTndlTGab1KF7B
h+5XNUkx5SP2dBHGY1NLjZmFyopd/FW/UFiCmYes0j5fOY2emHVoAW3bGjypcTwuZDLc1n5LrlnU
zGCc027MfJc19+hnFqsxuB0xgaISkGk1unPm/+L1ZTuUCudwZ7OdbZmkSVIhdAjlk0B5cluiZF03
6dYHJ5d8LQLzkuUvtWAmc8Hx978xjZF4nsFZrJzqjYruYSBW1bOdHZRI+badwf1yNjah1Vc+kA+0
6sFK2hnjpPPwnkDdHiZ3n8FU00PZzH/stvTVPEI7zZg85DuY1Vs6p0wVPea/GMZcxB4xcurtx9JK
Ood/7QWw567WTKQpZ9h7bS/3l1or9a+5hDZVs/8Pg8kZIPEe7q4bt121mA2UcRXOGnH8OULpqStT
XlltneMEK/YEsgUvS1uiDGIOFVj3Ywz/R46aWpl21i57tx/KJouzPkHEHZpz1zvJ2AusLM7ZMQwj
6eSBSkdjv2GSRkFOy32ttWKpFIDoc2Bn7RiY6Yds6XxKx9CcOcA5hFXtkUtepADNC6UIbgeDaBZu
EQYj0qAsKXgpl+f6xrG8E7gHQ/Bec944Yt8QAvDUBvyZJctc5NJqSqnPhEENsc5pbQWhZKJcjQ50
+P4vGJDPeeHlKPIrUj2k5n8kZpKB8lvdEITGHsxwUBS9eR0vO8uqUwFLE0yB0u4f5HDEUzeirZOB
1COclt1mtd+vzQuhZk43exyYjla/ApKgq01yQSFUQxT7CFfAWNtHZlF2JYTbFE5+v4iDxRKmwhY0
+E4YkYylhYb96vH8n4ZEIQjNnV1dcKv8e5MYYpthhrabw1kBwe5cm3gGcQpe2jl3P+wAV7Lu/CW6
j92RY2KBFMhCUBZshmQb087shWp5nMjYpMmZYe30CSwJEAgOMBsYYXwyRuC5uS6ZaGNh3N5f3tD+
nVmKxVq/d9vKJYsQGPArmawJFMDKk5cv1VHbVG/xH/fuqneRwxe5pllRA6UvJM98fwwOmo4vD5zC
OBkd6i61awVxoEwyrnEAjuF27s+46lSUdNEnv+bb7D6iH3TgnmBoZ0ZWraYtb3ou6VN8hEBDbf0D
ha5EEE8L8lgjOpkdjNHGVgtOAAzVtUnD5FYQRElrfasg15EodnZX0gPVwu1NGiv0qThG1lypbCz+
nyH8CkuczCu29TJpqWuYPLjnqlwGo++RAz+5F1LlOqteA7xxIBt0d2HJ97vzeMN0WFRiPW8/xKhi
wKNb1YY0yuPKbIk9TVBrmpnMKuezYBjMSsObL6cLKFfSvJoOmzTnEtH3Fl1BaBRtWWyDq4kGWPDB
GremQZXGaLGyfRpBZ0mhfyT6VM7zOPTLBgkE5GWZz3NBJHqbHwl9u2MezQQNzJca5JioFbUuCgX/
q3u8+RlfJD207059Ri4XFKlGI2NRpnTekPi2pm6Fv4RDkokdgdgesEwoJEwcb224MfYbAPAtEan9
CoBbt62eLIb4Xr0zMMWdEOOxhB5ClsKimpkuZ/TNvnubQ4R7ZnrEDlm70oLrZ+V+461wHtsYrw24
ajJJPGVlKFZCVqrnAfg68Z2Gn5Cc1jGGM6ZcuNkSRwZ5wmeFKxWSBXepE83J1FLdMqhq1l9AWXry
tAjGP/EY0yFzblKGUUiuU2HIlCDx+78ZCx5qViPlA8Lu1ZJMwIy8YD6/m2TWq7wfRZjwkldCwun0
8vAaQPBXAJNkaUSC4M93A8KJpzpWzypWSFBzd5zkgMCBF87f+5BdSb8uCBrSBfVenRAD91cg/VpK
NZ5ZdXYk5Xhy+0Ch5I0kPUMNZYYfykCkyRLsG92JpFuvoiSxk24eg5OLpzAt2Ylk1aTNmLVokAFi
a2Xo2yPr7ubG2mZzyrm/3yFsCFmsjx6d49EdP3CcHcMxtghPaimWQwaD9X9nyvHWV7Z5DGWnGUat
ET3p5ATv+pkS/gak5L7BxQJGu3dbw6Gtw2ru/46cymcoxqZ9q6OGsKivEPc6wTFcdD71FDZoWLfH
oKG3DoWcnTiWcUYdoDyZGF++lZ2XIK1MYJuRFONC1+OAl23gFPwrIGUz+kNfJu3UhqDo56Fqnb2+
94/PneZ8Ie4/ntyVzBw0iRj8f8ljn7FH9OLzrLYqCoL1h9vdimlXLSAGaSOOjjXCgMjGN0dAl9or
6kn8AxvGld+0/ZB6NOkVlOC0Pi+nLwh2U1tj7ap8h3qhuJEMaaSwTfKqVl3eVqg1efPRHRQOVsgD
iXnhKkyHFAqxC4bMzZOt0a0GErHi5jlehcSIUOAvpKi061kqaRpZeppTMkW2MLSi+ecYJZWP7xEf
OmPQEX3eGvVpA3KCswk+JIigDVVY6Pu+Lqvin1DTAQqlWQK9ahtn4YGtpyA494yf3z1tZGYELNIQ
HyH9yqeEQnBIsTiyqrKWu2f0PTdw+UiDjr3SSyhHVWDrFOHQOCsm1u1/yhzaf3Jrp9h4WPh+z7B4
HMKHvpfgcIxEFhVyKAmQw2C3/aKyzcW6mxIooO9onc8Zf0mexbwZoNICiOv+7knexoOTapUw5Wof
nWNtH+QulMFDu3sCkZ1DJEP7thm58kWLV8DodvQbRWk0KgLAE5BC/3UyGJS5D+L//PYVCxTHKn84
bNT2iwVHilVuZdFwFkZ8AiHfDbhaTP0m+jm/RWmO5IGI4MHub9uWXapsYm/ODh4c39X+w/ULpQSQ
icD9oENfhQC6cit4w/rsdSUV5HocEE9+Wbqsyx4lsCVMtFiTzprq7ufpWfLmD7U7uIems20yYtaM
b/BMrQ0rK8SHswLjrTL36iUJnAu1raeVepfm4RU9IY8rb1mzl+/PptfNlux42Iq5D0TAJH+YbTco
XG3Y8wrDwvnRjDJVWRMbfIpBcBk6hgU4mm/MbmvGY7E8OSiDIkbJT25WbLCjxLe0MjKrRrItMajT
7wLwgr1RGgoTtDWf4VfgHIxtrK+bjkXVrQb3owugvB9hbIeOl8NAVWOan+9B5904Xh2sbZ3ffBDS
o0TixccYGSXOqLtFYGJIDcDrQ/3rEKI8bVrpUmfvkVDG8oXJK/OcsAW9SpWu4WypEGzjr4MbgWWz
byqi28aWyXJq/W0LIFz9Zn38judlPUbQ+4oqlG5ohO825wHwFSXuKaJ26uuXeGQ4jOe2X6OnN+ow
42irRkw5ZChNK7hPBNOMn2+9/jmdF56/3h8ObUMU3o5uP2kekBBRZb9+TZgDQ6Rshs52Vf7PNbG2
t6QVX5pXLFLyndsuQPpgvXr5ur94enzlzpa/F2F/P7Jp42D63NJqjWsYlRqd35FbYLi2TXuAuR+y
gTLdfkfa/6hZZHCJUkltwLx5Jes9zSLeWQ8dRnlV3tG0HOaCkcMbe45kXZYTba8MIbEeykPx+LUl
7dBzvveQtQ6Dtx2GYipdWiAF/NG4B/1bkeNRQ9Soiu3RgROQxVhuyHHb4HY1neydI29NqsL4Fphi
ehWCnWZ3cvgaBlgz/095Ag4Y7Qgij7cPK9HvA2XuojmlfClQbESpAuLNFeO9KQLMmygGaDF/mpfE
Mp/JIP9QodpHXYYx7R/OoLn80DLLQigIOC8vN50589hSPU11bI9x02xlYrv0bRWw5Rt15euFK7BT
iSWusI6/JYFhdqblTWJHmltZZxnnMqe6vzN70gJ3lOZjPOtccaKLsJXTsX8sNHIacITbnjHCWUNX
rBnxaPYDkJOUk89ITJ/2XVqVi8brif31Z1FRsrItGiiekCSg1qOX9oCzo5KCFG/4gMCmUFHe7g1F
LVk+9rp3UH0LsHOpGUvaPDNJ/cywhpn6ZmO4z9zrRu2qG+hzAKA0V69KC0x/N0mSLj7IvOGevzXs
+rpCdNyEAr0DtwI7OLnRa4sdnwlgtiVn2dtVlJMzSmYhTrU52/49lF3M8dA7EIeRO+uGp04+iehf
t7vCQsreBCcI1LlZtrZS2G1MVBRUKpxK8cpM3L8i6k89Aoa+6czZ2f1vLX7PxVUW4DrMVgGlu2S7
sP7CT9GBN+hVhQAVcGZH0dAfl/Zv3zU0TM1WQgfgc8Gp4eJlaEhwhRnVZw0JVJv3DFj7VFlSzfzX
Gohb7NgI/MYBBRCp6rwB5xM82uFAy7j/cKmxpCKcPITWa11vFnafp1XnhmYAQ96zDACYMH/2e4/6
QE87aKOy61PGmSUJZ2lAqAeyJRSVoV8P3diVSVTHZoiuXmTJJVvRP+eSpjif4EKVs0ARbWSEXcqU
l/TpEUOlj5HGzujxqEWJWOCERzX+nNS2mhkJbi3VK/Rxzsle18gFuXHA8ngNcU8StDkHX3IdlTw5
8Uoo3fzYHPnRUdhD7rJzJj+FPIZ2gzCbgYvsLfy7FobfZk4O+xqfSch/xfFMjSBRJ+q+yIziNhNi
8y6cojv5S2eaWC2eSUGmhHFaHTrfeFGTfJA+6JNtCePxF7Z9X8+6/RitMX8WuzQQaRFOfrgSUEH3
CmbPKWxNAW3rei9Fm1gEBU86/+kHKgG4+y9T/I29VGlx/wLOck/D0utPNYRzjm85TOHpelwUsELI
KLqaR3ZRnS55+ZZuSS9yjAqVPUc0xWdk92r2BZSsDeaLnXdOoeCzayQTLS3XaPb9AG6eBsGcTaBl
WY6pCbBXHoKtVE95Vm1a7nR3pQpOHO1c9xQ9hI3dCliSrhaBCzgRMuNw1Kc89ilIdylasX/J70Ap
Jx7pgoNpICqAzthRGi3Ar7sjY6SH43Hs2HMKkybe/W24HPKy7lCKnN9Xd34zIIKZdPe+HVcGv+Qz
H7ixn6TP04zNESlUXn0s8lk54uNHUR847bleGSbsQ6fY44jofuRKyKBDvK4gJ9A7MqvkKtuW2sAR
bQt2QuIr+UTvYioVpcl9bIf/uWwjJd38qoLtsyaGM2k2J/DwTGzAIBCx5rFj8C/TuGW2lqU7i3hX
TFL1/Hc7PKllAj/Phz7NxnH51RgGfVO9Ojo6p7aD2J8h62T9T7kzm7CAj0TYSX5hhbKblLxRnj+O
cXtn9q8IzyH12fo8eUVmwQGPvF/ka1kHmgyS3nekU5reHeIJlu3SWFvCSgPKwpG+kQ9mY8y9cHee
A8B8BMoXacVQGVKjvR2Gvd2qWBIdE18UunZLpB5pUmw/a34qUXmCzhnQszOK9kdEoXDjm2Hwz+e3
oVi6QwkaaLf9jK4pcrme0cVa4hiWz0MOxTvuSqCONMPkO8I9kWzEFfaGe+aK0fq7atvCOnwnxVlO
cvas//+K3YBdKe3b9ItYiCUx0ryE6t9mHBqSDrkm+YOgRhZi8vtf6T01v5wrmVkFzFzjrxxuCJ3j
aAgd+7ZJ9EkEVkYSUXdKaYQnsNxQfsO4MXD5CpmNYA5pMY8rR3r+ufg4VWTdST7Y+X/YTIY25Ymh
XGEBuBA7iP7CkzBlcV04FTPYqFKQ/iSjlaITboNARGcC9XIufKKP7mBSxZQ21lz6BfT8h0R8MP/5
e7DnFAu/GXoBFkGMMJGQXwU7b2fIPjOa/H7CPDIXy5D5I4v7mz/hQjhEWuLo6mT0NmvhDMfjbSbo
Lu58pl6XgtVFrzqiNatYnlVAPqfHow6b2Kv6Y2aK/PezQe0foiqtBGQW6VvqnDT0o1NL/5XEDAfb
ISBrYcrppjLa4MhdxtZxl0ruAjwJM4yFiuOHIrVYFve56Ne0iMbYafhQDqGPFcvHdP9Kskx1HMLS
whV0868zfWAW4nOpXkV/6kPccHZKZn4z7glIwwgnteSof7AqiIJB8LMnSWOqZ1xJW1UdYGiRE4ck
W72+wjUczxuFP2a/qCtCUCM4Vcjve2sKgrYwx8kWCGDs0411KWaaVc9WdPwmESj3xrivFYkUwORF
MD8JsskaYq7NY97jLYVeAhc0pcQ8kLrO2Nr2d0mrMdFmOYdF/J4qrmpx6XcJURMazgTy0Raunz6r
8Uy1TR3VvKxjvqEzyHrPiFq0PoyKC1+yTscJRUPzmaQsCCUsyzWvgN9LbJpaICyMYUO74NBWcx7M
KEMXjoOKVu4jbAFmQV0zDx82ihy8CZSEdGjWzhWALbsLLGnmGmHz1rsBd3UDa8pSqB0fvetvVSBP
s4IGDBIvfJ7YKlxVunRIklwI4lLNi/+2RUx7uh9q3xFV4j17zQZyNXOVfmqvCKlOfpvjiaW3kaFR
oH2pTbyIiZmhHrQCckd9UHI7nd+yU2MejpdxRbS/Xp867wDaDEiq5Np/3WcQilliGnDjpC/rbA6N
m16p9vA4mXNFIJEoHEvFSpfEB7Se4VIv0ZMI3Qywlh3+3DwK160H2H5QudqMxLKuQELTaLkChUgl
2LGuwVP5Nj56GQ0Bd2f4+RQzubhI1qY4xiEdb46gaKPjW6fipJ483X00fQLkCMIuTWZbhKtDb6eF
bdg8c4TREHdEXv1UJ1n0r7s5pzHHl+uYMoEP83P1KJNQzYcSiiFrklBpLnEigLmpBx/rnB2MX7tB
+NlKpx1ig0mFV2ygEHCpOOeSwIIo6aUK2UkjVzNrASupR8tsFGSCok3SIl2oXx3fckztflQKjXb0
3lR1dt5WEPmNhfwK8uCtxzopJ1vyzUlx1z+PeB40VrqkCOwuXBXHS+uZvDcNzgOzYlFXsbLO2wcy
KgN8gIzvjL4P1HMyaQlwL5GESHaF3wvhJ0/hd6xXKFiYC/r7Fx292xEkiEdGHCyoLLza75i5lHZi
GGn60sdRsSD9nYJzOMWpiAHXsEQFXOF6D2rwg80YcxtWexm937XyGhAvFSAgnvC5bzX9YOmO1VSO
92srg9kLiqqlAKr6SiujAqVnKpOLPydqllp3SVUYpedOBFmDiHRq2eHJjZdWGwEzKi7O/syfD50D
nTFRhbmNfqbu2yYEX8ACJkLjC/QnqfpQ640oC62sdBjkK69IIUlq2Dn5GYVtjCZe97Fgn6YI3q2W
8tPXVdI0la0i0yvPOxgqsAvPhCKWGvtpqJRmm7e3JX7IUA98kNxoqcotT9Pf/nB1HIeV8sesvuum
hXkQeY0gq+7AD2n8xDFN/VkKV68nT9tGZWZDwD0eWFvcEkLtd7SLFlxNE9tZEfpgNsrlVf5HmPlj
XozWnlfacyHG2yog5KZaukMoP8T7jTjUg/eSAsNrSU69Q8V5XS/JSsZjiJTmLCaEpIYhF+8bYObT
UPbge2Yvci52USBVsYj10M0Egc1FCOPIbvH6261AGFOgDNsZSrc1NIvTU3fBg2cyrmnIAtGQalqc
+G6FmK2brMwdVMweqOcklUblIpItFvjac2pjv5jUI54Gllwwq4Y3J0hSFj1zq8n47YTi79f1uxQ3
tYjRfa/Esqc+XPh1xd9dZsB1ezbWPoX7up4N9DLJRjv8GHNrn5zyuwLKA+1SWTELdZs0tJ6l2g2f
XUB8Cmxo657g0OZ0CHj0UnSK2cNjsuIjDGWj3oR1COB7wKUbk65piwFo8NyRFR18dFKKuHFwWRiB
8PTWPJV95Mk75CPx6ltbt1O4bhtk/V95S3OQBIIAkF+MQqIJRZST2zMJXr38yvJIf4o/Pi09jYQ3
rntn/uw4iBOgUFLjXiUZA/wscMqUveBcTszzB9ZRRSzFlGciYv0Dcc4a/rpoRmJLoAq2E2Sj0mHU
muhLDR+VkrKiVisdr27EMN1uhdrCO8tSCgN8vd670HHwMExrtq44BYi5gCvUQ1T48WDK7tKP+f0U
yHVYQ1Fag1fVzVpTWGeew+zG2xAQ2xhb7Ra9U1XuSgryqRmrn4LUMi2gUa44qS0KsiajcRftNcgh
V5jhDfKbRKCxDKVA1WrRYysHxy3Lf729+czvBqFBb8Lc0M4HIEDHyz3Xf9Q6mfjmVdIfpj7i3dmL
dyWY7mU2LmkvDpwFhl5fvMC1ln7LvM5P/MuWL23Qf6Uu9tNie33fILwwN8LDApTncKlQA5CoPctr
EI0bg4gfPaWbokaayP9RuTEgciewl9UFSOrW+S2IjO4qfqPEQpRGVe1iYbR56u5m0WSyisDaTN47
HlqzL1fx5WyDoOwABimHybVHnHVZDNseEqyKAG+rDqXWAeXYYVPfmuxemQ33cMkgAgojjiYP8joX
jDu30Ex0ZCYnYBg7brw7HSLkzJsJZXkj05IfdVsElzR9S0v1B8cuEq00wYLiToHrKGGRQbV6vMsb
Km19PhWsFy25mzTmZxd/syiHa5aiSIEuK8zme09S43RKxCvAP5ktFmCBM7eu/iiF2mkRS4X1tMqH
ejHTtTsg4nBvFMDPr7Fxtmuws+obiDpvCQ9hnx78icHEoDpsysLbq/h4f/7+uQmNsaOySwH1a6dx
JUB9Gubx9b+lD5ovHRdE2oGtMu9umhc00Yjb0CCOSTkMOeew4rcNF4lWJPuM5YHufmtOTmfqb1f0
LpvRmufkskaAmyCboKR/ePG5+v4J9o+IrLn/EBaKYStOY7M8L/0dXp9bWhFevqEFxYxy0GHyJ9/2
kNtEdt85zeTGYYyCTx9cGCxgYrdiMB9nml80CTTaprPoyFVmrX4Aa28hboqIvIhdx9y7e4poMOAv
+MlXnIfAmIua1X6xVHsV73R5J6mSSQz+A8Tdkx9F14Ai/14dUmPR1j4A82MDSplk9kr+wfq1XnjD
iKSd5etzrZVQRwo3gN13q8Ayu13yMsRRY0OIQU12l4xLUqcon+tlDQiy8uxtj9ny+nFNmsRVQ6Qq
g1r5dzzKkVH2DXEhhE4fyJB9spdN5m3zhclvEfQPL8eyG2O3z030Puxun/xUWd+AmVE8jNJ+l2mq
efcQF9eZhEjxUlVZqczAj6XNqQgTJcxY20C0HBd41gpwrzaHCLXkfRZWOXCgeWkTOmN7UrAbOCwx
KxwsQQ82Kx1DbD9WML1uMw866K7LSTG2WArKyZa/WtZMMCmleQB4mlkQx+HqdXVBR5SyZFrE/lTX
GJE2P7fueQP8TcDG7iyoxbyz/WqfrpeZCpbDMUh18fh6T6/vT6ICd9Tzz5ZImLI014nfsLqknN58
9FVM88CFsjd+TlHd/rNIZsUndDruodIf6iP6Shv47JMi1ZyfguQbIGm5IpGk9FWByRAbHGwiRl05
MvlkmvZfoYttlGcga6mO+34tfetirGApxaYQY0LPnKsGISoBBF3Zsph/6ilUJn8xLE1D7j2+tWPX
juyfuZym8pBMlUXUgqbfgrT2ZV1uuI9K+lVSKSrIbQZrxVyQSdOK3/7BSW8voXfUurKQSwLkIffs
UrQT4wfgt5nlfdN/uHoIpFwQ2b1YH5/ta3WsRLwGwhh/WU3vkFQljshweudfHDvgVUZeS20krnij
fIRbzO8L3f3qKhnbpIkHHBvN5bvESggnX01lzr31ltJ3Io3iXQSe2J1JVUKcsST9FrFszFzYdVrc
LorikGyg/uEILQRU3zjo2u8D+CHqqPRLiFqU8cfSnZXNZALp9/0J5Daut2UsEAB8YiS4Tdp9u/gB
7K+d/zfr3DfB0+0JiXP598msNkZurrDY4Bsv5VnkjdeAln9bv2c0aIYlYfrYkaqOL88AiTOyTT00
MHkqZmR4948uLcW+V3YU+tE32sWEGJZs5ubG9eoZA48DoJECExmn2SvdNfc9Rx9Zw1T6gGy6t5gx
wt0yALnSo7wCcSzlvwteCuUIPWunYpCqtPf34y8iXJh4n5SPsAqBodMFQMF5qbzJ59p8TpGQ5eF0
PPR0ts0k5l4FErtUa3+lNxFKsm/AuWVsP9YeoCsfISNNUid2zLJfUC+mv0uHRj4JPsCLH7LLtu4j
v5SZgy5/sOr1KgfDzeYTIw+Fjs2/IUFU2nJhn8coSMQqIN08t8VVpjjwc/1+7Bsa5w/MBpKcrmqY
H5LEISaxYX6e811jxDqsF1R2Hhq59EyRh6R5qCBC862KPGS4JcRS9Vo8iPKAHvtZH94QN5KM+l+n
+OtiMSf6MGJHHtt8/MTNT+jsE1lc6Am6XK/cZx3G7vRJm69NLFxQLDsNhCj3ktKBWqFS2tyUqs9i
1z2b0BRkCT+silcYAjyKyV5CyU7GyECKtWDySDl0kg2OrmlklfhPUrMCDzwqssm8Y1SgjJXWiQvx
OL0fU1f84/1nHKL1wrYjnq7eGe2qsfj2nwpzmrxv7aKu8KKDQJtx33TWhv+HK+L+l3tKF+5qvtoB
FpBbl3j8k8kWDunEhWAcCj+LPkiqZK59UOlJfU09TVqNN+3LlkXVVaP1WtNhcNLjjZQHQVrF/25f
4gbyRuikYwCEbssCHUd9uYapztKQ1Aq31o5y1S4DwGZtyS358kx1x4/+pe2pTVUWvEYS8whR0ZTM
+p37HQAILHA30m363V6YOu9b+jRxo/KK+sMQ6uPr859g/2UBw20aDe0w7A9D6nS6KXKV9+TUHObT
amAjNLYwsh3brTZG85nhhSs72Fr07vnVomrslf1zlhPuGvIXrXHPxo6ggCMOHCYUBUy4yMiNgDVl
bx2SGRliwmvPQaV/ApEJNQfQhOiCVKeRvIaPhjhMpx5G6LsaXbEMXIcS6/TciuoOU14QOfJcKqSJ
RWlH+Xn8QkE5bzI/n3daxXnkozzPHl/kfLpGv1kcTZwvCcXmDKiYbfxp3KTnEfsiP0Vm3W4lS2Nz
cBkRFW5ahPS8TBFOoWJObPj0rhFBske4PY6CWDXqCrFb2j1q0Z4t9QzNRQje+kL+y3efRn+I83yf
iwoo1cHux15f7QZzcRdEsotxbGXguPlio9M3ZNhh4aapQitc2JbnWWgS8fYVnZ/DdfDHvIAjgbdG
V5JW/G/3gkPYOC1jQTKv+h6cGjZCSq0YrYH+O3B9HWOHz5c662XAFGDu3LtKwsE4XxQ/G7l0El5s
FqeuRL+M096FDOJZ77Yy6P3kCFGYNoxJxniNVFl9+KQCoaDvcDL6FXUzjrDKLPmo0mqvxUsYcaDM
WfZ3TaHZsC4OC3fHMAkKnMioFSDXAw4hQFV1g/P7gRJHqtpztEkG/yQIVASWSdaX2b2uJYhDmc2/
PISWXiy4/uWb0kX7V5kHERHRDWn6wpSF14YS6zBps+nkbTs1cCD/toduBR3hlBV8Q0ZrKvY44Ycp
BSFP92vGsADilcQvyTRtDIodAE2TqNsQWXEZmHs9B5wjx/rS8NL7rraorSs9UWDQg8qf2sUVBoGo
4K+o/pjhxFaIBzhg3aYMlDhmDkygQJSZfkDihGoV8u0ST128xrLDP036sMrlpzWKhQ+MuP6QvTT7
SHGeQtEGknrz4Y5LxjZuR16O9ph+qQuYGK0wefDyrsfo/1I1lYk4IscBWxnRMRr+GBdhWZUlTqJN
4QLhmfE54vt468cFTqb5HxMx4TIDV7PYjo0dIm2e8LrHFrXRhJ+URkAegxdDJ9RbsMi2S0+mRzJz
mD2MLs+ZpOtbMegeS1ttWcXEPanfwt84QlxxbDkLgLBd3D6ibRzmmqRHptkpTblqbZEDVwYKqYAO
Sf+WJygzq9d7O8PNjiOdV1enttEOxNO7Wk+hnVpePBHMFzM2tC+/WY7QEQdnnvEMA9x2DBdmu/op
uKxBgAYTJYgSbl6XHe+MH5VE2xhLGUsXfaSzARlawlaf0NcEqlVr6V23u+sH/n5lhz6gfMkR5BG4
qvDi3FiKd+cdHwvHpX9Do/ABmRgWF15DDWrxkpSay1KE/Zcv0TLU12cJKds1RhnOCqYV54mPAD/u
mVZudVb71H0AbxegasJUTaZapXALTStvB4F0ZrmITZxxj3SOYXfKd51S2XFm/zuHrxtAKN0Eq1+U
vL6/XIt0/9sAQWKOJt66yUjtlW7bwzNrnQOJpaiFEluyA18QYbrvuC43FWEo7yjszYIzqjMhPRxt
5eIq5oy2UZtqKlcpyM2hh327zXuOPyS32LBv5KvFKPjsshi9JXdxpYKxz7AuJNVPIAs9dlEhK/U1
94/M2fDGGOmQdNrEL8v+r9TZ3jpks5Htpx7TVm/zf+bOSlXdc0XW3t7uwg1U9ZmFRob78BLeGDaG
p/hMUVK3kv7bjUzM5b2Su3ZGWAq7WdJLjC2e2qmRs/Rgv4A6F5zFIOauEfsjLvM8lGteoksN4jcL
6HTF4whJQanxQvi6Xu3Vny9RQYPsfwPXX6/02viOpkbSr4JBOZrWFk7H/s2b3JbftdRHqPN9wsZt
+ahM0uhB7e1CVji2vMXcLSj3LGk2Klbn1LHTWmuDkkvfAD3So8hyhokSd/VX0ID8ADhkkd7E69/y
WtXMmvwcjuYXglvrZsG+eTe5TAGGWICBu0AWrg5ZJur/j+J10/4JX+Es8eO+LCMIr8SlYl9WuC8i
Igv1nGNSIqoV6HQFO2RV2C/tdkUxQpsVUc9RoLuw6YSUGjQvdaQy8esiqPbVvMiw0Xnj1iv3XHjC
wnXDh6hWjdjLHnzHzvhhC0mXfj3KLJh3/vWnRTtimIq9HpXXMw8EpcbXxBn9HQJENK6v+eC0+Uda
GeWc7VeQkiGfXIokJXzOpynoXwq0qEd0pwKcNmBqArJ8VBP7cxJxeFvytNr5bDK1T70jjPrmILmI
vfympnJ1YI7YnnpjrXgNil+3EPOLtDvm4SiG94GZP89cJ8ycWSYTxHVV8t3rwVEA03dqbgo+nsKl
cD/9fjYxwicXH0KZZ/enDfHAfyADLYFLs87XY7UG2GBM+jo8wWQxXogZQjpgL5dAdyxRSWqkH717
k/eKdCZ3YuVhEYjCz5A3DYWy1UEo9R1IQHCWMP66tmNIBhuAKpnO5WFiGAOyXrTbBprWvfGLw8UG
a6YOuoOJMmcmGh02UwMmCnYBtwFaPhwE1VH++YplKg9EDpwdAmH2GjlaGVfqU646aKvHDDE42Ozo
6FjeS9CHfiTt8crKiEFp14O5eQBXBWpBl8wbmqZDFuLHgyzrcEYxdZsnCo2oOKLpRRxQStPm3f1Z
NFa8PacfDhbf0N/1OfY/EyVZ8HMEBeKf92Jef/+qF4M1vV4cfsNnYEtDsgeSdOJ4yBf45vLCHVJD
tOTWvvFYF4LXUvH4FtykzOWXj09vsaKkhXh0OXQZ4K/ZzlpFMoZenPHnhZEepETxaaAN9UF2ES4w
YN5TNBjpRYB2e+aJ+n5nkdyU/ZjYPe1ZWml8Gkb4rm27QY3LY1aIiS6dMbu+ny/alkIOYazSMZtM
aq2qq/c/LbNsN7D79qQopdHH7fvKoKmPIciDwgW/KVBzE3Sh4BEgywO6Hr+aG0P14NkvHxYBw+z7
Wo/Gt/n65tJuFDPjL4PmXztltwAC6GY0pctbxWBuEQbFJ22cWAlBNNdGfsiIyHB6G7+bzMl35ENS
C3ZkL1+DUYN1It7105/5ieHrKDHNiPjazpgj141Rk745NDZI8xI0HBCbIHzYokolT6EQxXCEGapD
eIHjLsWSKUtHEOFhO7QluR9pVstzGquPDweAblUumZfM0GuZfe9KgW4fnSottmkEhZfOUdTsaIvy
8DT4HSWdzEVsdNsh8DIK7Rz1AEgIwGkjyxGvePL+/mpjMAhXHXrwhz/yv9GzL+M+YQ1KAWhYTXyq
0+/3TZHvXHyOvQ+ETeNfc44kpxSWhHVqRXf+xzsEMRkullBkHXMIsyRachjZm8YSPu5wxIyKihoL
a0IzfWDMcm/pEn9MXWRHt+vL0ykpaTHtrWh9a7mvE3Ku7ekw+ysKtB8md1IXiqMSBef1b2DtxMh1
V6PDNvJANyIcqcJb5PcXVqNBkYW9b1bAmngdpQ+uN+TIDHnT4n3xWvghrl6zf7OHO3Cjt5Di/2Ao
uaSm/nCynwZzJeJeuvB69pHIsLrpdAb83uB9vnnTwKEWOx40Y3hXg4I4XpkXPDWo56tdZ4dNxzYa
s083XB335oQgdCYs8I5bF07g/6Ei71hQAjFGod8q88Srv0FaF5sSOA4T1PqMMsYRvrTfpRgNTRTp
rM3YPwDtn5jG75e3nvSDsAbzks+OtMOk+rN3myis52YtqKSiVt6tPJ7YzRg6QSHmtyRSyV6kZjvF
68REqFqC54yfn6ik31uerFo4JPZSTBJuFnk++y7xlRZkfjSsuDtiUswQXexgJn2Jou6nN+GkjEP+
3imkZgfnhJ4ERqNqRPV96CsNGWnPVEWnKUwvfJtEOhv7Mv/p0u076mleugY96yZg7j8lXi+WJHac
3TjzALZf5duxSyla+QtjkKn1u6OO8uoW3KwU1WGmF8y76fQUv4hDgkB362tjEJB96XWuNawad/uM
olEHBmpOe1MexdZTBzYM3IeLQqOH1E4Eqbkwrs+CvI15HTFgfdW1dVQsNsVLPmJ4RIHrbWXFjqO7
VG5xvNWuHYZ5HVLM+0K1QQNEmKOXUyP7lTZMVPFX4/+DWzERDPdcpLuL01U2z0EsuKNbgPLZ/y8A
D4nO2IDTbAzN/+fsdsPQAMLxnOml968P3egTgU6n6tvgq+2IrTDgo7pPrOIyBYY5drt63j1V9UFN
fCuQ6fNegTsPKJiRwV3lNEPbKQwqpmuN1WEfBx3cwP+fJuZUWg/V5Kp/hKz1UwEWDS3mo9m+xDS4
jXFJjhnFHru+1JrF+QAvhWITCQWJZIWwFpmZnrKBHuJdn5NNpySU9Eilf0M5aPDP8q/sCqa7nbbT
0xZR1x+0oxbfoBQbeVK4vxJQWFyqYV+ynzp93YVo1Lpc8Ph1e3v0Ab/fgCMKEcgZO/3YU0FYGPXU
AqH/FRd24MXUe6fjbbjmFLumwo0MbR0nfP5Z+z1Q3B3DMxMzkAqpdbRfkbDbC1wf5ARO1SpkCxE2
kqEfKRaCar/EADq4QCmd52rlQuTpFUPDm6/V2O/Ar5ifezNN+yGnxfNVfEVcyNNGYwSLm9HD09SY
0ftlF1cY2qRMm8j/EH6iEJJpY1lM6sUAFWzaWU9YOvTPJDKZ+lFlxop8mfUD3xB2w44RIo+RBYo6
Db628xSYbKD7B3odp4CGVE7DlL2QFDPnDxLXZeJ/ihSj1Fh/oSVhQGQhO7K05ReHv8opNDMNEKxZ
T7IiYNPioHb9buIMKNsPxgTASneW1Ih/tBpgyXXdktUzgWcLpvBLe5wysY88GEXxzkTQrPhDJsXY
wgWLRlBEyxg6SDo9beCM34oF9vmm7paSSEfaa20+fxn8XyTeYVVYU5UMmx0iwnMhcMwmL4eIV82t
p2eBNVNCVA0fYVncnh+giIa1Hkzw7F8Zzkm8L/5NOUAIveVUYuA1ukIH1Z0hayls6N7Xznd1RR1e
2UtigAxLf94UUxBLoQ2dBaPinvTT12vksox7icnd7mOYYyVk5aIl3NifEEMcJCUxPGI2DJRpfd3R
zCt91GN2JM15iMkAqygkD1HGBWufnH4LOJPr+K5hIXQFlxUrMM0AUtyQnArCQAPrXsP8hkLdNG7j
Rnqw8UhKSgC+5tc/UJJvNR6B/iYlGT/YRDfdskQAhErKS39/nYCMQUd/xXEljbnP9wdcNKdQ9CzA
cz/hSRTO+wXMSitFr0FpEAWM+JHspgr0VtqHQhFIVDJ+rrq+mCXrmVisXNQmISDu2nL5Jnc9/G61
+EUDaGnqRrUqdW6DLN14wffnJoFb6cCaZBdRplgWe/PrmTUNa5Xrac+PyEb0yRiYprDmahWRDEhO
pWDCsqCtSJWT6bpbWn1E4HmR+EOcxy+GpS6js9tAZTCAggYnkYitxn8VxF8F1ugSwnJAwh9dNjFw
6oPk2HijkK4ob6GqYYhCHW4n3TEPd+3L9SzR/D+FUEGF0/UKhREZoMk3FSmt/VuMpFKS31AnKmvS
bVWiYhrenCyOlsBzr1abO4TnciiBFy14Q8Jt+Kp6afdp+x0Q5SN8zr24Glmh2MubW3evRmEY9YFF
z06puORARqKqNwXpNVCi6GP+sUMvYwix9F4Q/UtkkeCNCq++6VTZQJDRJevUdb/CgaIAn+GvPa8U
mvxB8O8f+gYFC8PeBG+9T0sbD+DtkCAHS22H0GHk6ruz5Z6fpNQxU2QzKrgXkBUSBJOiC2GtS1Z8
6kFqR1KZ3vSdM3j9RVCnLXaZ2f55KgQA+h5qi1jiMx4R4w/m8z48bTt3pvOdkhlWukFz9Diac9Tb
yJQxQNQOoq7icOkLA1WiZl2bh34Yy70SEO8zpSIVVt0cGpsrPZ6ebeRx+dsGp3pirS58jOlJ9gE7
FZqk8RMPRWTjfzuhEMkIgRIDTLsP5yveIVLd37G0omwbiOStU/OUoWc3CYkj5IfBrnT7SeP+5cem
it7NC+oDGkT8OkvQGC7ha8uWAqPxxVkimwyHSLwk289ECpSlBtZXKX4EllZAG4iHlwumVCF7nH/t
l2dpZaaRcMa6efYnfIUn9xOukaRlfnvR4QSIIgWerQwiXFfy9imCjsErq8IWO9+Vb1JA4CauN2a1
lCY/AVarBCcR1Q67cJlPkyKjpGCCsxEPfhuB4leE+sR6Vb+1kKvVQ/MuGnhZssfwt2YO7plxLjCW
bTwlnTBfGsnBK3UF8YPpKgjy0f+v/lY8v+6QMBVbjWICmWjxzvp7wK01QRQ/+sezRjXQ02MLM74H
Y1ScZZBv8nW2e6ztFNiJJK9xw7mWpI17UxGsHf1CB4Xp4OG6SzS8BJyhBJ1j1nuRfENF5vplVN5m
Y5aD1mDHXniATBtZGKRm5uP651JoCXY7h+MVSavT2A3Ov7xk2d+2fNPAupPkoKH9CyCPY4LxTl+g
arTmpm+fTuBGf5GXDFWLbMD0sjRV3YY8l+HiC8qsIutDF6h3JoXaJfXYbo0Gj8xR2jntdYS+Fg+x
08CQaJaTQYjguYtjmvBAw9XnwuRXfiO/cIKK1jeR0bqqzLbCPDypR2sqJ7bsZFhc+WP6E4AitSAG
v0Rw0SHwbD8P3PSSRByMF3Mwd5zgZwsLJnM5sq1tJuncKryN0FI3zcy67Efrx5NMi2Rhrnlw62UK
yr7OeGmTeF2gUQ88+yr/X5ZhiZZKyUygMmx0LWpk/ZVZR/JwXijoYd68bxlwC9OMrPg6ROEe83On
aWZht7JSXKpLkDrg1ywR6jgzuVt0TwQbaxFs+JuZhngMWsLkvz5VpgW1yUpkAJMBO+DxLEp1P29r
bLK5Yb76MBdTguYeSCnFdgI8SVaebjw2r5Nq4PXCo5PyFdmLgCuzlLxBQy4M5/PGI4PEOWfAM/db
YG2bXyDSbDv1m7vwZ6GPMAmL306sdwG0WqKOt4x3ELZ1MTQKAXgtEnqHzGvsiYTxwzH+bVy/+3rq
2zH4ll2/vTCXpeIVF+MpfMnvV2R5z8p1j1sC7A46uhDUoMCzpBd7S7KhNZ9RSmc59ZYD9L7nu9ZF
QcRv/mIYV4XIv2GxQwN86gvltTPn9qI/JwH+MNU8OfzdAV7xOaignrPFoMlS+i1n19tT1X0ITF8p
gTSuRgnS44ezygTX3KPyw7YI4BcGf39zyDCCIAeaIZj5twCY8i2IL2JRqccRYRIIsu23A52mAtHE
a/BwBP9oimuwS6zzj0C9RtvyShDvbMZEOF35KwMJeNJ++rOPVJz0dcccEi/WlIJCSWVR8EGQ7eTq
LS38QSu5/uaXmhUWR+o9e2oXPpsSYYe0adxSKqKhzADIcyWuxbBtzwzNqJaK0xtqftk2Vm4YRiSX
MRQ+3qkoDsH5zbntzLokljk07IUhDWpl/lyQBGNAMW5ExoycGt+CkhXDyY3ve+BZPOMkPf9er7L1
OInWXfwsOwcd3nS0jYKZZx158EA0xs4JJjbUosVOHsZV1jBx2m2AGz56fyTDUrcTdQWACF7AC6iu
/U6dVgR1biu8BP+iTqgzGG0zPLbldZDLgeAIdoMiRrKCx4MnVo/UlJTZAFfE9JFQjdr95gSWJ1w2
TdyeHGid4Cwaj6+TJTLoYR721Zwnmtjo78vvqAFzd8NB/cKbtxe2ScYIOHxgH2+Nd/YxjS449dYJ
7ZUFmxOivQboiSDUOaZh5uylEDKy0fq/vjgFIV4GEVxAGIu60frwnnm6I8DZlkFEybueOEDlfXiV
3QEuHI2PlzFoApTP50rt8K7DE4O78qCUhDv4Wn8qG/OHoSO0UfutA+a02A05fLWId6CMizVjFUiq
f8PzDoBjcLsddybmD0M5JsZKD8QgKx8RWDE7OO5FJTD1V3UMF2rTQcDO6N6c6GNUEUai9X67Ugz7
se5pB5o8lAobOiGuSV57/DgGc8qYuv4YPsT1CY6wjiriL3UjBFlnxZh3PsWdpjCmLEQ2OZfPYmmK
4P6cEyiYfLpyBRTQHxA7CqnVYDJ+j23DFUWWMwTu17tc5tCsV3Xx6STKhxGGEIp5d7TGeJ0quzwo
xnKACL5kF222QK0OKuMe46ayqnliK7FDn3DgYHqAkMOI1lqaKQ4pM8/U2oxf0EsZaCYqnsQ5ppJQ
9QRAHWZApcXFivPz+Q+kks+bUH7UOGru4JfZAiYxhStAuC4p89nCviMWhZ4LSG4+8wnzpfrkaa21
brfk2xpTAmn5nGGovqfq8ysjc0ovl71K5KVoq6IRp5WXGehDDqt0lunqtBx4hvVPXo7B8dHGV+wV
+f9bp/5fyRAG5mQDtYjXqr8j+kJAlNPAMC/n0pss9f/ssc1eTBBwtkQL8hpr8aFUe4Vw0qOouCjZ
xqKjZ1fo64O6ADm4C42vgc+61R8lf133Xh9pd7FmtAt7bY+i1SoeUjDWWWdj8S8W4ioqEizEnYH8
WgRV35iktEAuXtGytm2DlPuXkwVA514IMqxxBKmy4InYTFoYhdexxIIgRSo30p7GN2jgKhgG9Z1T
rgzO15eXO0Yqybz90nQdZ8DV20mtILPkbFxAIAD7vL5upEduzCOXBUOrLb73tIiINQULFShksVlQ
kswHYmc7IwSXNwaGNegEbie9Mz5YpLq84Pl0ZyHZV+atMS5DFuk6kYEHGkCwsSoCyCisKwjpB5AA
2CafyVz3NQj3icilgfUpafOH5fHi5bGwQXgdy8tGW0P1KkHu0R5cuEdcJPgBYjXJ4fOn5kDlMU6B
r6qLyD5+/bz32bQSl22aqQPk9Tt+F8qWRrZQassZGsTbGY1iwDO8E6K6hUkqObStsfLzeqNNpr2b
e21qZ/5/3ucULSbG8qqkwhh1RQIQEN3/WRRoBDk8B2E/LR3HxvXThbukCowKlqD8RbFzl0LmV3w1
LWYsNJ5Qe2WPOw5lbSiYwSzDEhj4mIl/WvNTH9OXWARDhioqdcu+YUNlcIcI5m7fF3z9UQQNaVJ9
wXTZ2pUhhpV1VZXKW7WJCcf9OSNtbZjkxxa4khJoRv+dzJLHPZqWDAYW5dwVNc8JnZuuglEa1FQs
Qf9o/tvo51oPkZTfIGHcw1pQCchw1cgDMucGDeRb5JYjKiGW5joM5zSmPsSAPxQDjp+J/J20rJq1
bAORWuj1UP5jkvxOg5TRxAb82pXXUOmrO5TbaN+CDYJUg7tStuZy96HphH8OOqT3BkV4aY7eOUwR
zXbhf/wSf5/Yu6oQFv0yXtXmmFY2IhqGpFfHMaO+36ipBzew98LLuvIzRz+M+rmtXHKlR3wFcC2W
4g8FGy0Wnd1n9Qp/Yq7YqDEqUSq9cH3s7Gh0UuqCwVpfJV1ViRvOo8Y0NlN5lR1hd8EZyRAiiD8s
DHrrhOOXrVYZOPydPM+T473aXz1HSpZkK+MOGBlYxBDSV3V1oB0Mrs84qAHbDqYQh7x0sc/YDjm3
aS40afjZ8Wx40ORv1fSp5YpGF5ohM2tpp2ujHjs1VVtovoZn7aBv8wFwlg7Bh3co8AEKWAf1UEi+
mcxoUPBE0o5Ar17tnpb/RCMnr8dM5jVuUowS+OWtjxgTvj3otKNbUIMUDDkz4nqm9rBv6tPSJ6Oc
VBY7dEIXHmujmp+Gj1XUAp0bKawhpButdV8CIk5OvubrVZLd8j/JUB1ERB5xhRWq1CRqiEcbqpWe
vpGmU/VcknNSpa45LDAYxBPcqDvqZmgGeuKrhhawyCoZT8B+6752+J1UMSeVjb4Areejti9XcGe/
2fv/Zhh0i9ZOmBxOowlFDCStaacM1I1crj0LfsWCX81wOJ8Rdn/4v3By39saDsR/gOHsxk3D8T6t
ERQ6Nsz+bbg5cSm4cWo5xgGPG4M/ve89VCaTxhNKsYBmuSU/+oM+gxVef4etdKavoCY/QmbG6vLE
rDwvKOB99JEekM8y/UBOKq7xmM/oRakPg8Dovlah1OmBJXJadU2DpPcfV8Uc2dXD5phfVLIyfcL7
IYh/R2eS/Ss0IWav3pmjDDvOw4coaT9FGqw6vxSVlzcX9vtyoAU1jmKoRqvMt/eU3fV3DVf9HQJ1
tZdoVPlIZGsh9dsyybIOikJKjsqcJ5CoD/DA8k/oRm3y9/2G4+1DyzmIOR5Rj5F5YcnBZ5NwxI5g
g/QlG9sFpaNYckA1Vy2MKC62pZiQFthRhE/InQXZVPLngdKjEDWSj5F+FzCgeChVwtIpQnUAulZQ
0KCJazKKqQmsCKiABQZFdx1I4gh7IxQ1FSSJyZnubCKifJyw5lNTd6yB7U4ZqgFT090KENQyOII/
YIPdnPW5F4NQMt70pAgKarlPYXAdsTgUpiV+15BgwbASkS+trhOZTW+fvC6WDvZ1jtB8F13vEfsS
uG2P0f3OYPDXu0V2WsuOhfblw3WsVluqCGRXUdZ7QhBsctkD2+pDnS9iDPtGRl6ulKvSpo+cYbX7
T2YYjnC2VqW365eORhFBfm1neUf832W4lF5l7YErdTm2v8h+v9thl33tEeyLYW6ZJYHX8n7NaX6C
Hm03kQAOvr48az+Ajpvji5tZi0iHHN5t6lE2ELKtd8LqYJtBOE+Ke2Q71TtfwXm6+R/bdpQPJnZ2
YN+MvAOGwJunIp6I8xdIahkX2yXakZiOJ52jLv6839RgJkKY2Yl+sSyb39S+0CFc0XqHaUsJasNQ
h9Ay4+ofEk9E0pSunrijAikd5hl/P4fyOWVQJU+lA2dvhVXkPt6q6rXW8ueBJyCm5EbkFBBTZp0O
3zFf/nRK2dQrd9MnpRsae7wNydbXy3c/MLiSzu0XYMPl8Z7E5Sc9FsNrYl7IdB2RIPDjeYS+2X5X
XvdS1g8zvnr7/qJ1FGuM244lQJDUct+EqzVsfkoZVmRFJ2N64qvER6Nw95aUqoZJ9yDQfc6tJrEn
tn09dEBeLyCF8Cz96rrdEheKqQWDO3+MZ8c44P+6ukk+PpeY0kZcsry7qE7RQAJHMzkphixRss5A
wPvBz3hPOvwJEPlaWi2nGId5kInCAguMIE6/+Y+MtB1tbs9Sw7uRVcoQZtEZl/FIQvActS6/ClP2
wdI5UQ6HoDNLOayLJfN2DJNAxamdpIPGw7nN9L1JdcOYKdS7kx42Rh56MT0da+yQ08j4SiyxC593
3nM6RWqwSK9DdE3WwoTzVMjhtpgaPLGjRbrv60VD7E5NKt+5DwX8zQqwhO5oC+j96B8vV+lSNxyO
F80WAraD7tMU0VlXEEAzD3/7kegr/4ejChR+CwDM6Fy1uPkVulnFfCVEFaffMZO2r0nqgnfunKXu
5FLFYObbPd8UBU7H4AriX6uFOmwPkZAzexgh+vkeXFVB3YmqIkP11wn5+UdpjdpjQNp1PhRm7ox0
J2Rjcymp1d+/11ELC5bVUQUEYNPxhT8H6mbXcFmDXrlBQRuF4v7yFXmA8n8C0IraRlqTQzw8vWSu
We1u6Ix4k+DYeOZo+2lCr6+uAJwK1wKggPaWfmqgjZ72NlBVXG81KPjf61a9DRG7jiO10wolYfYj
PUOarQcNVnZZh35xzBOjdZ7XXfGKsaNweSC2s9lKqzJ4U5pars7YU5zD9zQuwQNECTAr3jotpJqV
D2i/PWdCUx/IPe8XwKBdXSk73TZGcg7pBBUla34NI53Mf6l0guFCxQdHu71hfHqLIsKqjiVHOUTn
mbDpsPqJ3ROjQ1e6m5fxsDs2Kj5GVXI8J5xP3CVGC9u6XCxgl+VLfC5U3VK0Q6EYXvdhP5tDntIP
/rrQ2FHBhYOfRMlbyF5idOzo2JeXloo4n6ga/i4+s8ZN76oDYnd4JZazDylEQqj/FMrY25+u2Fz6
wPS9u2BCdmYdYie7ihDWB2HCOFSIxoKs8lAIh0AkS33T+boJnndJNXIoS6ICw4FTu7doz4M+37ZI
/wYX1zuOfXr7i4Jr+eoqT3uruhX7WQ/dzIFVLBrBPuwWg3/wBqghw6wwkEKOwz9KALarnT6WcHHi
xwGcAczeSk6PtdEwGxDrqDDd1AynbpD5ebOn+aM0zaeNkA4aKsuZDPerbh1CBT23DnlZDPU/fK22
/uSzN6PjB6hOwzFwB6ZXQVXSCNv5oJjKLHRdiHa6bbuOS+Z2P273thUBcjx6o/l+wnJQ4rdrgsme
8eVW4swWyJmsW4lUag0lzPt/vWVn8gbn0cYhJQHSMN+LzhLG1GVVBp8nVLfqlbGVdXX5Up7LICfX
PWscmFVQUnnryHibEDbjpNi75xImV9/69vBr2D9/m8tCTKhnvIdzuQwbtTQkul0yL0JLmjLOp+eN
hqVaj9k5/ni3cH3NId+Ud2SsYqeyu1SQPHGlxIMStdkfAIr+6rggmWtNBNjE8vMO/l8163FHBnLs
sHJutALf0jdu20A5HpFn4nmnfrYAjKYKojLpKrrJfNYZvH78wm7ZIkHc354VNSRuMTT7yst/t1HZ
hhrMU8AxVLVAYDSeunIsoX8YvVaAuDiaFebixdaBlesgWdHjyz0mo0Gil3JZ0DwEcuWelSi4xoNI
Gg2iFZ7gyDJzJmU3EvoagnpaGJNE4Hc+KglMV1+jDAPD50LLbsAQmQMdZZM+vnxzVT475r4tZ25B
BakK0XYLSjNw4law0Ajv5QRxaQshblbPUA5u3zKGLRgkwn/onqTKNFCxvE3tDecN5pwl+XMnz21s
gucWCIz5cTj0eRVKeOtrYljgUha8zGrw5J9xRbAWs2QzBqL68a8nqE6k30NaQWvFaZD+bAoAfkYc
oUHoPpmxj7hTGxTzM/CDaNH/iH0qnQXPVz/svKkoaadWn/8aA2m5HjIyFmpX8VXHSnLJhJ+9TKQy
oGSMYoSe22KqU75vVJJdG9dwPnV752dt5br08kzdsHOX/Dfpsg9No0s/KTodnn/mTxzNkBtgvzmm
YFyvWe0d7Teo5eOjLEs80Il6MFTIvdS7yiSzDHGMnJPoBUrmEnbe4G+Ryq+dbIELTfKELv+T5h6E
dFb34+Mv0VTVMN7CUvzBRBugxC2gfP9Kt4pLsGGVI+INJv6rjNnfy6aKpIB+LlMJPJnxKWO2r7PX
P8FqVNiI8zFhZnU+GH98LX3u8imFDC67qbuygaHYfPQlr+gx8GW5+rQryBVw/+NJLlFFY22kndmQ
5R+oJE8IOo6fa2QbHq6qBo7vdIGw3FCwKKlRSXxvrZTjitzgxlGqUDwVL2ns1jX9nT+iTf9BGN3q
aHRzlPlu1S3W5K+pF1p42TrKFAdNmlTlyEzJTWaEzmnUS65thXUCjiT9BxT2AZMJ6YdyO+coi4uw
xrOsb3SDPdPcen02uYf0b1YODAchJzGZZ3kbxp4wYvvm0rHJpBhzc2ybic1ctgidsGYeb36C6fGU
ZF0XFQ98W+knC4SF2jnRpjSNWAMk4IiMj1ziuHiaPcFprgAGIVfK93cdIkzFUtHvMD4sc6X9Rnub
K5t9BQjsNZpBZ40TKhZOZUP6WNJICAolynjBtS3JF+MAqKbR7BYrvGxityV2t4Z8Go3rSYXr1vtx
tObvVhY7axdD8W/Din+mgRG3E/TunVkF2QVP4FfR4MSUpS9aILrYhhu3agkEpQcDrSDnURPW+wNI
KUgnkSBi3yjWQ84J/T3I6s3ztbVWyfMLQNLNG/2x2dHnQUWpYSfpBzAx54tjOQ+QvI2QxCk4ytUW
gyHToNd0GslibetY1WOiX2KKAwrojO01WWrgqfKS1YQQsJGmIwAmR//TP3GNnS5ARn3/kOWPedwJ
Au7IHxB3W4eE7K0p+4xUmemIKHDyLDZ1BsoQZZLsPfaMdqjyS0MfdSZlzRfLEqy1cczJP0PLmozN
bJ3gFb4rMH3WQxaKjFT68LDA2Ue3wI4e4HQAv6Ksby29hDz5RMI1QNpfS8wqLTJkwAAWjTWlEn3U
yw41T5WYGQrF7VApVOGuR+4h6sqQXW0FvGk4dV3Ph0rdJa4mkIMwE2SNW/+u4zlS7GoC5WkkWLcT
Gbq44mnNKXbQBSDpQdhAWNWFXHw2JnbqyWh+WlHqmYuMoAYEPlL4B+e5PxteZUOmbXOIdY0lfGVU
GehY1PhaRd5JcGLTDwFo78Oxn6VXVjTpTvjE8T8NPcII4tmcxRP7q8U7Sm16s3R0fIzr5+kggZYp
KdI8WMZjHKnLe0kU0MK6g/+iC0n0WncSrtyndYQGN42hO5JELoKtS5s3JgOQyD07vlAg+9eUUtys
vLwJB5lTiwBrYzoo1foghSWhEksGSow1K7XPbB/KB750Rx8OS9V0/6wJOwP7pNkxLKKzGaKOV8gp
U1PVGlh+yMLyCsx+WGCJyeahfaTbEuZ2VQosPLHrA/Ge9G5LosKu0FWFChc45XVwAgbZw8Nk/56v
cAye7VFEYRTrWfr0nhnMNRwrCHnBKTwGl+FVNVuVUInFDINtua0xle7Ki8NNymON86PcpaPxiRkL
+ioYC4XY7uqMyD+6K4pt9LUtktiulEMVNzoqqqakGNx9EZvGb/aC5W4XXpbXvnIBESIPGBxr8ID5
g0yE/JIL/+S1VD78t9F/QFrIqvgDaRecBYbWlQ1b/3UWxJIg2bvEiUJgxPIoVbmjPrUsod5eFKNy
SNJgJ1o619BdVXsGMnBBvGWASSonYiBRujY95x5I9IZ97feYTz4N9RDJJtcRrPBI5c8x/X2jOfxj
irRCygOY4MVYY7L6pP0cwHfky6OP3Ax4EeHlKucwy7qJtRJ7pYyVRIuApw9UKJ7dC+VITOOaT5au
FiGBg5cpcMpPGCdpQ6fmoMAk1lfuqLk/Vv6vBE7t8Kk+i8uu0EdxBxpCXar7NoBEerPZt83+kUVS
niU5IQP9AXHE95B9vcq0+0ynvPcTU3KkyxY6QNrYRM6YVBJ5KulvClBY/Uq33Q+wcWnbfZqZHeCv
uiOqAOZ2osncwIeTHwfQ+G5CBhLTpHkCMhZaXQ3TQYehBi6G4Q0vCxgAnK7lw0IRxMi7s82STE3V
TzyIqE5xffJK4KH61EDYCS1PKx/B1S6TbxoW0x7kqHYiigMzri1eEJnl1r62OehhJKJVAQ3Dz1Zs
GLj8nFFmXXcvha6ywpbG8A5PRJchyIalbgTJGU7xJA1D6aAGpMihfyTfbRK9frskdDJqi0GGgwBf
FkkYwFFJJvMBETQXguZlG2U5imax3URTY26bbfvI0YSqy7ZiArklslTpwRkxMlK+uPDRLe4LYMKl
SHwrKY0BmpHXRxTTk8JLlgJJI3dPa2RwF7JM8Q4vHIHaHYl+aB8YViMoUe5XAmlqR9GkcZCSzCY4
uz1P69Jayf8g9T+z6xUlnhvbGgPtR7Swt4Sknmqf360caNMHxXg8NGeexoc3AoKwOsqALyL20sG3
BPX9E2gzhzweviLsaH5OnrDuacXUnkENKxgqhaDNeSFrbms3W7IfnkSO4Wkrw2MfNMqHxBDWveN2
M4c/1OZJ5RPTjZOb1LS7FHhTdE6P4aBYu/LNwaDhF8E/B1S8KMtqYoCXAGBVYJgDcf0sNJwMwU0y
UR3SMvF4EiKcMpQ7x2kgepV4PRwL9N9DvE5Tk0jPudAJ2Fsz7gwb6TrTh89RRtvHIcQokTwsPCcE
g688qafEIYFs9DG/HFH6gnvVfsb0K+c1jDYg4T5cMKeNUNSTKMl8Jr7sEcgG263/0l2kprt8n/VJ
1B+PwyF0LLr6wPA37B1KPKA120vRyty9tcrKsZoDaXkStJ7pqODwmKEhGivrM6YEUAIjMXyMfXTV
v73QqaRGtmo0pGQ1+bc3WgMLQAvb/kryjyJDJmtDZ2UFOrtFCb9blFF4paO+Jym3kp4NJs1wvkMY
6gweYkvkJxCKPXOC/W8PHNzt74yJsYDHdVHfwW/4o/DnTmy8v+rU7PP44Klirl0HXDzUOQolJEAo
CIoGfdBDFb34SVdgi7iCGeTqke5w3EjzE9ciDO9Stx5sDIFGL6rU7VSRmARWvJ5lujZ7vVRscTDY
B+5l6U/eUvQ4bWKONNvhBl+TnUEdZxWydswn2jXG7AP4PrSShSLVQzJPTTJvRujZ3PNeE1H6PiyG
9jJeK0G54p0VEYkNp4ZKDmVMjQ50fLSO1jKIXOyd05iIj+nPOyTSQCc/p1JPsdi5NwVplXIKr+E6
M8lLH/qKd+m3Ou0JIE8I5fsKf6BJzrPXW5f0iSan+HYYpAl4cQj0Da+WGx/S1/66Xvv8S5uAlP+j
0LYscz5HMvafaetsg3GKrxSe6s8lED+vp6agPZmoueUt4pVuixwsTm8ds3Bi8a3SixRbtS+pZjrF
TajkRWEc1XhsKDrDDnYGSuyfzGWy/g07bKESlfh1UV1rxEOHIagd/BIaXXJP1tRHgh29br+t0nnh
3tG7j6QY86Ztv5rASEiIBPMxqsKf41sdhLYuDW5Zox3fkgnTQD6bvdC2wWOAwmj02I43sVprXf9n
hn5Py2Rmj16qNNJJ/81Dw+I3JYaBpxDa9P32oxNl+g7OsYFaZuKwUNx/FHwVfqbjgc2jTfkndTOc
4JVowkWIg+OVh+o7/Wq+Zd28gaULRjv90e6sHBYVK2Hi3x7npSYcrfPBa8ieeqrgLVeVknNFnLBL
RajkA9q9z9+U11k4ROkyuQ6JJ0uSAsI9BA8O88Mt1M3NZUxnmlNLzUlOzf+vVyofLgI4VujfcOT7
vzr3VkLTA7/oElSDmFP9Tl9De6RZ1D7BklpQp7MB11tClqz/vtUKWcbSSgz/VR5EBlzXcDtCSqk+
K0fOqeVi6mvqw5hapIM8Ps0VUaUEp3x7AESWQPLfk7QeTU1Xib6S4fqt5FuDWA2gy8CwRaOAsC2a
jHpUWd/geEytd1P/zEQ3olT8j9I1jm9QWXriAwfCVYYxnkgt/FnGbEW2vR2lQQcFUhHbaFdUB0wX
D/5JO7MT73PBNN5+bBr7lGCxz2g9qknCdRtxfiv6BT1ynHwB/6AFwJAzN0ZIRV+F4ivFeYj6ok7G
ULrauQvLR3cVut77xsM1Xchra0ZvRpIuchzq/F/UhODyXzIlTp14JEKQ/0i9yyRZGdM9XZVk3nFH
EvG51biiItMwZaEqoOfnMJA5Byv51tdhs1tAiCxFXE9CHdzyJ4KgeKmpZHeS1gEz4TaxP3osDaXe
whWKA5bfklHYFFAZa8iklJLIjBYhZRATlHQxlZ4uRP9cIIjUnlWS+5aN33n/NE4ytRkZcsg97xfg
kuxE5sh282AqR6XX4eDR37mA23jOXGGoRas0RZ2SbkbF2ikNhs1ZH02D6NMnOivv8Fa40XvstXR6
cabm/3voBbw/ok4+K2bFcI6wJH9el4y46aOh76wDYx6enwBRk82MyK+tOB3TewaYZd58vM5P99Vk
DIw96YsunwGt6enIwB5R0BPSE2ZwP91kNm0Xlqi4L56o3B6i/N/wtzOL1bNjrK6fvT/d9I6xlSSu
cPbVC86lKzSL3Oi9jYG2iVKGP0AFHwOKDpe0yKHl3o/r/kK1dINCdktu10liKa1z9SQ+9m2rpqGu
Wxg0gOMPz6qNpeN6Zg3ckl2k2dARkeU59EAUSPkE+H8K1jMC9M7/EG2HSgtUuCLeYWPPvKzRSM78
ZK+7Vwb22eslrsnVbRINK4eqbp6LlapEE+BUZZ/nmBpWqFPYzWK/gsbQ3xxC96CmbT07FtXTn0Fl
G2y2qPbaMZP9OLXNteXWM9hfsz4bA+Bf3FMW3QxhI9F2vcWucphM6Izb3Ie/Du1Hx/0BQm9+wxWL
S+kt7E6Eqs5zaThkYZBUjYpmJJIOYlWlc8aGV+MAnYyAaw0U99QDGaO6rL6K1qsfrNSj+kM6W5uy
tWMXRdd802gpAAVim/mIbjnroLEZnrsFmrDe00W+3cDu/nxUeFfD+Zns3fVMRouNFCUlo7JhUj9H
ovo2iBN3D9YEGBTgIFSBINHP9NUJooVtTSKw81GfK6/NV2eUzv4nIazHGrU20/Z+sUbFlM1kMVO/
6SlMy2pnBgAHgDshAAzGyRzz/rFFJz9sGuWG6IW/1rer6q65ssm25UDz/h73pZwd0CUeXCFddn5W
ZxmCgRBSLF0MEnBz758LmPIrjvEOTRfGFORFQDavBaOpGQUEP829lJ1NcaLUd537AmKqlawBx2AX
VtlikbOveCCtTps7QasyDjpNvURSzBrhtlgDorqOj1hCHzxl298EuV4cbWDDTz5NSsBcS5hT8TUM
oxbwCy0Ckmsk92j4JucP995Rxt25f0VSDi/g6cbP7/Y8QVvQUCHC/J5YxnG9inwDpBvI9hGfhB9B
NIhhS5qMjNNXITfEL0lCpyA2wvoIlHwy+HeZtTyImyeWz12FNcRE32UP/3HsF5MNvkr2RrUVjHbE
VlNiIRUtvev6dZvWoe5J1+X1Jc/FhgyPqsByN/hSmbn3Yf9VS/CwO1US3IJOzfFNl62MxdzvwZAR
llJ7tpirirP2bFlan7Q6ZaQH3PQkC97CJ29bq5NcnwCLPw+QqmBUviV938dg6yhZpP1cRroaBFn1
TSTdT1BjnOTGnQrGDIEApm8qkmlIMIW5dmZaILodMOwsU2/W0UsiassTD4ua5g1uGdOnVBTngBHS
AfpVw0Er0z7P6eTVMYTilB21FGzIBtatwFNUVL2F1He+jxLAKGgv86X9POhEOfOKZ9bPKAhW6CLZ
ULFatMEIRc6LD4G1XFZSTk6IODfrDC4CbOJP+ribGRpblCm6B/lguZo5cG33vx65Xgg+9f0Jp4q8
w+pDbe63jG1Zhvrc7YzurF24J3Qn6yAvEDY0M85iVP4e1QznbmXRb10XQ/st/sQJbfTUUyTLJI9z
lT51NLHKk2T+2AWgdUXDtE7BZOiYPv9VeVBE1tBc/qMtRXwxNKDETf7jqxfRAKaJ7ZGGdMSsLjxW
BPMoqx+VcyvMqBMrgdPGuoRM+76diriqFsn7mgz7OfCd40cjfbAVGHr80NOS1pqno4GANnDqQsMK
LODifkaqv2pS14iYAxwsDFw9MroMP8CcortHvz0MyuZzTEJ4uJgEj5irsDd0yZ7M2Eeeub4HduxQ
+A8tUEkrKniQUXJo7esNmazClHazZk9OuQsHjFDxEyDXDt6XreN42oF/9PGCFzd6meZtorrDcxfI
Tcv51AA4bb3DMYFEi4cderytrRaToo67FR9QLe7hwE8husu5se2Bbb/1o2MLS2saq+gIX16ZylNm
g1clYfziFogs8EG2WElYkJCU3ih1X6C/wCFMupGae41taDGR5TJG0bnXH2jOgGwui65xX37sOtv9
5+99GM3rdbrrFdlbncyNaqx34u4g380DqBBmKsYXMEL/sSn+7ORFFx4G6J69z+KzkwxaeMOE7YSz
Bf8tzsceCvu/8VaPvOgYgSc4PwuW3KBHE/3aFJI66g4kKaaluF+M4UtMELwViaOYVbcoZmdlh5kX
tOIaCRXmPUfekFhv+zAmKgECBv8VvlZkRD3BJ35IDX1aRcbh8Y08aXANj1z2vH6HnGpgUz/Njuv7
J8mFRCU7OGz8EgekxdSsF5li4ILQxuarUqWlg+kOsI6OtJemPLtLBaaJPhuiFs2/gw0M94ULTxzY
k0hYOMtXZeSWS+TXF4QJY7Jp6pX7PcH925XZCnX7f9/CmZ/prmi5KTd3pntbE/IpcVwVWGZS3UYh
MxGSjYAG9yuFgW4bl0AkGY7QNvocSEAL1GtOnS/XvM8UK+UfUtK/FBRBdUlJQrB+NEnZk/9E+y09
S6mUOdLjv9Xi//dfnFWTXJX9gcssoDF6QuAaGYHQnpMLmJYg5fghVdU3WlrHqoRq/MzwJaE7/lpG
453M9qfwsrXE+OxQw02YLxHKw6Jd4YNtVyJ09GzLqJtc3y7r9fKsgfAPqnUIP8CDnTmo8HxhhA4W
Yh4TL3tA6L9VbgzFt0mkrIXrLn0sqdZWPXp3qxQiFhToznt+hiuzmC1eBEkGmmgPTA4ZDO9dwD/i
BMEtJEsxe+REZgF+uXz64dZr+Was+FuHtmUx2h+Kr9ksMvl9RXrUKYzOAjlnGx0RjhfoYT9hUa//
Up70qFWeAn6+8GaRYXkELFqAo0jtC0xPfjW96ASHnyLoqBjIW7WMGbi/x6PNTefPrb9P9NnvGEs3
nWYz9RCvEF9tLxj+48r/wppobVUk+wRIUBQiMkaqxaiNXNmUCZjkVuxVsaUkEJP/ehV5gFI0y9qW
2Ty32rPptWm1qh9ig1T/665XcfYLH6romnlLF3uYyhrfQmHoUzJBjxgAJAGSLSwNRvy/cW6wzq/G
IWrCUvlqcEjk4nu680BQ/f74a1WJKaVRAj3Xe7fvUSGzWw5hFXw1allYPNY0qB0YyByyBWbLe3SD
Z7OmR+FCL5LTCvnD2kFt9XmXq3agY6vauSj81Gfr6lHeNxb6Wm+6t4C/n5cpLJZ7ZKU46fzXKk1D
o+St4IiY7N+UiA+q2crpK6cpf1hkzUxNR/4gJKNjgHWk0NSSgF2pZHF3FkHd+FwAFGuQ/JqJi+m6
Ea+qqifuOx5FiJwRJiSCpWcDormw9PJH3xgtTCF95VHEQdr5W/c/eDsUwyxrCQk0VvMtnqY4T2Df
kf4AJORdorjizhITiP/duYzR5gSWwcZSW6lc0oGxyScwNmKeVdByxZM8T9/X37x3PU1ShZIsWb9T
TJxGDCnKsJ9x5Vio+QGJ9wzJt88GQ6kO/3b8dKCCiRjosCEG06ZBuHIZ5sXe9ILxmKlPmUkW6MN6
pDEOyML7dnz4hYZkySyaXv5JRJURyGlyJeePKgeGwzS02MXG9zmYK7MISTOf5o00A534Dh7EjiP6
OummkHFwTrD8WjtKkI41+oWSYrHygQcCuV1eSe6OC9gHCVgripb7L+RtOQdHUHzLKR3+JDOQ60Cp
58qc3tYGZ4uL5udHjwd3s12S+a8QI1f1tjN1mjCAAuDjoMM+NPzft/7XeNBlgGrj/NESrPZDpDig
UripW1jEHatHItet7AJu51m9K3ZUYGyltiX7LUuFAP6RayuJfOewmkHmW2wijPLByQIHFd+5Pc5E
Zl/Osj/gE6sXbrzvhpx4hn+glV12knjEk0tUm505XydQdMsUxm7Q9eOWvUoDNkiuhCQkWmlH6QkX
GgYXViS8lMWbWqRgqnX879q00P/05z06VQiZZqIbfua/7Krwn1aoHgq4Fo3GiPPQIgAU/o/2vblK
ScTNYFVpjpwe4N3AWk5tKUG2MjoLjSf7zRLo8nHKsxUDRhpeOgp+212ohQnpgEO2zs+av5LHy9qA
1XA/n1f2XwiCzHKulDAi++YpE9CuxRDxgjlWhZPMYv3wTmBkyTVdYxgD21x7iPKvYPJ0sV7hNLKj
QiV8Y/6wOHN3/PGQLf3iR54N4sRgZTor+AEdEXaIf2P7Vtv7lZ6YG/9lU5OCLaZVL7HGBC/vLImm
C2nFay6MU1AQBWgbX+xpdQbLU+g6NnZmqO+qm8b3FlAsIz5WQmJ+i6CL+9n8jYPQr9xqiconbQ8s
IiXO93Wtb2BXKHLEIhQzH/yd8ROsrOBmgrT4eI/WN4mwzlJxQozB0TjxdYiwAI40YjIfcW7RlHNz
CMt7QUWJo7GdoSUo1zbJ9ad5fPXXznmgYNk6fPynR+iTsZU8F4U9Yr5ub//8WvBWcwQKmrGqv2My
hOqPIIkRkkqShSbMzmz5etbEZca8rx84u/bcVKgqqqGi7GOGuEa9kZLoUvnmVF5E/isJYPDxPt8m
W9tVVzkew+yBMIX9svltEuR1Pcwea+ZwUnXnWazF4w0XNzkprHyPzaUrj9XIlPyOaJTRnEDdN7Zm
DrSJrkQCy7/fubC3aLW5QEx6z5zvJQzx2/b0vgBRLliRlgXRqM6kChgu5/vZMScD3gv/bsYwb5q1
JtLW3VghA97gFLqnDABT296SdxPeCgHr4h3drXtlr0Csk8zY/eQarlDee+49UFj0VRBbNs2F00ve
HatBjrvWeqrBYIJ4DOWamOnOPe+RbV9IhhBZ0gE0Wj6s2veI7X+qh98Vy1ETOmsVDBRU8fzOtbLf
ckfdNvKTZco5COqSkzyZ9DfymqxF821gwz57ApwvppXWoqrUZf3upULyte09kOk/22mgxhVfwj5Q
PYTAVU/XkoS95AmVnfoqudjxJhpez9e6npFpSkujDaeXfNSTjryGH6VzJuRtuU4+BeRaGQEnB/C0
lp+nY7mORNVB3cbw5R6u/gNZK0tTGayEzakyf7fGSOw6ZXEQkZZo+4gG2sWwDvRtgElcZwRJKXQQ
b66q0bVd/62nHSmQnQILS3AbwZtk1mM4ywY1pigZ8kgiQZO3yh597SGST8NA9aG1ZiyHdK7Knlb6
tcgKB4NwVNJCopZUOzmGpWqZk7CHA/McFzlOrDgRt/Zn4aSQb2+YTPG5eSJdxXDn1vNGQdeGHLJ7
AXaXD54HWq/sQla9E4w4Sluaz3tBSi1WtI8/QNQf3hv86/BCZ0xzz7vOUJL7ejo9P6uigyQYJyWc
fNYZF7g6WQa/qUwk2ZeXc2iJ8paH1a6rsMvfzxWIAv16q4KDkPXDfreG5DDhPLRkAQXo7/hCcQlV
KAgknem6osi1BXY5t3HaVBiLOpRpZofiCOe5+dSZrBCcHHny6iP+gxtmOgoIQ1Eix2XdKOeqS8Ak
Fs35QKKHyeMT30Om7cSSup86vZA0BmkSY0jfn/e0/Jsq3ACpd4qOO2Kj9Pbd7rmF2CiiqONq2Tz8
nCU9wrvutDj5ooB0vnC6BB/jvN/CvGLEHTYsu3pQeIvDTK2gK49tVqRYAB5biyb1LvdYoDUpAdiU
wdYEwtDnda3gTkANldBAju2Qh0M/i9U/xCOU4ecNpn+FqDaG5QuwvEkBp94Bu+YGQOlMXzMmqKoe
8aF2UWWoP1O29Pk0iFYTIHkss1A0sDNayGVDPpDz1fWcAb5X/NgGo7SO41ZXGPNpKOh9nktPsURV
AK34l80YX2k5GY1fbZ8P4ZnwFR7mxb1+SbgBbgX+rnEHi8yFAvejYKeTFh+RY4W6c5CBVtdr5P65
ruXh1Viuw3a3ROgG3kKIXL9caZsD87o2/0RJYZC8QNaxcFqCda162j0ANHWUyLWgcBZrjCg3M1Ps
O1UhUImMmeSNMIz1xEF8ltmWuhGDq2MmklduJHHYqTOeMs4/W+vDAQfgEeAomajsu0TKQIz4z2RN
yU1CWAE/a4XrTwdA7YLQ3ri1QlXspEBpBOB+P/Km1kaXjBch3Hh4ufT7QFBynpGpqvUeiYbLCil9
tO6whpikpSXk2Y5goC4j/VDMwi8hm8EltUFiw+SC5VW41CKrrqwsJpA7iQD8Xds1JOwab5cpLw3M
928BBlXZG/H9Yl+jQeZ1s3Yh/sd0ZwhAfnwgL0PN0j+yotGUIKWjG84Pp0b/sIXUEy7i/1UDYjYl
gCZ9MfoarWYKgGuFHb8b9nRqGFutYIWdpEgrNi3mpCtsIPR+2TrccyWKXpTV4nQhFGYq5Z4MHRsI
A2sgpGF01f+gcUNOG2H9tBB0s089w0QZrm4BsGXFLgpn+fJOXItEVCuBLVK7pux5/BE3n982S8OR
k1tZBOP0DecYQx+QvIPy1rPEnoRPwPx0OE1ZHGn2BxVoHYOTELk9B0fSjMwZDeErCYXtK0UANaK/
3YpoVAX4G4fYfCHserfhOpptahXEW+ahMgzKWvzkCCDyfeYp4tFDrLM8yIQR6RLsFuBuZurL1oO8
jEGhwsKcQsz0/xcqZ50DvPnZ7hwhRXeYwpiMbyC3+ZhweCpTH7sAQo93TgnfgeC1yrMacOCQDvoE
IGGTW9KYgWpoLLPLdGtSvx7FcrVl1DpOH68Jfkf4HP3pKXk3aP+IeNGifkiSwp8VJyOhLcalnKCE
/B0jc0PljgS5XUanB/oCaGrfx+dKkvFYPT7YdQO2y65YDqZ8oeJS4a6xLaW+ib33E2rjy+THfyFf
2jNw4K7Pvkdx2RD8Ce8gR6M4Vo69CKsjdEXEh/ub3yFddENWjA5K6q9W7uN8A2lmgRz4PSW6EAyv
RHbZeXfbI/ytGis4Ue2UcPr3XgohFc1bMMqwvs1OKnCzX5ZeJer+DOy0tAZLH0ySGrHxaqC2ldvv
w5XM6E0S6gp3GZeMCV9QG45hT6IV2GUvyxY3Ur+J59XbUFKHxOnLu2sPC8RrKZmwTLFnZCQoYddO
pIzEAChXd3z7FVRj1zf1K5uyPyTdpBTMgm1zZKvsh6ROaFbsdvEJKy47EfUziQQkv+9s69MKmU6/
/HLarWRUnzsqq8Ahbe7XmPwBIBz03i+QWi/ZQd6NZ9LroKFyhvQBRABdSzQX4OAFiskJkflHSkEP
1dGHdJGg67jaEpPfwCjwSHgNRI/qwzeXTEymVN09qgij0M0Wt78MpMEhndZEAzxsjH/JPY4Vay20
1vj5PimbNNKN6eXRDsHEQ7Szw4M3s3aSY0lB2N+yjEI71OhSp80RLyhWIgGh2a6bmujkAduQ8io2
2u6+iDRGgCzKBVcj5aOF1Fkj3xw3YKxJfktAhv6Yn2Nfn3clBpC4XDcjMVu2uz0Zpn/Ks8H7c8m3
M2zyIfuwp4cAcZAF7dLjaoSWlvJWsiGF6ZEUx1a0X2XkNDn34SoevXmSMlxa8SKjrgvbSwe5g/4q
Ux0+TRxFlKCXapFQC8ciLGba+qF6xKejDqLgtB9FBSENttyxJ29VjEhjsnwC9DHdDOJJz8BQVFQq
UqueQCGeB6Xcz1DTJ7hJAuDf+zFAHqyo3e+oMuT1QPGl/4htcSiANZhtXIbqYJUkVULRupSSpG2b
h2zwnWJyLcyAfSq+Aq6AAnFxRePgqSB0/jtTRilrqTv9/F1xLZTHQjJRfQoPoYK+nmchx5F1G0JX
e76E1LF4WSE6syNSxPLFwWykXN4zTcro1yuZG3EkQQ0alfaNgNOKv7Yw/VUtel6Li5bg0OC5GYAc
lMMKMBWgn75nzKEwzO/zYXqGQ2X7U5uYZbDIX2Uep+e04Q5cizjzGQ9kiCNXpfk/cLfC5crCryVP
5Ku9Q5xxIwifNKcw73Z/z0NuVWKgID+OT9q2qhk3ChXW0OLUEkBI0TeykC7xGzICYOcJWN9wTHH0
WAs1ccWRjI5zYrpgaM1wD7TY2sfRA7bQIoKqY1MXdP4OHmIWHPeVUHOJgkWQ6uDvyCS6waZMw/ri
S7veGi6c3a+XvgyLyDmYCfLQH6G+8e6gW0TLxGtXvy/pGSoAIrbefkSIZUjNsPC1apvxLR5+0erP
VDNz+ylf27mgTBkYT7oj+jFCP7ojTF8W42PE25RHDsCicdjge1Gc8HkKyfrcjL00CmT1QU86vr+5
YUU6nWvzzhXiCma4E/ZbpMmDQpMSGn7KWcWDg6uIQUFPN1G9lzsSUXr5yzaEQt+MW2vyPRyekVXG
jjhb+dg6NiuoCMhHDrWRh7CXR8jZXBrpprW0FN9DEFz1DMELFYEBDuetxH+xt7JWWqsklTOHSW/0
8aDO8kGByIHQOjrxzQ4yNMrtDc1J7n6Ps4BZF63fTJPxGPnlFhMNjVFdcte4HwYfWXaUiSkSFA3Q
YEdu08GpihNdKuPeBlmdgzaXuBaOSotO8Y4LWRxP+8ke5/6J/1gFK22GgDxgl7owlF2QGm1OY3DP
AvBlKwmLojBdSFjs5AyNOuvQT54ySqPeCZT+/AqFc3TWbN3kLnm8oPM9kdM4A6XubuAnPhzwkFvi
M060of64XTntyTW49hRr0x0H9QeoFk7AExdCkpZeqEg+9FO3atRHg4YAtarmO2BFiMGHvUGtBlWh
DWEnfRINreOr7ZcO7qtHzGiE2DYrJGSANVu+dQZVyp5/otHahyilB3SLHmkkxrSF+AgmzwJDNVKy
EnAkuQrbxEUShku3JE/K5vvgMJTHiCvprgNxRHEsLTMqkD04uh6hd5CHa5hbnmfRe5DQXej8TsDF
B9sfyCLSe70bkc+4Y7tjW9tommUU0eZ/McOOVkzoWYuEHzbShHPmg6WHCE3tKIA+za2qjrTqKfsC
M+QI6gHy0tPp55bX2bpturFdoUqj6heLAYsnpedimkuVX+E0rYH++m4ZKNa5uXm3QCKtdnsBFvCO
a2kz01mMKiDku89e0WN1/e+5BldY6eAWEsTCp8hGmnncZ4z5oC3oA/9XxuadIEF86O2vj0GYHiYq
ql8gHGvVUAu4xbCG6pEAFPoM/DOxTaFnAZU+804JkCKAKHcuEXcbcy9DvrvPqL/a6lR9TBymSfWp
vuqeWs5dxLRty8xw7yl91DA6sb9yJAPni1+LUSc45c/Ce00bAbTKixXXlBDtowAHyKaSWp3HPC5j
Z1vlkVr2QIz7q4Lzy+3KGxN1VEyjMR9QUxufCjbGrnDuZ1+zzSvP/wAIJlJsRolu+IKYOBXx4pWD
I/9+vtaILIuQTc0w8f1tdxjeaaQiDg/dnqR4v3Av6yDJ6uwsiuXuEfrfWHvp7crarrW9SzRzVvuZ
I3VHqaCOhiBKvwnVWCsDCe/34TrXWSBV0ibEMHYA9k32WDvxU2xmnxctOBoe+TUWtgYct2BKJX06
oL4kWJsc6ZnZc7odmemz6oyqxeIALX1J+YxqqdAdsznUVM7iZZrR6sRlG6VzmwcEPu8OIYyv6oMQ
aY2HEPMFEOmshD7Q33zoMfyS+nAddI+hMEhUC6vcaRE1tLk+DSy6Sr0OauwzOIeCZ7Bsdvy+tKgk
TsvTkkD715olefAsE3WcujY4PTPPvVghmXuOUAKeF8FhNb2Dwr/UtacXeAD22FBie1uT7Ev4dyQ5
FX25CXUpmdXEMZyvvPKQPFKBcSQnFn2xM5K7miEzCCME0BVAn0uQeb7s6kzPQBsFTkY6yyQf3gDn
s6GJprcVLWir4w9avXw3U6NBEq1L9nw0AYhfBg/qZhnvBUMkbzKBh31KBd7+In9i3uWhWfUgaaZM
svxBI+ie+uGYAXnjE56sEwsz3tKLjIfRZqAdRmKICmegnHlSj7QQ+3OTNbK9U+r4EM6wFRZIobHX
dByo06Ivi3sQW60eErN8f7UIjYvJjlSluT83QPKoSqUN+aR3m+xlZC+tEYdcTHp3kIU9JUTvXZ6s
9q9Lc5kl7yuOWBTkitoOp2vn0gYGU2iuBoltKnM/u5Ez5WDbGUAuDI+6mlqmTlQBuc+Q5dWD5Jw4
HFyXBDCofGs9X7pbxQwXvLzYl4OqeML5f6SwwJ5jvV8ha7JS14bNzKQfwaS0F3/Lx3chSRe1jL72
P6jxJB1E2toZB9eH8NvHTzyn8sgM6FHYFt4mYwoI3mrXYXzKx8BFMiA+cEb1RJRxzKtmscIvnXHD
41Cm9ihnAh+oPPMj1aeAhSZLa4a7USvFRcEy5wjpOMSLN4HtBWt4rgRM5vrhlucftN2eTSVm1z7w
u68XFaBdW9SKN1c2V/Bc18OMU2m/tqDDUxce9ljxvvvZLt73FXVgrnV8ob5xklngslyjA08u7KzP
Ads7swUuzTumog0aLy52fkhlIT07ogJ+JBM2zSS8uYyyHzpQUcVYG7dyCh27GWiiPWjKtrzCOX6A
4lGFnXZPyaYAcbCBzgRhk8A3kz+r29eF5sBKRJj1rHQ3A4WYnz3hZdyBemvv2F34O81HPLL0Nk3U
oQv3whvVAx+DEyF/ueiTbcx+N8sRPTUu2epW84N+yZpQ/8mlacuXIhZ2h5xvwz6+LEdehWV4A3cu
EqbWI8sx6Yj5FOiEJEKuebnWjE5G0NILc8gGnPYe3Jzvzqti0NZJbpVpqRrX0zZUCvIx6pL1gGB5
hpA0yDpAwqbny4V5Rqk0kF5hGOFeQBQaisQXzOWvhMsTIijoXmFwJ57/XabcwXBwHMTBO8BI+ld9
7SXeP7gTJRll6WyIt/MS5fWmKtqATWKb3ANtAJbyKV3AbauT21KZFbwhtnQVRF/7MtsO6bCnkvG9
YqSGUO8MorRNEaAKmx6JJBfkEVb/i783BRJswrWZoV4KzxJOm9hEpY3kaqGrQoDkG6WI9+AdP+Db
k+nKDteQP67k3MOGVwXR3y1kq9xKw7TrrS4tM7w21Vzrj5g0FNHlR7GHQZRGiaShhe1pD0mdS3d2
pdEd3IP4wlOY/oh3DeuGWTE2rfEFd0XfhIlV3nUZInHJ5Wr7eidRTYOITUZkWaJm7K6tyC9b325T
FIna4vb1gXIvDX4MR7xZfhZwzn7jG5fP8uSbsMinDwfpFcVOgVhBXoHwjSr0axmxyvG1FnBk7TSw
lGSFS7nQsuato7Bb969p0813VneVvWU7XfAItCvB07px25wHgidVWKwCsA8RvilA2OFf3QrpDCFR
vUr3M00Mbndbout8ueUbh94oFkIlHEIQpA642pc39ksWBenmvvjyG5m8Ix9Kjma9Igx9zvKUu1GL
C9YPEge4k7YjCwXyq7+Nx82NYVMGiGq+WXoyAGe7/sUEF9Odf0B+MqjJSoqgcAiMjpyHG9EQEvvm
v4pInHGI0iqigte+mYp2PgIiC3GlFpKUV2u2Dezo5jw9I/NV3EkcjqbHb9cLj+uFiU4zCO6HdNaH
+ZQCFIRM3WSke/0FprfnZ9DQUvS3dnSjA0GcgtdRF9KtEPpq6/09WXaOVc3qf6UA/4x7CytgdORN
vB+0+ey42XPY2p8yCRnBOlwMtIM5g/N7xBdqtq7r2QbkhKh8l8k39U+140AUMwlPzzS1yjBmTzvm
Lz3qZvqRwH2pZLQWoQ4kh+hUbp+fzOzM2JE11nhyBrgJ+C8CAEag2ht15rb63D3UuywDnYnP3Nm2
0l3+gv6+B/yamacuKnZMjTbHL6Pq5QAqZH0UImQL0Me9qfAfmcs3aBpihV1uDwmRzWu9DmsTe16Z
67DmaRzCJEyBRwX4aRSVO0nLsJkgPYMHuCCp7yzh/uL06E1ivzVHxmZYHgWMgKyYw9ijzhzcF3hR
oYXO/kKf1cHfdyd/18ysYZ/QtVCwk8FTp83TJg9DvbC7V/TCu8WewPqhiEeNHZCS+MlF8/nKduCz
TtIAhtdUiookZaE73sk858gTPH4r48ja/YiKL1523UK5LEkRhB4htyNhCVvFKpcUu67qN8YPuc9v
Cvdip2bjVFA6wPJl3lXz0Y3rE71r/uOuxcoE104/LnaqPru3CxyH+QnQ3qVBLInIq1+Ijd8OaiSf
WQwGsOWoa1dkgGmaKAQc3s8vnicF3PezvZvex20AyPeXtHIDI7SnZINzlXzwV6dDPjStkApvIbli
gmOBc096l/RLT1CzJdl7JkmnMR0N6+94tEZ4gYb5fGxcsYkr62WpInfLCHiulZBtmDzy+6hEfcZj
OMMNQeRkhtXkbIp4gaynMI0TduArmXb7UrAHfl0RIB8wjzntRJYEMVE61GqpGMSY3xiGOvRpfFs/
ncq/4ep0gVwr5BT5bH+6yfze4yzkJ6tXrrfay/DdfzyvITFxcKFbCRagNRFFzBbQOMaKIz7Uzv9f
4w8nPrhFDI6L47+X9/pSp99YwLIewlQ214Y+RoRX2KO9Nu9i4MtFWJuyeNSfo2i5iRJnleGkd1Cc
1o4HDM//ERYICVfZGPcWcKhmnjt+EEY5etYZXYirsSzBZ9HC8k9sLQKGFHy1MWUcmbg1FNOImgwA
p+TC5DiD0jYMlYphBdwJhGqYjOZM1E3pCaK1+6d8yVF+MpUKaJkZWHVKV2LPkU2L+HJmOi3QWYzd
toDEh1kExUnixqPNLHsD+Yc7bzGS6Al9DtJLQXsGahspIYeVGmE7aCjESYB/q9Uyr+gHdKnW9Uap
IwwiYMxP7wDjSejvsoSjcTTU75yBIr1UegDJCdyNEVT6JdXgXdt8dCOOhiHN7bfkmWRLE72ZzUbt
VGTlCZXkbJIbfVvxwjiG7ADIdP+nadyM31jrRrsHJ25NzMdADMDhFfhZlX9m0phr4t3+J6QxHbgC
Ls+PDu8WF/nYiN+XEiAAnom86J+muj/MKfUC4nHTbTdZHCY9S4SFPjQvQz5QBgLivDSfM65KTDVP
84W4FcEN+jSVmlY/IqwQIx+l9rIhjciM1WL/dFk5w209EkVEZwwukw6tOy1YLp12UCIt+1bKpPKH
1Kgo4pGDhDTOWjJdzECTHZfJs2sK0f6bhRLoSxTcxAwSgi7T79neOhLCxsVHx2CtXkmCRLaHFCT+
MkmjUyaccIq1WE2rY/Wb9Wwme6pGKDUJM1wzlL34ZqF470jiF7I1ND0s+UHyp24aeumAsPxY9q8e
c7Uj3w9vEu53yi3whOimCKF7X4y+0BUrjorDjZcpljm1ZXfNsTSqa/SyQuShEhLClMWaiDKixQhC
PMDB1SbViHT20XxkNlTLLT2XggbbOLI9rWE4GOx5nmEjCxBcy0d2yQ/0GY3D9xRzxrI4u1sjgqoi
EcUz4J0oxfaHhCYqijLFjJ2HF3vPfnvalloTBMxHgTDepF5enORnKzjXSWyoHMuNH8Ud1EoXB8JE
b2Qi7Gc0VLASH0HwzylAYG4M3ZAPXDfKa8OjSnBvlD7YdsAuoDa4oeSrdycUZ6eb8kzRakrokzgS
OlIdUB+fCf6tA6gudyPeWQxwVpOW/dcLEzuXDZf6BUjN8Op2co+bmhQRCSR5JJAQy5Qv0ejjLfuR
pc1fhz/3kpmwwOMY4ahwPj/nlyvB1taUTg7rWj5Pov8+nXTkBIHJZnIulpQIjhhUwQLT9CGm1bN/
6DeMjRZW+lv6LT04IK20qHskdlMje9ZzVhvjIsIcyS7vH0YvLYqwfXxJE4cgcEQxUba4eODq7jdP
RM1f8zgv+88OKImINkKp9YKwSRrivNEISyLaXC8hnIfJHNcOh16fUtT9oQwhwOHXEl+PkhYUIRz/
tz2XLilwzHZKBwyQ+cRwyuLznq8Ggzf3VVpeGs8IwKK0PNs6p/OVh69ecTqEDPCrx/Rn4ekJTK4F
2KbMEO8dQ2+SdSY61oSt/oUuAUdejo4+vaas3WdoL2eWbW4XRslxTZQhWNbUyHiKKYOONla1U+KZ
9zbiBy1giPNbjVvuxYV1dgNJ1FX/rqFWcYYCCJUg4ZEj0Y8TxG2j5+ZQrMJLCbVy3EDJbIEUQM6Q
lWjxoTZEneIcOay/IIGpveEAhFMPG0hi6cqTlQ2HV9Akw9Ki5JkUCDYeHyNxA3pzKlyElW1AnJvx
SBlA39EiyXraQrXXr2I0f7zX3QADDn+dvWwywNqIPKYdy/bsc+hf5V0bw/cP6ds7mdmf85KHYRKW
TAPuUsygIH8G5b4wzRELYQwN0mYmxx9K+KxNN02M+V9ucSQVkLGNhs72RKXM77sf79w+HCsr7sF0
kvzcxtlGDTZS4ei5XnclsJbyVrwacVkcBvG9M34HXHlhaKPE90a0Sv0rZCFMOCf9erJwmS2hU28K
tgsgU+BAU/XmKUzZTURVtS27zu2B2DJNtSj3WYhqzFM10JCNGaGEBMGK9yAXXFeNN0/qoxVi67sW
ayvOdWcEoK4x391QicT04Eo7Cp2tuk6RlsuUmC3wlGyuvTX10kfHupyD5vW354vI334c26wBWSHr
TWMucZ/bNlNGM5sf9gO2g5mVAxVYUXnNk3unjdbjdS8cb40jrbK1Gv9BlvyWwuhaqK0l+Bi3Rs6V
MK0at3JChvwawAI9KMjB7YRX5kDZrtVmFOlfpqzL+6SMo8X/hCT/oupXz8HeHFLl3K0uRiDO1rex
iLjDc3pu3p3/cK/XiPcQKX2gisbZ6JGt6LaC5eVB7QD4YiM5LByxl1iO8ijoGQHib/QCR1s+oOT0
weuXjsOrXLXmvr6HyYRkiCeQU7MuoMOccJlbzo26PDtWcBkVXe+ckCmPsQxmcWBNCuWjEWjcbhkL
dqDgtclmR6IN45vbm7/ZtPnRKIMUlsvCt/wm6myu1kCVBtFXffI/XvXJknjfjwzgSPsutj+BlRaJ
YkNupZGV+CqT38OaTrANvNeWozKjtzlZaUPtQXC/bhUGvD+qFYVzskmfTvgrDTDewIBPOYxfadEH
3ZdfDKZlZ5BnuDI30bUYk2tHv712dVt9QAXtNIkJhj7zxTnbaxf+XKNBjfrZRr0zmtbDUqEp0bv5
d/qLp/efy8lP6fEr9O2ZifidRwGe4sXSrywLpmGzZvOjLk0a/3AiOSIl4i1zO5oigJm73tnqKz1b
67/pX3SvdTBg4vWjFTVSmac159CKPD8KOu0FBjhDfqjGorQuJWkPXv+4QlSWdWT6B83HKR1GQley
INysS39AVvv56JapMi6Wld3ExFnA65PcQ2kWF8bfZ67bf/w3CveOQnWAx652rS5iZk9oIJzF/WRa
eKoh3n9O1KKu0J1B29Gyz7vYh/qGUB3L0Grh4doOvdxyiNb/SweMDuY3navv8fQ2ZuvlxbwPWQ8s
9FEorzhGy0hgrwoDF3VRdCCDPhWTBtuLAQMK6djEUADYAmlJbAM7ysoUhKAS9ewbEpIJEzBW6KkH
VdD8cLeaq6el/9BTWoKS8fBbIe+hoWpZx0otZujuhow5hW9yXO3zbmbOVY8EUHLYL0Vo9/q8AII3
/VmkukgVKKr9fzj8Gk6Vo1CI1zpm1wbUrIDJkjZjm5OY1BIidI+q0HYD098Gzka0BU6+pW7BIzcu
zEMdimy1gkl31e+uOoFhhLmlFDlnxtjgHuouopEWg2iV+pmTl6hPmV+MPwQOjI8W8boXOx2mgucI
ueUSo/FQO6qeRPtNx2GVXr2WjPsdvSEV/kXtc8jR6K3Icz61ymK9e7WLGyOIhgdm4/TguK+hOi4v
xX3dcCW/f+xt1ZqOM8xbbTgldkPgAooW+e73QDMXW/zxSYIgCegVXO6A8N1453rFx233sWs+XYIX
pRdFjnNiGGTomTDF9mXy43DeUCAN6e6ixYqmrIJuMoRczjAYN2yaL10OY3oYHiMcG6z/ERJo/uqd
W7NjqFIQ7piE29mx/Xzqq5KV39uG6waweVBAkVGlJ84XQJx5MAQSlBm60bCKt8EgtA7q1Tqhgd1x
FxuHGV+zxlSTeRyQpQtmfMeg7sISjEN/a1fw3F+A2NcYaPkulgUeWqRrAmP8aRICR2W5Er1q27hw
+o3RayjA2mlzj1GtWPaX7i5rqQtRbV8hgnUgjzu5hOGIHWwUpPkWJOW/6frj5XJS/4jX3yiOR0OG
UTiWzEiq/wBpDDwDxA/Cykhd+5tlQ77kv6faKGUsWiB6054lt7bj06eNDdJgeh1qRNwKUH/OnTsn
TVaszhvasH7LqHnaO8ECXIXMUiGGRVNQHVoLZtE9nfE6vbVm1hrKL/YQchEq8Ah4KwYty3sP4L5d
gGV9bKzDtTuzrR1TjH66Hpv9dv/QPukFlsBaD0AJ7Igiw4RaFZ3DQwfbz8dGpmgPn0Va1VYv03Rj
Qg3VzIYa5RloA/zeunNJsCHMiIV1EjMj8rWU+nhyAwQZieh9SMrwWknrrRWRTxH9CF2vv0WtfQQc
SUBhBGpzDowIoNcINmXAJGnqmFeX7/hdJsOvZzUwN5D/HzuY0XOQVoZFe3Ls9GdXnpcC6NqJh6oN
mrMzGzmhEYM7rrsozShFiov2lA2Kk35ch8OwpJG4poWfVQPDsxyPsIDY4WmXFDwsJN6gDnDb3+tT
0joIQQymQR8jITgy+EYySLJA6PB2sCOqFYnIxEaes1qdD/o42KV+Hgy3dGPA5sdsHTNrpN7OyA2Q
fbOxDcQ+ZUcM2Ps/SnJbrvR32rL3XqDo/mMM/Tul7CdP/H8apQnhKv5Wp2hn7MoBcmboQR6jml16
975jgaZ1G7pEw+88O41hUDQG+xLyX3eWKT0GeWohLm4aWrhhHRehs+ntjRhSZt6hjiX4S9iVSZmV
4YgwGTnUySYzzJSkNo5IEaEmaO4ixKWAs4paB9HpWfHl6D4O0SBgGA+5haS1usAif2zpJ0OexOwS
lhNz7bd9R4u3TBINsyAi+gVOw/jbpdHSlKyjgiqmkWHkUBxM3Xjuy6D2fINU0bxZ/Es9NYcELSt0
WiB+qODCfYB/FZzGdoVCXMy4Ul54g0HEXk0HWfyEcZHOtv39bwbYnsr7UA/qEHfg+/yvihTZzEB+
xmdH/2W7K/TUnO5NdFglWz5+Ot+T/5ZRpmFYwMy6f5OQG/mVOHJvq39jSkVmyjUNLwZrpfveMJY2
xNym27dsZCjgvFpOpfN7UuG1VfZv6stRN34qG8unqK8rMNqVWSFM8vx22y5UBlH6EewOVFHVgynd
pQTnRauOjMB4fR5up2FgE5lswsP1N+XPyPZ0c5MVGaI8mNwO+zEKey+pfplS4QolodI3jzDYVKh4
LWFWNyXvP3Bg24i7+S57u0pDy1d6B7LfuHBqkfdcD90f/Jt8U0bFPAIje9F86s02ax8CLql6LtzL
/E3eVLWt5O65rbkCai8VSScLanCJ3R0dP+lFTWXOzdTd76CQQqv4bSvdPbwKh+WHPYqsvpKYLTyg
ihM4gok7uOg/2+yV5d03+bBJdEFziM/m4oSe2O74qr6NhrwCmQjivyisH/fc3Z5U2XfI2v+3tW5C
QJFrYYVdcM8teF4sQe26jQJbsWkmUKGxlG1ZTbLUFkUu3C2wXQ6EIEUqlwlhWwD1pVZZKPuxzqGE
p20Z4XQZnZFme25FAGv7f62iMnW9RUmZKmHa/eqZotjvz0sjpObYtenD2f1O7K1E4wwrvBH8/tMj
yVA5GO6nGLDH70NLQInoRHZP+OMX0sYtHlYx/9TlEnvGh5aq2zSE33bu6Q2qNtuBUmXdvmszZkXz
Y4Z1WaOyhTtEsFih+nVwq6znKDpUyUfKIOEtirYczgfWc9HBJyoiz0B/Qqi71RUeS7vUYSLyYbHV
16qvoQIUj7lqjFGsXmS2Cbswing261Y4TyovEq/enrBii0LG/dQjUYCUI7GflOVxABhrV9ZHja5d
iuBSN/bo6fUDpNwyFQrQ0lyyflnwCGh5uVWkg/YpouIA0PEG++RwDPRTBtuv0icxKJl1mSUsrfFz
YRA1f8yTTAO3FhVeQ6Va+R9yV7Qz5y3BYsL/cGRTvDeacQNhxfmj+Zf80DfL3ugv6FI9C7Fv8L3V
EikMrm062hQjny6dLoBZ01yXi0+oyPKvSGBIAFQvjmnxNUhcPk5w3L7OQs8eazmwksmVsbB+nZV5
y9ic95+ee6l3DJH4+QX1h/5HARuEtiWRfPaOrcaz6NGM8e8ziY/sHIUSPb2TQVS5L6/2e72sFtQV
as1RwtZBkZ12/kDOrxdAgPKLMJ4GgQNLfn9Q2JcB+QCEMNC+Z0pZDc9nY6dlGcqYYayjZl3tamsK
0E652iX54zpQ0KGcdZBmZ528VItnaec2UAF92OuPUMv7pSdLdCl5govRO+GINP29CCrSkhLCgCHK
1yhuxjgjNS0hdwp3LyhvCW8Jk9g5xaG+wrWpwlsg2cR43Vrfj5wR9+4OOBQEZ7PXCM43bpcclyGF
xkROQWb2+WYrOpnS3RBsGhRVBOQ51IYAEkLdcSEnoxuEMicOHZriZu5kGLWaUQbrllfaQMT1Cv+k
nZXsQMstQ7RfJt552Rsdw4V9pgotlsEi0wzbPm9AidT3MtbJH9mBDjovzWtK6jfipp0UdhO4R18/
cn0RVfQzUkPh4jKaSNsKdk3olR9hVFYl7I4nth/uRX6NJ3X6Tc/n0MXGM+6UEQesIqwGf4Q09UyZ
8hAR8GiY/RNFxZQSkbANQVZzd+7qK7OwRA34JyQkwt/Zt6cWUK3rIJnCYNIys2jvp8V3OzK6PS96
0g+yC5s6Scqa6v9eMPbHJck53/DOIY/5RRT7QUY2CRkbMP2fPYjzYOPadIr7qOG4/Aenmqq5rDkz
OmJyQFE93/iihWStS7XrWTD2MV6IApl6O7gockPR54Ol3Uo18wZCb8yhUS+DsuqDNTB+VkTHks8j
cHUOFNdJC3ab5xPmxPx7a9KI88bNLOB8uCIdYGaXt03re1xWF46/zLOOPWDVHSOPcz4oAzEh3xHC
WGCsmik53AiejVmefxZaCknNYa7MLgLgWLiffYyqfF2RaBWMfOhm6pXXdicSbO0qByTF7qST4tqj
VDZLEajouS/3FweA5iKvGKvuqe4dS2ps1CDG+Xgsfe8wOpXUCjrNPNUAY4XX8o9EP+DoZWn1uNG9
nOpVnD07SCwt0UIZlTHo6NMwRH+VXii09yQgcnNw/P4AndMIHRubRibSdOYkNCr8LKxy7y/XlGqK
IaHDyCJ+cl1wuaOgqW01fTGsD3WQSNf8DB4Pw7MX+Wozl9EmCAC+jDLX1UUMVZYKNGfDiqVUtEh8
qB+BthdnhTURyqfx9GqqBTRFz2961OM1MEStLDNr7nl4gQW0TXVcSmXUdW7uCl/O0HnokUysYUUw
YD00cAHo3NvRnMXwhTFCiaxLXJhBr1N1DxGKnFwb4YFNk6BQKx2MNMTP9i1cuMLo9SUARyn74BgC
9wXrctzOIeuR6zFqo92TxX6zMcK0x9txMX1TLVUPBPeeVvR0Smv8ForpyWIC4/fBPIQJqbDL0nuZ
HeP1rlP813YnTiRaRmAQGAJaynTW+7PDtTnzYiS6He7U+tcXpD+H5EWfcXfa2rZ8NvY39nxfCcQz
RHZFpHndD4LFOkdX+JR35pLPFtMF6Rc73Y4GzEWDEco4L4YY/UyXAvIEstE1qm180t8Uv2jkE+HL
WmbdhwKtNARrg5B6ugjK4mHMiAkjGNpRTbroFX0g0swUA8jCfv1WMtayWukoNg+/JRh0boqEHoL7
prpQV4rJ656EPiKgFMQxtHg4IT90pCt79dE6mbVbGESrs2CgDcy7r3InotvzehIpyfYLi5vwOrtX
BQEa1Wc8TjkV7+Wm4ZeQCQ5nzIhydVWZEI6oM1IEK7ZhfdI5bqDYOYDYyBjf8RBK7wwpNtQoDXaZ
Trmk+2+0RZwfvlLtO4qwjHDilNIWhavppPBnOHV5sBEdT8Pp43jRTtCcuVyJNXOkS/WtuYjtxbEp
RkT6d8rJU4YHRZjMfGhmCQMnmvg+lBQ1ftZKBpIR8ID2Kj0AFPalI5K0fIBKZIrwGAvYRhsK3Why
GYKdMnIKxmPKE11qG8Ih3HYdN8/TS7tsaNgjt4gYhza2EGtIkQIl7pZsccHGzFHlHynXh4mfcKKW
GA81CiE7IYR6Spwo9Nb+zrJzVwLQ2XhrmTM5T94cKKvjcG3U/yqZvpWKshAmqC8ozFDr7D0rYOW0
H/dM2EnVWLH7sO0vhtbp0+uOUND346zHCJvEtPqr7FB5yLQWPa43/0EAl/P9vPCscJ9QOgljh9dZ
7IP+KTFcFgGcwNQ7eoESb4PsaOGtoXfkQiLW0YRr03DA86acJUecnSVjpHEG7zebVg0u4J8YO47S
ucc6ZLeX0YUwGtB/f/lZCxSQLcMi98OfdMyfxOYSxaSCnT/qMOWRKSZJyvboHVPt35Q+nYLqqVa2
vaYylfV+3hbr6DDIDvXvbH2Io4s5mxmBnjkRK8iQHfgEjy+/MphSVLpmM1TXbGL/mKBmqI49cRkS
4qUSyxSVLGdHa4q4nwsJqAp9W4wo7jm/XAD8QQ5JnI3TEIMFrQ6iw/ypFLiZ8vqisP28vIUvHxV5
jVFn3saqHtUi6SnGW5rsQBoYwNSlEYA3o+sy3YJJX7oCP6RSVqPvpvwKc7eStZWqXfVXfmsdzEmc
UnPv5aB1soTdeBa7oeOwCRCiwal0A4JTUn7SJaxL7fQ0Bf2K5fJZpWzL3sNrsp349oXJP1HzvNbw
bQSo/H1MaLz0wW8nt5x3KonMbCCyo5g3tFtjzJyKTxqPBqxF2uUTjJwz/l097HrJZgy4mKhpTSXk
PdMunYv78ZzlEICZGvwEr9nHmShTHXpsnAu1rCNfiCsj/IJa9iLtEksHUX7dGRySImnmfDVCDefN
iWTd8upsqQVzRIYXZN9LT60reS6srqqM8RJVdnRcb7SnMG+HYOs32BuLSvxyf7dLBgplg7XSvOA/
RsdgJKEwfZ/cs3rPcrYTnFBcJtwfjMq63gGXdhY3wbJTZluk1C+5QpL5lNBJW3yg1hSdnVxz3bR3
343S9PKMsdGq3a3AXXsgUaqIU1uEwgvTvnVQd3EzABEv+IycN56WFMHZ6WdRsjmk2CNg/93PBKTI
w8gmkG67oCj6HYf4PI4cJz/bvcxETm09KYYWFF+u7dFGPcxepdnoOnHP3219cied3Z77CHpcHprB
M2HksZJy/NiSPC1SV8S9ylBG7Bbnw8eFgq4XMUrX+zLVAlgTlUpCawXzM3rSmlU4o0Lb3ZfqrCav
JLf7N8s7n4SNdFqbqK5Epyn9/3M9OerrZjp5KkbEYFQYnk0IzkuaY7KMId4INtpcUZOZaftSLhXb
hwa5ufIPBwYM7/7Uluv+XPYXbMI29C6INhUCMPQqizFxWLQ4e9/ur+p+wducI2vtjC2Ti3TVb2Aq
DMqVzoD78YbaNKQBiYmNPiD83HTY5O6bzVoC5YK5S5hyBvp+Vix2V56WRHrMktqPm/EpsexV6+Nl
1UsJtvH0fcxd2vE1g/TXhxCpCsmnMVsEJIopXO3XnBmiAPS79wgAz2B9DE9//enENXZZtMyht5QW
qQi9wbblCp1bLNhbNojFidjh3fjMw/94POn1XcgvTPcXJFf+1I/pcqqLeqlvTFI8yT6YRSLvFth3
x6m7EHXxnyOCdiwpbbzXGUIszsBYNjn/psXuoyVCITVr+6d7hQ6fKQWFlD2a0RPMutUtdCGQoyfX
13eAPUd8eE/LN2VKVSAo4zgGCPFzVVjCZe+hze09U7mx/SGTiQUaMGyeaK9fyXOSYBYRsMxEpzOH
wR99Hg6ZhLZA0k45QF/uHnDtpuQk+J0XySUQBZXCFpy2V6ml0vLig9w9e/n3sRfzAdZhqNLaRUBh
wJG7vUCDnUHvNjOMoSa6LQLDnXRFS5Pi+1ttg4NLjwsAxRCjpke2Z0tJj0Y8dnnBwzezbF5nmm8x
N+BHgvxzaPRI/jmPzoNGZLEnt1aI0MedwcktHK5ZtEgv1H94h/1+9uFtMaHE6pEQ3MegnL6N7OAD
N6rlf8vlnc5fFtpknDKRZafydCwGLqsyXxQU2OhisDMD2Z1Ged9PXnjvPF5WzkDqGDZzyVbdKFFP
S9XgXz025yyqrhMnb4KlNbRSTGoZGYtLUHtVTgLqOJDtQ3O6Btp7HXHS9H22/yI1CVPK/Rgppm7G
mhujZ99pRvzZGViHAPlzG5yTPjFZ1Qgq5C6L2rmQwcpe9TsFSjaKdvTgC3iNKAAIYK9g45ibIgOV
aHiOJL27QukAQDyJOd8C5QoQarxo5JexKhsBDIzPXinPUCx+4zTSY6pcFHBcT65Jdbni2nV0ElSj
q7+w2pFM52YgwOe5pEkbEKKlJyJ63sPJE56qW0Gunrk8NQGBd90GGZQpzcD0s6Y6PAfed69ZGuHv
XnpyMvlP488mk8Rl6XSB5tQ/9c+VFucOVB6gMAvdM8KnchRi88jROgZS4OrAXuwwM3E+UPa7eJ4I
QghyMGDK8iNoXBnHF3m6of6S09FNz6qyTK61GntSG+Sw45gYEaVXlSbRqvIqAMgbxcEM0nvL3ZJB
9Y6dwRP+s6S+hoqN/yASKbdAgPTEwI6iio90fU/XgG39POnYsSmQy3pPXnS8NFclsj+YlWqwsU3p
JO4RQ3iV/Y2ZDTP9XvpYZ6GNC/lsc553/jqW0vjgVaTSnKr1JuA0ufq8Al6yPYY++nOLe2W2ytjC
EQhl3sykZYggYnPEyC6IgKyQHr1KGaFLMtWjsUIZ5S3kWNOz54teNtnLavv8zsyoAqIYpF78ct1i
aliGELJqXOiLvSlTRpZQPOmuvt5oS9zVgm2RC3Ccb/N49sXcMCOFNGBRXPBBqauGyoW8CPZfA8oh
G95kyrEGh/MqlDxEttCsMjtyxStTuF0IK4ixrtag6okz2AxgznuIMQmwhw5s1fHp0El5EMNwZAx+
CYAg0/mxrW4sU+L7UyuNbFkIDn10ea3h2XJY5NC03HfVkz7KJ+61u4UPA0ZXLCyAi0J2XH2NGdDe
Ph6K765T9Q+525uqz7zvjbMax0If6LQoUYGDWoVSWrHVJLhVKZ0TKM2nZ0u+SJPmQ8wZme+xRMWA
cvFauK81i1WQCeRs0R75NqfjcsQeFaR8U3ag169dvvidWBhc1SOatGPxhHlxqTA4/Y6HyJuK8dkF
jv/CKiArqoeip6DK/s7Ehcm20x4PbNDMdj41+ZTC2+vXXGzpMqlbF4CNa4/J/wQQYxt3AT+2ocjF
nRYqdrhQUYh9ouhiEpr9qtRHAJcPWjpmGnt1L1ywtnmoGZgRLBGBqf6P8DGq3A4C0FfrR5mB5qV9
p7hyHLoc+tn89zxDEgkGv9Sd12Eg8tcThnWJKd/FdHxqcPHEWy+zupoqim+Y5ioahhbsI+mcISio
MzXorZus0RXq36tcC57fNsgTWHrVvBfV23BS0cfVtWzwWcbpIoXDR4l4EjmtrnElM+VsKnECimQV
JhhDeDeJlq8G4TentQWhx8rhLKlf60c/OKbK3/XsMzLZNG26lPcU+CDXsuSCj0f/Jlg1VLMYUPIZ
YZchZHPBeFdc4tUwdoyXAfD4V6/Y0OAFzvB3k8QZKC52LuTVQuC4Ni28oTMxEhyuyEh/QuXFI9yN
v3VeYkxk//h0246g24Dm16L1mC7KmxflM6rlctu+HLDVB0ExI0kD4f1HK9WZ7DYW3Oo1nCaYOy3z
h6FmXh3Iq0zxEHNogZiFlFfCjhQCzQfVPJJrQgUbMn+/8+0eGg+KlzvItJnzDig1Z5Rn+5smZq2V
aVsGgzvtH8Us6hP2qMMnArYzyMu1Q9nbZe6b8BxsQ3dihDNgCzAsvnG8GmEIQKHfRdldiWTh1dNx
Vi13EDgBGmhpr/wE5vTbnvM0E7PCotcm5JfApLwvHFZTRviu/mYczwLgXb26lKA3S3IQ2xIhTbYQ
b/GV6oLvnjuLW2xagMNko2xpBX+o5fVLM8d4cL0ZsMVq3h8uvoq83nks4THOyAg5cXMJa3xmMInH
sPwczuCiExW3/kUGkKwJSXRujdWGAMgGhF1VZe8jG54PjHH/8JSKsItelnJUsRSoexbIw0zVMJaU
k4mmd6fV/Q0Jo7C0mDxGJsgM/nVIWHDBlsYbuql1iPZmNLwpPsAb6zHbqD/UH+7tzUUMTbWDj3rC
gWViMjb7nrdHqClZcIFBJM6EXsuE51YnoNihongzfh+d7eRYZMl8AKuM9MSyxC97Gsm0Gl2JoqtG
1FWlUXwQUUcLJ3RTG1JzEGtHSivR+HpsE+JG7a1EfvjDvJSbZooLKXAjNLnjSWhkUtEf6ZWePuoZ
c4emdz34bjfqH/x+XZAqHXtQPQCJONQVtkOda7rTOxfCnstRicMJjthfpc9yrwFSDOfJCEj0+/i4
wBK5ASwwUzcTETmAEwIzzd7nXnPONALYAYWsN/W695q2n5i1kJ1j2OlmHm6v6nxJGP4RovakB2G7
rab3U+IK97umA/OdDFO+Y1cAdVbX6bxAmvZEz9hx+Y8/sQkwdbRmw3mriWkOga4gXH0SrnN+6gk6
/sqHNgjFD3WRlgkiy2RsFlOxS4gFCJKc40aFVGxJjDzh5aVSwihUDi1doSmymm3BFuHXgRFw2MHn
RvX/juw5lIIbdP2xSI1hTY1y4auUwxEMEPrBNxTvuoK9p9cChABJOT+0Gt7UM0klEGIeXZaRiAvG
2PfDQICnuVXUzTkym9EAJFlLDfCCGZQoCzGNHZyFXf+SFcHqeKxSfRAAawA/UhP8HOrzLYojcL9m
tmZiyNdH46ztFK8xmtO0mjICmkqKX+AWOiwLluOUjrpLHLsFFKh9vvBUZGfPxY5X2ABs4Yp51XKS
J+NVDo2p8VfZ2nAbvPASwdSaFtEU3xEkNpbuYw6hIvO9vEU45a//qvcT/E/tN5RS4Ka1F3fabl/v
oXrjWd5ZmMVgYYAZuyc3/FcHpV28k0s643Z0IJb4HU6gWEonXJxtKC0OyYlRR2Y2Z8aQ+gEXC9mz
+HBdWNk+tIHDNEw0eu+011h2bBu5ssx+FcYQQDHa769g+11OjUPgYiknmNDJ9JxNcGXcyMFD61Rv
yt+Ys1DiU+QEwbdyE4XKY7MTK9YqmNvBpIT3zW2lpWx+zOMjW2syJi4nbxmkL0x6CMkuxjqJxTQ9
23CW4+RaAvC0v7ro64b6vnpNVG5HdVmYPLLp21awAnKt4COGx4OJoyfcbvGSBHUFyO9KFZb0LCQ5
VqGYQmjszo23H4tfVueMJDD5WzOE1Lk6flltGp9d1BBJSRsKWivDZ8qR48t+j8ZOoyE+3CDUQ/P+
6Opsd2MQF4bJv94S54HLz5L1/fY5An/J48KLXgDKoPIsSKpPNbeQPmeAmQ/if70iEFVnouiECgVu
43Nh9LmkvydW5xeBAM0QgVskh1hhCz4UzIASyNQQXg6WCO/NWj9R9+6qkOb+7jsbdwH4qw7dBNTD
hbUvcXRHhy3jwfenyqz6Fk6DYZ0knDmZ1587p+s7iItJV8Y63HgtkjtwWMsfRQ10v8/aO39oCQni
Jga/JkxeD9X9qBSnjAnyEQHIYAZSzthjp3A9jmShtOLbFwuwT+W3VRs04eHGg8qZEHPRy+gDoFx8
zUmzdnxtY/5Y0m8tY/35GorDWlntssKNuaEjmM1IS0Y/9fePvG61NCJbOZW6BmXnFXsbHFlwdZRo
P/wI7tnnddvMmHtNV1oBbTTCgAbL2CImkK3riwaAchqLTtw6NcsK2rgzB11oSzouqaBRFELJj0M5
0S/uhfqv1A/bB/9F9HS+R86Ux/Wd0sWi7QJHn+w64/VCSnMbXQmAvE/R5UfmPDTCqM5DF0OUFnqr
nC7F4XO3n9HALHJWWkMRNRCUYSuiymB4T/N3rtueawiIc80f6ZNOBEc6GdIkaoUy2kkMcHFQP4o/
QRfv5Jievpc+IpTeD/7kx0ULhDwsGXuNnEkhuCdk8vhbX2/L+9ZWtPPU3T83v5dHyuvhXnIKQs0P
hPYoXls+GTOqvcsXLOLSVcsjUn9Or7LsoQJ5fkmk6kg0aB2VAke5Fh94n5Mm8RblM48H/pBrEp2l
LqB+XCLT2gdsGOMMNL1XeHs0UU9O+CcLV+RF5YKIWy3LTBLR6R4h1zk2VSEfITKOsPTG4t0XWyYl
ANDLnDczbEderxFYPqr9r8BibnNdyToWK+V4xXt9Nan6mqmt9+QSA+aq5nyX0B6S60C9XxwGco0O
6MRg+zri97HZN1rbR9r2AT3PhrBtQpIyegkldacO/eEJ5ang788iGBEgajI3TwO7xGZZf0o5YhZ0
XJoJcInMzG+H0D4UWAjZ6ixp+dEDDuMkaaszDgtUJqM1szDMaQQweqALHgtI8dFqJfSBpU/AyrAO
ZHF9s8+y+bPxUWRNXXRj16KHIRwHXYJRAsLshDH3hOLWMoYB0QxQetwt7LPDVeQRDut8ugI7WyIl
+0KwzMD8BOG3Yq79jcQFjUy8zxa7WqTEmkC3xJZBnhtoaOoLHaa2MECQpM2xNizfs/3Mk513TvAH
OvSj364++dLRo6XuKgY3kO1IxOjBzxgVvVdLykK/uR27Dz/mcJkByTNs5mXQ9yvZtq2xxgZ9Rlav
5087hAg4N3KCs5gQ4o3E11DJhemFVfExIEK7d7DOK/2luHn+ZAwUSaJLq32SNr2UZ81o14vJ0Yjd
AplZmdm/IrGUuNyXEU0C8tDDv3r4ATvVe6/gO7jG8BY4QMGu9i2CEf5NhlW17vsShQsyxRrMh4hM
63LCvIV+yiQjlXB22zP5oLZJvMqHqiB1NZEtYP9tLGBwi2NRYxhpuEhb5IKtwnP32SvEKc4KBNK5
mwximkIOKzs8Q9MDei5AFRgUTX/ZxpZHglIcbXrw3UqPWaEYEClmBky0a9E69WUMj9bTrrsmS9/3
8h2VTIWoJT0MKcws0ZpcIa8aDxn+6gVhXr4/7k8pdo2gqb8SzjEo9UDyGVrBzWcZYLT8M9jmCDH6
kZdbocYySOTLVtOE+eNgYKO0C8eiu5pNG6jYu3H3fqe/W5z3CcnWd8fHE8jlViMqnUOHpRYzZRtw
hKMjFA/dlLNhNqz9CqfrmdC0UrwTZfEVOONUUkK9Dvey80fbW15w1d74BwLAY/bQx7LQsRWPJdC5
6KpAoQkeGZEa2LOCWsCsp3AVpsAYw7rWaKdl/72sXm34cIp53Ev91DpKZCTMeo7TF903+shUcMFn
rPc7ZYcLnrbTPyzx8hj+olFpOo4Y40OMf0uY7n8IKiMb2ajN+KsHWEb00E/qUZTQbnjP7pcLOJdq
Xz8D4fs371R1EGKBb5AmIylYimm3WyYUiw+zmMg9yWf8Kf2skMQa8DfIIT5MuHb8g0Zu/K3O6SHE
vcZCF8Wfm+zM3mkGzX+L+q0ToWfXfYeDLQkVUElMMUmejkTvq/GFQeOyzbfq306f9lMM2DA31I8i
Mml5/MhexLSuYHGcrczvQ1WkGK8yqlR6VHuIMEggsr9gMKrEA/GEmbM9MuB9KNftZHSViC7XGW6X
rfY2hCpA18SgBUSTVrvzJ9/TIsIYRaD2CLQn4mL0h6tdj7ASO7DOCOh8dxYgdnRNTQ5H7aqwTvmG
/91eemEzDNqCvDGePHtLjlzVuoqfEicQSvD/FqUHuRrmKWsfJbRkQEXbPf9pfIARjJG8MdjXDe4C
4f3rmSUhFLyqRLtXWxUaSDsF2Ifpmw/S+sHrAv8YHFr2wYpR3z/g+SK7Wn7ZpBAlu/Mhko43jn7W
o5jUndJ+NsaVMcAoLKg2jsTQ3NhF2lRR24dCMnALwkd7oQvogytJmdaQmxhbK+o3SejERlHojf9d
KUxHUrGAX+aXR1wykkafiJ7j7qcq/cQqaTS+mi1qjibjl3kgeANvdpJuoiabnA5Qv3H0ZEiNGnrE
QbiOX0SPJo4BY3SatBIsL7SCeSbGI3YULd5LEQ2PSdQ090lrLqcByfSGMyh+GAQ7sZaNs0iVm1ql
qr6uuqePjCGg9+DaRTM5l0oZOboBuzXgsD7nYHIYXG6VKAI4ou7YDJqTtJk4lX2hS7Q09cnbqYzc
aGI1FhqJnGB5xMF1tiitQSS1DiMBxCpy8cL82kb0T7UPJyCwdEu9gVJRQEfv3Zyt5PmGRsiKg7ux
XGQTv/F0Kf5OONolyq7geTnWocoNEPPlVWnEHG1ql34Tjj1UhaWmNK9csmnq5GRk7TBStDXLncb4
zc+rLUSDInvGvvzOZq2YwxAUyql1P9Csh6XpGMzYJCD67tl4aocubkzR+MkdNVLR340c9tptBM+x
ltgl1v6/eQSFZKLZ4j5V81o+8S7KJb4PrCvhR4/FxS3tTZRbCVgEHaH3HTd6HhLcGMU3NAyL5kLM
LJUmpaNS2Cdlcp4Pm7UJz1muyeMmJbc+xbxHHfuUFRgUrmGb3cfF760jh3HJWs5gsX2h6YDHY/hy
/MJSMcZ3zI46CTTGbTnVq5Z1hdTQ4M0WVNt8Pcf11/B/EkPf8AMy0tC5E/x+Fa/i6JAVka9SscsA
2o9Sx971ZJP5On1ukEm5OIejEj9oUju5hSJjonWFISKSHwV1qEkXTOx5BwWXUDGA9hJt9KePHUrc
+sddLlk8uiJeV8GldmVQpcSsPxMqpYsZWWeAbQkCcXB81SjikZ9/fDCFPvCNsShFGCDJrCTJq4Am
eBkP007IW/axMvekF9e4cFkpgMk8sktaNagENZ8SSanBd2CxsR/arujLt9Q+gj8PXSk15Zp2uBmT
vAXRhxQaht3UvXPkXZLNR0iRN6Xf+ZXNVeEDuQB9TTMYoq3Nsc5Hls7hcp2SgXIpIr1suTHLmVeY
iYC6Kxtizqqa82TfaEp7ZbJNBiW6E2E4r5LWniiA90+l1NUtQpz4VZGf6PVnM9FK3LvVLjhw8CPB
rbY3BVwm//tj/0QyBhuqxGdIyRjbwjLLsO7NtDCqO1yNEoH99EG+ZwOo9RSnu5SiTY8fo24pNJZe
Wpup/1UoraQefNP/VKVUNhP09amGTeS51F96P90uRTzGNMW5zA+MHOft8//BMiCcnbWTxwX0P6IO
aexOOhNDWLEbcSDmMdNlO1c2gYqIv9hohRnit8jlUYfbB/sMiGvAZYhrWY8zkE3RGMAjRXGQrXPs
FOlXawfNk6JBW/Qs73i6pK4zHS6Q7a0pbUOj2pJWbtNuysFjMmPq5q3iuZJ0i7p7Ay5uJkt9J3I+
XLNIb6g7ULWm3c1xTuJyzs0qHFqV9zWoNnUcqo/FXo/89LvsFGfL6PqlDdmoK3+01SUUrnXRF/TQ
ezI8BEDZTGZbMVoK6wMkzQX8jxDCiucBO4Zi/VRK7AnCk/zikk1ogxCSIo7PgLWRX6q5xQut0qYC
UQmwpURhSQJdJpjo5o/MrQgsrk9fNlCSDwzwf4Gl1h+3wtsZBSZ8VrDXxUkk9gwmbBQszb/YooNd
WIFKRZSyM0Q8iCLv0QOq3SX+TLSBDm2CQOtUEimOA6L2+9taY4GkVVxD0nyZ+VWDavy+ZYm7V2AT
ZHSJYI2EXwKwDja+u0bCU/Uke3Ytt2P3/Pt6i8KhNAOQdIn5JizSbIU6GahC0MDJS7xsJYsIUTBy
D2CniFG6RULwnRfMAXfh+/oSTm5508KC6SR6SJbjRv2edxcm16w5uKA59VmqZp//KqjDS2/BGfSP
AtIykOOd3b5Rlq077H9kMLYEUigExl8/Bb/80x85cv3P8ONR1H+PjBy+dHi4h43uMRHLWWCqVyNg
ZpbEMWN09AimaBdS0gzA/hkyCdPKmcOzSeb+pDBszZdmAI/ckAUn0JshDgYO4qZ0whgpU0OqoLg3
WAfVaTJe7D7uDRBuVqAcLGPXfKj8vwTsvbz3BhgcX0ZaTrC5+KwftfpF6QST/RN4fqDfyJTGS9Vz
5PSX1VfeCgj9/ernzP/qZqXNvejLJAS7/7qC7Ntg7k4JCVZopYCDV6Bw+ZxS6i5DGYUAYIo2f+Wg
HkC+yKHfZMYRa2Fh/jS+nL3/Q5aqTGG4pTNHs1ZONefnx7dwrxlSY+3HEzVw+eSlnVFiwHRhibSx
VJaOnHi20emG0vciMeRIWOcxw/QrODja8tVqP9fD7Uijq0QCZkHZxzblQjzU2L+yVULO8n0jNPO8
rKOwERgzPam3IHiHZB4tUpCAYzQZ5MVvUAttdKkMNNyrVyydM/fVllKmpKFmOoVJ4BeLEVY8WccE
lgy+9TvDfK8a2ZSTrUFRNx39Wtav2cR3v2Y+bboDkfOXaPXOzIKidrIaxBJ64J82v8g9vOtMnJvW
bjKWXyC7fJ9IOI9AXsO0Xm+pifAS7IPn5vk22H2rojCOMC8zX/6Pjo8gU69sHNQ8FMjFBnQPvPhE
VLMOsx1mNSSsQyBL7OpXIa+oxdhW1u8LAfOpMaOY+ba8jaqbMUexCkXjZz420pE8jbf3XyBhosLD
DU3skUDzWgI+4yggL9Wvfcor0KeKThEuGZbDk7DxlgjHlfbipeanyDg4Yc6Lp2W4R1awzekY5Uuo
gRWH4o58BjWchCHL0xmuQgz1WZuz/BW0oQL1P1TwuKtZ9zab0O+TEbosKFZZAbb/Vc6ho6moHprW
NcdiI/Des1kKoDurljCUHLgWHlwNCfdZHZVzBqw23TSQx9xrfDIAyXbyxMgH/fJU4aY53vbUT6xO
dNXV/EqHpBc0GPvoV33p+03y06etxb/wR8pKNIqTbl4Xed5SRUNq8l/RtEZKBOVFlIdONuvH/LEd
CmTBcYoO8eohZOaDEowb84+6d4R/drGAuPvpqf4V9XZNJxiZUwFR+aMS3nKMny4/UrGAC2IrJP0W
FSz4M85DxaWh1SxjwUQOYYEH7g5gHNgF4gH731qSy+mGSa5T3YbDCc0Uak6A08lpWWKNFxaKi8Lq
hWR6vlQ68dhxlwJxYROEU+pfAJ2nWq/ZlsOGdD8SdU9W6TRIvONptFzhI700SpG2uKV8m5tP4wRu
vKC+Pa6RbVU+m1+3w8zt2cauBXei1ufWgjqBwBcaqyROrmwi4MJkdOw1YIwUMJ+C1T/NL3DxdPm+
uVsOZGPcX9CwVMAdxYYZSZGUxl7Fch5op6BpIzPvuW01UUXi0qsQB4ntvTgXOvrQytYZ4avzJ1fe
gFdXvqnpIvp+eo6kdgVFtNY5lc9lfsYAedyD12GBBcxh24y/8KGaBGiQ23Yn5LpnhiaCEZCYCYJ4
DW/jCvecyvnoAv6jTZFLnHG8TgPblowijLFsWgf0PCX9JZlmO7ptSM1HNdBFPzHigAJRALi+t+PN
XVWvi9KTq+JDg3uD3bZ5T23CAcNzvsaGuFEo37p0txdmHR7r5tGgOGjEbgr1CmvDin2INAK3Casz
yeTH6DsayqkR0yIJlzTVhbmtixBOEVeL28vsNZ0FGiGf0/s5C+XgCnO69GeIvuOgfevmIpzrSn6j
iq24YFk1vReoAuxdccfrz2LVzhbJdsfRjYWiUrNHJNEx6Q9JgqPAFffdN3k4BI3iGZQLcsFnzdTF
IfC6h+M6Jwtc2+oSqQO5z5iy6BZXeLlnZ4IpwvRRkyMLDPl4WRYIZ7W1jrk5D6ecZZneyczG5Lcv
D/Carj8pUDp0w8tuTgNIWaCmfEl2a8OkBPRUy8V83X4Q5KMJ4QFe3/VL3NWe0zbx4A0f9bHM68QF
FoT8jEZYSEojhyOADeP1qtsOa5VB0AfVwyQGdnDrcgDGJyxeMJ9QrkLo1MvjRvtSfvvHlirJbp0C
uf1PL55ZXK3WsKSkDISApSof09LW+SKxQVGAvSV5wAzADv1BAqt7Lq6JYcn0//5KhY5ZCgwhwHmQ
jT9RumRPa95RMWfN9TE4DKBwKPjWykiSDBDxigLL8vJ9ejrrSMJo5lH7OTZ328kZH4oeupfcZTzs
SG6r1XQdoRsnwSYqlqMkbrqWFn6NUZXenjpVTP9xJSG0bDntQiwbwoMeRWfFS+Rv4eitLjgHnIpV
yxULvQDhzSZO0HHHRzk8F73NW0id8AjSh6L8xctz/qmjTK0aulkRk9pr7rxaIlg3NC2VGQMm46hw
B2TSM7LGeo2bDka/Ox56YseZEu3VHyFbN+gqHXbVLDFXNSOnZ/dPXtJvJWUPKHN9vS44FgXP3Xqt
A3znaaqvMzgyEmml9pUqiQLhHIGUrpZ0kUMnA+7O/ERohfEsB9muhLOiC4eykXT63tOKfq12ou6L
XS7dgxdFRKIPW4LKKH5g0LURnUaulFi/0TGKQyReVn9pwVME/P8DOkf+ghxh4PZuzHUMbPaZPmzA
0703vCP6XIlt5NO7GufrdDDDdx74iWluVN1a3vq2IGa4tg6hhEl+KApwrnn/0MEOyDYO5bydaYjH
H70sEnzCRBmA1+FG1N+ejJb0g3yQCas/Ow6hgyuLv80o52tc1cS8kxBRwMvTUbLVL1KKf6E+uLVR
Fp0O2jk9+A9wT0DIEA3Wf9+yDrvL0vvqcN5RhMelWeXDhx11mlRJYMtZgjhfXjn/HGrwEmfdZ191
22XkN8rEM5oSmkF7d1+7Og45OhqP+9VSWU944FDn9Q5c9wUB1DGbm65oaJtfbJ+wVp2g8i96eU1w
cBx1gGVX8WcJz2b0+OJ1NI+ZUevc0QTzxJBU1/2T4uNyyLKbFTKDTAWtaspmIG87xIJ3LUZJasub
4E8yTJVhoBOuI/IvjZtW1feB6IdVukt/VbJ0bj19hAdg5Bdy6LtbfG1kHDZSHH94eulvSm39Cnoi
b7FBcGjCWpb3r2GNPSFml13k6fDOPRQfva6+g2yTibVhD+G3uKyK5v5Ytt7cqiMGYecJoOsVBU1G
ix6/TftltHC+e/vJcxYU8uC8wmoX2r4C9NfO3Pem0r2I/5SQAvxfvF2IY8KwcZBi2ipavXDcMKOo
zsjnA4+3vzX735/PZ4xzG0sRh4uty1EAOJHsu4sIFZxRmgkvWmZk/99cvV99Zs4wtctPBh+yySDg
nQddJojMkcobeDpPi4fQfPO/Y3yAf9A5OPfZJDPvFfAo8iKWHjZYE3v92VJozf3k1R3N6emoG5Po
atbpwtIlmdPPmlhlQizrCo59gc5CK/iQDR+OmLHAngJNCZSfQZQhOu0Gz2+sJq/TbnL/T3yj9Br9
G+LFXSZio1fXGwJXU1fUsEQiHA9rqnEzCK/EpZIYHbHAycjYlP9vZ/xyylUPwGUTPfpdYoC0Uc9S
CapsXgSyTBY6Ba3LVyT28Wsdn3NK3zDxL0S9Z6v2s9egdvbK0cEkrUORnnkfE0H4C3yUKSkpJ5P6
D8BFaMx1eTr1ZjcER7qUNlYlNuT/GqkOlIB8s2hto0705cqbAxrlZT6gipxhqjQMVTFVVU6ZyWNU
zSBke3aeJ7Fn2rLQnrzoeTHd0Fvaj0a8hPL9/NWguJnemdM1rxBEBujJTSB0Osfqx+5OjYrfeU+X
A+O2kH8y6yuFGQ2cdkHKTFH7jpRDPlbD2to8/N4wPh4D0e5GQVXXeZ6rIIv+yWle02cAtZwl1OoD
3UAp6Av2WICdWeGgkdkeLdd0GkwfjhILOnv0/FfsdwKerziOZ89Sl390BxkAMGPILZFs+Y3CpF2r
GtKPZQ96rXBHzkX/cEMYZn/iCW9FF/OQql/Km1quaoiQYMPidBr4VvbHBQCHzKsmWgDUdFU6EI0F
JKn3OyBslToZei4ePDpXs5Hp6DHFGaQa/TZkkikR4COdmI/9VUUIAaGMiSwwsuWfjKJFt1hSKVSL
FmKr31x9gOH92T3dFrG4V8JST3S7CPJgRxP40Rsptowy3uDnosYZ0yRV3WSDTYAt0h4KQLcfJSbm
hk0ULOgSHJbnMR7dBzCrFW+xfANhlf0AxSLcn3sg6ycLiC9yhbu5efjDU/6oMR4s+fv7nr8FOp7r
7p5z5Qj9FfmjsV6eh/qmUMiwJ8PEcE9+T2hYjKQnui/JOc9sfY0x2m/d19mPwgxLBgGStblAUdbO
GOxyGVSdgxAw32J2ZIjff3nGgZ4FqWlLRlLZZ22dAA50MGnF7YdH8zjg0JDyGe/+zSZh/6+Nq4LJ
t3/6LWZN9YIuEdLuDs/z4uiSJc1oGJqcMlR2LMCy7jyIw1ZGwYIB8fGxb+ZFl6BNtOvOsvoNvrUj
FHEuomiTSBXQMKaCaTo+KPRe66OCu4K/IxzqEG+QTbbKBStPGeLoS2i09atpXFNG9S6khMTUFSKu
sel7FenSUdFmEnpZRKqsm9xGa1dzm7ABQlj32IjciZ9m8mpUHSClmrbYJk3my62co/CT4UPCNgZI
2PDSz7HVIDNKBxG8Ife4Zvl2SYEZJVaZRd8d1iJoJmhuUehMM9hRynsENydONenzziumTjHkRDwA
P6n1YFl7R2Y+Py+2jeWdm3Fxhu3m9c1dx8j6WTvOZAMcSyM+86wzt/uF+0vwAcuus/J5p/z5VkZG
ExhS7enqruixdSXHG/fipiG6N8eb2GUfkVhC0tGD7sQe/2c+/Bd3x1FGoaWQxb0g0BeGJHavqwrt
94+L5rKpP/24hRZCFk+FRLkz1HZs8AyNrbw/kCV4Oh3P81Sq8I3EsmxhkHjiG5lohLrdhmNgBgxY
+ChFTtZ4gFQ1zAmMeKewyANrTMsiApnZtKCZ8G/EdUp521r+FKZDSs23V4X0e99Ps4GBPKm0RZOT
m/Xb0rz9dx7oKdJ1qoSzadm0XbfX0ap+g2xRdMJT+FhOUkY8Omqsk8YMKJMzBCfsCsdscS3ve6MC
YbVasXR0Nl12YduYZXzRTat2i2Tn1rGYscihuRtSLUGC4kyTLHhi6dmhlY9JZVZZQmSloyfl6AEu
ggnH9exKI+xkkTcTzDvDe4bloEvZd35/vng8WGwqiOSXt2/jf5W8Eoe+CRFwjz3EzA7GT0wjAW2w
Mmqa9D7XuDNa7rcMh7cJsepln4UhE/103yJzpiH2WXfeW9s+KVb5woY0vNNBB5w/SKW0LxoLoAVQ
EI/bxKjGBVdvlKi/ANGXZqUYwkuZu00KhBj5HOtkCK1L8+3MT8561Jmno/TjdKy09/dwMFoWBuOH
pthAbGvCpZzDd0u//6OQlgYAetkLDd0prN+gM6/8jaMUHn4SdqVJ7vCPxURlzx6FLZTSfpPtorcK
8CPRWpiTNwYkeoUZwgoHBoys4kNvpRkaAK+29KBPRHEe/jjnMn3JM0yks5HlPQpJkf2149RvFEDU
4or3DzfTyS43u4o7hq8ytPXAXve2am1mztG9itSdOOy3O6aaKDeQDjh4HqZuuVU1vH9j37NOCh0x
CuYb1gWVuU9pC2tkR8woj5PDX9riMDPYl46r3y/+rvVgqQv1CSkskac61r/Tyl9AGb7cr8whVoJ/
PGA1MI4jRS0tbmD+CFLjGo4eRcOAdc9zGMA+qQjcvZa31hh6M7EMfXQeeXV16aXujCEIH2VZiCvH
kCEdvYPT+w0AAi4dEC/K7jTTt3fTr9FxfT05hJMnEckOoFPRxYQE0KVjb5cqla8FeVU9FUG38EEl
t17JWkihZPB2JBzcLUP3/2+hEO6TmW2yvKGlUTajkuaPK+U6z7f7zPsWn31ZEZpdEkGYn5/Qmini
TIG/krjW5GBLwekJ5LwTga2GziKwCeFJhUzkMH8X5ZJ5e84JNKw7YbhJGiATVgVxWQT+Zrb0pC9+
AsGOmRZE9TroqYx34E6RQ27A3TTpCETp0SZVxihKC9HlWqU4Vd0SWnMQLNr8EWLjNEDvQBJz1sO5
iYwH1YmkSaPuWTWRgwbhfQDHVcC/TvfRmZ2TyunCL3mLvVHQgie2MQcvbtH1XXSB29qJX71xbYHk
17DP8awKqCdlat8pF6fiLXLIzqKOagzEp3SXL+03zycZfj5AigLBBEl78LCIE2RlEIbrmt2kMS74
gEXb3F7Ry6+rYIL5mV1MxtWm97/KTl//xjuyObl3zd18iNdp8JXKWi1ZWCDHpkZU7dwpEZ5yIzGf
LTHY7e8yqmaaqq6fqhVPOLexpDXZcEsMPyL8lEKOLnJphEgjJrdt0Brk66DSQjeO3qk4ZU6WUeRb
zqRziZg6pIwtxcW9LZdEKsBI7c5n5v/5MauVG6GlkrrxWWLAc44di/vt3P8QL9mRwGeNQncO1tpc
06++71rUyjRzMwF+vUMN4sBNOKhtyFHSAcFOno+SIbioR3oTosU23x8x1apai50Y4NLEBUe8ZTKe
GZPKakZ7bYolHp3snrgqK/59yIPjEcyA2m+SWANeDueVnjypFjqPJQCwCpXHskrWo36v9LcNkyRa
+9oO38DPOiW4Vg+6o6hutkkUs5ABPW8AhZ3HdnBd32+PCtD7omJOGM08Hi9nFlFmy4X7LAxKPGW0
jPi5A/+V1Gav4t4ClDTF5JQp6rwOC9w+qU7tln+uoFryYYUg2dNJ9VxMZxfqrcnWXIRvIeTZYjuL
mtB7p2PreiUrqH1BBursIlvJu7wtFSebKSoe43jZqahQwUAYGGT/w8IPKHbHQeTZVrJULWmmGDt7
1KWmi7e2SMSCeSfbDNg+wCIHmnSh6DGXMx+fZzEYJ88MIZuFdVh2jjfp0iAw0XRFUZwLvIRQ9Bqb
zUDqj2eTWx5xR+2nNrf+EDitBU9FnLG99YwZLf+HH2Buimophn6EliP/UhTfspHP5iCvP5w7TZB/
LeLQYUxZVWLV6CuMSgeQTzCfdzP1EmJygvkWaCgvS23OtPnBzyrGkXTAO7jqpcQNZjfhPZF6kSfA
oqmLxqwtSbOBw3wNwLtGK94VwTTv1bg0ibIbfbToWZ85ydy3NRQHIGubSuRsqI2G8YKfZ2HCjZI+
6h7rtfGhRrz0rswyTie81VQnvrvt81JU5xOEsSOx2BtaoficcqVkbk/D19Yao7p+AikDTvcFBX92
jF+QIpq0uO4tuuW7fwgKQbLq3xg6w8U2xUfvkxjjH/4MPwIlIi2575Uxa/w3MFofajSuI9fHmHXE
98yBoFW/cGFEYuz93JOtHAybovYNbZOn0IDjUWHmCLOwszr6XN/Tp71rxenJgt5p6aIkRhnY9Adu
Me70dM+m39BVRvEMjJnX+V1gMHDecexOjUsi7qOsJmEccN1yRmAElfqup2i3aOlBzGTOcvpQPDxm
Z/ThLHgxgpeC7yesOUFOh59ft88xkjJDxFRoiHrH0lJaH5veJXUeWLPFxcv1ixY+sIkGr5dABN65
/xxP2sGjtS/jMKwhcgYqtKbsEgVzh7qROZfKPN767LYfgZHglUftjAfMN5PnPy4aJZHYxYPXdW8T
Osco5nX6KilvsLBuLpSqhJDi6pkF1db6KkAhBPNMsRIoYxcLD3l+JmPvuS4smkzXywTfqS5eHC2x
KVBBendhp5vZL1WnXex0qZ+RnuouQTk8pMP2dvejaNF1OsPuOgjZHeu/wswsHYmAkkdKI07IjLqj
bOElP7KnRKY0DfDgOop1tYVIjVYkHKFA1+zm2iIKoqiREMzCj6ojzbR4nj0IY1YTtfILE3pZ/Lc4
qPCdx7cwNBIOfiz3LbFpeDnnSzjLBdU+t6Ximg8uuSiJcpci1HUSTZcs5US2H/dkxKXTdkVi3pvS
30pf7EJ7bkT0yDKrbGtuGW73Iyx9PTn8f/YI/kln0udoAREhevq2pSM4rpmQSOTMGSZAArLZnDIQ
5IrGHDRqsegR2DJMSGFxYMoy0dVwwhJtumLUoOxFHw+j0a4/vpxfvNl8zkFi4uAeXm5jOd8nIc2X
4Sf7jj7+MVfEx6vq214rdIJohYn/xWdqpiLH/NQ3OxoJtZVGEPtC01+wLlHFW59SD668dWi7Ife3
jwzSsThTv5cEhDji//zADX6p2aPnlNrwS90MAMx7+HJvcgE2qkPgUqGB0066McRezcOGQJfGweZY
fSzgWjQKmoioPfzjCvIs1aXA+VsOyJgvBCa1qzl5Wd5XAZjCi0zOqCqoWkCsYYLP5qCwhW9CbHRD
Zt6JRtxuuPIf7c7gUiZtEAWgk9V9DWwxzqdKRLN7cXRvMtb/6t3/hNvCgBKIZgwHgvxjPbTvUxBv
VBMchcNi2lE33UqV4mqXUnJ/Rou9I/hKDjttaG9TBZjb9hQ8pNz3LQDbG6nIemap+t1kHg2ZZbNx
xTY3eNX9yrxMDdbTwNCjFpKJZSQdvAEpiUqf6jy2Gw/lERKyB17UNhXCwefX5Ie4PEc3UJaUFV2N
yVggWHmVtQifPuAUQMmY1k/QdTRmcNvlO4LPb+Jo4mzghE/XQtSt9Ma0CUHfAlgeXWo8BCqGXywT
lJxr9cmF9z/Xq3XqlgbVkel77VAx/uAXiEorsdiSDJOg+XP/A3VYjfk7DV9NAdXTNJyZAoOj2/Gs
PBQLleeRIM12WxZu36jNmh72YSN7ukx8a1rXjpkrYGZS4/6XamBWA28u+0g05b9UmdMcZVkUWcBk
Pl3nnjJse/Btpt3dOFsPNKRqHFQFDt/ptEYMyCnxjA9vUq+LkBAyktWjYSGGvu8jaYUod6me2BT2
rV8Tns5VxJYAtThyv9JYjtxrWDAGUF/W3n1KkX1SPN0/jcNPySoyJCe4bIyGs6aoWvrO79BbP98s
iArpvDpdnm/HRhMO5kTUEAnOetVEqwDBoIX2QWRRNhYlCfAXN2CJuyk8lDwli6GrB4T7AZTAH2VA
fKUvfKYzp1pasibi4iw33lvM6Qh638jhvkill4LTdOzXG9llCLLdSYnn3liN5kbk7rW/3fPa3q51
rzxKNbUJx+BNXIQAyhea3fjT9xNwgVzMHwzHaNSLLVQkkNpHxWuz/DPf4mTYn3pMkVi9Cajxyz+D
h6ClD7g1aK4bzZfv7oO++tAuBGY/YFAYIJbVVvWvTTcXVieMZb2oHIUeyAzlHUHZzafcOYWthkVV
ePaCTIY3K/wBbbi3GNxbuKQdZBxDY8VkNC0eAXIJNNkneZufcBVE81OgO6A7wOzMHH4gIVBJwmG4
OLxnxDn+CPsooK3Ms0p7HEunwgFFy8k6rsSq1Gn14i0ahd7yWHq5RlAEJSRxKqFsSs3Elp3XxjzJ
q4rmXjrqyeRnPrcto9gekDxapw64DDBmCVJxQA5t28ZmHctto0lldTpT1ruzuSENgG3AQhsaONJs
Z6MJyDlJ+i+eKjgfUyxUkqMROcSU6Ha+hxcTekYWECo98huMqHb1O3KQI/Fy8CRvEzqSugv3RN1H
mUd3X1GJMrbjY+uSfIF5o8MQsLKM+c9fyozlsJbeiJ+2C09wKxnAntIfWqGfBvpaoAdvblC+jhba
fpIR9gF4MBO6wiZOPSwk3sEfqm6MDDXZfTkfvBOwLsnysGJgc8bbNtv0LqeqNrHQIjmLi3s+k0Tc
3wEReBTXf1md4M3gF+0Xwf8GoVal5g+rqTOXYtRAwgYE+JonvcaWIMVNDN9/W68czryx9j1FpTSK
bf9+tqOOSYTH/DncES7hnZh0O2WWsKXYPu1WfKWnTY4TLqEky4ZdXd03ZKpVCQoSDgcsKrzAU0VI
/jBghq7YgOvBSceVRm0GvwsRjMmwjkhzuvqbSmGg4BaRn2RyFNNAwq/0FXXa5L7ZMA5yJTDyRs/m
jgYL0HZP7weFsvzvNg2yqnJKvaKUvkcOwNQuF75Yvfb13WjukqajSWX+CoM2NMVEL5zMy2yOXtnF
wK4pbunIsXkWDDqXvNCbFSsrQNqOcMdEMHdHzfJ8vRDTngOA77Eg1rGgC7X+mJq1lPbAj9a8O2Xm
/u7nXiTr40pnDBig4K7MbQCrla++4zn4hMAx0Ulnid6lF5Xd37Yt+0Ry05vcFdwAASiy9sXSQv+T
iGemE/UWs07g10EGXuNbxHbQ4RAgyfXxIfR9emOQlpg1+Dz05VefNejKymbqhZmSjx1EQopULGKl
oWWeN0SFPARuXWUkd1cv8M55Z6WCkhvNCeguPfcoO0uDmrnAAN+OI9o60NmC+Z8i7Huyi56UK/+e
KLnDTWlueDhtFFsFIYIt5MJ6lbktypVwbAcKJy53X7h+uRJQyYNqtiyMfKi0wp3HlIQYfSW1EM8x
M3K4ElUg/pXHmi2YBlMsW+uhOEYPZpgwnh2erpyhqsh7Z0q5nWZait/hRznef1n5qCKjvXMy7iRY
lu+SntqAcVJu3o+k1jXPqENG36ftYs+pIpJx2MDnPq0pqgU3dTV+FhI4HN0lVkhPoR29iTjWRCtt
KLEEFx05V5+mnJNooGv6VcWe6N93CB1SiMIn9vMqowqGn+OamEY0WO2v9yTJsF+t1h2UiLaRrUGN
4wUXswI/zV8npD/V6Gag+cgwB3gkbRTQfW3yTwwlPE3xEaSUEE9uXHIIZx+MGeCPhK3rXC6Hd4Qc
fDqfPo6aS/qZc6gzinYxpTRlLreGV5xV87TXW9nq+YvCxez/PYxtpZ68rcZMaBm/TPaRoydsK501
WSpL8Jb66FNapcH1prsREUCMVA/ZudnRQlJt6rIYfJeiKGiAeoVE7B3fPDJr7yhJ3LBrp4F4Qt3p
14BIxuPWav1M0d2pZDfGNAl9XxU0OBvic17JA8g/tTzJZc+1dQqdEeOFjEgTxx4HdNbOGGBR+njH
3TwfZi+2nRxO9c6TotfQf97o0TsbcBIf/bVBEpPJ5vfZjnNr3iTPlmFh+MIBeF2xb0l5sV7ZJA1T
upFecTYcCilKd4ByD7G2xnOjUVUIm1V3orlVqWxxWRINz1yS2unBKvU8FAkpIuiqg7OZdHMqJrjB
ZF2xDZyvugkwADWh/rHgUDDEfrKj+OALxMxfaUJ/25MyEjtm/+nORBGqx7xpH6CcE8Pox9v+e0fP
SXIzhbD15bc6wBw3F45Wdqx3qasjuiT0nX16ztCYlEmSeJn+rEXRj2XSNZwzlT2cluoeWnNcTN0x
P5mhMXcaMqY03SIs89i6MF5DTItCUtuDmv0Kk9xOQZHBgikLs0vkPXpsCgjr+F/nRTQ4HvQ9XIFK
FIHhTDUjBD3daB5JmQz2K1/ayf0gwSzeMlwNcgxSu3T18S1M4E7LKVWxhFrB0vpxFmrEO3FoierL
uX2Y+KpOr6X3BuNUyl38sf+UeBtBoLfmaQUvm6cWuL9vZi37Tb4V0CwwZl3zS1VRQFud5f7ZUu2I
ORR+LT8m2/hoi+1ZBdmCwp6Ct1nOdtLtpp14vHOU76yfk2KpnUzqMITxqHXpn25DRDRfglq3AOjq
Qj/+eq0cBKQNX0SCc3SFJ9oV3rJcl85Vk+pN46AW3jaWmpUNqd24PvVMBfFAjEwubZpeJN+Q+NF4
j/xpArJzX9uKoaESDouSFmQ4/JHU1xnRzPluRnZ+DBlXYPmVeKV99XbqLlNC/RaOU+WAKAKiCoi4
raRV2kSrZ/SqtYqA4OZxhUyv8bQWyXYbcvJy59ZZRJGra96blDe83NBvotNoJzcAChwJbRFrH5z2
Om6biLWT01z8FFIEmkvVfWB8OFLLtpRr4cDivSweLiySvdiN/lMlCermM4VrjasCa7QScsQS3zWn
n8ras9a4SuE+T/4hRd73aJZ2APr3xBpIkxW8+ePxEUIZbhDOV4hJkrz+vxhhAuuDPaW3JlhFysrL
dpp/ZrZgoyyX0NTNLKI1BU1WTe9Dsuzr/fma2RhIIhBjMQ6b6kPuRPHQYLED432NqDoGUH5S/RKy
Ys1DuEAfe7RplBruY27HHsMkeCYrSdJRPWKvLa20zZId+gXseQeD7RnXhNe0H+TUMRGZS3FT39En
OReXZUKLXLwmowRxVpmKtsWxZzoUwcVA1sg1eKRLnS2IlQvHw3yrPRQPXKeFcdDVmiRJ8FNWkbBu
Jk5jX4qFifmQBIKWwMY8v24RQV8eAAfr3DrAEtMrJEHEJoUjeqnpokC0NqAkDqGoJ1GdDNIkpZZC
cIZGorC2lNy1Yc5Ersxm6zMEhjonxwx5/+Gll+Ez5pT1nmjpZwdOt71W5Q9mcb6m52lPWdv6tHzP
kZ6vz1q95Gz3NLZKXeI/aZsBLDpQK5R7rzgkMrR48744XrBCNrh50OxdBL4rCTBtqEkczLkzcH3q
zd4mJH/6aATKWzOZEifxg6finNzc8DNuhHMeBmpLmLHjrNXIOWBIEWPobVVqbPXEA4zMTBoWMT4h
VdR6PptB1igZqk9PI0M/yGvmEtipylBnwvSywuVtGEu3csr46XCLEdthII5tHRqsiODx82DiA1/N
yOMa6CwcUScxweBHVcVCmAFrk3/NCPqbqmBbVxTsb2uVmXCz2JRx/MeOM3bxJWqSYg2twDkH5Qe4
JXuE56lXkdV84KBkHeFhxGyHPvMUNeaA9DWZe6rfVw62iDxLUmd8ci3KwKv4CBm60rzTDDEWdgXn
J/M0nM3pWkeookOjPA5HaDBCZE5jzOdckeLhrAYUpUOBgybe8h8kAxmA7S0Mu3xnkOA1ijDKyF+S
Yjp4464XxB/JeDP1c4l30FmMNfzWKmFa1xyRFzpfW2wOIjpUbXKjZn2i/kBVGzP84Xn1+41P5uIY
T7MaARAOoFEC7FspM9Mksbbsh5jJwfruturfzM/wYZyZ0I2niwIJaNjqxtbN7JIwqMogQWBg37Cv
poBrhxIXUhLQ7W8DVcov9vXrfRsKN4A/pv+0+sy1f5RI/sEew7Tuz518ezavI9XFiDCtN319u/RN
BiTbRlXRLi0XH7+2tMm3W4lrhIr0uexP386/fAiVWsL7YN15RcKyOX09ABo9zI4qS86A0uqQwlIr
6x+L5+KQfNOnCgCesIkRSPlv8s4wJZu4ED286cC9KUz5zKZuXuUKfPZcapzfZr5kSTEMXz1cSz5C
GbS/FtEH85gcIxyzvExP75RQ6uZiCz2Rx1KGwiG2fksPdATC3Tgt/kl49ZFu+srFPFe4ljnvajQG
QvVVtrsfFNXO04VIqrMcwYwbtqNjS0QvdHzK63V7GkJwp4ZwAi18mtGITXIYU/ftz8WnJ7LKYCvF
9YVdn0Acy4P195Iq1/D0QbyjkXIjQRK7FlJYGCVGqEiHJNecrJx0jd3Z1q6Lb978NhyJSzekIFmk
RwN5WnN84oFOulHcuU9geldkS/3uojlD0jK1b3Ke8euORVxfgbuWb1uMtpe2CjnStPJsVWixzsT4
5aiB5SCkSfSR2UlvrF2YFjCZ0316viUGxHyNsTWnH7EU4ewbsSWEa9vD1h7Te0BQK8r5k+Zg/fel
Lx5ySPRwQpcBQkJHCXq7ihfRk2PYo9XT5K5HjMuay+7nsKcfjSVOtakcWtqfBZ+nFO4s2ZTWeXYz
suQ/VDcXeoGMq1Go2Y85g7UUBhI122qTs2InJjRWDPGFxoqMa8qfllyDL7/rWp9XUVaSsyt57pYO
ze3+q/Bqs+FZoFO1/eJzIUAmDshMCJ1SeavnnDihOf+vp7GCFnGbFaL9MAcIyulwuFGR+ApraQSZ
Hk/dDvUyS0niDfkPd0HzJ3SiJBihun+4PjnnU2y6ONR+aKoZ9ipwScKNLwS5sclSq5BPSIkE6h3/
ly3Ds1Ex6UmAEQ7JHo5gh7XgHvmYB6YHkRAdEWSoHwTj7ITdMAX+mUbeHxg2RUigkNglgF+Htqxf
oPwOx3TbPn2F/A/0bA4MODJPYfnpbbPJ/yNeoZN7i9m/lHosj7ft7RJa5nYzr77Bx1c+rwQfLHUg
51OeKYVsRFc1I+rxw1M4liIkb1+DBXd7t2axKWwyNw/pnRZ8n7d2NAScxJLVpztMJMEvTHmNF6Kx
rrc7iDJCTRZoa7R9BwLdYiw/wUfhCyF18GpULzbr7J9ln4wggei/t1UCxzKDKYDZI/RY77dnT+yF
rJZHrvdQevzRwvkE1bjOcLMtWPrsLBCCu9fW7JLyWZBcDZW7gvxFFPiZhUj5+V7HZobko/bgDrI4
nP0YByYBUtWc4qD1q/aKYiiYRtTwf7+u1YY+qLPoVhr2nj79UFYkiFuyT5VODK0UdnHWQUv3LpGr
uajwAhZmehQm9FcPPjSXrbZZ/oGN+pT7TL/6DPxj+ZEWJGO8O11ubX39yhh7HwTzuEXBCyZSfpu9
LSZuohNtpXoyrytWUYvhUJLT/8VumV9nTtolEEajO5AuY1O61hpnBio2IHC/hkFPujh1WODO3otn
+tf8r8KhBxY/gkagZv/WvFS/QiTvw1JWTFAPXFoKyFhsIjMJ5bHobkBKDOPEnH94iCmRqI03f5aE
gvzv4BMBVaOGuYa4oG1YbvvUhGMh7lTsBND1pUjq9+STRVf2wKvJPDa1Y3urNhbAs0BJ4L3E+XxY
YEJuDlvOpvK0yUPoP4oLivG9G4C+Hg6C/rjk0QbkhGeQD+ULE/yWgSu0Wh0MQe4q4hvP83RPNDT5
8/AkUae4pE9dwULSa4vu9jTQ8TlLt+DYjgHR6mkz/R3AS8eOlLgS9AkHOIk04u6EdwUWgTYcrseF
KmBIfaZoXLW8/xfV/Rt9BF/uJKcCV7YNHroyXMWE3/Cjf2YbQsggXLBglRMpdJy7cj3Pka9+K2f7
2SzxHwFRu3orkIRCR2m5ofGz87XGFdcJJR4Y6EVOG/LPQ0EXksZywEjj4fJ6ZHqRwszxfrGwdMx8
3A1BesTJ7t1nxIbIMhGzl25ObWoTnKe2GKdvDlzZcwEz5UOHIzIo++SWSUUb4HbeqKCcYUg+vKX9
R2UtILJebmM0dE2S5mf8n1LtKS7M+qbz58/Jrb3tb+tp9D6y3ZRgh9o8lxjaT3SkGFFHWG76Lclk
7zCcpZalXdV8JLXh8AiD2+cBbziZ1rYHnEaqX6IFLMl8jatcLa71WXLCaljV3ixEUPwXMH5n4IH+
dU39oMEip7aupW6sfwjFMKkBahqKpzr81G692K1sW1e8FYeNdEpCZJHuvTtHijkIk5JxrcjQ2FQQ
UjbC+WPrZm887Z7fi4WaekWy0UhIbgRPt8FhC5GG6E1iq/RNfnWJxx7VrTVc7eNiXdfxR9oR/DSB
t+yTNHMvBrrwLbYcmos+n1fBPecOl7+ivoWcgss4g6L+ptkNotOXJW0aV8IUq7lvpLUy0rKkZ1tt
izi4DLlKiPt38aMaBVfNrnlBWJK7JOur741yXphJcJqquYL9jxgvCsSmA/yustXHgIY6hq2fn/9l
68AVRsmic4MplSfNWOjZS+UnZvIhcI+hzew7jqluMWYfKn05gi5r3HMvNJwkAPrDX6AcQkROf63g
jDZ3BgCpw1EFGFFanD1ZKYLa25jlXxdV7ZzIN18JQVhI2c4jDmkRz/l9afvjy+PVCbcAtTrm+YG3
m5vMhIs/JsNBTFuG/ZI2bH09CRf0TlXuLF6VP0ubQ34DhLcy8JKCkISgCyXOde4Fn9TuD5+BF3uJ
hBceY9mt8Do0TAEFS85IV1mee2Aw9RjilVXZcD1S2MDXsFa9ZuhQTXsIU8gxtOJt/uprzcxMBs9O
QeJVtxiqqNU7VglsX1i8rQYB1KxI1gTrwcldurzoN2JV80FANEWkVPSSd//qm9dpLig+AYN9yn8q
5UNtTJrqv7Si7juv0P3c+mZ9IR77IfPw0oys22Zm1gRCwg0CUZMhrbVQYznHQUizIyVDwd1y+lRc
1DWVqoNIZXQzOqQnjbTi7YOVUGl+3I/Bdv8K0ot8GKRtJvG0e2SBmPyEuFUQKmPKk3RS84JFop12
w3F8utDfmkEUqZSYXO/5pk27okKEZqlA+lCLxkbt+kJCUQZhuU2Z779F5VXuCWUKA7gS2iRT47+t
7Gaq1+Fpc800jvfuRMVgM5A9TqH+nPUX/BXz6Y6zzjewWzm3h8O+j8d6zWk24ntwjd7iEQei3LD/
07ZmHTdrHzeW9GRKE1r4jrs5sNZvRVxTcpeT5B9Va6+t3vWsRaWvUXIIJT6OxU+wJ959Xk2sQUAX
K8Urak9AYM5Y3NEQ3vUfEueKsYZ3+g01uB9sc8fCn12hYHxlPfUdhHdjsDhf3ym43ZvR9EizrnSw
cfQNXO2QhRU24h+6GtgT5UZKSP6VzBiDhRIcQvHvmcdRyjCd6bPs6oM2qO4FcBJ3zTdfz8Ngqtd9
RveJZIqlruKDQ3HtQvYOguXp6vAYRoAvffhBkS8NJDps6yRMQB40k7PIAJjmnt67QW9y7RkwKbVL
eDls1aGkOI+DaPCzyX7C5Nb0NiP38QPLMj33GGnhxG3PfxbJBmjfvzcFAMzy7t8z0qVZJahW5N1D
j3XuIpDvIYnR7ZyTXnV0VJpnlp8tNR+3/y/vBE/86rlVzlO8++7EOs41SxzDJ/BTcN1dARpbeWDi
gzHgO1zbH+e4gMk2e+i8pcBOEwajjsxsdnt1WqrQoI0NIouBdvlGVicwBSZbKuAgz6vM0kin2stj
PWCMeP8n9S4PMdBz9Y/JcVa0Z34sXsWPm06kJjCr47ajh8Vs8qUfDy9JGwTWpq/d7ej/0ryCT7Cw
/OluY0OjgQ1TELr1ia9gGQLFdmVQYcWgUdRYy6/Hr2zOVDQ4B5VPeGuQMfa4vvlk6fgDHHlcuPMS
OeVMGQUX4VrQyKvW1hKHMY8zkYw7hL5tXpOAsKRWi12O45kN4mPQiH2ZPV5K38lxNIJAdzOCDZ3l
8huKRj8F8IktIiliR+/wSKneQUoBAGBYwHFzT0F3y5qr95T1SIcWNUdioxFdFU0+8nlFjwDNBXO1
1REh8HkQDh4VJdMbt8hFDkhY+F0Zs8ZZa0nMS3u/AX+XWuTLMy213imrn5HU3gmg6yKtVXsV6ZZz
cJNToj2eVrvxH9hSSUS0rIyr5SZMXmOgVUcYcDe5300ERtSdeJQ4vU3aYW8+1qPD9fraWL0k3ktN
7dxkrPYZoVYuLUJxKvjxrfBcv/MsBxQrx/c4JR8q8SDSIJ06kKdTUXIMdooFEgbbnIEUxqUH5jnt
fX0oLsxQoOL53JdMH+nO6pmRR+ViA5Q4k2WIecKK0Ve1bPjCgHz7bnZpcF8QH3cwfs2or35406Up
rdqXSrU0AqbwSR7lotZTBiAy7+r4HEUBliJjMnG4Zu2eAwrw7FfEf2ER6vaRC8hFwBCxyDOEfZkF
/wCWTvfgUcu51nHiNY9/xmziGeuw+aq0Z+f7PiY44a5dQiFSt5OShQLQn5MzhOek49Dbsu++7VzX
mfLUv33VN6Z93qetYaa8DWhwLgyoSxagWYX4RnWvmivHP0n2zHuPg64YBp8ko9R6TLBY+RXhZAXg
XRFOo82PowOh5+3ogx3lWyhGlesUu+WWhS3q6fsW9W/BzJVKWH+mEggR4t9LHTLDowEgmMW2btyr
8h6tBBumgAsTZ7Odu54QLJK2nWoZ82d0mXlwZsCaRpNsaaoXduxykG+2sC4ZwimHprNvaDP4QygH
nw81qbX76pmS/SR0APjgz0uAcbXZP4gY9zIGgcpiI2UrgScF3NN29UJjtoLLexrFiJI9lWaDXWt/
5ePYybqLN8Nh126ji7vowwa8ItAQEtZ0kz2SQFB//9GwqmvxFeb33acflippYkdznDFRpBes+nj4
W/RckQurJ1RawuB4J0AX0jvg27WP1sc6hZS34bOHwyTSs3gnjUca3KIjtYqBf6y4Tbp9kJG0vyQg
f5v1AmV2nLVGBDnSOwjitySXPQ3mi22gkcskTOWX3tzQwOVWSikgKNkfiKZzdACUh6H36ph3Ns6M
nqzI3F0ESVpT6jBzbRxGwae1vH0b2V5OQQqqYjiQ5ZKYaxr7abOxd7q8iTfeVGYOsGuIy66dN7Ca
iat1Jwnx5ydYKbfAzddKLn52Abd8EDRrxO6pEZeDkUvrMFaVAO0V5NmS820JlBeRR1X81/DYAPG1
GwHjbf5RXah6Bacb9+t+v5cw/5siZ5L4/MEU2wr5mcerxXu8tf6Ek4wMKs9j7ddNfNLue9Qtqpht
u92mynRb2bvdt5+h2al7ZNg3gWozViQ+CLuJkDmIRFIjOO/ux4wd18PLGMY67qMpCX1ZeT4X+GLT
po6WBzH17byP4HRJicd3FCXrp4W6kfutH1J1f3nSqNc5xUxuzUGDzWYb5mHXBtPmnhblUh4mA8Gx
6S782TKL750RjD2B4Pzp4JkH7TW6I/JzNTa2wNqnBTlnBpaDO3nbr/t4Tlrt3R59XIUcz9sQoptz
G5ZTUW/mU3hE0UdArgAsNB19Wu4emjdQQ5nn2M3J8ZCoGA/WILGEVjzbIqgs4wyZyPIoyXl1j1Hg
zUwxKzGrwUBzzHDJDtBVSCIjNTZ0p0wYV/EkNgb/uCPOPPbu22v1pZ/Uhp7kLMzn48/ZuhdlY3yD
/knPjaKy/Q9M0iGuEDdeJYr8LNAtXi+nrm/luSWhac7fay+kDhBHWvU7/u75HrPtxSGO8agelrQU
CpCMFRDTZPiEdZF2/VCFRd+oH9bRuibvzvAIcCTwRQRN+WtArfcajOeYtC4oFKp3ePB/OqpQDcqv
zNanZpE2Zd/Np1Ymb2N4/auOjgoehA+OeDm7xZtpwMQPy8u99bsbIQKNUI8AWYkTeWx6/9hcLJy2
3R65bo7LjCodg57z/sLFxWFeYNULnrImmSyNYSek417O6vtlTekYk1p5ykvNAkHrrDEkw05yUAyX
1oA4lyO4QgwD0FXbGcyBJuQ9Cuo83CC72Q67iYzSK61EZXfzINUqd0AdlG2VAvuSjSb6ieJ3fLwE
rH8EP6C/9ZR3zcCl9X1qux85HirnFIH3/ugnPWnCG+KSHprYJKL7wra+xuy/ti4z73It8N7Hlyik
NEMW0tyIL8n0S1kIhsSHcKEqcWXSbYFBawE7g/yxCSUr5syv4R7eL4k84zHISiwRS8ckYkSkYWum
jxhuEsEevQpC4V+jvNI7k+NQ8aO/xWpInc7NdJAKAza8AYYwDcn3Ba6wwDH4o7RgzWalT66BFojc
swuVF8fwVLl7oK8CkttDg33hQEnWCDGm4S4abhlh2Cf6p063HT+ruHf+N/Fv8JdLiqbRukz4EMlb
cBWcwqf1Gpg8UZvZRFOmzrW4Vy/lrsrEyvYKiyIZ50OwSiFiBPuuaP7m4UUMDBLgp4UKF6Lwo2LK
dExZk4d74EalQVL1B3khRUADFQD6K6agUKqqwUojzN13BimMVV8WQgDo36DAsE06NMaZVnzwpe4+
77hhOsdrvrJe1gUOg7TcKB9fJ3R+CH/e3BGfFGRFhZ1H1ZTOmk+3juoBmwGmiQcOAlegyi3w0W/P
qrTN0MV39VuI+4/J/9+52FycpAwGdZmMg7tep+VCtRgKPhl+k/GMR+Aw9ZI2fFUweUADRINXaLXJ
y27/NaU8I20iSRhB9ID6JLE+nplrxp/UlWT/sk2N0PapsxnNwmFHpDhubiOMaJcGZh8cRosPRhMp
u13fJphxa7P4yFsGga7aqoLwOAQU3nwrrA9TWW+PfLONgKQsz6MjNqRv/ymfv8XSLE93+FeKEiih
Ad8Y8BQcOMV6zrojzLV3oTJKLLc0yBpWInIDW69rlsgBuwR0rPuqxYIUhufb/dVgfx+qS4aODnGk
h2gL5w03HZ5xrBAq2lmV+ZEpkNAPASsV+2uBa+AHTOBrgdnUCPSiVuc/QI/mPh8vPeU3Yx9PDd+l
/29x+KIKMcNbewOV02gsF1tmAlICn13yqC8h6Z0oDV+9+mbo7dp7wyRRXLSmGKGSTcukGhxa13Fy
uO+XJGq483hTRZ6epOK7frsXFVJA5CDmUPKLvhyrgyced4nt7ECwLrNZCLf6nyinv7+BdQ+i8K+A
5E7RxDxgXCsoyFxdHmzE8pK9cHUU0Ioezhv0Gsl8hYmacwIEKUOR7i2PCX5wx3TtEnAO3PdGDu5a
BDg+MfxETRzajLvKyvf4br0raNJHkmbaH/ZBLTK+6ij5bK4BIcpDRVL4YwqBArqec/xQaqYaS4xT
56Q3A5yOzQL0OcWSpsEdolTzMfOKX7SNFwW93zq3n8Jb+Sox2Xcs0sRUrF3xT/fDM56nXycnMDSp
VhEPM5/KSPIuk0A/gfILIa+ayV9wqbtHVXeej5IlJkj21g3PUKYdn0U35OYIYamEWkLNNqcZfhuZ
9ZTX9GA6OJk6T7pSdOw0DoSX/GRjk87zmKCCd+9IWCVghUidjigiEinccL/ExHlQVOdiO5tXJawB
RMeABm9tguOCSjU47IIwtbUFYzYSFIn6Z62Z+Ufe6NbKP5G8CwYznOX9kGARQRordj4Ip5lISWHu
R5xN+mnOhWs+ZvMB150mHbdLrCz2toOiMo+CxFGUwdiK7ePMJ8TWV9SX2hXe3CSUxOUDS8KskoAz
44WI1RhW+GILiz4d9pQPqxFQKMjYTGmg4LtxlrXbxrXli0QzA3zaD6t8uvcUVUtZHU79dI2JojCu
cJF0o5p4IxB+IfSs6sMUuuCMD53M4qkSsLx1OOaFA/xcypwU/uEXq8sh+EivYE59cSPlgSvJDtXF
VF1zcVDbZUtgVVVEsxOPnqnuR8HcOkAwkM/1PvQcGZYOIXRrkluqx2E4lEKhfwz+h7Kf32vLJJha
vi8dWpF6h0gh9pVetwdenjfL/LBa0ddUT/tjqusfu3d8/hwFEodRZR4GFv2q/1t0I/qGKV3O9bjv
lPzC33MLOGf6ugWprZVUT5epK3i0GlKum76ZEcRAdDX6kPzbqp110ZqQe4eRTkpxp3G9wgwThfE8
Ip09hg8zisnNIZhk01Zl/fJsM0dQIfxi6zL+qV8G9jrU0s3JecqPLUPvOnwZ5etusV+2azXfLZYO
lywU2SzSEWtq2BoSVppVZzlswdxG8yVs8x6Bn9nXG3ULPVxXvenG4+fBLlPMeY7SLEpbe/YL2iBT
M7S+SqU6jpErzK2xDquhxq8o+ZP4y3hHjyeFwtSLBQBTeBEKkjVKsbgEA16KkhD+NO01E8WQB8LT
bSGvZo6KkJdeGpxitjFIUSTDAtPagq1dwGZuN8UsDh3IUejf/hYkSZCyh0QhBYfLkSt5XQO2fhbC
as3p5c2Y3LfETIvrGTSgOy3A9EuECkEnvDBDEprjcwxmBHVgSin1YtnYPvUwCjJ21IHaqzRTbKWn
/KCOQOSqFA184MXziWWXBM54HyVozYLUnEb0iyr3K0wf+EAjIelBKNkBwxsXy7QblRl8yAcicXBt
asFT1Yv1ECT9L+HNeGnXe0IEloLeh3eWOVUpViFThN6SE8U/6AuTWuAdJJCQAPI9GHlJ2gyvHMAz
FQXFN5F2IzHiQ6gYhLzUQ1+fBpF34xzRcC5gNNvTGnqPXNY+NrhlDF6qZfv8H0nIXUVo6/B/AmdV
NhW94u9IQE+nKbT0Lefj5Y84sBZD8kQUK1dWV4lH5+0O//hAKlXZBddJmiS5gXXsLpMRo+ISyedb
pP4Dw1Q/jXs0rnoqWAbJ6Np5SEPanEBrrCQCHg01CwCVjFgEpsveFMEeanFXSrdaekMxC4+g2xQ9
EtH7GYgrmPWp4RTAGvbpEj9WMqkJNBJAhcrJxLdqpUhlP/MN7ztkT7M7wePHya7++d4Q6apUjkwW
ekpsFe6QnwtPULveZ5mb2W/2A6sHlY4PTWomiZYEqHvpwJLobsyJizKbF9ttjmVVuPeFayPB5Zo+
OxklWkrDAvJ9JUUMMdUXf17eAT5Rb9adZAKGbBRpYbvVZqhXnYmIyl4PxWWDMLoSCVYzLZJjxMPu
gzOl3fzSZ3WSeC1XdeZ88+9FW7LQTd1c7jsAmhgzVsqMsSMjDEoyP+swsKW9YArb0Cu5zt8Hv86y
KUbKE6e6unP/vcIFjpVjYsitJ3rpZ+GcioXnM/YAz+0KHvxRVq3SEydm3QLqMpgP/e6oR5dMYCvG
ovGe+ALwfEXgqxK/XKR19J6VW3zvfhdtUkemQqy1Mpd3RyI96n6lNPh8Vuun6cjP574RHx0FGbjB
EbyJ4xfa1pJZjylLwS+5N+VsZ5v9MFLSLq423mPu9Qxm9MAJwQ1SVtiPM66TrZ9LcowaQN6nozS4
Bpk0FlpsBcRM5RkwwnQYwAKer8gw6hduw1yDx+x0QHRI+3UAyYlSQXQml3RKsOnnGcVEzWPPyW27
5J7bv6OJ4mAfJetRRksyZ4fIQPJVYZeuyttSW5IO3JsbZUcIrOqOuabSJlIFlefS2oQ3YIP/zSHw
ZTIm0TI0SnsQ/apHLJPo82jFkozPy2Jk/dL8FZi7rccflbJKyyxFJFUqPwOayEv4nD0qbB7KYJN6
NyiWhzZZBfXOu/pMbgDpPCtM5LFmC+MmV1TcF4VFRt1kXAgpPH0EMzVq4/K+wKTAWWE5QBYXdp1E
5GtbHM6xUVOEy/8kMlwkbRHylM34AF6f55THa/q1DByUxGdGzI7uD8BcndVflsBABsxuwAm/2aer
7h8kOb/mvoyy9RfLBDvp2SL1souOo2URTpaVhaXx4SduvBjcfubIM6n5Qs89dhj5pnHEfKBFuQao
QBPrXpTsEP/WIHCKK41lP8G6R6xKsxoXXO/7laWnecLDdXlynzHBK5gcNEMHhPRGkokTQmMVZS3M
ZqRObt8VRIq2SOO170YoZjM7lm/be96Z6GCHayrJfMS9882ggi5aLD8MdxErGJRz3Z5lXnOjItRb
Z/WtM9OzscgGagpppNE5FCGh02BzWKsb86iZ2DzcE6qX2AC4h0cXCoc34tfSHgh05ILScmopESLq
GgUZkwAUxQZ6Ypeo8TI8xNRjGi0XW0hnS8Sqa5uJM791hw6UYypODuNWqXDDjqN1ZCERpjPaZSr7
ryVWCH8l+cODbHoekAfRJ8AMiNDg7wt9KRhPa2HFgjiCwd1/ht9rZYjWt3o50F5i2o8LzCLGf+wa
Cv/rAfIECgTaR2jOjU1deY9CLgho4+WkQH1YkLisGbgMzXbjYaVQ/q6QxfHIA43PIq4xLklA8IwL
zR4js13mftkDP4f19z51Root+ndR44U1OQnF2mUlK1/SAmsk28ZWUfff00ExdW41uml0lB0xK585
24/Aw3Jp21E3KLwsJ2VaZc0qfCL/PF5k8uUMSwTIp2fh2ImZtlaRBfdgYfFWNbRgscc1Ei6Xc1Ki
dP/Ic+4m5IqBLGTTSlM2BonO1/rgeReCMS9U77v/XCxDDV+LLqJv2hp0C8QtLba1L8Ti3Qa+3WYl
hg9azdR1pW14ayi5LqWHEr1dz52WwqIJUx4QQrhXepRvYkg9/4iHWxbXJdb1zvmvLc6Vf6wUPEx+
0FsowZOUQ5JYJhxanEKAzweyQw7okYwqVMQH5iyxU7y6dVsrhCUCPYCJg1giznM+SEMd0R3Py3Pb
46kRd2PG4vliG2qDf5clmGvmZuwCavvO/OEnXzMYQgj1RUm5F4Z//Riz9luyvAI6wKDq2oE3OI/y
WFVgF+U0NRLqViaUhS+iH+d4/QSdZjUvN9LuvZ9+0sTER7o1AE5bNoKN1tjV/VrsgXDtyHUoLBKY
idLT592swr8JRU/PRJf1vSj4vukdVrDIuQdyEC1AHbF8CG5W02EQYLS+dwfokmeJmftNUW+kVt7u
9aAkRBgh27WPLI202wkqfPhCl7q/weLLX6R6yOINbZpgBPO2hJhNy5WlzMs+RkCgHulcfVjn1c3i
AYtFRW+ihPmCzTSpzAOrd25uculEFef1JiZOz1CIwbgpnVSvyarjQWT9/qG7gHvTgfxjFtFy9ZWS
9ICOUZUSLem2pSO8/RXJ4Pqs7lUrXYe7B27CdEmGQu4bZ3miFER9ufm4JMwJr/UJIpa/XiKkkZ0f
SKKg2LnA6/AtJilWWRYLcxENR9CPfN2GgGkf/AEiGGHy0L1KwYDCp614P8DE9hgd8ZgGUMoLYtZu
tDE3WaQf0HgtVgqJrInpRwbDK1nzJ2MczDR1cOTkhxG6f0Tb5ImOV8T3JUvwTqwD/WHCDjggwKFb
SE8x6IewGQMb2zgdBHUUZ9CwtUMW0iqTW3N/I/4UNnhWGuE/lsUF4kmH6jOJKrqXhY0d5+bR00KT
LiVkoNjBEcwwWyNMwpmoGwU96PUR1Q+p2McDm/4NSSUntzf59a3qVFTCHxT5oiOrQb2t0b0ygDKv
bhLMK8CKzbSx8Ay2v/bIpkF6rVQBG9/shTOB6zSkwzbTZoATydABU8BYMxCh3wiThCPKa/DyMyXb
/j6ew8vQyfALQFp2uFJ62unN76jwR94fLXs0ZI4ULZXtKKHP1HokWMcwzzD0zOG8RmV+YUyPurx0
dXHPmMBLrZKT4ojlGFCjwdELk5AJQV4nAB8CChqwFkdnjp7Gk/l/T9bEhH6lBuOzbvPkaS6KF3a+
yGLBo8LH2NdT/id5PkJIeWMIW2Um86h/7fIw1FGXFcw1fPmY+B3f2DG526D+NgtqKe1TVNhZMOrd
Q/Vf0FBvhAqVYS9znyOJspJIHPk7tRUfyPdLcoyXWIvqjke0ZDylllPvODOT8HKmWXKuMSncxOL7
CzYTEexRu/5W90nLK/ttd6n4f9DLefJyn3gwhKHj6e/MxIabQCEk+Nj3AnTsUKsWGoqsIrYEcyPL
CVz4ucfiGHz6N+g28srB4HMGEdd8iXTMWmyOi5Yz1WJUV4vcrWwGPIqBmPE+79MVivUd1keEFbx9
r6bbkhmsDUSsdfMYFSLnvgDRU0VdpBIBlbb2ekXZCGbxOEy9h8ejuiYddV117+/1Q7Q8yYgFEuOg
FYU5mMNmN/CWMrerMvfCwbsHk3NWmd7EWGsjlmq7Sg5yf4QfHQlIgwb07FzJ8uBXO8IelmJeCUzT
aHf61QHy0OIVreP+3DeAqZdDz994CvyEdnPpvjpxI2wTC4q97BMtXk+lIBILWdenOr1gu/5fWMHa
rqhal1XrLh1iT3N+y9wgj45X35yQfl39VC91FJ+kid6HHyhFx1dyAxUnCl4vFi5NhS/Vg2EYh7J6
46X/vnRWa6CqCFKiuJmWknVte/E8kEPGlhr8iqkEA3ub4dASMgBudcoeCO1u2VE5wuNLv6qhW5IB
Etvvp5B0yGseEHn7d7lJi4JdQh387cgwdmaOgRk0gc/d0kdcoAcN7LjF/kaE582bM5jyKxikR/UL
e/xJZhHc14XaYo0KtRBSsPO0l4px0JIhb0Nw99gfITfcpbQ28EihxCg02NmwZaaM9dqcPQNKPsDh
BtQplGpcO53M/7MwyJzHGICfyFGmUhhj4Ie5LVJC/1Ix6D/IWh4bj6btBVR1Xb5WCfVp2o7ymwt6
I4JW5IJsAOEs4JjJQg59rC0WuYfddULDCfcszoxk2UlfIvUUXASfp3+4Ub9rtjDJt173TgxEA24Z
PjnyTVvoMWDaezDmp+unSz9zsGyvoZBhHhLrbYMezJRybBje1ZYPcAYD6t/4z7vxzNx3KGHea5W+
JF9m0oBc535KrFjf9NNrK+ZT6/C6Ac88SnProJQ8p0KblFE8qvCV3bVbI89mfSLQrVUQaaCccV+3
dhngVkylhEEaaV6fQI9y6kfVysOI7kp1VvRqjxDG3I6F78Fws+5iGbyM9q8s2Yn25H4U3Cr9hC46
fVVobiQGiEuavRonCpIaHWL75WlFaYCyzS0kU6sPsX6RirnQMcJkfo+YEt9c8bLRZxTgAH0aUGhD
wttlPYFaiRbGfpPxL7dHpWg7ztD1aHp0/+ZfaWM/iMmKWRx7Pz1F5lo00p6P2UpETsmBad+ACQjS
WVTGh/eB0Ia/eTyTG0ZAlTp3WBQ2nUq8nO2KfjOCrFhorIHp3xz5M/kqjo2vuu4WreE7ssevo4SA
RMdo55c0mjM9jeaIoprY6SU/pWkBzvdukoT0vj/u15sdSx5FV5hHw5aH4LAFgvK/dSY/G5mqZfeY
4smcXebVoR9fSlE3nQjSYgobtl+DPWhviiOG4mti+8Rlzm5SxRVuygSkA5NWXiKAX7o3fIltzSFK
3mEI4nkFcFLbZROYVaFtZV6RYkaaoY1MvcTUNGWOv0maYtUx7XCMNMiZ1wYsqWrjyRtsNCuS0e8P
+7rBo+mf6dGcXL+1lOpJMz/JDrdnAiWbXx0BTaYxmJDbbTQ4lk00fnhKHoz80eafY7cDy+6hvbwG
7+nDOiPihiQm1PhETdVOg2ja3s4g0DjKG0Vv3JRmNfueSyuPmSI/9SwvKJNWNH38C2puw8/au5MT
Je7eGSgZ5WY7stz4czYon/mvoCUehiuUYU8tML7R0FLUchANJxfY5KSF3BvXsxURu+5lGxGyV3su
y279T/6ejq6ziw0J7plX3yalLhsLo99K6Gcwa+Pc2cIhdiw67vjyYvcsgRBFe+tefDifj4POpBAX
21SXFXZIg4yxCli144CCfJvFirsfwyjFSTvJHEs4Lnw5nLW+7ZS4rHa4LAQqkK+7xNTVoKRlDRkN
Lu82g5kkoOa10bK/dAnz6azjjkc29ROML5lEUlO2+i6+s/8TNHYEfJ68dEqTZQnLx2So00grNtE4
YafMngbGgUDLV1zxltu8kfi39kIOOyZWOlGJZnBxhysHAk3ZUfNusgOV+oIcUvjwzdWFfPFQ2KAE
TwOE181grD++Hc7o+z+Yl6B1E5myP/PZGeRBSWqXYdDEmFAKPfrFnEYYhqP1MMstxp/tlfFUEbFv
R2U8nKqq5uCHOd7ZNeUQG0Q+ClrEalUDCJsxZwcmpwbhRRZxhXyscXJQG8FEi6dg/9J9XGL+E9ya
ep45gG9X+UNYizuWcO4OD1kN5Q7jnSMmxTYuYzChLA6b9Y73i4npMShnypqJgdROMed1Kg3HASQf
U1LmJQPiypa0p8d+BR7vKqnc9CRrxuMCqZHuk+q68i9+X2Vz0lZT02zZ7pqjS8hC19BiAaSw29Z7
jUe1fesYeF4cIbo+C1/95COYe0T49HqHnSxgdLQPrWtJf1FnPk7wSzQu6eZ5ExeDaPmfVx+aRn3d
0TgZl65Ij1BL/5XWa2/kIF1XPPHHXzm+Tfgg1g40Ifr1aEd+cWbHgD8MpnOUE0Og/y2oPe2cMO77
HfU3e/RG7ph8Ht/ijl0bAhkPZPF1CJbAINzYSZTRJFCsVgV39yMf3t0wj0aUK4pChTSEW9TOskQT
drIjKvaZgjvNoQRVUhxeikWOHelBTdaVUIRxRzHLNDABvQpeBvrUtaXwXybY9uLFFLdXSdc6J5Uw
bnVQGPYr+f2NEpoAw/NaW7cXWcDblbxsxon7VFsflFG/VAp/ECUz9eshX9/OmeRUkLPbILw6qT1O
6MakzR2kYLcZg6XkILcgJWq8qtCONxqfUM+VCcZqoXAQWy9nXeg/lKPnAE6UO7px2rXixT2deogm
0ZrR6KIE524jXUP/ztcWvvuAPkjDvnQm837o8deeRsjgL9sP1diaYQZDgJBLv6B6Kt11SXzx9Tmx
apWDspPxXEFWfkxlVcm7JrH9WiccrsjFVscS+DuybLjwOmEzQPfrYrpvYOzxnexqSqxi4xbIbbFr
5lLXBmc2Sk5Ep5yMajKSiQHOtbQ9KC3U74AoELcjwH1mo7sQ6juTkPTUMc/FKGuH+SVn1CcpTCzy
6WjXqr5vSjJegpP9R6IJ42RN4bLubSMdE7fC5DfHYq+Y2yQXy5clRwNJwe5jVzW7D/JGuqSxy0Xv
eWlNMILMjMRDXNzkrVhqWuLBrlqX/hYjlY0kL0aqfcZHu9BSls04L4Azq4N7F1ok6tN26Jr3ceGd
k8feykapTXdOooZLKPZmiqduB0qAOufCN3tmyRxpVoqMevmriZHnae749ODh94yirIw4kcPJcspS
IT+E3u6Z3YjYxa23ADZs468XiLovt3ujBgZLiVR/MZ3Ytt8QZH0tOdaPxqDmEiGuN/iGdrlBz1MJ
IvRGLJFHsSwTvGt4y3QUjCtaKoEmtlX7KVuciT3Im+1J2j5chldbOyy1uVfW0jWWkxK6lPCZ+iYy
eqnc0fQZYL2qC4R3YpweaBSkyxPNGy8M6e2rCJTUEEzqJRLH07I4bJSHwgJVRKNAFvyx4zuivnF/
mQqHAimumqiEeS/0MARNvGeQYfEo38HTOZhOeOxS+UNC1YOQL7/MEiPcgLSnzpWnhc55B0O3VnfV
gDmplSLSA/wgueV3hYHnEQGFqbwKzH/Sz/xuIcgAK6eOwssNGlF2SgcJpxmCwFPuA9mi9ZNnFJHF
XyMEJRMPcBhtspZrbvrj3iNR8LZEKpuk7AAFn90GDLb0UD8N+uioiRX3pBbkfQNw0JcxBMVFo2i/
yvQ0lvqQpWRiKWaNtK/tC5B2aaSDb1J/0f1TmJVc0od7lVFq0wbpW97KUcvTODnWdtgfNptDwbSX
5D5sI0MXDkowbfS31K9da7S7O1WOTM52Ic1HgrE26DP8LgKoeZKRsaI1nzp/lsOwPPw5siwhlSn8
ukYlzQ8nLPbQi5ROuzFvkMIdteZ/66tceeJc2Z/cNz6K2MViyI9XuoCduJCNsLTfI63k/O8u++kp
UAGnlXfJWDR4b1RaYq3V4EpjkSv8PEVou8KCk1wavbVWKRNK/304FuEqpJrLy4GYlgJidkq91co+
mCHXgjHFMarPdc7HvCYEJo8xEoRy1VXevTWu6ri7DH0RgrYDZzyhvjoLnHsXA2uujyFR6C8Yznjm
b2sFfi3mtDYVL3B3h84hDXErNKzF+LwUuzRA47nlzYoCniAAfxOJ6MCsPiXK5bVrSs1UmWyMimkM
VcdZaqBHeLhKv+Gkm0trjcfp38tEnpxzBNMkkUN3j0wE79n+dX/NMOU+CsB+e2FKxTjs8xiC8xZH
wCO9T4RrtRWzPWqRd+FYcw3qGqSy8eMruoarw4VXdfSvqkR3MJutZBs+npAraUbXN2BEcArINyJK
y/6i/1KarPLjswYFHpZHWkRnhtRZEZvxbOT/eZs9lyHdDSXlUqgeeRMnoQ0WDdyN4P7JzMDDKHHH
bcbKUrQyHt/T4p9lPmalsPSSHaiTx8lccl7UA6Af3R8EHkeZDmoILiXrGC6nW/O6cPtE0Jz76FQw
9mAKbDT4r4Nzx2AzeeUe2+KY3rfKeEDEByWGBJshmuEAuPjeN42RIF9sHGY36Cd9kPIC6oLZctB0
VbPUnt43+sXdvwS2GSCKJoLhY+xe+GKcBUMTp9RZhD3lkEtbd9IGl/pDpRUdXg3nUIC1ID7LrjWX
dCD77HER0NBlnHx8YBBaIUASCrCL5NopU0pIOaQjTul7U2qNNo+U5EgsCEA+Rqzyxk4n5N0nVM9c
cUO4F31E9O5W1JS2rqqKoUWbV8aUl7RdO1ZibrBs8NqGcTIun0s71kC9hkmwvtto9oxVw5ikm4Ro
5tRW56hhiyUfaleURKJgwf6EnE9maaLmS7R1Z8pGy2IEAneVgbYPK+e6UoeQHPUnry9NZ2U+IT5o
8Iu0cgN8a3rQXlC2om+G3l6kDMcsuEb4z5Bdy6FIQSA3YTNdzXeuCjfpfz2M6dPGrhKMmfM2drLs
s80UZFz2Vcg5TGhr5u/acDTmzyMu/7NMkQhb2dH8enyG1M7SIW6P4nK9Te2kTQdPbO6lZtGv1eig
ClqhqZ+YOgR+IWC8gj9lPbxFvFvjDv6IZfsX+B4NLxavpyJf8WCq2BuM4X/joo6Kd6b30YnJg7hp
gObMVvR4uaNoZpToOOaFsVGMkPK5fCNWH9u0DkykT/FpKD/qWkTofEyTOwxA3mOwJOCpzeJYqOfp
dfQYtwV0fCFWmhgaKhQQXydDddMtj0EBjO0Xun1M3JGrQh9/VdbAUvER/fmnLo1oRNSNqozAVvT1
rucvnqKRpPmIeUulP5wCdAf9pw3QYx6G7ytYb9VrGo4UTPgtDwRF8zVuBt9b3ROkUchylGg04F8/
jWYYGTnrNljMhfZy8mHJkkzztirRRsZ1ZsSgOeW6h/hXHL3V1sRgjZ8mQabDcl5Wk4ZB5o5D2i+H
zfx/x5Sf8kxNgw3BIUOVduL3XbBEsQ9xBe0b5jRbidTcP8p+9h0xwehWCUZCDOlQDrDyLI5AM2LD
7Fj/ongz21W/9Gws/3Yanld3EY+qUIqKNc3bKUEW9p+YICxeWZgUN8zY3x3jY5yM1cGX2hilvS8H
04ZQTOjyFyc7dFa0Fs0i5b/FxmdgxMSeKfZ43uBC0d23bYVwHdJW6Z+tZsdAFChGSGfsr5oCF8nN
kNuFdoVIDvlLVp+a7QD35Xza/ugxro0lAAhRERTLe9GIYYi87FjpwE3D+TQJhtXs5tz2W7B5KxeH
0FNdGjQ0iTGquS3ljVQR+EAar29Ixwp0R3SMo4Ky4pP0IwrJpJmjsp+HUTAdUm1VqqjtDgaZhmAG
9XsA2qaGPpapwBTXji9DCV20iPonw8VxGfB1JzD6ihHgcrA5cBHhUlwomM/kYVNldwylREQ4mnGj
fvhazD7EbsFb1H9PwJRx1I/Z36zR2V508Zewqi+W6BaEFD+3au8EeGa6ReNKWHhGLflvxQmYtywX
3Y1QZKTnfZPTMxVnaMMjiqGUL7eTcZLSxFgnwVzgAX2bvaIKoNpEtHskAVpa4uC+voyrj3NHrWEw
P7OkBcEbBqFzr/BFTz6kaLyS2GWrq8SOm6jtZxe484dJzfgllloAlIOsrAVKYFcvfMwhzPMViSWA
ZUbf68CskU2bN+S9UoaSvZY6V21wFlSqQFZjCU/mudE4p8s2zGhSutjgomp2MAW94yta2sXMRqtr
bCosJg2YJuM99qFlFA5n7WFS/DekTdAyQGHjN3waZ0pk5YryI4w6kHhsguc31Re1eNc3MHOsn0oe
Aj8P4Ekx+NP7VZWXG2g3qkVo0CK0cfq0JlhSS+LtHbnDXdOAHDiWj1sThlozCJCKgYtLnOue5luP
q1wIiabDaIxirNcOgDnZ1MzjmS5WpjZ8lLo5C+h4F+jZ9atAqUS8geJNVf1LQNqgACnHnP03+FYM
tNlW5AP2kj8SaMB5gcbI+5jrHk0oCQE0zsP8RdHBzIY7dxLXQ4L5+ZFf8jP/wKwmt+94uXK5j22I
PcPyjAMk2Z5hJFJvm0NMDgFrKPiPhl2YRiP8+aqgoUE8u5/GZh9pJqAOqfg6hrGitVlqawba78AX
eBM6GTBKsbuzkhvqhB+6hc0pP5F10gxOODkkAvSV0QgzjsDVRzYlimrkt3UHluRN6PGZx+9EW4+o
h7nI/e07g5VRxd04FPcti/6gHB3QYBS7XG6LcN5IzNuP4Togx+BCrfS/mj1XBHYBXVo1BVpiT+o/
t7O2pyERiRGN9qzcRtIhpeyJyJ97E8eNKk85xTN5htz1C/a7QB25Bveh9y+A5x2WxfeP/wGIfJLM
X6tGSsi8wrYI8bUibatbRYfyNNpstJHK46xENXcWfdVRFV/mB74IZ1Tm6MQixxwLZLGT0qKJ3X3h
3bY+8R1zoLzADROBT1BFnO2SX/cXHM2VZv/rBeDMem6VCeN7rqQG56utozQzhzoCIJ5h0zVN9cBN
lqZY7mZHbTCiSPae4jUC56IWxsWvLQSDoHmjuiOcFvWejOQdUJP60SdV4+SaoVJCQgQ3EQ2roiIy
MSHnhfTj6eiQ59abjq7gRwoXT0iTT1ClhD7ikBXgfpUArRFijRouExkQucxeIrcCJlp3FYY21q2e
NxzojDR/CJqGyWCPUxfgs5f7Pdv4BZo6ftbHfCU8Ac741hY5xT0DMm0W3MUVslbhadTmD/a1rbta
W//3GSHQeHkg1F/OzvjLcmxAQb7RNzE5dvyO3HXYUmHUwBeGEYxjhBWXN3AYhgirLrhGoWHEbZ5S
8YeXphZKbVYWKiTrGU8JGpVHugESsv6UX5vdPhlUElyONn/Hu+7jc4xK/1wRleJL02q/2MGb2XNS
uc9yQcrcygeIEhw1aCtBvaKM72U0+in6aKogNScofyoC0I8UZfS8ggfviKPcEQLiaMZZp0WJ5Dlb
I2IAjp+BCKAdHdw9Bdj8+SjyAUDipaaTAa1v1u6p0qXb/iE8ZP2SUebkpZPaeys+8anYOlj/ut9l
ZsNAmaB3qMXQdJbR6aXFW4yTpmC/ZLds6OS7Y+x/gc0P9wBDLfF9OQ4JqCpeJU1mDuWbB5b/KGp9
1lca//+IEfyOSXo0IqC0B4sGQkQx/zXjCBmlPjRw7ErmRkI+I8GVeKOwwAv5BwMIn1Ozlytl7XWq
l71q2mpHRHxEq4HUFA7x4VODAAjJdeIwBjun4FcMaF16rhCGTb0MvkCoLoNnNv7RZfohQgQ5MzME
YSXBuwhki3VBw7hE4CRfM1balSlLTqqDktzilbTAZnjlvRiLAH/v/S+ost/pr922bmcpmYo2xdqu
X5DO1DMDAKeqry6b3K32TI3s2hg2aktWTL6rwgzq9JPyhsfF8WTGtoPFdoFLc7NC5qL923gGVGHf
RbfY3swfErv4jZOZBwC3Wbttxfdj1I9xMLYYBipV/U7rczpuQ3MSro4GStaG6DmrdisjS6qSEUmF
rUj2JZh9jwRxpsmrVmUvk3WW93xzxJBFLMOHgEFrkJyPqpMilLxTy/weBM9x/QYdt27kL+uxf/yf
lF4yees+RDPHm8F/TtrjA4BeXpRtuAolIUmk70CvpuW/XgC2hlw94maeJhsBn/No8Co9iRPlfBJn
BSmRCE1xpI8JjHjHoffxeNZNMwHs6O1NFFGebwq5v/ogZUJ3cna78iMhEynSwxVXej6RSVAwo0Zw
vhRYxK63EJmbnmCJyozlYeRtXSrV2XEodgB3O5o8KjxoqFy5l/xeyiuVqRNEDqNOEmlQgrG3A5Dh
Q4yMSMl/1ju6TJJ2Hgb7BCxRaKpb86gZjOTEM7heZqHr0m+3XA2FYg9OrA9EfFuFnemLljjXpCBT
3zskNdAogD6LRuL5eXO6VsN+/RoKNuz4genvP34duMIAW3Vig5E6zl5S28ZIlSqwKkMy4Ho9X2uJ
ybh6DhfXkM3DksmGctRnKyYAEDQhUTdyCRUW3gE9/k8kKjDgpxzOnGoW0xs4RgnNOZYoJI2C5BqN
mn5dUOZny9gjyW2wlpGYgSZLLOZXpAFGzjbVJQfZWrHmmjNl7aehTf8AQO7V4ljivH+rbgff3q8n
kD00s0Yu6w6Q1LaR15SQW10nPzwlOGfeFTjLhBWvEju5//z3Btly1H7sHOcZkG0lvZFy+QzXzOpK
9yKQQZWQKRQD6/VaharWSG+IIA4XbHNBE6DlbWn7iQcVug6wYhRSCNN76EgNumE0rJ2k9SEn7pur
2l2MTaCQ98a5rCEcJx8hTqtMB7wW/kVJ3kF0JeBHREVWZvBC2zUGWiNaUC4tgVMMewEoo2DZRFD9
1rIL0r3Fa1AuQ6zqJP7pPd1K3/6DX+jDBkAhf61eTH7+hrMxNJGHPCdO2y/+AlKgmu0DGqmjKtqj
+j7/iQ8yGlF59N0x2ZTWUG1jpZaTBjcqPgmH+a2CLODp76LAWNhK2+/HzyO4gQ5rKEU7UQBtwSUd
1t+m6EK+OleIXVP2vShI1KYy0oE5YAp+zVDGwjHz0RCOb048hyB7Nd17IL9r8youC23pvjCtPRK+
MJl2s9YxDQ0SclqwZ+2LHJjFlECu3sVsXeD3XOC+N8CuCGKxJZjloLym1cj4LODzf77DwpKb6gq2
cwSkDv96+/8jUBZKSzhoWcftF+DMG4Mj7hz1c7ZJzwaMVTwcIft8Hizo2WuaE8ibysfqwvu2MmEV
RXrZJMn4TrQpRAQjtiCiXGBufXRHHUauJ3ExbPKLdJW8Ryv+Nz9Ujv5Y99kkioA2lM41tfSLn0gY
myscJwW8iR5I444/k5tQ0k5wF2PMZLkyjF3yFleGrw6zzqj+JVjktngwubzPwUWR/b1waHT2TgoZ
2pTPYUGg8vK1sImg8hpsaWFQ8GtjPDNilcy5BkTJGbbuja3JzDQ5pPHcyeHk0CwK5zBrhkmr6Gu6
r3Gwtiu5ln6fqhriaKKuPyHSlGO5TYKxO2OsX8Nsao/TWtUCoHs1Q4Nn/CzlD/RXPNYbJ+98uUyp
CHgN2epAhn5OYQVUPpz/xcq4CHc+P0OCPCJzesOxZ+vF2qIFx2DjlWYCup6ykdvyjJci2pByoHge
67EAVGl+x6Yb8zfPvfsKdUMht9FJBeaRN8n6hGkmluq80ULsP7yWdWVm25oQYx0TxWb0c3/VQZd+
wLwAPHKBAePFYRe86Fx+Akmw2CmobVWqlK7n5F4eJPNJzHbuyPdH09dTQpyIp/sMfOgZedv+PgxP
N+2fl782t+VziFB+6oh2FvR9i10MnAM9RlhNnhKuBAkyzxBBRo31bfzVp+TLiok+7XtFftIizzKR
h8aFR3xO521SfIrnAOxOxetODJwUNYSY99GPsVHBqUJj+oy1h+RNBbw23+6jYJHEGYD/RS2NJU4Y
loXvQBI5vcOIyrSu7ERWu7rlg5sKFM5NlO2yXQwUzX+34SYND0FkfJF9JKb0OH+jeqexhlvyHvXh
2wXFtFuCDUIP6pMG8trpeMMW9UAxoRrtS8BJ1bsn8N86W/UH+UiboStz+mcHLbrrwII858+OGprs
JibD34Yh6KiHsTc08PJwSC7MDHvhpDpuT3jDTBKIQVRhm8Mof8QOnY40VXKs9Y+FOMAn0VHHYT26
HtJPR4n9v1ciAqdSs6GVvyM6SgiizS29l5NkQXJoNMi/zH4aYmDlD/UCGVg5vVtq/lcf92mAA54W
mg0mxozppflIGAEu7sP13HoUk6U7+4dmRdfgJ9lsyVEWvqjKE4DzbpU7+K22sZ8QD5LEt5A97/q2
jX2k6fzgtViig7Hn0SgMifhteijF4njfspyt6tyV4KsvOXJiEVU0M9Vs34x+8/R4aJLQt8oJL3li
HkQGc+XLigrQ16x+X5/KaXcxOkNpNPMc2Qx9ARZssFD5GIS5xyXxuOyJ6sPlk35BYncHhspMGpcG
rRnxsfjNFVJ9F6ANs9qUqJHtt3gzS8qO+lYBMFYn9+fKR2bE+1Us36i1gaI2+Vhv+/YY4zL/L3gV
G4EE2X1GT6K0VhVZXzOFJIPyYCp0w7aYTCpkAZSXae9W7sWhfxV678UaK+0/dKe7oW/NLL/1Wy2C
bRPkABggWfbXxQuRgxmeV0gG2c7EPj7Iu6pFNQ+Y4+nnyVedn96wPZ1RKDF6deJIjhZGBiJgNbyb
7k2K+RfJN0MbE+qJak1ilSSHt+Swj2A4i+jfmQRx7N8ujN4PBYrG4fp5T0WjmSOApZvpGKbxPpS1
OWd9m/NuE7xxXMrSdkkOalCk5jkvIBSy55tmpfws0ZrxfR6SXWszJgowzj+o114+2epS9GWCHD1s
knCX0nLaoNd8oOyLSOFS0jW/w29L66noK1Fr2h/jJ3Xd391XF7t2AyoiwxPROzKBh3B+CS0fhOn+
03p70OSCmCCmawVy37LX6oAFW0mdaR1G5zeNkxnqkNgK6ZfqsqN/F1VHnVHE8vUhK6FHRigpKlyf
+jY/oT/TTw3bSnINzACS15lIUF7SBixeetZxqGEL5dwcpc4sujQe5kNJJCZ4z/OY9C0N8pTfFjtG
XtUChnZXknu7r4YhXiF2i4eg0CTvoRjr6W+RfO0/j11YmrmbNrdXtg/pkzF7aLpMlnziBpEVZgWD
G9ukCkq/Huof1PgI0ep7AYrHYv52EYnicbFyAOWbyJfTS6kZ2x8JXjVLfcoVOl4RqoojRgcqnIp6
FOS9xCrdv7X7itU80rIDwE90HobVLaXqm4qKzPPgI3BlCOqvU4c7f+Q8brwCqpvnXbv61SXdrZCn
5BDI7t5I9rrzYKfmL+CCIYij2PNCBKEy/MxwuVCL7iu7hvY3aeuKdX2+mAf1ueKNZ+CQ6DAlw8wt
YlkX80VSntU9zzLtwQEQdbImSDLYZf7eJj2HYCBvrRJmMQ2dY725PCr5zbAC26lcketf5Vf7KCPu
/j4gB8FwhvOqEgKeL+Q7Ckvkg4bPnERmZ8dH8b/7A4/Fb7o4RNM65vdASQ1QfyYZWArLnvMVlcvB
OjvusM/FXZvIWGgEQtFlsfgFONQTVg2irTpKpPcQX53RUP019YVE7H2EKgrhPjNKOqGiH38rBupP
cz+eYcjhNiG8V14d5OSsFj0dhRKtugU9x4efas9sqwt4Ph4aHqzy6Z606w+/RSb4jY6sgT6MiQD/
Gs0WzyT1jOlzDhxBaMFsZTwzraG8Hr49bssglnAbm3eXHCNMA0Qk1DKS4ZThbUOYPinqFp9StGOJ
7aG6pbbyKgBsD8Ogc1+e7I+8exnxuFzb6abUDJfOodmQ8svC8OwcEY3ZIegBjnGmBkwbhbjP2dQg
BrNIfmQsBsEwe/ODNT1QJQHvWR6HbEvErec6u8XKBqAMCoU2X8r8jG+d4M3xdEjfTsQeOLraT+Ve
qgUOToVaEYpQ95o3qFG4fmmRIXXuUA+PXy4P9qVWueqGRRJt12Avn/anziykwAF+cVyFBqjbny8V
4HUSmaYTgc72nVaxsiq9jrBN8tyA+YfIAj05c6K1T6Lkedxg+cXQj9OGBXnmV2GsSgdFHaV1H1dF
8idnId7rJE/IGTQAAd/JT7v5P6qtaTTyJFVphSUckYt6/BrR+gLhuLFjQmhp2rakuhwISEkwPzz+
1iXm7fQF3PpOiT9CdNuDrfb5hPlvQZz0fkoCQLxqIRFzKldNkg9EIaJaSKRDMM8eh41rW1BXqxyK
KOO9VY7jPuTPm8/VjQIjgwjIzc7DOLjO8P5uyqml5eyx93uFutcfW9R8x6jBc2BXNzTOH3F9FefR
Z8GIKzxsA0wZ+XBMsPEnEbTJnmz4cc5y/T+/4aHuO9VWNI5rCSyAZN11Vd/Fmt0aNaBt0kZpKLPv
rZ4ztkBlCjLnpK7HwybbhRasGhwex9u1zj9j11I6FIXl2uVTddJfOM8/RHX4HhkKFKqxM7bzWTUt
fNqSOn3CMQJ+nM4CicGKE0BoIJY4MeHTzU3d96D9Sg5jfmtXhLbM/32YH/UPoyJaEcZGyi2ZarbP
MlFxPnmFhGeadtT7AMiWcKBDTp67VW2AgVFE2qC9Z1Qooii8mqiclvVwldQO5KLC4CKzH91o6ZNE
0P5ihlcB32I1etsSBvCEwBWKMTh/DanHgsNPdV6ndWBMBCRSdJt/atvzTY31umy81CfxxiUNAuZJ
2npy99VIjnCK72yGbT6lpvnLL30JyjvEfkaLKrQncTmgIVnoQIwVW77uoQ0KCOT/oZq8OJlXXguq
cdwDDRf53jxZSGSkbZPAVyQ8EIV+5zhkbetQSa9LTPZdyWukIk50eWDr0aC++fHj0Rzd+wg34jol
kRnwJHILAalgG3dvVyxdqLDWwBNOz/Fr+nbTGEn0gCKcfbu5J2sJqB/0xruujOOR7cg66BqMGOrx
0o5wzQbORvYs+p24atb1YAB4PxiSQZHQK0CVBOIsYSXCgirghiJzCpD7uIHmmvt7Pw9QR69fJGBp
b6fucF5ZSPQFqyr4iJB+Rm9rnRHRtYAgharW4RNqwN5pNIN5mKjbN0nAo0k6gwMOgr51p4vM4G9c
wabiAuMCBXKTMe2Bg/dpF6OSYtj1l2SDvDhis+rsKp5cE8mfIgnKieeKMHAl5vwca6VvDo7k3ZO0
NyzPXEAe8zsCl5A5uGQDzjHYdEbtGcrDU++rm01XY55/uG1DVNzY08maZiUbZ50ijDFURO5ReYDi
fY46oluozjZmMLI1Dr3FR3IjmIR5cnSDBab7EG7BtoqZs+Ni7P9A8vFlDzziPTL1Glhf4Y8zFpmk
kwIdUk5eH/2hCNmu8KQQE/XDI794UNsGJZqLzZOf6AgfnHyJAwqqs8xfiUah4d/i7TKC6d6NEG8D
M1uYOPp/e9BaL9clDiCmPjHBGN5FH+UqrKvzbXzfT9e0+V070/dPyO5ZTZ+nwx1ucEd05pSimnZh
MAD+1dyKXnX6lk4YDaD9ewI78oO6wt3HoNgGTvBtCJ8GP6+wlBfzWcsFWXnJMBAdlIMkXZ9woHAP
970LFCe8yyJ9g3/UsbCWMF8+TQr2g6Nz3Pc4qRiNWzsX0Es5cN1sVTTCYv0ccCxTI2L5Ke0Kt6qg
5KkIdIDEdXJ31iyMof7Ntd/Rz9BQIzS3R5LzkVLOVQHFAuIu9P2tlt6gfCIxYmQy2tRMVMhat1dq
Z4WOngp5iihSesRQYn+MeRKD7/rQAIJV+4FcUYCiZR+IGZf1JJD/5HCgr17sAmQAOmDM4YqOa0/Q
7bE09VzCV9kWREDyq9BSIg0mrumQDaA8n8uUPvZrWLt6JpdUEceG+whNaEgPoq1hK+mja6F/Tq+3
0Wo/TPMRNQPaKXHYiRtixc/0SqlmZLx3sdyph48sPWh2B7dNCHwOj+vAcVseD54w0iFaAGCheCf3
GXJejqSB3at7evUq3iG6IIQhTEtqzWs5v3aX+W/gM2V6J5/+uYKYey8PJzfqNfTlStwt80qgVoOX
13sQbdQwqspySxinqVz9vSqqiDIlKGyS9PBnwqH7YsvVNSScumal2kVxaJdFDshnXnvDuMnqTQuk
v90m4ccUhHGxSJuXH+02A2zv2wRuGt5490XLU9pGghPOlDlyU6mQhrapAwHRabV0l3ubd20cAsvl
BrYjPOALly8/lHWnIHG/Yhm7P14C4xSeWbzueVSZmfCea9dklV+3zbEF4LSdaCEi/hIsdEA0fWE3
WqEPeJ2TQVzLVeINvtDBns/stiRABONdLqke1RIYKrpYw0l40uBbE+aA/aGRrIdNeTwulLAczcTJ
AzWh/Pn9XMSeg8t5BuPNA5+jOSgnZpj1Z7ghAINGks09Tp7rQYuUHyFX4RWhggLJC9/7/jR9fYpz
fFYvS6HwJZtPmXtO59VrKTx7Kmm0bXXtw1Rypi6cVgqSCLy3OadTDvtHA5h9vYCrHG0CG3HeTbWU
SQUH0v+sCvM57WSjUfk42VPYBVl/hU6OEa2iNpJdgrz6M3R4kyCqoeOo8K3/a8txy4aqlPNz+31w
88ryqNZC0kI+nn59EgDRFaLyuQjwiWzZiXlxmXx8Yi+HfI1Fvj6slTy7std0urpqOLOj79MIA1w/
80RwThQqKVcb4xl/+RxeTTndGJB3ScvtXii4tqP6abdpmsIThw8nVXUqwjQIqK+wGxo9rrq8g9Is
nBP5IhCJzpOf5Xzq3HyO3pGBF0dWllamDvjC+B24LkNHptJqPXBMe5IbWt4Uh64XOwPX8x056I7J
TE8+GoRUo6tpEiqMN2BkoTQ1KTmvYDwwJ4VrR6FBervLtZpY4jxKmyp1asulSOSt1FDlz1CYfl6W
FlCXcXGv9N0NzkAN3ysO/FavN9rnTM9GxhGIL1P2hNEmYCQx4aS2MHhGuhfNTDIEo8yCzQEf2CaF
lLIJAzAm/IQRkOb9OOMAWwKgE9bghe/rJ3kBrQop9QhPz0IpmMvKfZi5NX8Ux+AfEEjola3Id8tz
zs24djYtUUSDpPMTBAywgTqUPbK6HzawUfe9plnYyr/YHS0R9L+syLQbX16S6BQYMtwOo3mmSvyT
v9rjDhMwVChGb2JG3pnf9ycZKqrtcTHP442DYELGQaXeE1mSOk1+XuQ4Kk9zJNK9azEUK9kRMWz5
mFimSmYtKp1mA6fBbJRRM/l3jMTKbp827Y2yizGixHShDE0c6JMQwVHsJHMNM20cD41lBs2uyWDc
auYZ3A4KwxiZVybGDIvuk+pAucEuwsXV7U406Tz0OIb0vUVNGnGE9Faoq7UQj+oId+NC1RxSKv5m
iMZ8tyBCzuBpWu/vzTmSHt/LX/9mVrJPmv4QksdeeWyu+bbkpibH8RCxyM6p7LlzCtaJxde9GcEJ
knDUFvgkHTaF9AYIJOVlpghWRggIBuHqByvYS6wUBws8RhkmwNMGxvn6wiidwG707TdGkLVV+QCK
mUlyx96Wk5CnFihZ7l3EABUmjptxch3BbuepFZqsK+4Jow2VU+EqzsPv5ZAjy9nkexSyEZG9jH27
jRG39Ng7ZzNn2i3Raa7ivjad2MCogEJ0G6fi98s3sfePVRjSLV+NywUBgI36InkAb5Pcbqlgy2TY
znCvhz+qHNgeTLu6IqH1lp25dGhSra+UJ1nI2C5GQUYy6bRvAx5Ws4Kmd2Nctz029izm3B1I0f0Q
cOs13SwBUTTh+SdF0RtrcLiIk43v3AFWi5W1In99xhBvfSgGtzTQOgWgrOpgzK9803IE3nV8uVJG
b/ciZWgCzd3ZViloUZ53p/W7rPq6jsjbmwjX324N8EFE+lWu9MeYFAXXDfZvgZG0mvrUrBmxQWfh
GAxT2Cs/AtoWLWgSXJCzUOCCCyESMQn7Nf9mgA2dYHFUi/eDh6us+e3JK9Yj1j+RWQJt4qUU9QWM
83EMjmTBygPMElBLN2H8By9wxgFew9/0ysADvlRGwT/R6AURTR7c0hc0FtthC9qPN4Zs1HzpVYXE
fRAySPp4drullMNQvtk3eg6IB8u8zS6aQ/qqSncCyw0TDMRngp/O3byA/b0k7RfGHxz75Qc5E9Oj
/E/rSecXhkB1OAJy04qwLD8PSqZ4+DJ6Q4QAxq9cbO5WpRMpP+c4ge9cwnGwBbUYJMJh+H5goqIO
+x/S1N5imCw8BeDb21qWx8XIfE01SoP2CCrNO0bwO7puYa1px2jWAA1qGERKGlWQ01NUIOHIceUM
RfdlPaznYiQlIOW9vZEMdKT13DcXZUopYy9L2tYtiLLgYQj+VPTERaIfHLTOMy7vcVByxD4AJ4dT
9Q+7BI47Lt4njFt6EgR9Mw1aVwLgJz6oam+CE/MhIfElshMu02mhU7VjjJ9s6hoVTCbaWvcNcKSG
sa0Y1vDII2KeyJOED333pYudDOh1AENHoEwuxdUaztXuMRG2YF6l2K4iAMhyNIsb9TvwglfGxwtJ
eVJPVLVmJZxeo0VQJ+YfX3+DeziQK94dcQP4cAQ3/Po6nnANg17GG1BDnCA7hR5DLwSG/Gcytle3
MHDpiQLRzMaC67Jh2M/WT8IZ6RQDCL6qGLD8KZNX01Jnx9D1v7uXt5S1IydEEakzP0i/+8tqp9nX
FnsxXd/w3h0grtDTyc3oejvvEFvAAvZqiqWyvobi/KusVOcMZzTQlxbkPwQ43y8jdAAZ3TaQ/J9x
FrL0II+i4RMcgcOSY2PaKCLkDBCJtURkBAnjSKTG6tjSYCddiz1oWE/AvxxqkKnMlCLZjWG9WteQ
+bXq4XPHXCNbVN8GrW4jwlN0FcwFPiwd2OGT6R0uPgLKRghWuh5uwh8NvIM0Y07tqGuATobY8/dW
/d+KT1cqdb5sP70zHMDacP7XoanFdmuMIsRNQoAzKlPBgWk6RTvCuZvWTC7ZLRAAJnmwyl1R3Gfe
13PtFZTtovDJGQ4V/vqZFL+adfvdEn86xAMOuh9Gvf5oEggBQ0iUOtyPDjFtX7Ngxwa+7mOaNY7k
OCpGmEALkENtca4mS3oG8N5Y5P9UUmlHGwzV083j1lgFQ1TuvSdsDYuvQCCOWzI63LPgc0LQ4PSH
KVmZ8cg0n/u3Ny4YCrCSqhVmTlm3GzrlQwL8RqdF42quPgKdtlawqQR/zCWJs9RqWJ9PSNsQJJdR
JP/8EPPiha8yDhVUktGdrHQ250Vrrn+r3TIXpl7MzaNYzV6TmsKnTVGg49tB3BFcj5K1RVhOvHTE
pttdO8RhcayQC92fQP+oRhxjEA+bYDsdXjOVrY+VFzNsbEgAa/6t2PyPbJCeZ/4Sz5UH1+ZCc2Mc
RRZH06rQNVKcrx+OH630SKW98mSpXu4qnkxDiVJ9arycDWggcld+teX4olYglx87P6v8CR3B0Fz8
UDWyry8i+Eltht53O6VwdngrJye+tJLpvwT1vtRAfJ1lPP178PHAAKsLQT1SHYDYdGf3tBp2TrEu
EhKo+XihGMcKwCqSsvHryhXCe8lg+1Xz8cIBmdn9tCRmT4+oIyl+UeWCTJdsKOvzv2uq28QXjMVe
66czMspl0Ur3nEkgXml8O7Z15XeMw0N25nQiQaIVhdUN9feJlQyY3bZTqKQPmD3h7LMD2WueWzaq
OdPVQEIvuImgvd3UFrcw3Dqf9Pmu3Kgl/iFhhVbiT1i/otq8NQGouaJA9eaBUz+7Kfb5Fm7q0tmp
3DwuOfK+xHZk3DDjGYL5Bs6qRinlCIbWWV7Zn3KXolO59tUC2ppX4JqHcy2wL4709jZgl+uGqC6X
3wW53CQDApO4sqfviOr/5X35/4j4sdABfdObf79C7mokgIHMC+qCbmd4IFnFVpTfXk5m/GIgnrOo
wfuP7ZUGIdfXAR2JZjUeKM6A9ufxGblN63znvzLdnD22Ybc8TnGqCxXVeAmxRTNRCGOBk80iA6KJ
Escy2p3Vz81cpDPVg/7vFuSp0StANm5HCkdZ+mPzIAO5HE5tAgpZejjpv2eWRYw225pnzwjpYNpu
BhBWXzWMq5h5/wJmnmjJq/LcTiCxEO7GnKKJY/T+//eASAf/yn9L6ODe0OmLGC56sH2fkjHvoFYw
CmHqISp8yPkUWZTy53azUS/cPqRlV+TVwRKUA5LZlijClefeXdIU/vUcHnRPLvrUGJJAdLCmAvn0
D+YkqhWTNtBkDOugQYPHcw0yJBx/EzpToexBTLVcr//aBtctVsPs/0uZOIvkChsIDV//MOXqIxf0
i0EL8tjEL55vmTIMpjoor8sSpJbv/olF9rajFl7Gd6o3DjMHSfcSUI+dxh85FXkNXyiGdnKoWmfr
UtFQWXlJj0c1Y3sIQueIVZM/Oypq/logznsqN0X2UXUYlJm/vuaajP/RDLKLC55Awj33HbHn/+h4
xxlZcfn+hP09vfX7UU0Sked0vG1eas8tFTzRvqPfnk6ss0jzbV6PFNFRBoZjzHFgFCIt5I/fnN4s
UrgC6wAAWEhg2MgXcYwz2WdAYjDc5PgOzX20+sqpUpxS7hkvUjLERZz/ay1NBnHpbZiT6ywCSMhO
G/mq2XJ3yooUarRGB3PrK95883TUdsOlA2WzyOC2ZIVDPG6Y95G3DwRGxCOYWXZdDNp7t+k8xw1O
XiGUVe64C2XITYgfAP0wzcRQOStV4wcnailnCgw2nImADbKXXb5JYT2p4X+Dsjhik/GE/7XteJTt
WuX5aEq+v/z/oj7njQ9jQAxACtUqfZJhqPzi7Fsbop9Zt83cMKvLeHDy7jSXVziIOQ++QLQvecYl
YmtGmRWWwkbUPxHXwCQnPAj0WLf80M9hNq1rYq+Enq5B8WmDZhRNe4kZOMACjmq/3AjC39hoEf4U
ESjaFlFv5lhuywViPCxqQIvSxNKesr9k0fnHDrjmzF56fPgJFP2WHTGShJHEg9mOgXNUAWcJa/2f
qnZgUPPT38fPV9VQGFvAos/BCFcQVXlwy0BlnycSVu5wf7mjzN11jYnwfxOxmpvOfrYqu7ZimQ86
H9NgKxf9W0lhJ49GlZOPvFkS4yfEFDqvrolZQFKI1hQaQfejw/A4zBx2VaiY2xzehJhC5GXGoFYF
ULY/FO7VcBMQgiK1tzIOwBp3JLGjzmgMvibW8Me3W/Ov2ciq6kfzpYvHmQRRnj37bNcfn7u4HD7b
UMpl4vyAsSiNNc+VCKavYtAxc6aCzWpcf8GCER62xUriWT7lCBGNmpxMqFWj120BKZbceOynl9so
f3AtstEslsvJo2u2TxR3s8Nknvm6BUJBwLLLKhtB3JVMZzS8bwqqZouf1ovxIMeTofcZvpa+scL1
LTzEI5Mz4IJuVP7qSAAxk7srspSAde4PFNJqPnkne+Pv80/yqzmrTibfD2/2nmsFC9I0s2GLGDCJ
Oje38IWNlgUn7k1pnjHAMuyIy/cq+bc5lXPWn35XZ/GbLKkx3I+YqAbDyY0EwW6FIKFCo7UOLF4i
Yt3x69SzN7GEYj7w8pXXj81LbjQUbMpP0N3LFgW8LXwHxlk6sY5/nZbJr7O0lGPlgxsuvp2FgG/a
416T28MVFd5qzxhhacUcNjYjJAAvcuEUFahFdFiKl6selw0cJPnV9ycRpPObWe2scKdoKFfX3DX9
hhL8X9XDer7Htqugqp/P3ugSotZrsmGkFOSmiLCKCVQxJ0yECCKx+sHfIsoq2/0Q9bgtfif/0l9n
lbEDXvEWO5Q9gmTNGIUBv47XQVEfzWxKO8rSX/8W3SNJqiJrdhPUoVGYM5DA86t1W2Iz6NZGgbsw
2LD5n5o4vkwZA4roj3eB9ApxByPAKdOWPBM7NGTx9NGEvPWqyoN/iDHR5Y3RSNRzSd+RCLuAx4Hw
oQj1BtmG8SICw9thAtabNWGuAw1g65WwZon1Of8B+kzqL58wKxQOnKPneL8+4WqhGKA4v3/fYeP4
c2iMbaTUEV38ypVWOS0AhdhWsk5++5iY29IASPmhCoJXLo13bY4EkOLHnNImTOMFsrYyLI2ArEb7
+naHR07/MPfUzHJ9UllxmbUrnusTi1vQe9xavfQgWZgjGUJLFS8VxjN3sgGDDwgKadr7ADBw+C/k
T8b4iKVNqK3EkUNQvr65SAJTORhXEJqg3XbXK9PjHSHWZx6KVLz5ic8BCPdVLsPdnRzEFFmQuMzm
eRQXcaVhoTTa7UEZenROCoa2r25l1lHWhGPVRbc7O4KeoZrfWvp7kqrXHGcOiMAsS38MKoLiB8P2
2wD25N/rMWLYy4waBOuKjxOrdAqMHGGvSmadJ1cdJIpJdZ+C8EoxURHwFjWAWRYllUuRWZ+P2qCC
5+4vk+sEeAh2UTmhMHsGXYRQWUraaGJ3YJem9rsEPe9bumi+qHewO+qfqx3c8s6aDPBmOnGz0G0a
qGYomtmWqKD+TE4QSq5iCEOWZ+XDNm4f3xN1ccGDP6Gxcvm6lrkyNBzt5LwzZ6XuU2LsdW1vtZEG
AD+yB/+c9eH7Sjksn7IgrVjQPLFuRxa70TmHfrrsoHu/wUV62GAjEEEFThjWq02BSZxlJXcEpbQ+
Il95DwtIE0gFj7jmFC4AHixRVGSPcH+v3d+yYPjvaurYucEmZP8ClwnSteQflewEubeTWW4LiVBz
g0DoX9QvdbG5sOYtm+Fr+BZKIba59FQWxVQ0DGJa9aAZGZhUSSVwsIz0gTGcFno2lB1iMoEMEd1e
yDDB3YXMnig1xgWs9LTnBgFPfoiMu3kuioqiUdvbKFXW+HyIQe5PEUMEGJrPijjL6snywgiZ7IDf
hbOMTkpsk2gT2PV70qPIzl+jQwbndBsYIsnnkzR3SU4DSdFKIlPYwnwgaDskrpOZL5I7iDGLVgPc
7GKqxYkwIJ7uyNUddM4XpDpdhi6qE3DFZnOuWvJYTczy75YWt+iV5n5URLGREHFapRHmUzdasBw7
z1ApbmtnrPxMsyEw+K0ckyEwsZ/oFX/VIC0RNfmrMrrkFIuQVvtGPfQ8co3mNwGQZ6Ld+6Jzw1Kp
l2UYutYIak6u8UX8pccN6zCeGsiIqaCj6FPZCx6sCnfIX2hBgfXjNfxH1s6F4pdMxFvjKBh6u6Pt
PxvAMIU4jy1X5C9saDkb0rmLcdKCbui4aeycS7JHKgLK8nMJHkKxTM1bnqwOGK8dNx809L/fQj6v
Zvju3Qk+q2+9o1wAjGOiqs2uthfUOHbAcPNRWNBu/7WO4u6SwDgmXrk6kLgba8t78gBuOGPLdG6j
plO22mRGZU6z5D8UUgksSQf5dcgH8kN8EQLq+H4BoaeksjvB9bH2YOY9Bogtmcq/u2DY1j+M9SmL
SOxIF82BGgLWr9cXLcWFLRn3SsE1Q7sM81txWL6NN0FNLEsYFCgYvaK7OlfkxSf9kLtiuzObh/yj
yBVXwTkEEKI6dXSpBM2odmgSUIidFIs9Wi/57QXYFyzJkXWigIKXVVg+7Z2SkEPqDfVROANMm9T/
G/kyTnfdllF0BN42lB1AgxIXobMrEaBPABfmYHeBJekWRJsmnZGX9lslJ+HVbOjMSlIFX4aIhBh/
IHJ3NKP6IjU1HvOMAKP6SfmZPgc5PVzJvuSdBnDlU9EOp28C7II90eRoSci7YusQusQn8Rr1hDRL
zpEql5cU0TrEMkHxh7hGaa+LFFDujB2UXOmgKI5aA0EDSA7Pf6CDj9aW5XYlYkwp5PE2kkEo+d/u
uEulrip4TvdZQ//e9iymJnCH+4Al6dZtF+vWNqBCqXdg7zVrJB/kx7rhhUX4chxGQ3ZPj+JfA+ST
1juAcsBPx3R50XhQs5Jr+q2yWilPYs/Fs+A0Z5XBYB8utewgrFlr0GPIc3uFgS1cUXuBUkXr0AQw
YRfRfW5rPCkOsHZr0WoGGfmN8hoL/YimmOk8ICIpXvPsVLvdkeM3PzNz6V4tYc30RBweyQ7coxV0
7NL7GsnagyGWTtc16gLYlMIZqGA76pE/sg2QWUPM+/CNoCLCaF2hj/Dfm2oQk8unttkYOIdlG86I
Ocxmg322Gsa9KrAsgLyw4Fgp+hjIyjP1Z5G77LYBlc6OUZnuleRNNiWEbe/FUXknN3uPHzyGhYOF
saC6Z1aM5KMAAL72nX5QTwFfmoF80f4czliLxJwCpDaffDI6o6KMCcQuiAiIdkbCY0wnwAQ17ahp
XVOMryQYQqS8WWxK284CmbbFGna9WhczYNUI5RTjo3Nels9T+/+iLimMgOLYCZhEws3NR/EMgClS
ZCGcaDl88uJPrg2WUyG4imo2VRwEj9pAArkVvDClA6Ct0PnZ6Twza2XpKTl9wJawbCm+GRLpIrcD
A0eGqlIQf6ybzvLTM8s9pUdf+xkyH5T3xPEbFjIFa5u2W5/ETxgjTKpgpSoq9zV10CdxEvHVo/JB
tPPAUH41Uy6wiEWFhKpmC8CpdZ6rVfF1CiYGP/acvJaZGjR1ID57rVmIqxJGyaB+AaVIv26CWs6T
RIoJonrcZCrjSsQOQmw5AKk3KWKBXGMun5bab74SISMlcRSKfwoYi07RY+8YeeRY+RewpFDQhgUa
RWi9NSa0F+cRwMXoWwyNNuvqxqpAruXlawgO2rhMybg/8sVKLxd34qPwv/jIzgr37nxcf0BacVcB
8gWWAyiDYVBJpj6PEYXAqmmK5eBD2WR7Fc8w3T141w20KBlqF5g4y3aoSYXTcC77d86Tplxy24Pq
owNIh5sj1r4eaifg1cTLzE88LGOcMXTsa56slK0oPF5w7M05I19v7s0JLBzKexvQkOt1v4vQ2VCQ
wP+U1wXmfzLmnK+G6KXJF3OU1ipoowk4afIXEbweKhsulTah4I94/NXuAN/UMYRPzjM0Emasvhb6
cjElOpiUu7H4HvOrc1GlSAlbq35BnY7/aVlq1kK0fWentL//GB/Zr0U2Vh87Z+74u7U2k88Tl7gv
nG1XqDxVo6UGaIonFxDUg1Lb2UcsIGrPf6SZAZ84DhsXS5sdnpmr+EL/gbj/qBQjcyr1wFQMs7cj
MFbxQSfEgNajwmI7abAHG2StuubqG3t/81Wz9pNX0kdxnJkFstRraYadXcBNRBYy2Ua6sVnRXfVd
KEhuKSxxfLbWmpUP+6CRWPBiJavI1ytwBMREA0xaGqv6a31NYQXE85fdGC/tD+KYkshhXjL4AcyX
tfSWB2IfL7uWhNoWV+C9Q6n9NvYlpEQlaljNrEVL4ZHOxug6eorg3vpsjUVRcnzzqCwOkWa15iZ/
87Zsgzu6aHH/BagJp9JkNdFESM3dugS6K9A20C17Oy6Toa3AkizmJ0oj1RX5QREyJuSji/0H0Bh4
nD9PAoHZdAbsZZGu54yAx/8zC+U9j8widy4ptHtyXlx3dOMaKV3cqD3SP3xjX+XgLZNDtQswvEgT
QaVLco92repH2cgC07XYIvnGPqY3dIase3vicOJUA4/vAmUE6NB+2oucpK6Iz8eGcTMFHWe+OTNB
pKFoZMgHZYhy/Cgc1ll/nT85ZGDMBbV7HMQgSV1bh4+MciaszsX9MQTVwfdUTNKSEohQFeKFJqGe
s17+GL1CtHrlveHGl7FC0Xz1SdYaFuHA8HA9evFa6mdXZYLrD1yCXWyq25F/eQkEfH35B+l1V7tM
g234A0oQc5hAeMRnS2teN+SwEJyfoqOo7OdZyTtCDh6LjxrycGfSNz1R5hN+ZT6h7hO27bh8GHZZ
+aVO8jf8ToYcH+j/5IFUL52lV1ymUnBPv/HJ6cRWx1of49HOIroTPJ8I2mCXqheb6eO7ic9Idqyu
8Gk5Ym6qQsRLPF2RA7Xd6OnCVaAghLjR3RupHXm5jMk6fGfKk/xQQXwE+94MM1/YMEvtF/talaDM
+vdAYbj/AtlyWAPmRvuRYSlzd+MtaeErJFe0r8pfbp0X7AZO1xqltxldfIvcvCZzZMhG8gTUDURm
hoAzJlIH33Q1RWLfEc4fNbq8d7weP7tz0JikycuC4T3n1HjiPy70rIF6xVBF0Xp+TZAwpiWxZQ4O
+9GYfGOQILJKbKMvXb97yqVvRgFsPetjxpGCGFqHHwdqNun8lV3yjn5+0ACyrTwtE/sL2s1ivo6H
bLNl5WWflSk6r0aSyNiVZosJrVXAbQVcTrjf5ZV5fPBNfsSdOAb0ly6Yan+LLxw3xSiUIkxbWbAn
XLYOFBamq9f8XF8rMIm/hjBAv7z9A+3HIzh8qs7K/5M9n25dGqwhCcy4JHBl6P+BJlf56rQkEXiZ
kVsQC4koU7BQJJNyaC7zq+pWR3xF4siDm/UEwkaCMa7CV5zCDb7wnjNAuwy/D8JVZ4D1sIfmaf90
1YLvFtRD6plKiDdW2QpWjZTTc+7Bjp22+EmCedw2ED34nEmlOEYJT8XYx/OHGRKz9/hD3rh3g1jw
J7XMYPJLuTRYMLyt82VsyqgbTU2HZhAAOikjm6Awgino4vnANRtkdKVNyXnMzkSLvf2Dv/BhW8px
HVty0S7vwp4T4ywzgdY/0aCSXrPK5LMIkBjSJ+RRdxTHhXTvEp0PqURjJ3d6rurzqaJb4Lk8cjxf
6Z+4PzuhX6zD1C24g0IW4QoxlGe5fZgWZBcOIUmeYWXQW+wSMdrQD9LgUC7llN0kc33fUFLINpjZ
OEdfZWGnTBZsCPx6iR1x0pYpjxIzh2b7lnQRFy0w9VqWw/Dx9GP16RFQ0keAYYAkrtNVnzlU4+DX
ILvyKcAOBj+8g4zAATPZ9RspdzejACiOGutt1/OAsSzJXPBHNvaG7p2caQxY7Sbmk45VCoR6fs8P
5b34Os7wUmhB8Alk/ymw0sQcUAlz2dlp6vf1NgpvXnIJyw4IL97BTn5QJ5/7mpfAeskfASGB2ydN
grb/Q4g8wLqxiAtY8U9mCwy4ZKdOn+2vSbphwiaEGw/aJV5tkPZTg+j+KC0Uh9i4O5yP3MfSgNFW
sKcpvSsRpGB/To4I7hY8UBwtThbzh9UNoBwPERCD0DHMh2D8DaYFsvOmqZ3lLYtymvStqHejwFcc
dEUo43dBth3r9qWP4GBo7pYmYObnmhv/b+34TZMxrhUpJ1wp6yZ6c71NsukcJZOx7b6xaFTzoQVO
GRAB+PMGDtQpgTnNgBBcSJ7kqV0h1jTo+QO7Kk8TzIQUWlW+qQw5y/BmBZ7phFjohRcG6GP9ar2M
7W8taLtUSZEfnsK6v+o2HB/hZUbGpjMbecBAu8NxYJqOu30exgrLGbxEePq8ZNRohorDOE+M1ktx
bPnR/txqWnJljfw5ZTL1aXUOlSUQ4QSm05qX0dqmRlBvaDVYbc+9NMBWjQhqLAIE0T5EdhuX5eHZ
dbqUtjLPyzV9HiWtNM2OUNnrQTZyXuF+UnYiTHtp2jD0BvkLgtMEMiQEWba4yqC5p/uklNi8cZ2X
i+TreXDWz1J0gsFViZJstFDMO+m1S2E2HN+VByTvPamce6ZGMZjxpZQu57oloeJ1DarfhFRh3v3x
23egxViaZuwU7OFxms7YWObkfwGWalMpVZy92Zcy7zjBrLN1VYVe5GC/2E1XsRbDSzUxtB6XXrV7
VAx6Mx/yPNxhEC9IiWCx+SvCOj9E6N57WBElRLNBUh2NPKDL/HQ1Kq3LomgxpXbt/ZwxWK0W/ZS8
py3wTP/iK+z7IQD8Epi0v/8I+K8HDaVz/nwYNy6ePJS8JPolZZyw4zDcZBckBQtqEkmUMyTmpNVG
e054VR7CmIlI33WcfzpTIcL4hiwtU1OZeELv3Sl+9lskxvHb1fGToSsILcpYIA8svd1e7HuNFZVJ
T83IsB5h+T7ZN70BWQA+fnnH3AenoeiZ5QPZlm4PCiUJ/UT8a56W1kVzVfn4I9BT0AnCJsLx44kr
J0h7SUEwop0h1Y0Phh16y305PgJnjE50Of4iUT6ILYx4sNcWdH43AhJlv+dSa0wtO/ibl1tGUSVv
RtLuTpDcwRx9V5A6pfSjQydmdlj1zY5Bretlx6AuntSRtv9P0CRSKU41S766h2bx/vKUtdG/hGap
cBdIp1UMfZ4UOLauXwiRMzUydljt7Mk6B3Ewzb1cOh/UoB5pCuwDWTrexCqwZb9Ruws9/Yz8aH41
hy5x9Bl6KHVkhVy2GFSd1izsP5CIz2UyE0xRQj062hSbgwFBp5RRM5MfaI6189Ur6tDYkV/Chl0C
MNqPS5R2dZjE5l1IW3/CrXv1l4iqTpGlFy8RiZR90msKtoOQPJXF0z0ToHKMG75RlhpeX9bilXId
Po/+VQL8gZ5GlGqRMtZW3BFuMu5NI76fQ/8Hs0vTXSkohbIwFKrBkdxhBVn/RpP99JR6m+N70AX4
E6hZQ4LndmQpzSjgx7cQdOyhz/fO0zlYrmJPkNyye+/1qckOE7z3HHMm+M44A/TfcstB3pcJB6Ms
8qxn8t6hO7H2RTyjUxYh33NKqYjyXkq/HKmRw9KL5oJA/mBaCOnsYyhVoZOyvDHbusWe+3zIOZmT
kzY7P6oXJZ5q0MqKN2iZV5tOit+X16D94WQ+zWr1UX5qi0GBDo3Zbxb4aaIuQnZj5kg++8WFmhEA
3ro2rvly0tyAhGr4WdQBkgxWwxu1f11iyUe4bSutpyXhs6cwq7xpkxxgWM/W6PgrHEKpaeeMgmOS
kGWSCY9qe14x0avx7ZzCaN1UGc7TCaMRSXvMJSiF0UgZivhCTIySoD5iPDW4m19FBbe4Oe30Ziyf
Bm6hPbVJLTOqnqSSOWJ+Qfw9R+AkVjq+XjtkPy7RIL366QSd5jBgauDMIB/RRkDQWQH/i6fHxur/
GBl5E9m180Gpw12j9TdizNjDue8wEThb0/lbFFiygP8WvUB6fme43VPW6FWTDTlZFEHIOC3BZcwm
vNfY6XkiSEbXJzuaCvTSRRzz1i4RP2clR0hu1IY0pd92jCnhmPb7SGVf/RzivVoOHCSt6SFdIOCT
k9XLvKP79qbNaNuoai+CI1C5jAbQfZCAgZpgw/FcmWTY4TAfIjG/9gWKT218ESIleN8rLf7k8yM6
oXzb+CqoAwpJyod4vtVN7EWEQvzNY5rrYgmjzrc/YuFwCPEWjlBW3/llSMXOx6rzXWUuw5ioKH6b
mFJJB27RmuisbtKQF6pB3PV05q7qyZOufzu+u+payZftbDJgBnZfXgRO1zIhmayGKPJjX06qbMSi
lmK8oS0MZgfB28OKJUqZ+DpxxyvSYdLUbCzha/+xDGbCGH+1L0CuNDLLN/uPhCDuaQYAJB5q5Hsr
ON9w2fW6Glolcy8tHHA+9QxOSC1U8pQrYWbBxMeN1o+3Vg1LKGTqMKHaW2ur6TuJrce8d7MZh1m5
nn+XuJ8BSsQbXWi+E+JAJHKeWWf98O5PEMFly2/6PTUzsSSDleoOyLG227ndkFzpLVeVy21efqe/
mLoRCXljvDFNPMEKSigyazRM3yeysGTJZ3h/uuL8dDXGvLmxjx8oTtkRtvUymqcNN6ZJIEsGTZCV
ceIAd8p4zVmp00iFoWcoMeELbbCYeUxcDZTaoOEjo13+al/H/1gkTyLH8MGOvctvq045zXcjU6xV
9csnPFCws6Vpmcnvd+mcnI9/KaBLDSsnlj89tGvKM/1fXSUOC00boHsbRkj630em+Ly1/rCadAce
ouquVK3YKPpvHPKE4wR3PfeFih1iqGi7Vl+M3qlI5mOV/Ty3wze5p1G6frTJBlZzpOTqflq557lG
viSM3LXr4MRka+txJVP/C86AQTxLL2g1cFa3BbR/LWbHPS4HsRvOUOH1/NM0nC0cvEh3bXUFJNIL
xBfz9t3xNaDU/eLv5+VlGAoVxgdT/9ipLQL1OAusBNhN4r1WumBushBVznzSxoqFnjhoSLk9CKcu
1x+fPOfL7aNLUDLDTNKp2r0dU63oNdCqJ52ow2T0OJ4uawdMD1P05sHMTX5ScFhXGt354ahGDS81
PQy0+gIAVsUhl3eiqA8v7ZkkmisbCT/UAFM5CoWnZtoCA/yLH4IbLxqmDXsxsfw5EzJ6i5mvhevE
CBzGfrN2BQ99twJ/oyUJEktyaVtxt2CBD44PbkyYmhy3UCSEwP1q9P9uv6hHFevRyIbq1O/8hWb2
j1XvJFupSU7rHBTLlgzTo2aQ6S2UVra8RwQtTynA3XeHalImK8B3e/w33XTOLZEW3fHO4tWKvVq9
S2x6itinJlSxFJV9D8TVLDS2jeXotywvn0dbYey2U30FAstqNQTRK4IGu86hriFGKZ/EaTfp3mlg
MLEnPBrOwYyWvt6gS+KKJH315E72jlhfG3IQGJbn9ZmHTbN7YeQJN6UfaeRMtTwL0tLolpxGf0Bk
5KZVl2b0iWb742rJl88oEnjs6puIsUeyxi8xxhhtrT12nfgsUVVDoe6T89MeloAuK07ByXrWceqe
B+rTcHP8Z1nIqqQwUlj20T7F9o0lX0JmbS/QYnwm0NGB7spIA8SLoV0VuJ0Kgdkvq18lEyaAt+c4
K7feg/oWa2elnwxm+F9y6cr8lrQMQAPvU6CumT7CR6d8UUt062Sm0veKNcKOku61cXBONGmIgnRH
TWvnuDYoRo00eBwBmyZNyfvPOLd9sjQLQy3PdqZtZecCBNwKeiVFmVr7h4aZREMGlKdYPDPyC3t3
auG6yZfO0RVlDSDJJ5kYTkUi5vPXnM0wk+x/93YZB8t6ifKP1ayzRlKN+O1LwoqPkttpK241VBID
+cuTxmqnTDSNnMRrpFAxwy3dlWqljO2IbUHGSkeN9QAzGmk7E1FTjIjFT5AN/L5LoRujQD5YR2eJ
eu25Vg0JJ3yYZmMBifFJfyjjkTDvV+CAt+U17sOcZqyiBZnc/Z2KG0exN+NrUftfhF/yMvObLbuy
QwHnlW+hLbYv24NitQ8ToVn5AoTUKjyY8HQio5yp8Qi0x6zol6iv2jnZIRKmgKLX/Ojm+nowYIGH
OE5mpb7sSgU1dQ7huJ2IUEF3e7q70IvLclx1FLmDSQORuKeNGRENhgb0cFvJoD7Y4y+tFsBNxFV6
xs6Z+awuFVDTPpQ8UUp3VXmr9kpv8/CbhfbHjxSZaCDrLQttL/bge3+2al4ipzPdf3/ogyWed8MV
0er9QROHB3Rl34Al1NKPy8H7k0of2p8X+7m1ToaQqxDjk2JlDCtMTzZATe7AiBUlsfMQ//O3+5IX
69wAbG1xpTOq2fgZS+EIzvpD2LJ5taiXe2hnnwYMAuWaUPxWr/qsnRJ+TptvY7TjshML4yITwgPd
Vq2UFxi4jgBpGfhPsfu/cSd1qls63qZWyz2uKqtSOFoS1zHkT4h4ZFkXLgUfF1BTN5DP18Q8WD6D
9yj3iZp704u+ca293ZT2ShsTKRoFD6kiq+ATmcSjsTJ9EUYF+X2PAHGMkWOn1QA71AMgx3XwDE0Q
Rcu97L88eXH50Wv0YE+KOaLcW9bJOM3xblCMcJbw+0JKjjsJ5yxYMZSNj8T3oSkQ9/XelYInglHa
sRC5smcXdK1ZXDJjxbSuAhMl6E2zGCxpH5rtE7NxljyF/4CVA/QHwyoi/sARKoH5bkzj2gu9V11Q
qbuHJzDupeDEfwlsPcPccRl6QC0MtnDJmPteYwWOMaP4cjAYmNy+32/YYbGoYFtHwyHx8O/z671o
wfmM+R+diSW3mxAu4gZ6B+T6efYmYT3R+/xkvMZ0y3rJ/MaVImmM3cmjB3GLIl4M+eUo50RBhIob
Pg8Gh3DjTdjsPJlRfkYxBO/SIr9FxpC4xkmE0IM3hqcel2WRbhCtzN+Ll2KZOEybh0tzpW5maih+
wbuH6ASh+PBl+hEUIPm/5p/f3krCcZIEcdo0Wl0aVMhc2yh8v21UVwkBqrn+X1VGGZ+3qcurkEhc
sBVbpWiEEQWqLNlyYJSNNyiH3IGK8IR2Bqzu8KTkl/H8G3ABKbmL4l01VV6ujcpqsITpoXVMQ2wp
X9IeWqYj61bl3PQAdbUk3nogpFDlC4F0mcOvX8XJGfFfbh753A4WH6xUV18hCg9Y0IeRhaiyoBg5
PL82yBMTsm9WfwAHmeHWAWsxVABTAvIFcKmqVuLhiZGM4cVdW0DXdH1PGsMqAgR/TEu1zxWwR2q7
CfiY2pCL7yS3hLazRkpaVfj9iMntrfP8kUO8JU1f67qLZYUxYnc4ajui5BPx3qrMePT1rZIvh6Sd
5pnnO7BfCs5ImXzQfuAJoY1t31W5R/mpKkD+mDq4T8B0LFRfA4chBD25JjskBWKtDMI45qhac7Yv
nAU6PbULSzhB/vrYdn7TULlfUljNw8W02pN0qEP9v8NFnfNAGavroclkx2mx6GeUg2Cqjdky+tMX
2k16H9TU+Wu8hTngD+xy5FzrSM7eeyn7TRzMXMDhdJ2SvlHrASc6qppSbV8UWXG9lVhcefrGFYDM
/qjIs9+f3zI9vBmXvluxdV5UJ642EpPgTIEBLphuoue2zj13HqBWjCmvZRFTSt/hrCK/MYBH+3rT
TpT0zgdAZiR0YeAzSECPP2kx5DSKeiaKb7fqynwesZp/Y/xsc4Lz19dxmbG6+VXOH2EQd3NdRrTx
mF/TBon+vUyKirVtOncajrzdThc+mh8gp0hsSPpApSwQlNhK7h5TbbcfdH96BRyFdgWgZlytT7u+
SwwSgImgVl+FJfU02aoS+sP0SefJe9uEoNas0O6vP3w7myLqtdNyOmKQm0Z4osjyX+Jt+a6kLWcy
xtG3bxA1oU+DUo6vJMu+I0OGyfEhDOw+olqH7QC/uQD73KNjpNLUXX+YB8D6t7ki8sT98WkA3Zv8
HpwBl8x9CLtn3BAxCOaYX2gXzQRENHmWNRHVpC8vodwsHja/x1g8DDlt/6svrsZZ/5x7wZbqoA2O
tLNx/m/xfpMGw8E3CR54mvFSEdkNBT73JUcNMKZrRONhK9EwOVG7XUalLXVw2VmFQoqLs0YdM51H
ItFt1rknx64mdpKZ0r5NGdhrBiKUceLh96gf3FVTIZwZXqslFqYHjbVdhOpFJ/ZU5idGG1JFbvLS
RD79QXemF6sKtV1dF2Td1Q1DA+rPMwtH2T8Qcu0ggCS/j7zdSAka5OYszCFe40W2XlqsqYx+Pkc+
ZonbH4LkfQT/BAMIgMRjjpoqsMoDxAAxhFRqxM5DPCAzJHO/1b6UwajHk85FruwI3Sx1YdcW2Ak4
lXD+SrFkR0OruM/9aGO+B6diUbgzUy+YK9FUxYvhxSLlH4yVEXe1jKQK7gpMc7ZrKQSTl/Wp0aug
nxB1j8Lsd127+dmhyNtw2ufXr/5NFwRpe5j066SQdxebJgCu/0gQtv8DLjqHUpCNfSj3vqLzbQkb
e9TtP65HdifnVMyIORA6rK0hNfHicgN0WYcu4xgUJDkWNZr3nfrjRR/rjJ3CipmjCXA0Rey7jYXE
aPyqAD4zEPYm8W2CtpsSUUuUJuvuDEqieOvkUPW3NGCtQYQcQkLxX0mEOYPLqXEHpZW1jngc0/J/
zwd4DPERfeDD38d+LRRokODX7hzUtymV4SSBhd4iYUkgx/LLWbs7Ui3LNqATxMkZHEYxfVZMvFQN
tkoduzl8daZHCujZdSParWp3rFqXxaA0jV76sbti85qIJKRKdoBymb3hksni5piP029nUJHRlI4O
tZFZUc8jyuJJHcj4BcBlYgkjoeu9DgAEax5xn8oY0bO0bh8jJxh4iFetk6dqKois9egoc+uZhUYh
NGQsjuLzrKoiWa42avp0E0Nhod6x63qx2QZhOanajyQEPOLxzN+qJq8LZ6IgfdURXLJis9a05ExC
jKzH9guxAOBOHqMzKJtcmgNVyAxJidblCo9TRZTwaP/zKYuZh2rDfBLKshL18Tx17s5mo/XLF/Rn
bRDI0YxRlFvnAgfGvquh2XNJHsQbWwYzdCgjhMr8BfE13502agCdIimL5ooia3GxpVxSwamS531g
M20DWK7Y0clJw+LI4RZM/nlkDzYy3IsVu4VGtyj+tVOzHOpH8CluJ7PtcNUMb+bxL3IsTkvx1Pb/
WxwpsHws/AcdGayhyOvv1zUdL8hHt73tFdkq9VnqqUm8d722BfYn6XqgcmeRlrIk1jpQdcv05Vtu
e8HvaL/b7vG9BuH7wSwrDgV0G1npF+7SIn5WkjTcwsq5tgo6BlLwOL4zCgbIplJx8qqsoG06T4QV
yS7zT9vRx140KqEhOBX/LC+TAtQkIDaZZ6MMRm///SizgYXmS/XZolO6AUYf4CSMkLGsZm9zNLzC
3J4DnCBYWZtic31aWfsbukB0lGiQZ2z0V2GVerBAuOF8xkvwdJ71wsZo9AZ42H2hCt2sIfLbl5mj
KI4q1E7f6+gndqOqbGyfJYf7xVFAy1IWc4UhEbesrftZipE0b69YVdx3U39kxM8WmEYk8zyGs8Mp
ZR6Cxc/+ZufernIe2kkLJus7ClzQKN5lVjo/n+LA5wByk0/l9bRgQhuL5tLeCkWJ0c4MqvqghGPu
0MKXo3EpYAcFUAv0+fnVi//WdctC5qyMdkod/ZsjJ/CQPP1oOdW0GCM7NBsM2MpxY+Va+CMHOYtK
ZXLr3nyiT8RbIv0pIpPe4VlOvOqlSYXMuKan+eBVyLY9N4UmwY+UWu+C0/uN0ggn4Lf3haraOeR6
UlfrPv5pXOM2ainQ9Gc0DEGf6UX0lYitYe6KL5epJpWwc/AcAmDfD9XIkXI5yLdMRFVmbphNZlRZ
Hgg1eznFAV9JgarnBnyAVl6lFRvbFejjDF37PWzsFAD8kCH68ia7FKRe86b5Q49lGgd4jQporOwl
XtpL1fYS62HCQjDGCVyi1pS+xMJ1chXQSJmqij36FZ0AqWyDyLokmByJA9etBwSzBNp/LbGXYzV5
czDFXYwXgareyKfUpAU49BJXu4klvraw+sYPR+Eqgg1SGAlEl5WeCGzQIVFWDA+HMep0g4qImlM8
O/aPJEuntk2nYmZczMHjJ4vAompXdPiMEZlzAx48YOSPgD6/yBPzWHfhYJdlNAqOPgmI7sKa62iB
kgnaL0PYZZIyloGr/3b/Qs0n5u0UulA55cMbY+hiEskR2s3wh6Ja0GsIjSdzpJhahIps1gvyrZ9t
EEQuvLVQAwjPoQSR4CFCYM/0NZLOd8U8PZcY55WtlcPmPh6F9JCQFZAHfcWfgcJA1i/8RkwpYDEn
CQUBvsfcRKmq2M/ulZkCOdmLGys9h/TXQmCepBMZWp8YFhhQ5uced16V0XpGyuSflmjPoiqLsI6a
ZOAV3Xpsh1VE273BGPEkPLOaSmIqNkF3Ch1K3MIZfpT8cZ63z5RvGsgT//9y/uO2CoGb2TcrUFl9
OqQPenZe8GfoGxrSeIBGuhSJrQMGEGkriPll+kZzK5kcfKi6Vp8c0J1wDDxK4YkebxoebsfxJpKr
8445sQ85PkMAMlqkuL3gZwLTePrh4EjHI7qdsa0MtbK2XFN0iWKoyGRMCmWagw8gOHa7QhkWUAGP
UWNF/ra9iyqSIZ2TuwGN599tbGRpl5DXQU0hHyoAKUp5Ph3buPp7GL2V9kBLZe7r3lWsLXsagiX3
aIxKSzFbyAKP5ECLi2rQbZaeAjJJSWGyAfIWyKdxDEJ0MnX8LUa6+wGKo7H5w4+Qo05JTmYEeQEk
lPJZEb6YRDLtsDwQ3I2ovT5r8SzNpDeoWuerdBe3U2/gb99YgyIyF1Ny8UXz/4+CyH+tvANC14U8
/9J54HEGc68oOhVCEJ9b94r+YxSG5rKUjQ460nsYXA1+r/9lB95Fkzq/yNYORwYh+uyx+V9iyDLW
j9gP/U2yafQn+/4HvAQ6ZPB7CrRFlUwhr89wSG5nWdHEJlPWW48GdPcPRgcqNmDtFGkKbNoDsP26
axp4jzGC232Z+Umiv+HWOAG9gSdTVKXCwsXlU2zzFfOdb2Aw1+q68k+cCagylmG56dhBBAMtgQSf
9yyBIk5xGpLmyRYXV/ALjZxGmKFWvlaNtavIUP6h43l3XQcii04TDk0Vn1FAX7+Ve+hBqfveT/lY
FZypeg8NNgAhixkzKs1wJo+gahO3Qja35xlXEAqtdMvqd3kpzUXAki2f0gnHp/WcA4z88OU/b2Ox
OB/uY3s2R5TtxfAc8JH4jHMoeCjt5D32UK68t91OHnbp5lgdq93ixfMJivk09D6F/JOQEpYM6DCK
LxGfFRbXvW8Vah+EoTR4t6RI/qwi5k3C22pmfjyEqdpVu+QiI6TJMMjsSIhga4bMr6XwEWdrt6gg
zLezejZ2yRnT2U1w6OF/6iVQTZsOgHJqQPFgugaF37JtIqzU3IEj4iu9oaTWM8m7ZFZKTLah6WQN
Nk8xFdMv6FCdnWKJ5GPc7uXBC/XV95N8xXRzeNZl1HMQJfcz8BYgDX4bCFKzVYmg9kiD3gv/A5bS
qHVV1fVNg71h9b+0Uh4CjvvwC2p76xGebZzukEmqPDwtdRhH58JhEqw19XC9IULEU9S3bwUkdxkE
Y4h5Il36boc71o9+g8x0zYvJe78+j4c2szT7DgQoApY45uVJysEx9WpsnXvMVTUX18S2q+8MrwJC
9SVW51PtAwXSk9PE2A5KxKSR71A7w3FbWG1LqluCRO92zk1+0TIrGM8GIYUBgnYzNaancsEARq1l
/bfVRSZjObp/svnGA2lL/dRM/rtr4zNaqJuFxeTAzEzDf04LQz4zsWpktAKEXT6hreD3w1E5gemI
NRZRHhWOdrMQ39HKEg+CSm+HbzaEap9GUQuvaBmp3hIMmlDmO2pMed/u/6sQDi+FHkfuGD3oQjBe
NDDjfKkPMDsawLqTTZvtbrxDezAPEb/L+JN9kbl0VxcLVW4cQGEmlyRubBysu7b+c2NVjUaFo17Q
5/cfy4vIy3P5haEeWk6MKCi5kOU0uGPQp3wVHpWr/DR4fN5k7/f1wJge535dIWx42FOahQfsCmRp
CJCrtX3F4OlQTqYXOF15ywLw9fEu6If1ZuLUymR1pFV0ZQnD6PXLzt4AaXyVYkeDdcsYwSRiv2Rc
QBxJrRa26Ld7ocbRb35DXu9SFrHJ0gNgxeyFJQYT1tdTe2gU9WhKh7CfRYSRhhrw0U6B8O6vsqlg
vribB8rYKRSONB4M1gvB9OIZgC5uxVQ8LB9oMzTN7u+wgf5ZL4UiQ9cz4u+ClIivNt23dfcp2DU4
Gu4Ddyy9Cu2rv4ZCcFhK/frHCQvp72pmOctT0T0KLwn/0iWaGjtKTKBg4Io+ipal+jkcp41cA2MN
NQDk1IFcgDgUfHvRVWrQUqwSUf47sMrNJ6PidZKdKH0AQg1Hi8wIwT2H/YY7aJ5jR6ICSB2nfZGz
bIzA3hkGEcYEHxuhOm+lopnrNG+AYNwfOuqkDkpmp99nEZ1l5xUB2bnL0kn1fquQGoZn2gTg5CH2
Qr9WO3MhNR0pBsGtsoFLiUv87NlIhVX1Supr/3vcS1OJnVbt0DCdthWfaWElldNKJIjUoPoHWcii
OWL1VVCfdJIWM6McL3XmYkPbbDPJxtOF2lYKBdh1BBsR5k7JF7f3QpsTtwzG2dAaiw7NAV+vu2EF
zgXiYTMpH4gTNHC8ZiY40bLsMaYReK3ArrZrJ5atq3i2xndjLrujyuuS8hoKYGTWPC7MtOH6Lnw7
YdRuzEO2T5VcF43abhYjFgUQKJYhq89bSjqfzp3V6TEqlnUaQ5WD/5hMscbC2oNfE9Rw8zjRsLUG
GZ28H7tcyNP5cdUb/cgP0gItYuiUQ1XDFyN4trNOQUq7IIRQCrNNF5FGkq8Nos2+OCzMmbeLatjo
4GqjLiIBXJKgJtOK1oIbaKpteimLVfuVHP463vhkYI0xWIvUvznWQXFKNKjGNlZj49Yt/6CikvI6
/SOWDoJoUE+YQ0xaNOd7acGVycn0dFonsz3kt3Z/Nfc21MHTFjfK8hqNw0CW22/ECSPLzZo0uU+U
R48DlRDWRqkr1MCmAzJNB/nYPoxK+NR2BPMd1yQOsDVDLzIZu5GJOKWv6KKiLKlcw8FvxxnXSFeA
NKIvQwyI3iCil2QdRVo71CTjQJrDADkx/BLlQcN4hEQC2NKrFhn5D4KkutWfXgbRsuE0f/J/9+4k
b//yNMjezMTX8RLcBGeZ3w861LoXPi9XADfr65g2Hxq7DQd5Abc6ssMCuZ+k9WI3c7XNYsZHBoxj
RGMav7Ir95BT8r1p5bjl1LcApi00OsDAIfdK5dcHW3ckewTbA8xEucvtsLDQM4tBWdzI1yPItCcz
x0v7q1L5J7OMLwg5jVN5bXFesj/6bvEZzempy3qchDa1DL5gbnpHVd+deGASorf74ByXL4CgoWie
gi2OPsnKGnl5Bui8+n/h38YF6PyTokFfFaXrEmevpHRZNBZVyN9hzxLJfqlnpOWhTnjGlrJcPd23
568nTkrvAs0MRzhtSyTKJHrOGFXRfpTBoalTKJcWV7K507llvIvWz6VFZkVVRi2pBeNXgFuT3uwo
+uCMpmFqL8638OQDt+7l5GvCpJvrR/9usE0X1azkjYMKxHE3V0FC1F38c1Rgt71Xjqt5IeIxesg5
PbBY226GyHBbNGBkxemFvupy6nlZUkmY7jiUx6wDuIEYDXU4zDVkHRAIQ+5xqMNlePRdvFPlIwCS
IKmWBFeNpBx6NwpHyNDaBt6hUrg0p7PP4ET6h18kX3r8HHNYNpVJkv9hJppFOZxtYxr7Zc04D5Od
9l27UZcy3vDEHMnpR7uzVxA6U8gpj2cmFaCjP/qj/MpqqtZc7Qp+52YU13cNL3hZGSQLDTaXDSU9
0vSV5q86gFY4YtMs3vOlQd5CXl0zBRvq7c49LFq6To+jA8qk+If87HEX6rSPpdqnzfoVEA8Gav4A
tl8E5WWStETtUhXj5i4lWkMPpBv5p24zFIa8mi+Ny5AuNIOzO/chIlu5MCnoW4y8n3Y2MgWBskmg
IZljSekB957L7n1BZ8q4Th0YpLBCbCHbx8QlQaJN2J10RMJ1MEq5zdVh260P/Y1BPtmiyJ6LHflz
IJT8ZvrBKJvc+D9ZbHDbw55nVuEtK8FUuUfSuDvJ8L25GkvkikR/HQn5g+rBbw+B5wyyGEoZ8l2L
13YPJw/xWWXdh4e77szV/1TU49zqnWXDqW2VMfd9ODulTp8C4hETpZc1mb68dVxRshJyAYoWRW0f
SRwRQpAm4yYw3vo1oHc5gt6Se/DzL84JfOo+1vFM0DV2mBC3uYqeEKGKkB8WLFUH/UjELXGy/bHi
Mm8SgV/jP4bmYjmVQvK7NentdKdT/dbSaGL1hHGT62SWJYdsBwaRDxtmfrJFpZzijZNBHXhxAGZE
/9PUif120fzRL8FrqCoAI4G4LPX+lDENoCwbfWFNY01wrZfavWMgDZrZmJ3V1CANyo74yLxyMpUB
D1QegrAunGHkDidIWu8XUFiyCv3OCN2ZPZoeaZZfhlhx4Ts/Cb0YAReZFasT4+lytD9g2K/BC2ql
GoqpfII6Sr5MYWAacIi7YxS5aW5IeBzBjh9rvqQuYsKxtDQcbeEYiG8Aq4USv4doUbwt5qHim3b2
ZLn4eyqc72h9KG+6Z9a/6HwSCIjF3AYiCP5ZRjQV+gYxK3i7EJ86w9lXMQ08l+9wnzUQutsz5FVo
8yXI95cGm5SD5sfVfMCP33iR0nNWuqwwtfroAdPdNdZyekFZEkcY9JL2R/oz9k4vtQM3jWrXh1dD
pRUaB3yShJB5XhnV90pO+5elwY2lfaoDPZX20aPbWSyLeB4PNWAInYrW9btC3tvrjRLN8ud6TYHR
QgUvfDz+RM5WrZOZDPsRpFH279PBEvqBDkoR0KAVN4V64shGc5gGxnK0nHoL5GMFIG+X0U0VUtMR
pC0H5gE3WcKsyVhOSACk1TcnSFr8ieK8MXwA4hCeV/fkY15puVtOwK3de7gh3CTnDHqnin6DkF1Z
87WI/nhFE6s2svEmBJ+LjcGqDw5AqH+mf4GAIVa4BnMOkurHMftCLAGAEqw8r8/z2JZmVZtsSKrE
HGSFS7+4tqTzaUERJRndZ4UwNCYtq8f3cYjCwCdOyG+HGyiATNEIAVNqWZ2dp0+gQAs7cKbNhFV9
6xs4ctKud4sk1jEWcbvypL60+nlmjcpNNAzelzAKVmkkE9Rw2qQK0aIxZNpVItVI0sHmwb6B7DFY
Qj3QTaQa2L2gY5ySh56EyQNkM9xU1vezLbuexCVAgxeQPmi1bf77UCMCbY5KfSBHD4kNYOjVXSCG
GHN+TBtCkPmu77+patcStLpjbZHnLKmTQpDUchwmqSk2Ux6zQkiTFwdnnHG3cG6iGZU0stiTVQpq
9C16CIJ9TOqNaLwoV+Vmgwa+wkFqDcszIi1l8UKfZndiKPfjBjqS7zQ/hB5+BHX3fY3H3WT6GRyU
541Ll+gHujZsS4L9/LPtFZKrSKk7lw4w+Eok1Oi7TeTD9aBVBOKtIb/K5lDMd4IJ+amRkMt3P68W
xLkWL1K7InAk/tg+c2DhBa1B5yu/HSdlvn8DYXHCsP+tLGqtGwfd3F0/C5eToTEfLPPe1iObyIil
Tibtr4BH2nkN6FbEJ2hubXaMcfWz703MUc826IwH67ocWSq4Tp/a7RkV+J49ZlW39pMZM+6ZDWou
HHQb8Tdf0+A=
`protect end_protected

