














module receive_if();






endmodule