

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
N0hMcXbI5hCFMXvbzZaWNMXky7Cb78UlPrOh26mC4IyomLPXkDt4pohvBi74RwhMjj/Bp6A1/EjU
BW4AL9d6yw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
O4cgU289ETKimPPpC1lQoWfngvpNmR5tUZAEw+00K8UK2gEeqXn1hb3g7AZENGEwMii7hns4XQy8
DXQ5xw0Yp1Lt5kPvabj5mKM1bMdX8dvR9NHP3g1Qjd7okAVBl07/JG0NTnpHDOfWPgdIKiG5gomz
/inOtmJ9dyw3SQwornQ=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DU+IJVy0UCp9Ru4O1AHH4hAsURQvG4KWjfdJuBdXBn/Aw7vf76lLrDggWEsh/tDsD2w8gcTI1KZj
gte8Qz0RBjJA/tV/Q7C3IGP9sKs04WbpHeToWiLkJhGVSOi1cfBwcXqun7kk3rw8tbtRvnn4LLnQ
VVSnOUM0P3u3t9b+354=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VU2OWBPAFdMWY9YsdLW9vHBQultKfSyqJgSm8GFxf210g4AV7503RY1sTzcwbpKduWx2mEapVrlR
2+Drhdzv1Rts/cH1vI36ZrlUVzIXAPfly2Vw/ZI3vZ8ecksIx4K68q0S13FJLdHLryPXLuFGokYw
gCOZnAxTuOQQMCgsJA0iDJVXFdmLXzqwRYBXguqf1r+OMVPXs57gcwlgVB8r2wrtRxBvH0uRcmEd
9XDbIcnUXETCLhyRgVVpblWBh8bZbcQBY/zZZ/sbyAPD6J7Rp8CEPhLVVCsK4EjNey5PsDgo/izg
h4bUKLC5eF2W7tVckgp7jyOfw3DgIr/wn7RxeQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V2G0fgDEE2OFe05Cx8OR1KsgdINzVEXBIBadpSnPXIoTc7xRwAe4/VP6V+6MXz0QrLZuQHVAj7G3
9F/ijf7v4vM07B7zCCzqKWXPOd8bPZE51/A2H7Mt+ilGqjbh/VKLmxGs4hilsENWISKVXeBdKnPY
gj2HGvaphMJpBpJwjPAKBmbUyTX5Sd9nNIMzcSRJNulwiaiEOrABFlrZOI+c7bZY5sHmVeOtg9CQ
vhwpJiZDt2xEUYZdJ+nAzC0+NS9jg6KFWoyyUeNOwHZC9//fhh1MCUzJ0nZg2R4hBpRaxLZstp3w
PM0at5MBtCkDuhRItVUmq9A0HtCUCEmB412P1w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RN/6I+vbSUSbgQKZutSOM516q9s9JryaK6V/qqxo3gcYd+gU9W/srRAx8TWXTu0WbgzNnJ4y7Myb
hqdFZXcfJ/PxMgXPrrBTM9dc9q6Om0xxWrgSNxYalV3KY2vgAYOZai6mnccqhDfT+ZicibnnsYmh
yf5l9IBMwTbxQ9cpGytJTrr0jtjFG8izeH9CEj3vxYZQ4tA0TFJhsFvQhk2xXEnWnEBhTQbSX/B3
CADhGzXitOUqpBt3ylEkYkNM5wRAzze9LtBQhOCFWc4AJq4+3/P22qqco2g+VSDFNt7Sbc/BGwyj
q/3tdC0FZkEZB5DXnSDvgc9OVq2Fggic0aDyNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
R08pqCOBZZThIBK/VQ6MGrQnes2zFXD3Ek7OjE0CzTsoBXe+vwmYnBae1epWEURpF4klJsbJH/83
kORCigHNb8Pr6xb99Z/85jXFF9MEZ0bQgt1y/hMD0wcwIuvHHowkoOXOKd6ZGJzidg9L4/rKsijn
veMLws0dQqzRgrTg3IJ8ZhqGRR+vIIyYNKEP9+p/fD5KX5E78RJapkrxUToDamMEBO+ZpPY0wK+H
Y1M7hk/+ek1X1cGkLNFlYFLIDFb3gTOuT/li5ReiXpxOdkKcFp1Z5C5oaJ1R7azUG8MN7VSt0yiz
CvQRtH28BpJ67aocCoJyWGfMxzB5KOUSs0+BaipCzaxyWFs+kTDQvyag74U4pzC+59EKWar5raVN
kU6/aben5yFlUbZNa21witsbJjyJERyok0ygjQ5xir6UmpOCRzQzCEgudalqMSlZhzDQDFjMJI3u
qhZCOORLDb7A2kcFRaEfZktDnrDXH7gPgSO3aoZ/B40ekmlnGAlvxG3Cz3Jr+VGUtxNW45jGmA+1
vluVgXhCAu+UT1MQYH6dud9WwrfvMXCDMBQZXF9ma1R6vjiBd2EG59PuF6WwJikbhtLQyikLbtSV
q1UShNBnghG351sQAOQTG5ruTerKbnkaXP3of0KeL35WBTyfcrfHD92+nsckqrHSxxSU39aAlHgP
pMaD1P/eNOURUpny2ZFSL7SR56VSx4SiswzxOXbNuAoGp4EkwTntYRH4+oA4Ld8mriy/v/WmGqxr
ttr39UpDRgh46kqE04ynHLCgu76TARZfEStWE/DI88CCQVyVLhoyDOveykkPAd0RKZjj+ZOP9Yc8
s0vcBtiXel4Xt0l5emXvPqOsR+8d9e4u4PepvD8uewco6hYN60se/SmW3ACgIJg7WCawgh4SN4ya
MwEHuWrWXNamURxGl1/A+ekdM9B/KcEVmXayrOj6hyTUyzSFMit2diuJ0zLob6LcKV+WvJNjLnOA
64NgdiWlVwc2/O4KCzpq/tcJvf0mOhQUNDriObsG666spGZHtxW54EaUeSn/mQu0ZpUKoLwWG57a
NOdc2mg1WPGIDgkI8aUJutvtoTVWXoWKEYLI5pHSIsASOtog9H73UT5J7m1Ih2wpDQ+GnassSLU+
kkyM4/9Qt7zOazEoYqQ82lmCgG5gEST/+F6QQqk107fn8gho75lvAFp5f+A/PjmSdP/AxOJnGq9V
6hVNO9ggO9MqT3f1uuIWfg27eyFIJu5FpqRxk8FjDoP2RvtxsH45+wdX/mTaYEyjmBHPqyu31hzM
9t/Wn3Jm+ttD4zPsLyKaVQsD78ggoRKGLf8ZxfKTga4i/agEG6nWtItZKyeqbiWgVPOUL3ShMPsR
gCMGyJ5SBWRW/p43WhOud1HHpGWsEAF/S7mpT3cgBp7kuMpS1WBfQGq/5HL2XKDFYSKzy8atw+Dn
lGrjiIhORNZOOFhb2aDL3YHa9FVss3EOBNYHDpQgnLZQppjXPzYtW4M3wt+h2yDnn71R1ZyKlPYp
3j0b+Hhquj+iZfG/HhkYwYUvO1TrcKO4C0QzU6NIuRNLnRk1k7nGhW2q3skZNVteE5QIIvrc8iFV
VYFPcY6FlPjR7p7i5yhbDScV20Zy3+wPdCyih3/TXsOEZXA0I9LthjQV673YOzRzgAykFiCcJQ4D
UJO2O0VJJr1veGhHvReto4ecSmk6YiMHiOqFo6DiwTI3OGGXccHCUU9BnhAWfEl6tr4mx1/nr6SD
9ztD521P1DywPsxI0wKtSX4rvA+ZQzoF39xiP0fnTN53RRCg7d/ul43DKgv0dOL0cUZ2DD4Gqd0X
9LVBrUNQWJ784UpZRymlC8PJRQ9C4EnjFwEwRp7GzEjvdpc3RFzo0JF4cxRyzlG/dxm48eNTogmN
vybJAbEXeuK1nWkLr+P3J7eUeaQ2Kn0Ek9q4xjWPBJkuSu+uGLasJ252luvf9FIm0pKGQVajs4y8
Fbft56mFBhdFrTw/NNaRcWqbrYKVujQ8cqVZKwcnw24NDOPZWG9WE6cAa5BYQli5uwE/MySgz7I9
HkdAFTR+EaLmeZm6bA0nMlnJ1Fy2nJb0hQASLmrlKV0tG4szeZdYlUNsFOHJGmwz+XWMNEd73B60
9irK8bMkKpoXWEVi5wcG+G8GvhAZHs8dhcJGuTesDd0mJNTgaHPT9A07Jv9D55WyGz+oA/bdg+rt
bnigSLzcJAwwTN3R4v5wzau5NR5IYdhGDHVXDv1BpB928Wla5xX5K9V/SoplPvfRmi+rdqAlYKQV
uTkkck0T/Nw4q5iJtCriKtObYwkVRuCkZnrGy/5I8whsUopB1Vz4LKmRbRedd91mUVnqS7WPCqxU
r2HWZcEUpCNnG5Sy/52RbpZeg0YO/Ht1CZPB7n5GKfWsQyQzRSyYyJwxGAvmnr1IqCT4lYRP4MLk
cJZYNk2j47UZUlHJHGa+kzTIP4nBohJsBOvxqjDCz/ibzWRMTvHa2EkTXh8RgI18f9GP9KIcb2mu
bd1tQ1AfvBRt6NjiWJVkKDybK81Ro/k0ra0oTMrYPCuP/GQ5QCV/lFIb6qIjmJ6Rx/TOzHNLTuZf
ieUgEu9RFLhJWcyGL/X2kErBzjRLVIKTTKRDZSJQR8GJnrgBp4hq0RiEYKdGjo9NzQm+lgk2E01V
RG0bneKz+Cqo0RSFAR9jOlYF+DNYQTuBpfqReNGx9R2m+cI7Vt84NGdib7ACRAIZihPIDZ1K47sH
yfFUNjv20L2JkZh6berjZuIY/sk8UY/d1lO22lmJKhbNW4fg5WBcKUHnO34QLn9Hlugp0Fx09YPy
T9RczPCiTChHX1Z49WBa9vofKj3FOS2T53XMtvXKe8t3el9Jul1AZR5XFXEJCw3MySJivKqgiobz
e536Z6wts/pNd5HT8FfU6rZNXuRCS8zNeo1XqUIHnJ/Bq1t0DqW2aGlFCRMCFP0RJp4RtjXUaiWn
bVlIUKV5YzxEN/GCYqtGOdZ/juAHpyVXosS3V9sE6C3XRa7RYdJloGAz0RMjYFDi8dJLH/NMDU4S
kSshB2VOfnvnpq9EoJyU5CIUILFSD6IiF7iDZQYhFeTi/YSc93WcxptvZkAmI3JAHvKYfyZMthBG
5GY2DrnxUN+QXVNb3wqHCMn90OfyprXUrr8AKJnUy7TrevPPjVUQ2RFJMEH+IQ//+2tyP67syxil
Hvy1Oe29Na2QL6ipJWPTMEKkUiIt+Sfxk6WqrRyq5mdWIPk7C77yB8YnrQg7h8tSdmZ+m0kiwBvZ
fgtOgg51Z+SsLos6dd9ggasmB1chnER14upM9k+2fXBj4sPNqCJSTifsQpbtB08IUjLgdv+Uy+C5
ccQLrgB5vv0eOqwRNd9CsBhSyqhaSh+UqzV8OE0FfSHM2+zhnEoI84lbGmzzJdSfbEkLzm4M8yTw
ZvHobYiB23LdP+Hx8MQ9TKgW+KdB4hArgb9gzI8iBN9f4HJjklCw2h27a+Pcw1AbkZ/lGiQZ1wgo
nDs3Ld8fOn8uOBV788Zt8KwTO9W0uQpA/P0r2BHdJbodsP68z1zFJHILQdbhOgvwGZ8mwybPDPe3
TR/n1V08chIy6kaf2R9BVZs1F2c7vTS2fV9lIpftSoUfmTJCdsWWXOz946MynJiJ2KZXikEUagU1
ldamZ44a2hRaf+oQFswvmPjS/b/hSvZ2gy+vyxfTqB92Hv4yTpTDsQr8ZcXnxrk/3rR8H8yDVFyH
m87DbBPFm6RBawzobl0EJ0mjyTbb/RoKZlA5dsuFMHYUe68CZiW+61gnlvwTccVe2QvjfUcF7Dxw
HqyKoUkDYCTCx7AqCxk+D2hASk8vT2Q2zfYQUDS1ZGVEnzeWvZfMo8T8aiRSd8fF5NSje+Gf3cB3
fB1DwkBJJI2JS2JeJx4fB/N36bHHH8PJc77TPf7WrSoBAP51wLKzJ743rDlHYj+brX8JmTdXvv2s
a4InUjpcWSAWmFVF4eKtK3O5N2Af+beNJs0ZT/MzTk2IbdJxsDFKz3gSgz9EPITbEsP10+8at2qY
bwnC0Zw8fhA/UYu1QUfFLwE7S5eSwyYxX+BeUMG95C3wVvY+dk/3BEcXDUh1YSCHVO0oV3o3W3rF
JU2MxtzWfmhIp2ITHBSqrSVUYHg4aGlvTc4HWx/6SbxWo5+/uYeF2UMgZOP1cxOcL4WbV/nzUojD
iNcjGs0VHC8UUA5gJ3pHB4i1+l0pXurOr2KmrfxcBVZ7rl9h1y/spSh33FeAM/tGaPannXHCd5oJ
5or4cqz/3FAUxYH3sMD9SnLz5CNiauo1wXq+XHT/BKpqTLfyYSCreohLWM+WbcEfvSjYck5nGiBp
yX7KEx24Yv6Gahwi/yFMfU5kTpmLNB6Qz4NuUiU5F7YqRfeegzf/LRdvoqyFYBg4ZaA0KVi9J/sC
LHx352CWT7G3i9R+kPDm+/gAL0mIXhIPZLB9h5hSXREAdZneIYLYTVuKy4amqmZ350osJhsDiiGK
0XHEiElEXrpFNvZ8KmeJtUZj8fwZSTNnGLXInHClveATm391xeF6m39A5zRy8Tv7HBbDoD5KFocm
vhhnejvBOqJxhWqn0ckZrUlUisl01XzIZpQOwowzWyutKSs494Vz5JRFARhwSUDSSWoPyeb6fxYb
hx7dY8beBtuEqVQ3hKMT8aapcd8Lx1/9YWgOOYvO+kFGzYZG4XPAu3Mo7FmoXqMCpC9HBoXc1Gbf
iDNkWXXzXUvCI7PkV7B7JkeWc3qqIjpUgoFLWm7SrGlrU0LFzu1sH02A6NogNCk4nmpIAnh/Kjja
Y9T1eGbtaVpfrUXigT+TfQdFl7nW7AqYt2f+FCM+N+5nHNqDP7F0Ak/hrH7ecAuwxMMfkCT0u2JZ
/8PKRurtJys/KaFmkelYgs7nwGemsxHzsmYZ45/l6TdlSVUNhAOZR+D126eGm3Ys7xxU13R7IaCO
La4ZQFvX+lV8b6RGnQBcWZhLiCJSSoFpL7S7IzebKPuooXrE3rC+aedm+gH9TE9wFIXuGDYvGCjv
iaT1by2btbzDvDvJ/wBxl572764m1jRA7MkjN8a135XShYwT/GQNalayPrj3FI6IJnRdZTtdOBZS
ODGbXkl8TVzanWtH2l844X2P5S0rsA1EMqUouL0JHmt5ytxYVTgGk4Ep3OOujVWGK13HGEEq7arC
pjTHZ9VEF6brmqs0xPH4QiaevE3sFONKBtfzXjB6v3pTvE59LLKvTJ29iXiM/afjjcGT3x5QCi6N
ejot68JLmEEFAziAEXGBDey9GxicPhVB+47WiB+x3x9fqsVGaGSgujU3Exzy3EBoWl9GZpFcj7i3
h/7IuomcazHJ1dhp5DAUC71gAL7t7e28QZy4CJcgY5L9biSTGgwLUQp8HvF8jeW5Bx+MMm+IjF8P
s+PxU/I09kZguXRciG6OVs3FWGMM+e8ZKBOmdq/alCGRIdZPC48A1AiYnmCYC7vPDb/f2FXoZWVR
PQkFTQ5to7dfuZz3QrPp0IuT/dleJ+y6X4pzYkLENLOGrY/3AdwsnJjv+azf2K/KQyWn/Z11ceNX
v6AJAild7hY0I1IUm7KySCff2RVD1dyrK4n4xegQJVlWIeqrLwLIfx31cnorCBNVYCz59MIJNq1E
YKAhS6AtiFJxgioWMzrKzaylB5a4Y0uPb/lypc3qglefofNnLbxuIt+qShJftdq8iZBDXJyJoBgv
u+RGgjN0QzE7iAcLUpr+c5Cmdh6++2lcEx5BuE3kIV71Tyi0Bw3DBo6OcocJM2m52+wVUIILmGCF
0WHprikTBj03OFQ89oVpj7UvbzSPsXJ8kPQsElc4+FFAOXXfQavxSgPemlSW46HUdvd0Dpde5+hX
kGDdlikn9YjaRqhoiBMp2ocNtpBK6ngxbT29Np2+NnYe3/JRcVgWMHuN//+E1SlRMRYfhUevR8Uf
UfGyDJ8v3aEKiXqo86NaUHfvN2L5Hw8OHQxB68YPaZ1Cb5Ilz/83gJhv1QCRvdU+DayuPUGaeobW
VZdqf2K+E5fY9ia8wUGGOlTtGKoumxxqTdpGxJmx/TfHqaQAxyHVMe2iYyQ5PMXQZXfzC290yrhQ
s2jIBqfkE9I3yqkVPLpHqr5oKF32wQpv/HhzyJ+moNoeKRVTUmduxfddq0YdBa2gZf7lTOL+996N
Nl1xZGUVkoXhkHmpaKzNTonqzS0wfgPeBPeQGQMi0IAUGMxhdDMLEc2LPrgFykk3bkDZrr3oa6TA
TvH+2yvn6pW6vvnkdiLTmjf8CYc7tt/pR0Ah3dVF4fb966r79FkYWHNdy6mOvRQ3k+nbNyEpu4g5
ynp0x83/fnC7uCtkK5MWpPjxgZ0A37+uR5cDcLOOIo8FZiguaZgYW7u61a78voZ6HCYzTsZCkLFJ
BhEME6pHPRBkKF2Wn8Kj9ML6VBgoTcyExGEbrPKxOnvISeVZwdySjMmG1X7ZEDlK4aVScQNDD4sj
UWpUHs4fO+CvVnzYDOSWX9ZV44uAHFnCZx/Kmy1PHNhdqNlgYGB78i2IOh2HhGe+PgkvOnAmhbp4
6aYU+CwIGaXTwBAs7dN8wOumH1Al+tUsRGuwD0EX8f7Igx+bhEwJtbsfrwGTEZs5VdqhTjxIIJ2j
hmNkehUAE9lDs2oYe7OoFbzB0Jk+1qWxZKOzEQRA6rVI5t34hCZJZ8xdf0tW/m0Epm2HJJO6YT/V
8sU86+rj5oiO13CEvcp69rkf58Omk9wyZuSSDpLyGbuMrElimb6A6Ri9EhuYuGTCEBSo7t7c0fY7
9RJtgMGEk2QOG51zYzq0MBWgAgKOuSIJNu/PIi1mnQfyyg/eoZOGu+p2JJCIcQgkt/mW73BvWjXy
lqahunoYNtPl3kyWB9gXe+/gnu1M9yH6jj/R2by0NEe590Nigw2tdPC0pCezRNsBFgo9pBnVpnif
hvqK5pV8I9943eWXfaFUIMxueNOhVXlDGt+9rHu1HYq3JCfQYkxExTOAFLYGAHDDgyaOqdRqcGH/
qXhw4BJP6VNh5t2DZwD1sFZg9mWK2Ph8untpQGU+AZgI3nqyPgGBmsNRSwCseSc0Rd5Vdh5q8mXK
Aj5n9J6iByownTlLrD8juALFvdaaeSS5DVORQ6fu/ItNqrmLd0di3h0nFgTMW0GRph2d2FBukd3F
qlGlBCin6HN2GLC7yTPNPSCHBT7thCdvszHN22y6v3kyLwM2gBzIxheKVgROxZZOLJLg0maM3KfQ
R2khrmznjzdnVdNomowgKIkRf9wJw7X4FZ+lC+jJelaI+LAr9AHBmA4/kpjfL+EJF/uwvF2dVE1s
hJwX6Sx81YUJ2Hf1xyjm9AoLZjq+DfqSoZ+UHUJbxUNCMxyP3A/0Kya2N8FP8jFV60uOxLwIyVAz
zuDt21gBUCDESHJRJCcRnYhEldnY0xpUqUoc3zQ3ODB07eRH68Ryt3OMKzhOT7IGIdX5wbNV3ZBv
Sy96Dd4L1i/dL7TdhGBFNo2yke8/c+h2RWMZAP54ghj2GHeaD31cjYUHsr08M6tYYC8RMSmWh7aF
o5dOgfFPkcmSzMF+QEsW860neEUlVsUlQuk2+ROzLGFmFJh0QHwpWJIoesFNJSSg2VtEmOqvC7xH
/fx7uAPvfCoFQA7Z7McyC+1oJMjTvzm/BizN9meaH+kFhuJndfOv4Kyk3QgOTFmdoU+L0vPw/9Y9
alheURKFjyUJUDRRI4kYViEw04AX2m79OufkbVugP1WRXlR2w6vS9hcvKB3munJWpM0zze8Iv3GE
m7g9716AIj6oLIV5mmzXD7aAx4M1AEjv6rhsqONWMrQ6DRv4k9fsIhabRjQDSzQw+oPBCLojuC3s
oAgi2G47N4KYss9KMQWNYKPfLl6YmTMsxxtUt7k7CtOiDN0j0FQbBofn9Xe+cdeHDWDzMzbDOvDw
7WztBu2nr66BFHKFL0RwVEL/VtBcp8NGQuFKKdDBtF5hdeyGOKdAl7fKCjFeeVHxeRdEf53GOFHS
VdGBpoCB1QmJ+u09ndYN5uILJD1mX2eNM6ixe7U+XO+/sF7i+b90Pw+dz4yL7WA07QzWc1Tk8rco
fxxTch03oP0IeR0CjZiBzRu2gLv2ZWRrkNgV+4LXqSK5XEMniGEwa25laD21KLGHWJ5o2aZaJXtZ
rCytwvV+OxiyldbjJhKJCErADV9g/yHdn4DMhqm5plnGz3L/zYJJr0ujl8UbxCm4WF/vsif1CVqI
lVzDvLhJAFH/RpH7KVy3KAchOQ7rVpJJ6WqnzanseqQuAoBQde8jH0NjD8mZg4tAVKwqz0IT80yl
rfCMq+tSRR0ALSnt+cV8bXhb51qVUBIC/cv5qFb2JIf5Ii6bzbmn2XhYy1o1mHaYbxwMQKXOZVtQ
pCAhSVdSReng591iI52XRoMFrMMMvkU/9M3HpTxHmAF/aq8yn8LvL00QvgZIQN2Wb4ujVsCGs5c+
+U7u61doZJDiicMUewLM+AFKLwTePw65NsLHxhYKkJekgQ/xRGCrsvO/lWj9FBK0ncMXMrLVK2HJ
2X8repV+fP5PKNAvi6f/NVCqJ8OspJRusKayoeSAsMG1BOP4e9k8+MjPUaDaJZ8MsUgEY9D016mK
Pw0Nys6sDLXPTAc3utjAnFkmY1PIrcHvmhsniwwpBOxAi23qi2prmSPSdHkqR6nBsunxNHXDHBGc
DOQSj1W8nIAP50NdcYXnhCdXsRi2BKW19i8xUEsbEJOmR2+oej/K8ZaqG1uGZY4qzQGLXHvpbLPD
ctvr6/jRp4xsVSKc8Fbf4T0fez2odmGSFhBdayrlphtaEkP42A9Z5/1oo2IygoQkZ+ddHHC7X2ig
be6oZtxbYtXYcyWwZjeLprOXXl6aJ7mu7sEcflBhTVqm/JNPvN8rr6IrzxVrR9RuxsBSTJfZhRJp
nowK2hHzU50+1dG0hLBDHMg4hdSfcMnqw4gCVScLYiWwy1ytyplPRqktb9Om6sSmomV1vvH36Cik
2+J5AcfI/2l71jRPFtY2XTRa5n5ygqsakPswL/yd5jyGBdQFkdmDvYT7GLtvyAw5s4W0JJ5Jp8+y
qrSXILclOSv1TFyJamETaFA1wisd6IJf5g5JSZmsEUXuwU+3oElT/bliXjjaatlniIi5oV/hIPCP
ObfttIABfWCT4epKO4thAFl99677UaCBpmOlvGOFffFdmFcCUcN2vM46ExmWYPLNzMiGMth6YUyI
t0FCYsQSQiGvE3UBOFesq8WMLrUXaQKuOf3LQTJjXglKaJM8WRlHwQuQl9a/c12bN8PppwvIA9jN
LQ3HrjSILH56CD98S3cUchjgMPA77If5UZkgkW/32pnihZ5kF/FwoyZIi8MjHo0MLGRfp1525AEw
e1rne0sZfd2ashg7IjZ0GJRTjwFlq3v881NhxqleDYwP8G2NhztZtBGyCQIVijTe6bcm/E49KWMx
P9mwKs5CRIhTEWFc+H4Kvied08/mRlXGibgr0G0t4gMdX7woBZJMFL7CQdpATG2LTSlTVGg0iZw7
KMKcFuR7JLdpwZ3LOqI+P2j3Wo/1rvviaHMkQmRfyvuHgLJtUNrW/t5X8OwZ7Az19dULVEieInvJ
ZF07B793pk+wUUPLYso+yAkUHfjvCIhTDDuAFMxiwmXVt8IXOFlNoUXwOZRt64ZPpHfP9jVKIQzP
qtyT7ApoICV8MScHOnoPAZPwXH5xigtVN+RpELB4RWCfofbhtoz92r5M9L4cw7E9ub1nMxMaQ6Bg
qE2/rR5fHDdCjeB2Fw3Hie/Gbkk+Vxu71CwSOxrt7iSA4PyShs1Q6sP4Fzl7h07jUWTY6Xgb0EcS
tppCTJTIqRCGcYmJihPt2IcYo7OUnFZhp2S2GDIRwafhI5W6pSpczLCwz8zx0Dk+nqx3RUowgNrD
Ctgq8GLt3agNJcyOBobFoSWYSFGrAOX1H6piiTCi9c5F/nD/qGkqLQ5C0Wgjc7jqcng78fT+nwH9
7NtbzHVQ11N4PhJyhoWtbc/8/2proqflwnwzqFan/KvxD+DPwk1uzXH/YwfqdvISp17gD+ObIlf/
SZVTvZLM+xQ7R0CIF7zDwa63Tx7pV0WVZXB4QEA3l33OfYF5ElAwdeu2cigNDJiErrP/dwVkgcsg
83xdAS4V2Uw1WoLapb7iW68wBGMHH39y1SsGfzJtxyjtcRyhwCmM7lKQ/s79wQZsjeDPkdjueSNw
bDr7BWAPgkTp9UutdoyLX3s5JvVI9yxhL2zLkZ4BsWtocempRzCcPf13/qS/W3r3OHYLM7woSUL+
wp9LvVuNrxDFAEJMk053h8cvXkiUref2cGvE+G705oUB1UWphD92x/FpM+vZrh0xaca/l7SPhveS
Xog0/1yFPkLuR4xchLUWRoyGur1PPtGW5J/MT6cZYHCkbv7nt5EBfbb72ZwF4pF2LgesRalUY8yd
cUlrVyR1IWcjI8opOFIsFPoudzEwlua3gn7+mbuPuhcLb5MYluY24ev8jUKveBX1iQWurxE6roqj
tdZOYzNiBekwoyqzx50QGVcI/k2VF4iqSlViaNGnTnMbZo/PyGCX/TyXtcWW1+5hU7CQ+oREbsZQ
OB/AQeKC5UXWXsQGZq611Dwzh1HjpMcqQLeJz7mg2jA2sz4HJbQjK1fqfC8IdAiR3NlEqqJAUEb3
dZtDNLPuHuQ8xmHceMuuSjLuFb5reGPQ8N6ix1iQyGlv7MvqmdPHaSF2MnS13o4fgn5Y2WhRvQNb
qIjhQZsArnFxXlztyj59mn/ZVTFwmehB6/Vd9tb8r2kYmCcFiDXAsncomzJcx0ge6FVdSmc7FyDv
JQ+K+l7rBaR4eVgn6MbYWQrAm17Z3vy7Q1Al2o7VBNwHxPyO98VyK6FplZHs9yPR+KNeA6ikE6ay
DRWEPvrvpT2qYa8Hlac7gN3Ld8I0uk9Je7Y3pSj7OuWkylD65lBVMFHzUU6S1TCKVpGdcoAubF0m
NXLfLtH/siVCU8gqJt4G/9DeLSouAxzLVivNd9HI1HJqQ2f71H3mxKwvBzYOwhWIRHzoS+HgqTcj
bc84LvOFJjqjmLMtbViL6EcXBYpA1Cz4Sh9M2cumsxVg4FAUPkD15frHMbsMvc1VRUo45C7avNoP
ep9efav3JwEqWvM9lv1igIHcbMJrDJh8eL2JqzGgGCFQcEiMbAkPyHrdts2N7KzfPs8LSBdiMwYZ
CEF8nLTNdajJZCFnu3rnNaZo8yOFuTZyjfTdKakEwpq2NO72KbLg1db+HtwIZ/U2bFTUpV8j7q2C
KXRBQ8jDmsxN/vN3HetEB/beEpERzOl1iSMcInd/B3GRyenDG4rXXqwrdZK3GarYNUIjhvR0aZ0O
/beYg5J5Qsuy32C1kfljOxdKCIo3kU3qXbdqzMB4DcV0x6hlDA2GeuSOuCP0nPBHbPU/EzIFrA7e
eW3olF+4mV+e+othUEyC7fsVqJgPm1GZLpAQKHYGh0JmGcJi3YBmOnZ1dTuxN87LrCsDMW0wsNCn
aF9m7r6dqBvRPKMzLO5pcF/wk6vHzWvapzCKJrmylRM1y59uCzuTGk8i3w0oOhI7ayEPbg7fY4zt
ZnukVH9qfD/dOho9kbMPRPWTzSceFgc5yZEZq6t0kWDvx6Wfx41i83GBuVOrkleFJbx2dUeU8DCD
E4fdj5+roe4Wv7WFZO1L6EANixQc0dQDWA+P2LZk2zT1WyJRl/DVVV9a13aiM8r0gxfW25h/vQ+K
t/HudCQy3gHSuuhXz1VYefpvJWQ2mzg3Uvo/3HzKZojtMd7PApfXKVvtgp3ggYHojsHE6wq11tKB
U72xn0X5TEAZJHvPfah1MXLJb2OKK6SPm5O+PtQoWbzfKI6v252Jz4ZM0xviyH3Iv8DO3EPnV2g6
M9kbXI3uKZhuKHMzuhBKRXiGLmMVdB82GE16LnGHa/dpNdHgCzsIRoFBAy6ve6Nw4uh/8GfvLDlW
KDyNBCXhfTcaVhm3JT/gxt7lNx0qozzBVxngVhHlD+oyIEpN5T5snr2G8YNuoilZWudUMgkshSD5
rtPFlQykxgkmHT2mEAZ8gMIDeUH2KfrLXH5cgRYB3q1WtpK1Mn79r/Tq69a0P8YkUODtpCPaN9Jf
YvAUijU8zIV56NUz36xQNpfq0T8q23fl+nG7nfPPiFiP/IeS8/a6p3rhMNhvk65GQABBopfFaJTe
EBgc7kzNuTRheYb586Q4pelEDt2IxtRooydq2rmAURKmNtMYqCyPFmLov5cCdTapyWtrs0Je78+i
VJCg0DnfQGLXfkTjlv7KfVpyw2h7VortCfHq7FJE6lonb8SWYHU9PLlS0n3LcunoPa4bA/W/MxJ/
PnJRLiPPy9h8Lm3LmkUO0tbgSax3IhftO9t8Kn4DmZrbrD6yk/FSqoqzDQsWtUwwoNHK3xtOyqHF
zMqNDP3iBO+m0e8ynxu+iXOGX4i4yOAfcGbHzKTxieHeCf/3eVsyVI+xb2Hq5pSpZ2f42z551d7w
AaH5lqbfjS0LaZVmsLLcQjhlh0Boc6+AF9RSpkm6d6DWDZpdyz6hv7ONVjk1COsVHfaHhbhbxsCa
Av/nYM+mNrwhw3Re+hsZ+M9ZCeTxadgEJvNki13S+RGKfp1NvScg6oI4jSgVnS6eSB8vMUC73rB6
eeYPbPJxvllHfGDupV+5r6q9+fSI/W7YyIrPjBDuJfCRB0iLHb0aNSsRXUD+kFWxR+kdug6g9Ccr
289RbMWk06QdA6NC6NMZf/lOnnFPWzG0jaDk9ryVU7F12d/c2P1RgTKWFBrWfrEWQJMInD2MNxj4
SqnlZscgJNP0vb1kX/7sW5TZOJcLx4cTXZpE4dbyjyjk7D+fYCG98f6T+gWRgcAJjNNYIPu8pD/f
Uoc3EzpzBqlUscwkyM9qAF8lOXdlEpa+YdfJSljIYrga4rLzBD4ghdCLcNxjfFy3yeaSw6HPau3n
DqEc3cULEAkjDEEamWR+8O9f5reQjM0HPs9w5GjknrGO/4yb4lJFNxb43FrgMygNM7T8qRmXehEO
eKIlWZWJtSmUizpm+l9cWQ2tW2EnLGoxNkR83fP5nyjctzXGPKuAst3S5fsBJ2UXmbgE4gH5121P
zw4xMtIwi1CTu7WMy0xzH1ZuZ+jqZ/jw4F2b0BkQeHGtWIknpGnSxwyJXPFmFP5zIVpA4pp5cWdP
nZs5m5msf6pj2WHMwLmbtz4i5bHWUekqbl6I71EO5ays4pHSlpygShXxAJwPmyL5h7vSryjDz9pp
QBJU/v3jpfXIYnocdqfG4o0lqPTXU/3AwB+AQCWanBDNYI0q3yMU/5wL1yJaDdYH44j8YsMQ0hPD
9Ohwh00qirFUUg0lohWCW/5AXWheAxKv3sXPoGMT6dYsaRCKit5mQeeHj5zp+iCf+nElev1SqCx0
qtONPEYZ+64jSaJlgnhNvhodWEYoQ6dc9QZ47dn3U47KNj+oYC75LWAruRL7ShZOYI7tFk1IsUt2
X3ebR09IEZPczuBsvEPZtH0mNX3NM82fkbRPTG5w3ARYKct9EemWPbccnhn7YiHJxobVXFxsBHN9
UDz2jgMXgYeqbzeQAFmHEc9bVQA960ZCGiF0C0ObMLZvxPt9x3V1b4pjle5N2k/QabUBj2DPnizn
EyQ6jNHtPMV6vktDl535lK/dYCR55lOzGoUvE3Vqr4jhQVwPP1bCZ1vJavvwWYH4nf9DVm1QB7Sr
U9PmzMWNMgi1HTq32LZTOwUXhXJycMCocDSrpMdsn3DBDmBcpcwZdbALCq3jAmXW35uBJPZK5v2L
2UgDVL8YEEeL1yrZda1yDfI+FQP4iZtRAv6lwj6V/TLPrw4eM+S5dwXgtuYs+KUtY65Zjb/SFBOd
RD0YOYlrAiy9sR/AHDEf4dsROySRZLiyxrKSPWEDLn/m2EmqvKt0fjLA2eoCV34rhJ0zzSdDUtd+
xOSHmRDaXnT8cYzgWxjKqTcJt1ki3X21mngY3LXL81vV3JcnyGq9a1t0Ydxc9yXho/KC9YeWhwrm
BxdkewnykaykAOP8aQ4pqb6oR5VN1LXt/A9rHuvbvap3Tom+N32VN6r8GG1v5TSus30SgfiXldux
Qej6NtwGRJqDJKUpbCz20g3QuUN7qDZJ5LXuW9SArIF6Ppl/Q5DuKaDbTxNhoaE7wl9zdSbaMWtF
WyyLRjjlyTWNaI3Ow78tBP+Xf5bOyf2faSPu9xykP230A3jBhcmCn7lKpodbwWBpdp0d/wIMdxaI
5a4eOJPG5xiowrDF6GlGNFZ0nFEiyusbzhahJF5bN15EpvXjcAhWDk0adSLJ6JvLlXTTigL401Eq
5VUAao5QMQ20Rq0mCw1mdMyl6+SC295KoVUXfy42iBHpA8SYOFUDOGpD3ZeAD7+dNaoR+3BAoWQ7
W1/yuz/N2Rhiyv2pm7ClkAY3LWm706acG9z9ertV+yjPq5ForBCf3O/Czj0XylzPYrBVcQv5GTve
7IkPeU3JvOqxEFGzZu+75knJlNE7ZyKrKmHbuHJMAht/FcNgqqc9KBYO40ZvVz7eR5yrxdoIU4ie
iOcLW218K8Wc2aaajFXLOOqZGp2jlInjQ94iipq7i3eZTLQMwMCPGXQkjei2CQSl52u45R5Bh1fR
njYaeIyaWN/cp39rMp/IrvWdxmWYFaKh5yRB6lhj5IHWjj+PmjMSZIOzsonfQX7u6VvHK+h9nVLX
mbFHa7gNsF+BZRJq76XH/JJStgkQAQ99BGBeqb7LENwoqAHgcV2bHLS4no87gy4QG1QtbdHFxKnQ
5KwOFLPfx9Iam8AfCn+IoSfjO955DeUMg0mn7ysednqBSdD1ZUitcKlA25b64e3Q5KCY+YCp2MUF
TFwMx3Volq6Nmw5DlZkfjfQBoyks68luEF2PWURG0Zq/Zk3iB/J82pK17XrgSKphccSc2gxDBnab
r593jtupglRm05o9MmDXo2sQQRhOOthzV25rLZ8Wyq4FCd9ib/Ntp/LuUWXCOFlfMhgnR/tVQKaZ
ocVvC5I/J+9+aek1iB8Bb9iMWVFH59vqpFjHS3n5AEfK3LgBslGl4d3WKXTe59Mkitq0FEd4N7zH
30SX9gjv8+31CxobXl0tEaN7QWCqcuSmueISuvV7s3o4qrQfrhbwfFSP3ScXO8HCMAIR1b1STh5c
7PuVd4ipyueYdu9kAmTZgx7a415a7dy37RrOo59tK3jFwtbH7iLbO1rMYmp03xQDOR1ZFyY0sVtx
fcHUI2SrmROXDPw+xAiG2QLUVVD7vPuz1FUKan49B+435tK33QSI2I7q19dR/xog5IFFMwzQ+f//
OC5cmjZ5+7a+2KAn3mu16iiY6G3oDo3QSoG2Gj0JX4ojH9WxAssnFmkXisJWLY8qYLwRTD6DEHy2
R/xtGnZVRhFfCqqM3cVxHFYvxqkbCS59hluYUEwa/NZXxIMPqhRfNY3gtTWOMUErJxUH65B6K958
TB4SAL+ICbr85Y3s2JanC5ah4H/kR01T3g0BfhuktPP2pZbRerCyAQxVcyc+pL4EwSS9HbPQf+u+
F33og0RA0UtHvpRGQzkrMaeKn+EdOjcPds3eTytI7XY9B5joK3i492nAIsXv/iSpuRgCDf0D5K9k
WraMf619BsrM7DK3qJSIGIJ1Qrfur6lioT8Hh6xPRmDtSvWNCLBEQ1feoF2qB/yLl+6MJQUQ/jIl
2FLi1ACYD7tyJIdVMwa/kC2YIJtn8an0WXluuCeAYyJFlQPeWh4Ad6KwjzKuUGiYKdupZYXatbB7
LLVqfvilJXvgL0Ojgj9OLsmdvk1KMnX9Q17NTZYxyBkEAnxZZvxAcU6tAi1RmCMGMXkn/lDBXhls
WcVLyFVllgIHVXl9vWHTLi8JScxTO5TYmNu51wsGCBVSp3eB9HpVXPu+hlRTDEsSv0UGePKMPWbV
+KpXF1U/IWr6jeFh6lQIDkY8cmMBuHUCcEEvTX+DO2Cp3/f0YpDeQc6KI8n+PBpgcrIxLzRuxLrV
Gv0vhYKK2b5AoOe+Oag0+zGzJICd6cNeaebvKJQoGbO3iBXMKQ1lN+myJD7ZUpaVpomllZMi3T5q
lU0VRzAXs+Anjhi3i927R2m+hbleLR05V33j03QSSMr+Psg8djYeY/CMJ8k+oOeTOHS94mgl8wko
sR2zXFvfv1z6/8TIKg4WQaW5i6kpml77rDEKAMVwyQwXv1uuBHwSnZ0ljy2gyU5XUuY9xyMmYeBV
l2FW7RAQC+yq26ohxpGoSosvftRRiis9Z3fuEWnfkLVY7duugxEtS+TQH+gVO6EU0/4hd4rxxyyo
7sFzr4VXRHqWQ3GdrUwrqDrklu74oOCWdCkgsx8SsFjFwlegKQoxglGxwKeIQvZRTQKY6yWg05PS
RPP584vD1rrCiYSwtju44pDGXTSoyJGb9tybtflZRyphDNb6A6kWHaxweDd/z/Q0h46i6U294Q6B
L5PhEo8pSNPAkYlGK6z8ZH8BnnkkbSPShWfPe+I+h2Au1LTlz8rC6cw7MDZCHydiQCkVKbURS6rs
Ixu8RR06WVtvPlyDCLZ1UGh1H9Q3pSezoIWcd/zuiG4rA8zaiuDTDolbmy7vatNcSBv4wouop2AK
OGnLDWpTo2VXGwMvnL3/8j37eW35q0/0SGOmbO1yGlNadSEOKiikKqR60x838+kpmm98cGaHSxWN
4/KDdbQ624W+laaVBOkHC6u7V0HI7GK/EbKDtqLn8THtHcfWORnqfwehZUvbH4y/y2hZzRLm5l1U
7hl+WNTunnfcr11rrzryiQ7T+C6RLl7lvUfqKub9M9oxdRCIC3FllMTS5yCb07KytPd6+C8IsTvi
DhBRSBf/sbaoH+xTW9d9/H35TOLCBHAp7B/Itguaj0HoECvrqdjkz9K9TbgVdOTDmrh/lCuhJNYA
oSKSTtVH6kkJ4iSQ7fsk7t5bMIeLG5i36co5OPjemIKdW8WRnvsrdsDyn+FtAR6UF0Q7E+7mBEOc
LAeySM4t2ADYpM2t5g+03tXKEnKPGGQ70D5xCU3SaFlIshskeWraYkSpWxVFM9FfQnhUVsxvhjXM
fa09RgbDs8ceyHFN+hpNlP4mEoXOLoN4dpQuLSmLbKu6B5ixA2bkFTzpyxHu7OUPenhnH2lgW4+B
MvmoeOIDaO1qliNdTsZfLULYGMmtxdV1izBHFzfoUJ9UTGD9xQqsfiXx55XW3waTJV39KRYi/m+w
5T4pZQFdiXDCcAwfgGCtubI+4+2r/nWE2Hew5c0lXqOA1HUutkBtLtrxoLb+5H05XMBHYBNH4YjI
BDOh/bHNEt3ybh+4htL3DTUnsUkeESLpcS0Gl+KdjKn047qrkySt+OpAX9SvWoRbGqsliUggcHVV
hAp5+rsOJOzlOHixMFuy25alJ/8awSn0zO/JwXBhqjGZBhMdnKekESj5cNN5KYCpUIy+VyxgRonH
PpBSBietFXrv24uWm51A1nZA6i4UTLwB5OnDUscyuVZ9RqXCPZ4389xYFxpSkqhZdFS7GrPAgk/K
06/BKZ2NJnhJ9BYI8XeTkZgstc08jyqUzx2brxLqvFx8xPtxwbBPkirI8NToAPO/gKvixyG11Ixz
PFEzhdH5KU84QeoS8QuqzXF8h64TI1b29eVjDbBSF33otJfERuJV0zk2qr1+Y7yYPkzX1CjJBV+R
rnrjpVviG/8pAEUWNA2mL/4LTGtHQOrURfXzdNtDupS0tKHJ7YNmm4znpQqGN0QdfMdrKkTzF59I
Ev0V9MooF0kIf9ppuXC3FPW7pNqaQ4DMItAWc9jw+pKqUuOnKj+MiNdFRR7yxc5Y89m/iwoa+GTW
0eRZbOi0yhN10RRAqNfNwNRT51vf8bMI+Puio5/lxSuc9m7UQhEHp4F4tCzUMIdhQecEn3letIkO
WkE3j5H1Uu6THrj/SMmL55nMRAiHPM+/XeKDsdnQ5y2spkHlHC+bQjXITwADK7MY22gTatJt9kmD
BIU2voodEL5sAJjuvmDVvHDLVf0+eqBsCBD5603SvDD/Uro0WpgLkAgTwwmdLlErgQWtXdDswD3b
+7n344ZYNH7Rincb2MRpMaoCoLRVF7RRNazx5Q9WRDourDq5ST7gi5dKIDTq8aKcJcYTugmG+gNs
sOSpbbCYbNpCAyRZw/jpnn1jYbCxDI9TLmFEWCBezTweL4gPYHAGPTWLfylA0IucRLe9d4FQvzUX
cm5MlJNufpSRK2KgzPZjFhsW30/FhkV207RDyr46iqD2JezUMxGeJh8EjMFCDITUHIpGwBKN4lki
hI+Dhk5MXwO4d1JtSwwCcA5zsf8E6JCgJKdAkRj9nXEy3kStGLLqtISprqqbTDarhZZKh7zoaLOk
RQVodmKpghyuLqg6MPBNgHGjxonL+Z9E/cQjZJh2vr4EPg5CsJZqdr8s3WbxncF5Y4AsPLePsEDx
q9QOi+0IpQp018uAKlIMHY4YgaiQ2bbbg7mfxL8y8dEHvFDf/QGDIvsKGsg0q+F6F4D8DNunnlJb
Xaty4LiJ76wu8VTFPiXZUoIZ9JVSTwz8r2YbSSRE+vq2RbwOH6ccTqWWC36hsY0eUJlhoOin3E1m
sxZdKq1wlkLV+/JzLO/WhZ9kXG1SUkpx9HhSwiWgdAx6ecmjhbRuqdpyjzNPTJbz/PRz/iyxRBhL
e1TsO7w7GYfVA3T9fH2QclPInGMCXMjqfW4VJV42cCFFWYSsQEh8ykxOWGDg0cefXHvhS5Ep5xvA
oKJje43ItDgtHaVM+AIGl8m4gFDj0I456yBh5zbGiSv+OU621bRVIfYlrAojKN90w3/OaODANsbL
TH2Nq9gA0Zr3VRGrwjtv2V3qVYPuvAQZsgNu1TbQ7QF+i2siY0+JFQHuE61SEuxgK7hilgLM0UnC
rP5APHjJ+0BwIXWth0H++pY1dZrnBf7N+mOH4RUsr7N6cKqhpJrT/yECLm01Olnpi2PoPoqjF+zN
U9cMLor4IUmwOYNio2DFvo9l0qAyKK0uPBu+pmZMY6pb4Rxpks8stiEl13JJhXyCVi4WGanPHOgo
QlrwVz9mBcljyFsFza641ZWdl1VRv1IZFg5Ft54dtlnclPbFfIgCYc0g6Z0KrNkS2ggR50RVPocR
b6+C1bBAF0I24eS/NeStcGib9/fr+VhHJUtkKNS4uXQpLRwLiykACYNIGSasWOfgq01MGnpCWh/i
6wik5yhkIVbEjUOf4UMn+2FgfB0rkZwcUc/cFoc/65MfDBlZ/u7A2XS0Ejrl8o3Lsx/G5bG9NHrJ
k9YKsc/UOlhyWG679+PHS8uTVzlzXGONQhyjVBSJadR40Eul2CBDI2U+DRaakElX2aiDc2wxHPIE
3S3ppUUmQAeRe5CgAY/tlxSrJILYMGwDrSa6+UK2cjzi6LA3NJmItWYpoZ+cxOSYmDwpFnEF5I6f
xh1cuzQa1lEDD/pFIM3DHTujoYZBZZ8sxaVZ8StPjTHlWOAJkA1ancy0ONXCj3/EsaLo07wtpTUa
RVwNBgq31I4O2pUkpEObZ5bBiI2lXEPX2JBCNF7vtJB2ZRfLvZL07zHjbsCpXVrBkKGn7zWPMfAG
IJZ1S+LdPw37DtkWIdVf5t4Vi3lFKtVYeVt8ZV+jl8dZk+TlORPFbdy9GbIZdFGZsius3HEOd///
huvZJeJbS2eGQqUUPY9qUF9Ug0DqJ+H73z8ZTU8e0mJxuBsCXp2yfGxPWF+rUQKZYnAkR04n+igt
cIZ73FLWu67QhYjlWq2DtxlwmtedB6L8US8U/K3fmsipd7Pui+jZZfIL6oxEzjIduSVRwl6MQlfk
alg3dWcBh7KU7VlxDM5mgLCx7CUcNsVujvbBtfPasBLdVOMcL4vjFJKLTzwDr3isfVMzwCgzr0qk
WoKymLs/KpRbkfI02DZN3BWz5P/dLevhoPYFds20mLt3ujzEjHN69x8vuwcfmPmBvnw7WUmZArnj
sopEy2ZynRDCHxlfEAeQUFmjZpzSWOKgVbeYoq8UPJ4GgWzMHSUvUJxjN4JqGvVcxeLkNm9mRMfX
sVj9B7psc9hZzbz/5to7TJj+Dj9SA+ZEOPk9AuzaHV8xLFIjexUlC0uspjLDjHr85fGPCcEOGz1t
WG7aR/cJNWTa3hyoulvqkUyNQLMW3bE1HjFaxccRgYWpSUuV39dLW62hKobr60k1IYnn1I0qbAh3
aZAixGCRTuKWdx84lE3KhJ7FigsgpeFQqgtOHhFP+lsfzFH35ZL1Cgz/ZjRAVcIlJCu2j9VncEdx
O546dqCPEfVF9TZocj50szoojI5auiHBLqQ6nNW02iYcsEQ/f7ZHkHYMtAAsNIUEFDOiP7lN7gjR
9QdpeWSGtbStk0srNzvvw4XfIpAF7Z0WUwuQP+cIB6CloE9wx0qbBtR5p7sAy9EPFbCB0/I5F7Kv
4khUuP+N9F3Ae9N3kvogj7WdQcDCplYyJMLy0K6PFuIvG14jSQ8y/6ott/2E3j50QteFyVK5WPCD
z5twog+mSnFRzPn21TmRcp7gnolRGC+WgZSwv8vVjm/Mf8FJNE42vu7o5NGDVoUaItTmnSwZ+Wz0
J6gn0qYX2ozMYxMCQeFvVr6lqBes58W3pUH5X3c7oDUk7SlRPyavoL+IiyNbx0IUkGDng6yhaWtR
8aJXUGCDCjkUTofZsi8vwqddYZZJpG7CITWYD/6tyKPwHjwnyzSoeVNCl343kx9y0S7qNWa/M2q7
iuUb9bhsMeiyYd2ul/qJWBGJA4H5sTOwLwIWOjfrH4dfF0138gf6Z+nLn/65VyRe52NTJ5B9gvBI
xGETIs7tLFAkSICFDrnebCQ8ZOcIynQ1budMoUEsu+ukW5ng6mVp2bJtDpX4kz5isVGPRSPUORxy
SPunFYrTCK9GOOVscATabEaOtu9X3+2IjvcpVC0NMHFKTOMOGhG/hc/91Desq82rdYeSml47qSiI
AIvXBK7uG9Kp/yZb0epif2jPdLQDtKY4hbp3DeEyqrRfDfguVulLKVkJnDESJRX3Ie5i394WjQ9+
J4014Zx6qhE2kPxVwD/l3NmcZeXsp5JYb6BmsEKUjF1SaRoTRhCXded1oSF3pOwbRVOMzz70z7kN
dLLrR0a7KYzsofs37xUTtp7UBflpV2S1srBjh82rGss1F5jeZnDZnHEAvYd2CWiPLppk+9DW4c1l
bfObt0zCSzA8t9GiWnSCMKOCjjoRLgYFhxMmDG5SB91L7LflNX7iknYpYer6EiD9bACVxsGRSlX1
YfcML8btFF/l1oOX9ia+UuT1qq7B59LSl1HxgyD6ZgcBNj4S3FRpQV1/02Q3H/x7/79Q/cENL49U
7cnd0Ha79tOJsrI8LY2FWxelOCmuPVxTpY3FjmQ62vOQpABGHSsIMk3F0mpOCygaNB8gegKcyB9V
FG4wjvEIBDOUDBYh2w06hPscI9znTqnaYTdxRc1P5+gD4k5cyS/SRhquxBIE/e3kWLRUJNpoaAW+
ptU8x9Ks0tfez3m5/KscDBN3tzIofVMVZkeWgUDtVb70Woc/LRUGflzGERrm5xtWJTDIhWm7Z3wI
pjI2dtT2nZ5Cwyet+HjkykPEEs8dJAcMhMtNZunYuxiWiRUWcl9VGltW+0Uj4aWXpgorxRan+uKk
HhfphkBLWX+dQHehFhU8jF1Fj9T9hyvw5zEFTRY3IxNSogfQXnFNJibJHaIqQXiPusQRM3BAY65g
ybfcmywNnk6ekDMHVGnQc3iTWPSyKjPaFvDqLRykx1tcThdO4K/L/hUAPjyEmGsm9ruX94s4VO8T
zg6BbY8M6qxQbhyVCqIUe2MuP6HzppyYq7fCvQ8MpYz//kycOYW+eRR81MVzOiDfnUSL9R1wIYOq
3b6hyKBFXtFOEXpSrL9hJkg7wJeSOtl0b6Rh2ykdPmeEmGrx0OyXLeUlTpHwukS+MCSzOtOhUz/2
a+7Hf7rPJM9AGmj9Q4YFAKwKr/1PRYHMl1MGrLkKmdoPZihpw8dxqpnoQjjGDeGF9my6vtMidZkM
dhcBO2Rebf4gF/5ppXhg+ozPln4rvMi0j4R60YXyb5M+rc85xfK3dBhWCGFW3AbUvVuKeum5qlLC
Pk+mhcezaINZOM8NyidZRuSmu8sGhSryEn8NxBflhWS1ziHgyYWvBucGPiSTjkRMDxQE/EKFl/fL
1KxD+Ov0/I7n/erILEalqeYWxU7kssqGBelrSrGcOJhA7DH7RmuJ+iDOYni8g19Ox8j1hHUeIV+o
yNMTPuAuAGVXy21ZR06aGXCDMAGghbiRmAvIo92pWCAe8PbsOoZi+eBQW+h5mvmP4Y1Wl0ZOgdDh
B9gCtr3tw7j8OF2otj0GVqsYUiMqF7xKb3zqE8+F299vCy/CYhvUomf5Pj6VSbhPkKnGsNSQ491a
MtZ07zYB9aIrF9OG30cjfXur+SHPN9eBypf707E8Js5Lkfb6lzbZCzZcvW29YMq1iaJpK3/Ec+k9
/kLlhZWBzk9e+NEkuPPTRJ0w1sVtgc29Rb+tg1cjp/XUnUFg9zefBQppB4h5KuOIE3MjJmuM80rv
8ryhwofyisgZdbOpgjVPSOH8GZCoTVpZS25L+OMJ2VnHH9eYJhLkHrXU4qLpCv+BknJTSIkX//V1
ntXi/l54vwD+Sdh0vm43u9R0S2Zumv9j2EW4V+zPm1Ngv2HRh+U9Wfwijjyi6Qw7pi/H81lbYxRa
lgvFN8DHHfhDniLwe68qrUgntzneD9lxXcEcUlfBGIXPjxzyrwnehebySYtvRveL9O1+QxxAL0+l
liBFgrUh7gh0kv845mwhGxJvr/5UoeL2/RyFgYOYUQjgZjQExFnBq8mQbd4B6kopGIYqv/xcmRru
4nO2IfXx3nxHHiJWkr/vsM1OTM47kyQP4afupvUozd5mh/41zehNH/wf4GrKqtIWYUukn++QIQ8Z
Mu0k/cOj9Ki9/hdGt8uvLTJAA0Mjl0cfDUG2x97cmoR86fvkZ4KPyvX45/jl8CPfhd/7d4mrf9cs
7jGxu+6n+A7RNHPp9shu2+WOaYGT+s+tD39fRYL5Sm7nSQ9CXYiiIy56lWlWlA9KRm1AyX8+RXV9
DNx5yPzjkB9+/vaE1UElBhKeeuN2xDv40P5kV5nGwB/bcNY3P1iNoumnnwqMYV9JAPgIIvgPhvEb
GuUMUTS1zElSpftoYTY4sM6zFyusYIk0XQihOanD1arq4956EO+Qi3hwKMbs+T170y6TdayP5PkI
0GP9kLrzM4q6eJsFe5VpEZWtMq78GwgWc+dbXzjajEEUYWKkDDJWDEWOOCZxKPs5J6FDF0+feYcT
8OJPJuWZ9Sw7I2Vp/eCvipMGm5032ZvP8IPnUTcL3HyWT64hd8hRiq96OG7UqhkdCfnkoeQbIPvI
fjyw1Oba+yn54iLFKQbtbkcAkNvmzX7RzfhYnpWFbetx1bRA73fDJqYhZ1fJM9rhHY8prjvLLSmA
7zxppUssAAuW7RhcmtTVUulOXJjhjW6uSFsuw2nPBgb0f3LEtkz66l/eidSbMR0B3mtwB0JwORyW
Uz5R6EZdPO8/pMFD2RLKyOvZjmS8xy8lq6rP/N3liCTncVIbxoHhNBqoaakmRe8zAwiDC6v5GuOM
e9sEcwjCv2ZJKNTM8ZYa4Mcg+RuHY8Dc/A9hCmnGFUsoE1lmWpdTX64IjPMhYu6prUt7k49c28IS
Y+gBToT7X+DIKZw15uKOPJ8CvyV6ctxuJc7eMTgP3eSKT3bkAYWrXhKCLCWiF9KrqWQDBAW1+ooL
qJ2NMHWGfHMzZ4QYiRcn4JwH5PljXDUT3yWx/19luENfsIWqNujxx8u6HWBptsjp7HdOEGgz3Z9K
YhHVOG5+CbLNeelUW1THHZaY3wGRbYCNks4/aLthIa8l7X3fbLnohQyeX9wVqzVpTX3WekRI03xJ
tW1IwN62NxoALSUAt1lAo/d+36EZTFz34tnooR+pdY3CceUBs2HK2dNveuMHhESOLSgMambfhMgy
rxFZ0dpyNfy82amHy8isZhSJeBKEWCunvgU7huzHxKOx5x+lFmoVMBHBw47Uz2i9Ze9UG8H0vVjE
Dx711kCi4rgoakDzLxFjCFLJhFV/7gqrKweeYSjWbYb4Ox8gho2vOgXzXBniZwbpt9tzcTX//bsz
1SnVuMvK829T7GuS+2jzYmStWPwMNBWhb9GKxm+rpzeJVd1qMDGVqF5jRMmNgWP0pvAtA2AlMeGy
I8RPytig6sIoYAP73dwqN4FSAZyw6h8IClHAQKv/CXS4ovnRJmn41PVC6T4/766Y1t8i2Fpw2sId
iNuBLfohRXIivdgt0LUbFNnm74BWOt4i6UP1ERq73w0SLvvG0zUPxEEVoC/lNVzF5P4djpr2Ti3/
4nmQbN07bjs/bKMfcuVRunz58grL7Vj+XKrVQsc8Ch77Ig6PhzhCakHCbBSCvmS2lSTP5/ChA5C3
LzOubPuAcNS16o0tNlCHIcTKw1ufvc74VMVIutZN075Z75+2RqTjQ3Fy/SA/DpqgfQPVNxH85YOO
GJrUQQEBb/tHo96m7Z4YqiIENULi5TnLxzE+0eRP+ufnecLGaqZINK1YlffkLQhvNRazpLBkwXe5
Xm3Dazd/pa7l2TfcDFYzZoOtwqpxGo8dc5PVoPRPxcVOdfK3YSuOK7pqIw6sB78wL+BI7vLjvw7h
yMjmhBDjqA3ueIaDq6WANFtIfSZC85bcR8CrQjrtgWIAalzd+V7UaD05rfzB75ZBhNk0gXOow7x7
D3ViBKrQY1vT+8djugVW2Tz5oHzqq/bDFDbGPfXN65MQIJYPUPCq6NrjOKqmTlpWSxoh0EiX+FfV
2NzUl6Pqe4EnueYtAy9puEl/baHqzdIxsoUu31zQCIYYt5XUbLaI9rvr9cazSYd7Kfwax5+9gRpE
siRFr85ju8/g1+iq1+J7VR/2yqYGfkIKPO6tgmslplDzQ4G96b04S10VPTauVqVNgE43vFIW41Yr
PWFzqvhFJKnUtWeIYx8icKWmQVC4Q8ML/JIMYYxuAE2N3ZM2PP4shXZs96FyJyyGVCI2LNyNL37x
6aESN4gcCJVvrX0lqweYBKuJmybcHJ7K+hhnQClBsnUlxNjP1LOQ73dkVrO+LOows7Re/piCICYe
EnWcK9B9Kf6A6FigXzyAzB8VbGoqORdLEV4I5JWumgd867GQzrH+rWoqefl/cPFo9amwMgEsW5AE
JfTSCyk68hOzYuNMwLbbBYDHxJjRN+NAVlCCflWE42ZjJQWWnLzb9sMMf7D0OAycW9lEcxXLancg
FFYU8k0qrxLqJudPkXSxJ6shJkDZvdRbuB0kuc40OKbUzrNMuq8vWxX0rhHIAs0VxzCWGjWPTSpA
6FchPJhfdJEPppkF+waEJizT+vxcYoQ6h9SMABzK5Ro6zxE9TrMGkyd+QYF6nM/o6Q75Jv5+zx3x
CYT2AhQSDQwK7x92PuYUDSDHxRJAB2cu6/mazNNvq8Y2GSVQ87f6X09vXvLfO7QttJ0Ikm3YKZJu
JgFp/xE8mgTYsp1zAxkPYvGsjR7qhqETpdJAHLKVGhbT09V1Oy4dAc16N71fd3Y+0NbDfhxNDvh8
4Xak13t+ZRwnlbDjg0xbguxu4DALfYcYT4NU9VhmPPFCvPtyHhB1UbxGFO20CPpe2//DjBzX8zTw
ORSsnYl6rHgFmnYNvXtJ3ylMrbdwJCi+GerLN3BCviZMXS8qyX88l0RZVvElgzzSYq2XWBTfzPoy
iVssXfCxri02Zgtk3eYEZRodV8AVteJOP1HAlS0S53Hm/yQfSJWIC7PMTsagPlF9cDEbYCphPvsR
i0g2DqEXe54kyEdzvduF20J31v0WkwGP3U8HI5n1CXUKFRbC0szpx82BRgpXgO8BQCqGJJtvNvaW
HcPpvGd0YgsAnYvHRTxkYYHUqR3jnCxJvbTVrR2VQnD/A7Vl8D+pIIoE95Mjef24iCa/T9hEiUem
D2NVK+4VUs5EFyp+WZ0o4rHtcwFbaWiACZ7GxyqpmOaqzszDw0VZe6+RQLWf8/rrt5Y3CwNnO8eq
pBkA08fvcTiUzzs5umD1QKxyZ45WuH/48Hrrn+5zO8BY9gBicUe7Z13DFda92IsUQHb4BH8YUOIn
qvz8oWMA5E20KITygZGej7UQinaqN+nMAXAknvDefvfetwnrYbtK9a1AW5XYMYW+pmMo9HZyWkC8
57CiGV61dPssrxpFZW3+VNoxyrINp/QpVmzP2kDy22LRdE/gH9I1mzKrkc5I416kc9p/Um7sHQg5
KG9hpiK36CNuK/hxu3NlZhlMpAnMUJ9X4c9CYRRO1hDYZYbvgnIFQ8jNkiN90dwwIVItLrxhv75h
UlzyQvybUAAU48ex+Q5+oWfNZdU71UArYt+vLP0ulFik6h4ntkvvGRwMQoII314Dl54xFNRjt3QM
uLB5uqBLl4hFDiaw0Ub5HyWAQDQtUCcWwenKUZ6Xr03JpcVh+u3ScEwL6p/LJPnJzVIHO8fmcsHN
Z0GpVTN5lWOfsm9tPumfZXhPFZ9qk+Zlfc+MIqQjrv0kvlmSVSaeQXXze9xgDln3oItruLIKJOD2
czsRf2KoUQqvqsqzDfD4EyRfJudK3tk3EM99a9RMfXsokZ4XIGPS7icCJsowq0NvkHqkNbuZGm9T
8AvQQl1kfjakSfqPOnfM1WYVouJfLKM/Fd2bD212PQXUZmcZXLJnShCCY5q1lqvxI/bMdtXLoUxq
vbuYbsaAkFmMUt0dca95aJu01PSAOiPc6Y1UPdpmXMaND7zwNA748wp/kdYJVU7wZbHUk5uiOG5D
4gcD/3DX7Cjc8K5LdBwhd7JBJW5AukWAcPKYQrFpP3oqGBaJLBDh9ZlwPEHVuXaiuuzPc5fazzQC
fVtYC4cg5Q==
`protect end_protected

