library ieee;
use ieee.std_logic_1164.all;
package nic_Type_Package is -- 
  -- 
end package;
