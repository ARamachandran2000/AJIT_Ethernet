-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity AccessRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(3 downto 0);
    register_index : in  std_logic_vector(5 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity AccessRegister;
architecture AccessRegister_arch of AccessRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 43)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal register_index_buffer :  std_logic_vector(5 downto 0);
  signal register_index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal AccessRegister_CP_0_start: Boolean;
  signal AccessRegister_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "AccessRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 43) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(4 downto 1) <= bmask;
  bmask_buffer <= in_buffer_data_out(4 downto 1);
  in_buffer_data_in(10 downto 5) <= register_index;
  register_index_buffer <= in_buffer_data_out(10 downto 5);
  in_buffer_data_in(42 downto 11) <= wdata;
  wdata_buffer <= in_buffer_data_out(42 downto 11);
  in_buffer_data_in(tag_length + 42 downto 43) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 42 downto 43);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  AccessRegister_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "AccessRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  AccessRegister_CP_0: Block -- control-path 
    signal AccessRegister_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    AccessRegister_CP_0_elements(0) <= AccessRegister_CP_0_start;
    AccessRegister_CP_0_symbol <= AccessRegister_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_sample_start_
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/req
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_sample_start_
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/rr
      -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0); -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_sample_completed_
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_update_start_
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Sample/ack
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/$entry
      -- CP-element group 1: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0, ack => AccessRegister_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(1), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_update_completed_
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/$exit
      -- CP-element group 2: 	 assign_stmt_77_to_assign_stmt_95/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1, ack => AccessRegister_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_sample_completed_
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_update_start_
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Sample/ra
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/$entry
      -- CP-element group 3: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0, ack => AccessRegister_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(3), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_update_completed_
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/$exit
      -- CP-element group 4: 	 assign_stmt_77_to_assign_stmt_95/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1, ack => AccessRegister_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_77_to_assign_stmt_95/$exit
      -- 
    AccessRegister_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "AccessRegister_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= AccessRegister_CP_0_elements(4) & AccessRegister_CP_0_elements(2);
      gj_AccessRegister_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => AccessRegister_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u5_72_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u6_u38_75_wire : std_logic_vector(37 downto 0);
    signal request_77 : std_logic_vector(42 downto 0);
    signal response_89 : std_logic_vector(32 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_94_inst
    rdata_buffer <= response_89(31 downto 0);
    -- binary operator CONCAT_u1_u5_72_inst
    process(rwbar_buffer, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(rwbar_buffer, bmask_buffer, tmp_var);
      CONCAT_u1_u5_72_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u5_u43_76_inst
    process(CONCAT_u1_u5_72_wire, CONCAT_u6_u38_75_wire) -- 
      variable tmp_var : std_logic_vector(42 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_72_wire, CONCAT_u6_u38_75_wire, tmp_var);
      request_77 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u38_75_inst
    process(register_index_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(37 downto 0); -- 
    begin -- 
      ApConcat_proc(register_index_buffer, wdata_buffer, tmp_var);
      CONCAT_u6_u38_75_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_0;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_req_1;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_88_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_89 <= data_out(32 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_0;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_req_1;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_83_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_77;
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE", data_width => 43, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end AccessRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity NicRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity NicRegisterAccessDaemon;
architecture NicRegisterAccessDaemon_arch of NicRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal NicRegisterAccessDaemon_CP_116_start: Boolean;
  signal NicRegisterAccessDaemon_CP_116_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_179_branch_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1 : boolean;
  signal array_obj_ref_203_load_0_req_0 : boolean;
  signal array_obj_ref_203_load_0_ack_0 : boolean;
  signal array_obj_ref_203_load_0_req_1 : boolean;
  signal array_obj_ref_203_load_0_ack_1 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_req_0 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_ack_0 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_req_1 : boolean;
  signal W_rwbar_212_delayed_5_0_208_inst_ack_1 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_req_0 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_ack_0 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_req_1 : boolean;
  signal W_bmask_213_delayed_5_0_211_inst_ack_1 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_req_0 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_ack_0 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_req_1 : boolean;
  signal W_wdata_215_delayed_5_0_214_inst_ack_1 : boolean;
  signal W_index_216_delayed_5_0_217_inst_req_0 : boolean;
  signal W_index_216_delayed_5_0_217_inst_ack_0 : boolean;
  signal W_index_216_delayed_5_0_217_inst_req_1 : boolean;
  signal W_index_216_delayed_5_0_217_inst_ack_1 : boolean;
  signal call_stmt_226_call_req_0 : boolean;
  signal call_stmt_226_call_ack_0 : boolean;
  signal call_stmt_226_call_req_1 : boolean;
  signal call_stmt_226_call_ack_1 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_req_0 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_ack_0 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_req_1 : boolean;
  signal W_rwbar_220_delayed_5_0_227_inst_ack_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1 : boolean;
  signal do_while_stmt_179_branch_ack_0 : boolean;
  signal do_while_stmt_179_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  NicRegisterAccessDaemon_CP_116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  NicRegisterAccessDaemon_CP_116: Block -- control-path 
    signal NicRegisterAccessDaemon_CP_116_elements: BooleanArray(50 downto 0);
    -- 
  begin -- 
    NicRegisterAccessDaemon_CP_116_elements(0) <= NicRegisterAccessDaemon_CP_116_start;
    NicRegisterAccessDaemon_CP_116_symbol <= NicRegisterAccessDaemon_CP_116_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_178/$entry
      -- CP-element group 0: 	 branch_block_stmt_178/branch_block_stmt_178__entry__
      -- CP-element group 0: 	 branch_block_stmt_178/do_while_stmt_179__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	50 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_178/$exit
      -- CP-element group 1: 	 branch_block_stmt_178/branch_block_stmt_178__exit__
      -- CP-element group 1: 	 branch_block_stmt_178/do_while_stmt_179__exit__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(1) <= NicRegisterAccessDaemon_CP_116_elements(50);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_178/do_while_stmt_179/$entry
      -- CP-element group 2: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179__entry__
      -- 
    NicRegisterAccessDaemon_CP_116_elements(2) <= NicRegisterAccessDaemon_CP_116_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	50 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179__exit__
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_178/do_while_stmt_179/loop_back
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	45 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	48 
    -- CP-element group 5: 	49 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/condition_done
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/$entry
      -- 
    NicRegisterAccessDaemon_CP_116_elements(5) <= NicRegisterAccessDaemon_CP_116_elements(45);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	47 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_178/do_while_stmt_179/loop_body_done
      -- 
    NicRegisterAccessDaemon_CP_116_elements(6) <= NicRegisterAccessDaemon_CP_116_elements(47);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/back_edge_to_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(7) <= NicRegisterAccessDaemon_CP_116_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/first_time_through_loop_body
      -- 
    NicRegisterAccessDaemon_CP_116_elements(8) <= NicRegisterAccessDaemon_CP_116_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	45 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/loop_body_start
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/rr
      -- 
    rr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(10), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(9) & NicRegisterAccessDaemon_CP_116_elements(13);
      gj_NicRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	20 
    -- CP-element group 11: 	24 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	40 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_update_start_
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/cr
      -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(11), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(12) & NicRegisterAccessDaemon_CP_116_elements(16) & NicRegisterAccessDaemon_CP_116_elements(20) & NicRegisterAccessDaemon_CP_116_elements(24) & NicRegisterAccessDaemon_CP_116_elements(28) & NicRegisterAccessDaemon_CP_116_elements(32) & NicRegisterAccessDaemon_CP_116_elements(40);
      gj_NicRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Sample/ra
      -- 
    ra_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	22 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	30 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (29) 
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/index_resize_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resize_0/index_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/scale_rename_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scale_0/scale_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_final_index_sum_regn/ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_resized_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_scaled_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_index_computed_0
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_word_addrgen/root_register_ack
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	37 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/rr
      -- 
    rr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(14), ack => array_obj_ref_203_load_0_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(16) & NicRegisterAccessDaemon_CP_116_elements(37);
      gj_NicRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	36 
    -- CP-element group 15: 	43 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_update_start_
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/cr
      -- 
    cr_212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => array_obj_ref_203_load_0_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(36) & NicRegisterAccessDaemon_CP_116_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	46 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Sample/word_access_start/word_0/ra
      -- 
    ra_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_load_0_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17: 	42 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_Update/array_obj_ref_203_Merge/merge_ack
      -- 
    ca_213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_load_0_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/req
      -- 
    req_226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(18), ack => W_rwbar_212_delayed_5_0_208_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(20);
      gj_NicRegisterAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	36 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_update_start_
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/req
      -- 
    req_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(19), ack => W_rwbar_212_delayed_5_0_208_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	11 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Sample/ack
      -- 
    ack_227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_212_delayed_5_0_208_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_210_Update/ack
      -- 
    ack_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_212_delayed_5_0_208_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/req
      -- 
    req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(22), ack => W_bmask_213_delayed_5_0_211_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(24);
      gj_NicRegisterAccessDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	36 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_update_start_
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/req
      -- 
    req_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(23), ack => W_bmask_213_delayed_5_0_211_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	11 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Sample/ack
      -- 
    ack_241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_213_delayed_5_0_211_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_213_Update/ack
      -- 
    ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_213_delayed_5_0_211_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/req
      -- 
    req_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(26), ack => W_wdata_215_delayed_5_0_214_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(28);
      gj_NicRegisterAccessDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	36 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_update_start_
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/req
      -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(27), ack => W_wdata_215_delayed_5_0_214_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: 	11 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Sample/ack
      -- 
    ack_255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_215_delayed_5_0_214_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_216_Update/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_215_delayed_5_0_214_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	13 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/req
      -- 
    req_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(30), ack => W_index_216_delayed_5_0_217_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(32);
      gj_NicRegisterAccessDaemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	36 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_update_start_
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/req
      -- 
    req_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(31), ack => W_index_216_delayed_5_0_217_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Sample/ack
      -- 
    ack_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_216_delayed_5_0_217_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_219_Update/ack
      -- 
    ack_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_216_delayed_5_0_217_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	17 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	33 
    -- CP-element group 34: 	46 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/crr
      -- 
    crr_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(34), ack => call_stmt_226_call_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 31,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(21) & NicRegisterAccessDaemon_CP_116_elements(25) & NicRegisterAccessDaemon_CP_116_elements(29) & NicRegisterAccessDaemon_CP_116_elements(33) & NicRegisterAccessDaemon_CP_116_elements(46) & NicRegisterAccessDaemon_CP_116_elements(36);
      gj_NicRegisterAccessDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_update_start_
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/ccr
      -- 
    ccr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(35), ack => call_stmt_226_call_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(37);
      gj_NicRegisterAccessDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	19 
    -- CP-element group 36: 	23 
    -- CP-element group 36: 	27 
    -- CP-element group 36: 	31 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	15 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Sample/cra
      -- 
    cra_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_226_call_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	47 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/call_stmt_226_Update/cca
      -- CP-element group 37: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/ring_reenable_memory_space_0
      -- 
    cca_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_226_call_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/req
      -- 
    req_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(38), ack => W_rwbar_220_delayed_5_0_227_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(40);
      gj_NicRegisterAccessDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	43 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_update_start_
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/req
      -- 
    req_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(39), ack => W_rwbar_220_delayed_5_0_227_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: 	11 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Sample/ack
      -- 
    ack_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_220_delayed_5_0_227_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/assign_stmt_229_Update/ack
      -- 
    ack_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_220_delayed_5_0_227_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	17 
    -- CP-element group 42: 	41 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/req
      -- 
    req_310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(42), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(41) & NicRegisterAccessDaemon_CP_116_elements(44);
      gj_NicRegisterAccessDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	39 
    -- CP-element group 43: 	15 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_update_start_
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/req
      -- 
    ack_311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(43)); -- 
    req_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(43), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_Update/ack
      -- 
    ack_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(44)); -- 
    -- CP-element group 45:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	9 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	5 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/condition_evaluated
      -- CP-element group 45: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(45), ack => do_while_stmt_179_branch_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(9), ack => NicRegisterAccessDaemon_CP_116_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	16 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	34 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/array_obj_ref_203_call_stmt_226_delay
      -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(16), ack => NicRegisterAccessDaemon_CP_116_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	37 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	6 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_178/do_while_stmt_179/do_while_stmt_179_loop_body/$exit
      -- 
    NicRegisterAccessDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(37) & NicRegisterAccessDaemon_CP_116_elements(44);
      gj_NicRegisterAccessDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	5 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/$exit
      -- CP-element group 48: 	 branch_block_stmt_178/do_while_stmt_179/loop_exit/ack
      -- 
    ack_323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_179_branch_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	5 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/$exit
      -- CP-element group 49: 	 branch_block_stmt_178/do_while_stmt_179/loop_taken/ack
      -- 
    ack_327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_179_branch_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(49)); -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	3 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	1 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_178/do_while_stmt_179/$exit
      -- 
    NicRegisterAccessDaemon_CP_116_elements(50) <= NicRegisterAccessDaemon_CP_116_elements(3);
    NicRegisterAccessDaemon_do_while_stmt_179_terminator_328: loop_terminator -- 
      generic map (name => " NicRegisterAccessDaemon_do_while_stmt_179_terminator_328", max_iterations_in_flight =>31) 
      port map(loop_body_exit => NicRegisterAccessDaemon_CP_116_elements(6),loop_continue => NicRegisterAccessDaemon_CP_116_elements(49),loop_terminate => NicRegisterAccessDaemon_CP_116_elements(48),loop_back => NicRegisterAccessDaemon_CP_116_elements(4),loop_exit => NicRegisterAccessDaemon_CP_116_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_141_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= NicRegisterAccessDaemon_CP_116_elements(7);
        preds(1)  <= NicRegisterAccessDaemon_CP_116_elements(8);
        entry_tmerge_141 : transition_merge -- 
          generic map(name => " entry_tmerge_141")
          port map (preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_index_202_resized : std_logic_vector(5 downto 0);
    signal R_index_202_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_203_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_203_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_192 : std_logic_vector(3 downto 0);
    signal bmask_213_delayed_5_0_213 : std_logic_vector(3 downto 0);
    signal index_196 : std_logic_vector(5 downto 0);
    signal index_216_delayed_5_0_219 : std_logic_vector(5 downto 0);
    signal konst_247_wire_constant : std_logic_vector(0 downto 0);
    signal rdata_236 : std_logic_vector(31 downto 0);
    signal req_183 : std_logic_vector(42 downto 0);
    signal resp_242 : std_logic_vector(32 downto 0);
    signal rval_204 : std_logic_vector(31 downto 0);
    signal rwbar_188 : std_logic_vector(0 downto 0);
    signal rwbar_212_delayed_5_0_210 : std_logic_vector(0 downto 0);
    signal rwbar_220_delayed_5_0_229 : std_logic_vector(0 downto 0);
    signal type_cast_234_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_200 : std_logic_vector(31 downto 0);
    signal wdata_215_delayed_5_0_216 : std_logic_vector(31 downto 0);
    signal wval_226 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_203_offset_scale_factor_0 <= "000001";
    array_obj_ref_203_resized_base_address <= "000000";
    array_obj_ref_203_word_offset_0 <= "000000";
    konst_247_wire_constant <= "1";
    type_cast_234_wire_constant <= "00000000000000000000000000000000";
    type_cast_239_wire_constant <= "0";
    -- flow-through select operator MUX_235_inst
    rdata_236 <= rval_204 when (rwbar_220_delayed_5_0_229(0) /=  '0') else type_cast_234_wire_constant;
    -- flow-through slice operator slice_187_inst
    rwbar_188 <= req_183(42 downto 42);
    -- flow-through slice operator slice_191_inst
    bmask_192 <= req_183(41 downto 38);
    -- flow-through slice operator slice_195_inst
    index_196 <= req_183(37 downto 32);
    -- flow-through slice operator slice_199_inst
    wdata_200 <= req_183(31 downto 0);
    W_bmask_213_delayed_5_0_211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_213_delayed_5_0_211_inst_req_0;
      W_bmask_213_delayed_5_0_211_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_213_delayed_5_0_211_inst_req_1;
      W_bmask_213_delayed_5_0_211_inst_ack_1<= rack(0);
      W_bmask_213_delayed_5_0_211_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_213_delayed_5_0_211_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_213_delayed_5_0_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_216_delayed_5_0_217_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_216_delayed_5_0_217_inst_req_0;
      W_index_216_delayed_5_0_217_inst_ack_0<= wack(0);
      rreq(0) <= W_index_216_delayed_5_0_217_inst_req_1;
      W_index_216_delayed_5_0_217_inst_ack_1<= rack(0);
      W_index_216_delayed_5_0_217_inst : InterlockBuffer generic map ( -- 
        name => "W_index_216_delayed_5_0_217_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_216_delayed_5_0_219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_212_delayed_5_0_208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_212_delayed_5_0_208_inst_req_0;
      W_rwbar_212_delayed_5_0_208_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_212_delayed_5_0_208_inst_req_1;
      W_rwbar_212_delayed_5_0_208_inst_ack_1<= rack(0);
      W_rwbar_212_delayed_5_0_208_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_212_delayed_5_0_208_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_212_delayed_5_0_210,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_220_delayed_5_0_227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_220_delayed_5_0_227_inst_req_0;
      W_rwbar_220_delayed_5_0_227_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_220_delayed_5_0_227_inst_req_1;
      W_rwbar_220_delayed_5_0_227_inst_ack_1<= rack(0);
      W_rwbar_220_delayed_5_0_227_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_220_delayed_5_0_227_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_220_delayed_5_0_229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_215_delayed_5_0_214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_215_delayed_5_0_214_inst_req_0;
      W_wdata_215_delayed_5_0_214_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_215_delayed_5_0_214_inst_req_1;
      W_wdata_215_delayed_5_0_214_inst_ack_1<= rack(0);
      W_wdata_215_delayed_5_0_214_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_215_delayed_5_0_214_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_215_delayed_5_0_216,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_203_addr_0
    process(array_obj_ref_203_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_203_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_gather_scatter
    process(array_obj_ref_203_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_data_0;
      ov(31 downto 0) := iv;
      rval_204 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_0_rename
    process(R_index_202_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_202_resized;
      ov(5 downto 0) := iv;
      R_index_202_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_0_resize
    process(index_196) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_196;
      ov(5 downto 0) := iv;
      R_index_202_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_offset
    process(R_index_202_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_202_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_203_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_root_address_inst
    process(array_obj_ref_203_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_203_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_179_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_247_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_179_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_179_branch_req_0,
          ack0 => do_while_stmt_179_branch_ack_0,
          ack1 => do_while_stmt_179_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u1_u33_241_inst
    process(type_cast_239_wire_constant, rdata_236) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_239_wire_constant, rdata_236, tmp_var);
      resp_242 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_203_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_203_load_0_req_0;
      array_obj_ref_203_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_203_load_0_req_1;
      array_obj_ref_203_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_203_word_address_0;
      array_obj_ref_203_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(42 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_0;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_req_1;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_182_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_183 <= data_out(42 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0", data_width => 43,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_0;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_req_1;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_243_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_242;
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_226_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_226_call_req_0;
      call_stmt_226_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_226_call_req_1;
      call_stmt_226_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_212_delayed_5_0_210(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_213_delayed_5_0_213 & rval_204 & wdata_215_delayed_5_0_216 & index_216_delayed_5_0_219;
      wval_226 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end NicRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ReceiveEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    FREE_Q : in std_logic_vector(35 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_call_data : out  std_logic_vector(35 downto 0);
    loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
    loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_return_data : in   std_logic_vector(0 downto 0);
    loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
    populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
    populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ReceiveEngineDaemon;
architecture ReceiveEngineDaemon_arch of ReceiveEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ReceiveEngineDaemon_CP_1621_start: Boolean;
  signal ReceiveEngineDaemon_CP_1621_symbol: Boolean;
  -- volatile/operator module components. 
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_ack_1 : boolean;
  signal if_stmt_960_branch_req_0 : boolean;
  signal if_stmt_960_branch_ack_1 : boolean;
  signal if_stmt_960_branch_ack_0 : boolean;
  signal do_while_stmt_968_branch_req_0 : boolean;
  signal call_stmt_976_call_req_0 : boolean;
  signal call_stmt_976_call_ack_0 : boolean;
  signal call_stmt_976_call_req_1 : boolean;
  signal call_stmt_976_call_ack_1 : boolean;
  signal call_stmt_994_call_req_0 : boolean;
  signal call_stmt_994_call_ack_0 : boolean;
  signal call_stmt_994_call_req_1 : boolean;
  signal call_stmt_994_call_ack_1 : boolean;
  signal NOT_u1_u1_997_inst_req_0 : boolean;
  signal NOT_u1_u1_997_inst_ack_0 : boolean;
  signal NOT_u1_u1_997_inst_req_1 : boolean;
  signal NOT_u1_u1_997_inst_ack_1 : boolean;
  signal NOT_u1_u1_1007_inst_req_0 : boolean;
  signal NOT_u1_u1_1007_inst_ack_0 : boolean;
  signal NOT_u1_u1_1007_inst_req_1 : boolean;
  signal NOT_u1_u1_1007_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_ack_1 : boolean;
  signal call_stmt_1028_call_req_0 : boolean;
  signal call_stmt_1028_call_ack_0 : boolean;
  signal call_stmt_1028_call_req_1 : boolean;
  signal call_stmt_1028_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_ack_1 : boolean;
  signal call_stmt_1041_call_req_0 : boolean;
  signal call_stmt_1041_call_ack_0 : boolean;
  signal call_stmt_1041_call_req_1 : boolean;
  signal call_stmt_1041_call_ack_1 : boolean;
  signal do_while_stmt_968_branch_ack_0 : boolean;
  signal do_while_stmt_968_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ReceiveEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ReceiveEngineDaemon_CP_1621_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ReceiveEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1621_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1621_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1621_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ReceiveEngineDaemon_CP_1621: Block -- control-path 
    signal ReceiveEngineDaemon_CP_1621_elements: BooleanArray(51 downto 0);
    -- 
  begin -- 
    ReceiveEngineDaemon_CP_1621_elements(0) <= ReceiveEngineDaemon_CP_1621_start;
    ReceiveEngineDaemon_CP_1621_symbol <= ReceiveEngineDaemon_CP_1621_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_956/$entry
      -- CP-element group 0: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_sample_start_
      -- CP-element group 0: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Sample/req
      -- 
    req_1634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(0), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_sample_completed_
      -- CP-element group 1: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_update_start_
      -- CP-element group 1: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Sample/ack
      -- CP-element group 1: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Update/$entry
      -- CP-element group 1: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Update/req
      -- 
    ack_1635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(1)); -- 
    req_1639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(1), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	51 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_956/$exit
      -- CP-element group 2: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_update_completed_
      -- CP-element group 2: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Update/$exit
      -- CP-element group 2: 	 assign_stmt_956/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_957/$entry
      -- CP-element group 2: 	 branch_block_stmt_957/branch_block_stmt_957__entry__
      -- CP-element group 2: 	 branch_block_stmt_957/merge_stmt_959__entry__
      -- CP-element group 2: 	 branch_block_stmt_957/merge_stmt_959_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_957/merge_stmt_959__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_957/merge_stmt_959__entry___PhiReq/$exit
      -- 
    ack_1640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_957/$exit
      -- CP-element group 3: 	 branch_block_stmt_957/branch_block_stmt_957__exit__
      -- 
    ReceiveEngineDaemon_CP_1621_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	50 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	51 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_957/do_while_stmt_968__exit__
      -- CP-element group 4: 	 branch_block_stmt_957/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_957/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_957/disable_loopback_PhiReq/$exit
      -- 
    ReceiveEngineDaemon_CP_1621_elements(4) <= ReceiveEngineDaemon_CP_1621_elements(50);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	51 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	51 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_957/if_stmt_960_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_957/if_stmt_960_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_957/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_957/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_957/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_960_branch_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	51 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_957/if_stmt_960__exit__
      -- CP-element group 6: 	 branch_block_stmt_957/do_while_stmt_968__entry__
      -- CP-element group 6: 	 branch_block_stmt_957/if_stmt_960_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_957/if_stmt_960_else_link/else_choice_transition
      -- 
    else_choice_transition_1717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_960_branch_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_957/do_while_stmt_968/$entry
      -- CP-element group 7: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968__entry__
      -- 
    ReceiveEngineDaemon_CP_1621_elements(7) <= ReceiveEngineDaemon_CP_1621_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	50 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968__exit__
      -- 
    -- Element group ReceiveEngineDaemon_CP_1621_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_957/do_while_stmt_968/loop_back
      -- 
    -- Element group ReceiveEngineDaemon_CP_1621_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	47 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	48 
    -- CP-element group 10: 	49 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_957/do_while_stmt_968/condition_done
      -- CP-element group 10: 	 branch_block_stmt_957/do_while_stmt_968/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_957/do_while_stmt_968/loop_taken/$entry
      -- 
    ReceiveEngineDaemon_CP_1621_elements(10) <= ReceiveEngineDaemon_CP_1621_elements(47);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	46 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_957/do_while_stmt_968/loop_body_done
      -- 
    ReceiveEngineDaemon_CP_1621_elements(11) <= ReceiveEngineDaemon_CP_1621_elements(46);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/back_edge_to_loop_body
      -- 
    ReceiveEngineDaemon_CP_1621_elements(12) <= ReceiveEngineDaemon_CP_1621_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/first_time_through_loop_body
      -- 
    ReceiveEngineDaemon_CP_1621_elements(13) <= ReceiveEngineDaemon_CP_1621_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	47 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/loop_body_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_1621_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	46 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Sample/crr
      -- 
    crr_1742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(15), ack => call_stmt_976_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(14) & ReceiveEngineDaemon_CP_1621_elements(17) & ReceiveEngineDaemon_CP_1621_elements(46);
      gj_ReceiveEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	25 
    -- CP-element group 16: 	29 
    -- CP-element group 16: 	33 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	46 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_update_start_
      -- CP-element group 16: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Update/ccr
      -- 
    ccr_1747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(16), ack => call_stmt_976_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(21) & ReceiveEngineDaemon_CP_1621_elements(25) & ReceiveEngineDaemon_CP_1621_elements(29) & ReceiveEngineDaemon_CP_1621_elements(33) & ReceiveEngineDaemon_CP_1621_elements(41) & ReceiveEngineDaemon_CP_1621_elements(46);
      gj_ReceiveEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Sample/cra
      -- 
    cra_1743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_976_call_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	23 
    -- CP-element group 18: 	27 
    -- CP-element group 18: 	31 
    -- CP-element group 18: 	39 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_976_Update/cca
      -- 
    cca_1748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_976_call_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Sample/crr
      -- 
    crr_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(19), ack => call_stmt_994_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(18) & ReceiveEngineDaemon_CP_1621_elements(21);
      gj_ReceiveEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	37 
    -- CP-element group 20: 	45 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_update_start_
      -- CP-element group 20: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Update/ccr
      -- 
    ccr_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(20), ack => call_stmt_994_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(37) & ReceiveEngineDaemon_CP_1621_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Sample/cra
      -- 
    cra_1757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_994_call_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(21)); -- 
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	35 
    -- CP-element group 22: 	43 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_994_Update/cca
      -- 
    cca_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_994_call_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	18 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Sample/rr
      -- 
    rr_1770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(23), ack => NOT_u1_u1_997_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(18) & ReceiveEngineDaemon_CP_1621_elements(25);
      gj_ReceiveEngineDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	37 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_update_start_
      -- CP-element group 24: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Update/cr
      -- 
    cr_1775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(24), ack => NOT_u1_u1_997_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1621_elements(37);
      gj_ReceiveEngineDaemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	16 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Sample/ra
      -- 
    ra_1771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_997_inst_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	35 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_997_Update/ca
      -- 
    ca_1776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_997_inst_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	18 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Sample/rr
      -- 
    rr_1784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(27), ack => NOT_u1_u1_1007_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(18) & ReceiveEngineDaemon_CP_1621_elements(29);
      gj_ReceiveEngineDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	45 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_update_start_
      -- CP-element group 28: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Update/cr
      -- 
    cr_1789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(28), ack => NOT_u1_u1_1007_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1621_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Sample/ra
      -- 
    ra_1785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1007_inst_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	43 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/NOT_u1_u1_1007_Update/ca
      -- 
    ca_1790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1007_inst_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	18 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Sample/req
      -- 
    req_1798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(31), ack => W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(18) & ReceiveEngineDaemon_CP_1621_elements(33);
      gj_ReceiveEngineDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	37 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_update_start_
      -- CP-element group 32: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Update/req
      -- 
    req_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(32), ack => W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1621_elements(37);
      gj_ReceiveEngineDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Sample/ack
      -- 
    ack_1799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1025_Update/ack
      -- 
    ack_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	22 
    -- CP-element group 35: 	26 
    -- CP-element group 35: 	34 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	37 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Sample/crr
      -- 
    crr_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(35), ack => call_stmt_1028_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(22) & ReceiveEngineDaemon_CP_1621_elements(26) & ReceiveEngineDaemon_CP_1621_elements(34) & ReceiveEngineDaemon_CP_1621_elements(37);
      gj_ReceiveEngineDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_update_start_
      -- CP-element group 36: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Update/ccr
      -- 
    ccr_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(36), ack => call_stmt_1028_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1621_elements(38);
      gj_ReceiveEngineDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: marked-successors 
    -- CP-element group 37: 	20 
    -- CP-element group 37: 	24 
    -- CP-element group 37: 	32 
    -- CP-element group 37: 	35 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Sample/cra
      -- 
    cra_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1028_call_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1028_Update/cca
      -- 
    cca_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1028_call_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	18 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Sample/req
      -- 
    req_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(39), ack => W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(18) & ReceiveEngineDaemon_CP_1621_elements(41);
      gj_ReceiveEngineDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	45 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_update_start_
      -- CP-element group 40: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Update/req
      -- 
    req_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(40), ack => W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1621_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Sample/ack
      -- 
    ack_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/assign_stmt_1033_Update/ack
      -- 
    ack_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(42)); -- 
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	22 
    -- CP-element group 43: 	30 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	42 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	45 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Sample/crr
      -- 
    crr_1840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(43), ack => call_stmt_1041_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1621_elements(22) & ReceiveEngineDaemon_CP_1621_elements(30) & ReceiveEngineDaemon_CP_1621_elements(38) & ReceiveEngineDaemon_CP_1621_elements(42) & ReceiveEngineDaemon_CP_1621_elements(45);
      gj_ReceiveEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_update_start_
      -- CP-element group 44: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Update/ccr
      -- 
    ccr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(44), ack => call_stmt_1041_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1621_elements(46);
      gj_ReceiveEngineDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	20 
    -- CP-element group 45: 	28 
    -- CP-element group 45: 	40 
    -- CP-element group 45: 	43 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Sample/cra
      -- 
    cra_1841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1041_call_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(45)); -- 
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	11 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	15 
    -- CP-element group 46: 	16 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/$exit
      -- CP-element group 46: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/call_stmt_1041_Update/cca
      -- 
    cca_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1041_call_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(46)); -- 
    -- CP-element group 47:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	14 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	10 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/condition_evaluated
      -- CP-element group 47: 	 branch_block_stmt_957/do_while_stmt_968/do_while_stmt_968_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(47), ack => do_while_stmt_968_branch_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_1621_elements(47) is a control-delay.
    cp_element_47_delay: control_delay_element  generic map(name => " 47_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_1621_elements(14), ack => ReceiveEngineDaemon_CP_1621_elements(47), clk => clk, reset =>reset);
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	10 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_957/do_while_stmt_968/loop_exit/$exit
      -- CP-element group 48: 	 branch_block_stmt_957/do_while_stmt_968/loop_exit/ack
      -- 
    ack_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_968_branch_ack_0, ack => ReceiveEngineDaemon_CP_1621_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	10 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_957/do_while_stmt_968/loop_taken/$exit
      -- CP-element group 49: 	 branch_block_stmt_957/do_while_stmt_968/loop_taken/ack
      -- 
    ack_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_968_branch_ack_1, ack => ReceiveEngineDaemon_CP_1621_elements(49)); -- 
    -- CP-element group 50:  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	8 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	4 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_957/do_while_stmt_968/$exit
      -- 
    ReceiveEngineDaemon_CP_1621_elements(50) <= ReceiveEngineDaemon_CP_1621_elements(8);
    -- CP-element group 51:  merge  branch  transition  place  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	2 
    -- CP-element group 51: 	4 
    -- CP-element group 51: 	5 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	5 
    -- CP-element group 51: 	6 
    -- CP-element group 51:  members (49) 
      -- CP-element group 51: 	 branch_block_stmt_957/merge_stmt_959__exit__
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960__entry__
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_dead_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Sample/req
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Update/req
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/BITSEL_u32_u1_963_inputs/RPIPE_CONTROL_REGISTER_961/Update/ack
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Update/cr
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/BITSEL_u32_u1_963/SplitProtocol/Update/ca
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Update/cr
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/NOT_u1_u1_964/SplitProtocol/Update/ca
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_eval_test/branch_req
      -- CP-element group 51: 	 branch_block_stmt_957/NOT_u1_u1_964_place
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_if_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/if_stmt_960_else_link/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/merge_stmt_959_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_957/merge_stmt_959_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_957/merge_stmt_959_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_957/merge_stmt_959_PhiAck/dummy
      -- 
    branch_req_1708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1621_elements(51), ack => if_stmt_960_branch_req_0); -- 
    ReceiveEngineDaemon_CP_1621_elements(51) <= OrReduce(ReceiveEngineDaemon_CP_1621_elements(2) & ReceiveEngineDaemon_CP_1621_elements(4) & ReceiveEngineDaemon_CP_1621_elements(5));
    ReceiveEngineDaemon_do_while_stmt_968_terminator_1856: loop_terminator -- 
      generic map (name => " ReceiveEngineDaemon_do_while_stmt_968_terminator_1856", max_iterations_in_flight =>31) 
      port map(loop_body_exit => ReceiveEngineDaemon_CP_1621_elements(11),loop_continue => ReceiveEngineDaemon_CP_1621_elements(49),loop_terminate => ReceiveEngineDaemon_CP_1621_elements(48),loop_back => ReceiveEngineDaemon_CP_1621_elements(9),loop_exit => ReceiveEngineDaemon_CP_1621_elements(8),clk => clk, reset => reset); -- 
    entry_tmerge_1734_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ReceiveEngineDaemon_CP_1621_elements(12);
        preds(1)  <= ReceiveEngineDaemon_CP_1621_elements(13);
        entry_tmerge_1734 : transition_merge -- 
          generic map(name => " entry_tmerge_1734")
          port map (preds => preds, symbol_out => ReceiveEngineDaemon_CP_1621_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1046_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_963_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1002_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_964_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_984_984_delayed_10_0_998 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_991_991_delayed_10_0_1008 : std_logic_vector(0 downto 0);
    signal RPIPE_CONTROL_REGISTER_1044_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_961_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1037_wire : std_logic_vector(35 downto 0);
    signal RPIPE_FREE_Q_973_wire : std_logic_vector(35 downto 0);
    signal bad_packet_identifier_994 : std_logic_vector(0 downto 0);
    signal cond_1018 : std_logic_vector(0 downto 0);
    signal free_flag_1013 : std_logic_vector(0 downto 0);
    signal konst_1016_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1045_wire_constant : std_logic_vector(31 downto 0);
    signal konst_955_wire_constant : std_logic_vector(5 downto 0);
    signal konst_962_wire_constant : std_logic_vector(31 downto 0);
    signal ok_flag_1004 : std_logic_vector(0 downto 0);
    signal push_status_1041 : std_logic_vector(0 downto 0);
    signal rx_buffer_pointer_32_976 : std_logic_vector(31 downto 0);
    signal rx_buffer_pointer_36_1005_delayed_10_0_1025 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1013_delayed_10_0_1033 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_984 : std_logic_vector(35 downto 0);
    signal slice_1039_wire : std_logic_vector(31 downto 0);
    signal status_976 : std_logic_vector(0 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_972_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_982_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    konst_1016_wire_constant <= "1";
    konst_1045_wire_constant <= "00000000000000000000000000000000";
    konst_955_wire_constant <= "000000";
    konst_962_wire_constant <= "00000000000000000000000000000000";
    type_cast_1036_wire_constant <= "1";
    type_cast_972_wire_constant <= "1";
    type_cast_982_wire_constant <= "0000";
    -- flow-through slice operator slice_1039_inst
    slice_1039_wire <= rx_buffer_pointer_36_1013_delayed_10_0_1033(35 downto 4);
    W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_req_0;
      W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_req_1;
      W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1005_delayed_10_0_1023_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1005_delayed_10_0_1025,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_req_0;
      W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_req_1;
      W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1013_delayed_10_0_1031_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1013_delayed_10_0_1033,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_968_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1046_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_968_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_968_branch_req_0,
          ack0 => do_while_stmt_968_branch_ack_0,
          ack1 => do_while_stmt_968_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_960_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_964_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_960_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_960_branch_req_0,
          ack0 => if_stmt_960_branch_ack_0,
          ack1 => if_stmt_960_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1003_inst
    process(NOT_u1_u1_984_984_delayed_10_0_998, NOT_u1_u1_1002_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_984_984_delayed_10_0_998, NOT_u1_u1_1002_wire, tmp_var);
      ok_flag_1004 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1012_inst
    process(NOT_u1_u1_991_991_delayed_10_0_1008, bad_packet_identifier_994) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_991_991_delayed_10_0_1008, bad_packet_identifier_994, tmp_var);
      free_flag_1013 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1046_inst
    process(RPIPE_CONTROL_REGISTER_1044_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1044_wire, konst_1045_wire_constant, tmp_var);
      BITSEL_u32_u1_1046_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_963_inst
    process(RPIPE_CONTROL_REGISTER_961_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_961_wire, konst_962_wire_constant, tmp_var);
      BITSEL_u32_u1_963_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u36_983_inst
    process(rx_buffer_pointer_32_976) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(rx_buffer_pointer_32_976, type_cast_982_wire_constant, tmp_var);
      rx_buffer_pointer_36_984 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1017_inst
    process(ok_flag_1004) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ok_flag_1004, konst_1016_wire_constant, tmp_var);
      cond_1018 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1002_inst
    process(bad_packet_identifier_994) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", bad_packet_identifier_994, tmp_var);
      NOT_u1_u1_1002_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (7) : NOT_u1_u1_1007_inst 
    ApIntNot_group_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_976;
      NOT_u1_u1_991_991_delayed_10_0_1008 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1007_inst_req_0;
      NOT_u1_u1_1007_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1007_inst_req_1;
      NOT_u1_u1_1007_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_7_gI: SplitGuardInterface generic map(name => "ApIntNot_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- unary operator NOT_u1_u1_964_inst
    process(BITSEL_u32_u1_963_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_963_wire, tmp_var);
      NOT_u1_u1_964_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (9) : NOT_u1_u1_997_inst 
    ApIntNot_group_9: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_976;
      NOT_u1_u1_984_984_delayed_10_0_998 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_997_inst_req_0;
      NOT_u1_u1_997_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_997_inst_req_1;
      NOT_u1_u1_997_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_9_gI: SplitGuardInterface generic map(name => "ApIntNot_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1044_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_961_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1037_wire <= FREE_Q;
    RPIPE_FREE_Q_973_wire <= FREE_Q;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_954_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_955_wire_constant;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1028_call 
    populateRxQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1028_call_req_0;
      call_stmt_1028_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1028_call_req_1;
      call_stmt_1028_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1004(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      populateRxQueue_call_group_0_gI: SplitGuardInterface generic map(name => "populateRxQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1005_delayed_10_0_1025;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => populateRxQueue_call_reqs(0),
          ackR => populateRxQueue_call_acks(0),
          dataR => populateRxQueue_call_data(35 downto 0),
          tagR => populateRxQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => populateRxQueue_return_acks(0), -- cross-over
          ackL => populateRxQueue_return_reqs(0), -- cross-over
          tagL => populateRxQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1041_call 
    pushIntoQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1041_call_req_0;
      call_stmt_1041_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1041_call_req_1;
      call_stmt_1041_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= free_flag_1013(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_1_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1036_wire_constant & RPIPE_FREE_Q_1037_wire & slice_1039_wire;
      push_status_1041 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_976_call 
    popFromQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_976_call_req_0;
      call_stmt_976_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_976_call_req_1;
      call_stmt_976_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_2_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_972_wire_constant & RPIPE_FREE_Q_973_wire;
      rx_buffer_pointer_32_976 <= data_out(32 downto 1);
      status_976 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_994_call 
    loadBuffer_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_994_call_req_0;
      call_stmt_994_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_994_call_req_1;
      call_stmt_994_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not status_976(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadBuffer_call_group_3_gI: SplitGuardInterface generic map(name => "loadBuffer_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_984;
      bad_packet_identifier_994 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadBuffer_call_reqs(0),
          ackR => loadBuffer_call_acks(0),
          dataR => loadBuffer_call_data(35 downto 0),
          tagR => loadBuffer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => loadBuffer_return_acks(0), -- cross-over
          ackL => loadBuffer_return_reqs(0), -- cross-over
          dataL => loadBuffer_return_data(0 downto 0),
          tagL => loadBuffer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end ReceiveEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity SoftwareRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
    FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
    AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
    CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity SoftwareRegisterAccessDaemon;
architecture SoftwareRegisterAccessDaemon_arch of SoftwareRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal SoftwareRegisterAccessDaemon_CP_1875_start: Boolean;
  signal SoftwareRegisterAccessDaemon_CP_1875_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal phi_stmt_1055_req_1 : boolean;
  signal do_while_stmt_1053_branch_req_0 : boolean;
  signal phi_stmt_1061_req_1 : boolean;
  signal phi_stmt_1066_req_0 : boolean;
  signal phi_stmt_1055_req_0 : boolean;
  signal phi_stmt_1055_ack_0 : boolean;
  signal phi_stmt_1071_req_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1109_inst_ack_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1109_inst_req_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1109_inst_ack_0 : boolean;
  signal check_num_server_1185_1075_buf_ack_1 : boolean;
  signal check_num_server_1185_1075_buf_req_1 : boolean;
  signal phi_stmt_1071_req_1 : boolean;
  signal phi_stmt_1066_req_1 : boolean;
  signal check_num_server_1185_1075_buf_ack_0 : boolean;
  signal phi_stmt_1061_ack_0 : boolean;
  signal array_obj_ref_1111_load_0_ack_0 : boolean;
  signal check_free_q_1176_1070_buf_ack_0 : boolean;
  signal phi_stmt_1071_ack_0 : boolean;
  signal array_obj_ref_1111_load_0_req_0 : boolean;
  signal array_obj_ref_1080_load_0_req_1 : boolean;
  signal array_obj_ref_1080_load_0_req_0 : boolean;
  signal check_free_q_1176_1070_buf_req_0 : boolean;
  signal check_num_server_1185_1075_buf_req_0 : boolean;
  signal check_control_regsiter_1167_1065_buf_ack_1 : boolean;
  signal check_control_regsiter_1167_1065_buf_req_1 : boolean;
  signal phi_stmt_1066_ack_0 : boolean;
  signal check_free_q_1176_1070_buf_ack_1 : boolean;
  signal array_obj_ref_1111_load_0_ack_1 : boolean;
  signal check_free_q_1176_1070_buf_req_1 : boolean;
  signal check_control_regsiter_1167_1065_buf_ack_0 : boolean;
  signal check_control_regsiter_1167_1065_buf_req_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1109_inst_req_1 : boolean;
  signal array_obj_ref_1111_load_0_req_1 : boolean;
  signal phi_stmt_1061_req_0 : boolean;
  signal array_obj_ref_1080_load_0_ack_1 : boolean;
  signal array_obj_ref_1080_load_0_ack_0 : boolean;
  signal array_obj_ref_1116_load_0_req_0 : boolean;
  signal array_obj_ref_1116_load_0_ack_0 : boolean;
  signal array_obj_ref_1116_load_0_req_1 : boolean;
  signal array_obj_ref_1116_load_0_ack_1 : boolean;
  signal W_update_free_q_pipe_1093_delayed_5_0_1118_inst_req_0 : boolean;
  signal W_update_free_q_pipe_1093_delayed_5_0_1118_inst_ack_0 : boolean;
  signal W_update_free_q_pipe_1093_delayed_5_0_1118_inst_req_1 : boolean;
  signal W_update_free_q_pipe_1093_delayed_5_0_1118_inst_ack_1 : boolean;
  signal type_cast_1127_inst_req_0 : boolean;
  signal type_cast_1127_inst_ack_0 : boolean;
  signal type_cast_1127_inst_req_1 : boolean;
  signal type_cast_1127_inst_ack_1 : boolean;
  signal WPIPE_FREE_Q_1122_inst_req_0 : boolean;
  signal WPIPE_FREE_Q_1122_inst_ack_0 : boolean;
  signal WPIPE_FREE_Q_1122_inst_req_1 : boolean;
  signal WPIPE_FREE_Q_1122_inst_ack_1 : boolean;
  signal array_obj_ref_1132_load_0_req_0 : boolean;
  signal array_obj_ref_1132_load_0_ack_0 : boolean;
  signal array_obj_ref_1132_load_0_req_1 : boolean;
  signal array_obj_ref_1132_load_0_ack_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1130_inst_req_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1130_inst_ack_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1130_inst_req_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1130_inst_ack_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1135_inst_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1135_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1135_inst_req_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1135_inst_ack_1 : boolean;
  signal array_obj_ref_1188_load_0_req_0 : boolean;
  signal array_obj_ref_1188_load_0_ack_0 : boolean;
  signal array_obj_ref_1188_load_0_req_1 : boolean;
  signal array_obj_ref_1188_load_0_ack_1 : boolean;
  signal W_rwbar_1166_delayed_5_0_1190_inst_req_0 : boolean;
  signal W_rwbar_1166_delayed_5_0_1190_inst_ack_0 : boolean;
  signal W_rwbar_1166_delayed_5_0_1190_inst_req_1 : boolean;
  signal W_rwbar_1166_delayed_5_0_1190_inst_ack_1 : boolean;
  signal W_bmask_1167_delayed_5_0_1193_inst_req_0 : boolean;
  signal W_bmask_1167_delayed_5_0_1193_inst_ack_0 : boolean;
  signal W_bmask_1167_delayed_5_0_1193_inst_req_1 : boolean;
  signal W_bmask_1167_delayed_5_0_1193_inst_ack_1 : boolean;
  signal W_wdata_1169_delayed_5_0_1196_inst_req_0 : boolean;
  signal W_wdata_1169_delayed_5_0_1196_inst_ack_0 : boolean;
  signal W_wdata_1169_delayed_5_0_1196_inst_req_1 : boolean;
  signal W_wdata_1169_delayed_5_0_1196_inst_ack_1 : boolean;
  signal W_index_1170_delayed_5_0_1199_inst_req_0 : boolean;
  signal W_index_1170_delayed_5_0_1199_inst_ack_0 : boolean;
  signal W_index_1170_delayed_5_0_1199_inst_req_1 : boolean;
  signal W_index_1170_delayed_5_0_1199_inst_ack_1 : boolean;
  signal call_stmt_1208_call_req_0 : boolean;
  signal call_stmt_1208_call_ack_0 : boolean;
  signal call_stmt_1208_call_req_1 : boolean;
  signal call_stmt_1208_call_ack_1 : boolean;
  signal W_rwbar_1174_delayed_5_0_1209_inst_req_0 : boolean;
  signal W_rwbar_1174_delayed_5_0_1209_inst_ack_0 : boolean;
  signal W_rwbar_1174_delayed_5_0_1209_inst_req_1 : boolean;
  signal W_rwbar_1174_delayed_5_0_1209_inst_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1225_inst_req_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1225_inst_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1225_inst_req_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1225_inst_ack_1 : boolean;
  signal do_while_stmt_1053_branch_ack_0 : boolean;
  signal do_while_stmt_1053_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  SoftwareRegisterAccessDaemon_CP_1875_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1875_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1875_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1875_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  SoftwareRegisterAccessDaemon_CP_1875: Block -- control-path 
    signal SoftwareRegisterAccessDaemon_CP_1875_elements: BooleanArray(166 downto 0);
    -- 
  begin -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(0) <= SoftwareRegisterAccessDaemon_CP_1875_start;
    SoftwareRegisterAccessDaemon_CP_1875_symbol <= SoftwareRegisterAccessDaemon_CP_1875_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1052/do_while_stmt_1053__entry__
      -- CP-element group 0: 	 branch_block_stmt_1052/$entry
      -- CP-element group 0: 	 branch_block_stmt_1052/branch_block_stmt_1052__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	166 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1052/do_while_stmt_1053__exit__
      -- CP-element group 1: 	 branch_block_stmt_1052/$exit
      -- CP-element group 1: 	 branch_block_stmt_1052/branch_block_stmt_1052__exit__
      -- CP-element group 1: 	 $exit
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(166);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053__entry__
      -- CP-element group 2: 	 branch_block_stmt_1052/do_while_stmt_1053/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(2) <= SoftwareRegisterAccessDaemon_CP_1875_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	166 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053__exit__
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_back
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	164 
    -- CP-element group 5: 	165 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1052/do_while_stmt_1053/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_taken/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(5) <= SoftwareRegisterAccessDaemon_CP_1875_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	163 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_body_done
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(6) <= SoftwareRegisterAccessDaemon_CP_1875_elements(163);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/back_edge_to_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(7) <= SoftwareRegisterAccessDaemon_CP_1875_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	78 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/first_time_through_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(8) <= SoftwareRegisterAccessDaemon_CP_1875_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	157 
    -- CP-element group 9: 	100 
    -- CP-element group 9: 	122 
    -- CP-element group 9: 	115 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	89 
    -- CP-element group 9: 	93 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_root_address_calculated
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	157 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/condition_evaluated
      -- 
    condition_evaluated_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(10), ack => do_while_stmt_1053_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(14) & SoftwareRegisterAccessDaemon_CP_1875_elements(157);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(15) & SoftwareRegisterAccessDaemon_CP_1875_elements(32) & SoftwareRegisterAccessDaemon_CP_1875_elements(51) & SoftwareRegisterAccessDaemon_CP_1875_elements(70) & SoftwareRegisterAccessDaemon_CP_1875_elements(14);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	163 
    -- CP-element group 12: 	123 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_sample_completed_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(17) & SoftwareRegisterAccessDaemon_CP_1875_elements(35) & SoftwareRegisterAccessDaemon_CP_1875_elements(54) & SoftwareRegisterAccessDaemon_CP_1875_elements(73);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(16) & SoftwareRegisterAccessDaemon_CP_1875_elements(33) & SoftwareRegisterAccessDaemon_CP_1875_elements(52) & SoftwareRegisterAccessDaemon_CP_1875_elements(71);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/aggregated_phi_update_ack
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(18) & SoftwareRegisterAccessDaemon_CP_1875_elements(37) & SoftwareRegisterAccessDaemon_CP_1875_elements(56) & SoftwareRegisterAccessDaemon_CP_1875_elements(75);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	102 
    -- CP-element group 16: 	98 
    -- CP-element group 16: 	120 
    -- CP-element group 16: 	117 
    -- CP-element group 16: 	106 
    -- CP-element group 16: 	95 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(102) & SoftwareRegisterAccessDaemon_CP_1875_elements(98) & SoftwareRegisterAccessDaemon_CP_1875_elements(120) & SoftwareRegisterAccessDaemon_CP_1875_elements(117) & SoftwareRegisterAccessDaemon_CP_1875_elements(106) & SoftwareRegisterAccessDaemon_CP_1875_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	104 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	97 
    -- CP-element group 18: 	100 
    -- CP-element group 18: 	119 
    -- CP-element group 18: 	115 
    -- CP-element group 18: 	93 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(19) <= SoftwareRegisterAccessDaemon_CP_1875_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_loopback_sample_req_ps
      -- 
    phi_stmt_1055_loopback_sample_req_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1055_loopback_sample_req_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(20), ack => phi_stmt_1055_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(21) <= SoftwareRegisterAccessDaemon_CP_1875_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_entry_sample_req_ps
      -- 
    phi_stmt_1055_entry_sample_req_1917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1055_entry_sample_req_1917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(22), ack => phi_stmt_1055_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1055_phi_mux_ack_ps
      -- 
    phi_stmt_1055_phi_mux_ack_1920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1055_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_sample_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_update_start_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(26) <= SoftwareRegisterAccessDaemon_CP_1875_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1058_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(25), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(30) <= SoftwareRegisterAccessDaemon_CP_1875_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1060_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(29), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: 	125 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(12) & SoftwareRegisterAccessDaemon_CP_1875_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	98 
    -- CP-element group 33: 	95 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(98) & SoftwareRegisterAccessDaemon_CP_1875_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(34) <= SoftwareRegisterAccessDaemon_CP_1875_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(36) <= SoftwareRegisterAccessDaemon_CP_1875_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	97 
    -- CP-element group 37: 	93 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_update_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(38) <= SoftwareRegisterAccessDaemon_CP_1875_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_loopback_sample_req_ps
      -- 
    phi_stmt_1061_loopback_sample_req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1061_loopback_sample_req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(39), ack => phi_stmt_1061_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(40) <= SoftwareRegisterAccessDaemon_CP_1875_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_entry_sample_req_ps
      -- CP-element group 41: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_entry_sample_req
      -- 
    phi_stmt_1061_entry_sample_req_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1061_entry_sample_req_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(41), ack => phi_stmt_1061_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_phi_mux_ack_ps
      -- CP-element group 42: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1061_phi_mux_ack
      -- 
    phi_stmt_1061_phi_mux_ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1061_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_update_start_
      -- CP-element group 44: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(45) <= SoftwareRegisterAccessDaemon_CP_1875_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1064_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(44), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Sample/$entry
      -- 
    req_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(47), ack => check_control_regsiter_1167_1065_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Update/req
      -- CP-element group 48: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Update/$entry
      -- 
    req_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(48), ack => check_control_regsiter_1167_1065_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Sample/$exit
      -- 
    ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1167_1065_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_control_regsiter_1065_Update/$exit
      -- 
    ack_1981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1167_1065_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: 	125 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(12) & SoftwareRegisterAccessDaemon_CP_1875_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	102 
    -- CP-element group 52: 	106 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(102) & SoftwareRegisterAccessDaemon_CP_1875_elements(106);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(53) <= SoftwareRegisterAccessDaemon_CP_1875_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(55) <= SoftwareRegisterAccessDaemon_CP_1875_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	104 
    -- CP-element group 56: 	14 
    -- CP-element group 56: 	100 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(57) <= SoftwareRegisterAccessDaemon_CP_1875_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_loopback_sample_req_ps
      -- CP-element group 58: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_loopback_sample_req
      -- 
    phi_stmt_1066_loopback_sample_req_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1066_loopback_sample_req_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(58), ack => phi_stmt_1066_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(59) <= SoftwareRegisterAccessDaemon_CP_1875_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_entry_sample_req_ps
      -- 
    phi_stmt_1066_entry_sample_req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1066_entry_sample_req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(60), ack => phi_stmt_1066_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_phi_mux_ack_ps
      -- CP-element group 61: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1066_phi_mux_ack
      -- 
    phi_stmt_1066_phi_mux_ack_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1066_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(64) <= SoftwareRegisterAccessDaemon_CP_1875_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1069_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(63), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Sample/req
      -- CP-element group 66: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Sample/$entry
      -- 
    req_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(66), ack => check_free_q_1176_1070_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Update/req
      -- CP-element group 67: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Update/$entry
      -- 
    req_2024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(67), ack => check_free_q_1176_1070_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Sample/$exit
      -- 
    ack_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1176_1070_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Update/ack
      -- CP-element group 69: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_free_q_1070_Update/$exit
      -- 
    ack_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1176_1070_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: 	125 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(12) & SoftwareRegisterAccessDaemon_CP_1875_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	120 
    -- CP-element group 71: 	117 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(120) & SoftwareRegisterAccessDaemon_CP_1875_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(72) <= SoftwareRegisterAccessDaemon_CP_1875_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(74) <= SoftwareRegisterAccessDaemon_CP_1875_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	119 
    -- CP-element group 75: 	115 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(76) <= SoftwareRegisterAccessDaemon_CP_1875_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_loopback_sample_req_ps
      -- CP-element group 77: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_loopback_sample_req
      -- 
    phi_stmt_1071_loopback_sample_req_2036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1071_loopback_sample_req_2036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(77), ack => phi_stmt_1071_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(78) <= SoftwareRegisterAccessDaemon_CP_1875_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_entry_sample_req_ps
      -- CP-element group 79: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_entry_sample_req
      -- 
    phi_stmt_1071_entry_sample_req_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1071_entry_sample_req_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(79), ack => phi_stmt_1071_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_phi_mux_ack_ps
      -- CP-element group 80: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/phi_stmt_1071_phi_mux_ack
      -- 
    phi_stmt_1071_phi_mux_ack_2042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1071_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_sample_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(83) <= SoftwareRegisterAccessDaemon_CP_1875_elements(84);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	83 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1074_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(82), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Sample/$entry
      -- 
    req_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(85), ack => check_num_server_1185_1075_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_update_start_
      -- CP-element group 86: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Update/req
      -- CP-element group 86: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_update_start__ps
      -- 
    req_2068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(86), ack => check_num_server_1185_1075_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Sample/$exit
      -- 
    ack_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1185_1075_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_update_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/R_check_num_server_1075_update_completed_
      -- 
    ack_2069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1185_1075_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	9 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	149 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/word_access_start/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/word_access_start/word_0/rr
      -- CP-element group 89: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/word_access_start/$entry
      -- 
    rr_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(89), ack => array_obj_ref_1080_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(149) & SoftwareRegisterAccessDaemon_CP_1875_elements(91);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_update_start_
      -- CP-element group 90: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/word_access_complete/word_0/cr
      -- CP-element group 90: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/word_access_complete/word_0/$entry
      -- CP-element group 90: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/word_access_complete/$entry
      -- CP-element group 90: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/$entry
      -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(90), ack => array_obj_ref_1080_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(92);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	158 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/word_access_start/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/word_access_start/$exit
      -- CP-element group 91: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Sample/word_access_start/word_0/ra
      -- 
    ra_2088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1080_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(91)); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	163 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/array_obj_ref_1080_Merge/merge_req
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/word_access_complete/word_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/array_obj_ref_1080_Merge/merge_ack
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/word_access_complete/$exit
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/array_obj_ref_1080_Merge/$entry
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/array_obj_ref_1080_Merge/$exit
      -- CP-element group 92: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_Update/word_access_complete/word_0/ca
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1080_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: 	18 
    -- CP-element group 93: 	37 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	149 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/word_access_start/word_0/rr
      -- CP-element group 93: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/word_access_start/word_0/$entry
      -- CP-element group 93: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/word_access_start/$entry
      -- 
    rr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(93), ack => array_obj_ref_1111_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(18) & SoftwareRegisterAccessDaemon_CP_1875_elements(37) & SoftwareRegisterAccessDaemon_CP_1875_elements(149) & SoftwareRegisterAccessDaemon_CP_1875_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	98 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/word_access_complete/word_0/$entry
      -- 
    cr_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(94), ack => array_obj_ref_1111_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(98);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	159 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	16 
    -- CP-element group 95: 	33 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/word_access_start/word_0/ra
      -- CP-element group 95: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Sample/word_access_start/$exit
      -- 
    ra_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1111_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/merge_ack
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/merge_req
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/$exit
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/array_obj_ref_1111_Merge/$entry
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_Update/word_access_complete/word_0/$exit
      -- 
    ca_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1111_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	18 
    -- CP-element group 97: 	37 
    -- CP-element group 97: 	96 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Sample/req
      -- CP-element group 97: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_sample_start_
      -- 
    req_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(97), ack => WPIPE_CONTROL_REGISTER_1109_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(18) & SoftwareRegisterAccessDaemon_CP_1875_elements(37) & SoftwareRegisterAccessDaemon_CP_1875_elements(96) & SoftwareRegisterAccessDaemon_CP_1875_elements(99);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	16 
    -- CP-element group 98: 	33 
    -- CP-element group 98: 	94 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Sample/ack
      -- CP-element group 98: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Update/req
      -- CP-element group 98: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_sample_completed_
      -- 
    ack_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1109_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(98)); -- 
    req_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(98), ack => WPIPE_CONTROL_REGISTER_1109_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	163 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Update/ack
      -- CP-element group 99: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_CONTROL_REGISTER_1109_Update/$exit
      -- 
    ack_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1109_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	9 
    -- CP-element group 100: 	18 
    -- CP-element group 100: 	56 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: 	149 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/word_access_start/$entry
      -- CP-element group 100: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/word_access_start/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/word_access_start/word_0/rr
      -- 
    rr_2169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(100), ack => array_obj_ref_1116_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(18) & SoftwareRegisterAccessDaemon_CP_1875_elements(56) & SoftwareRegisterAccessDaemon_CP_1875_elements(102) & SoftwareRegisterAccessDaemon_CP_1875_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	110 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_update_start_
      -- CP-element group 101: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/word_access_complete/$entry
      -- CP-element group 101: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/word_access_complete/word_0/$entry
      -- CP-element group 101: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/word_access_complete/word_0/cr
      -- 
    cr_2180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(101), ack => array_obj_ref_1116_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	160 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	16 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	52 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/word_access_start/$exit
      -- CP-element group 102: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/word_access_start/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Sample/word_access_start/word_0/ra
      -- 
    ra_2170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1116_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	108 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/word_access_complete/$exit
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/word_access_complete/word_0/$exit
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/word_access_complete/word_0/ca
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/array_obj_ref_1116_Merge/$entry
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/array_obj_ref_1116_Merge/$exit
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/array_obj_ref_1116_Merge/merge_req
      -- CP-element group 103: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_Update/array_obj_ref_1116_Merge/merge_ack
      -- 
    ca_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1116_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	18 
    -- CP-element group 104: 	56 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Sample/req
      -- 
    req_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(104), ack => W_update_free_q_pipe_1093_delayed_5_0_1118_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(18) & SoftwareRegisterAccessDaemon_CP_1875_elements(56) & SoftwareRegisterAccessDaemon_CP_1875_elements(106);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	113 
    -- CP-element group 105: 	110 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_update_start_
      -- CP-element group 105: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Update/req
      -- 
    req_2199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(105), ack => W_update_free_q_pipe_1093_delayed_5_0_1118_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(113) & SoftwareRegisterAccessDaemon_CP_1875_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	16 
    -- CP-element group 106: 	52 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Sample/ack
      -- 
    ack_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1093_delayed_5_0_1118_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1120_Update/ack
      -- 
    ack_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1093_delayed_5_0_1118_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	103 
    -- CP-element group 108: 	107 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Sample/rr
      -- 
    rr_2208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(108), ack => type_cast_1127_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(103) & SoftwareRegisterAccessDaemon_CP_1875_elements(107) & SoftwareRegisterAccessDaemon_CP_1875_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	113 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Update/cr
      -- 
    cr_2213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(109), ack => type_cast_1127_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(113);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	101 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Sample/ra
      -- 
    ra_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1127_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/type_cast_1127_Update/ca
      -- 
    ca_2214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1127_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	111 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Sample/req
      -- 
    req_2222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(112), ack => WPIPE_FREE_Q_1122_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(107) & SoftwareRegisterAccessDaemon_CP_1875_elements(111) & SoftwareRegisterAccessDaemon_CP_1875_elements(114);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	105 
    -- CP-element group 113: 	109 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Sample/ack
      -- CP-element group 113: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Update/req
      -- 
    ack_2223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1122_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(113)); -- 
    req_2227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(113), ack => WPIPE_FREE_Q_1122_inst_req_1); -- 
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	163 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_FREE_Q_1122_Update/ack
      -- 
    ack_2228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1122_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	9 
    -- CP-element group 115: 	18 
    -- CP-element group 115: 	75 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	149 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/word_access_start/$entry
      -- CP-element group 115: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/word_access_start/word_0/$entry
      -- CP-element group 115: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/word_access_start/word_0/rr
      -- 
    rr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(115), ack => array_obj_ref_1132_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(18) & SoftwareRegisterAccessDaemon_CP_1875_elements(75) & SoftwareRegisterAccessDaemon_CP_1875_elements(149) & SoftwareRegisterAccessDaemon_CP_1875_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	120 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/word_access_complete/$entry
      -- CP-element group 116: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/word_access_complete/word_0/$entry
      -- CP-element group 116: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/word_access_complete/word_0/cr
      -- 
    cr_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(116), ack => array_obj_ref_1132_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(120);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	161 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	16 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	71 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/word_access_start/$exit
      -- CP-element group 117: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/word_access_start/word_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Sample/word_access_start/word_0/ra
      -- 
    ra_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (9) 
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/word_access_complete/$exit
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/word_access_complete/word_0/$exit
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/word_access_complete/word_0/ca
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/array_obj_ref_1132_Merge/$entry
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/array_obj_ref_1132_Merge/$exit
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/array_obj_ref_1132_Merge/merge_req
      -- CP-element group 118: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_Update/array_obj_ref_1132_Merge/merge_ack
      -- 
    ca_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1132_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	18 
    -- CP-element group 119: 	118 
    -- CP-element group 119: 	75 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Sample/req
      -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(119), ack => WPIPE_NUMBER_OF_SERVERS_1130_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(18) & SoftwareRegisterAccessDaemon_CP_1875_elements(118) & SoftwareRegisterAccessDaemon_CP_1875_elements(75) & SoftwareRegisterAccessDaemon_CP_1875_elements(121);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	16 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	71 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_update_start_
      -- CP-element group 120: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Update/req
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1130_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(120)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(120), ack => WPIPE_NUMBER_OF_SERVERS_1130_inst_req_1); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	163 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_NUMBER_OF_SERVERS_1130_Update/ack
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1130_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	9 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	125 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Sample/rr
      -- 
    rr_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(122), ack => RPIPE_AFB_NIC_REQUEST_1135_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(9) & SoftwareRegisterAccessDaemon_CP_1875_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	12 
    -- CP-element group 123: 	124 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	144 
    -- CP-element group 123: 	152 
    -- CP-element group 123: 	136 
    -- CP-element group 123: 	140 
    -- CP-element group 123: 	132 
    -- CP-element group 123: 	128 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_update_start_
      -- CP-element group 123: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Update/cr
      -- 
    cr_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(123), ack => RPIPE_AFB_NIC_REQUEST_1135_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(12) & SoftwareRegisterAccessDaemon_CP_1875_elements(124) & SoftwareRegisterAccessDaemon_CP_1875_elements(144) & SoftwareRegisterAccessDaemon_CP_1875_elements(152) & SoftwareRegisterAccessDaemon_CP_1875_elements(136) & SoftwareRegisterAccessDaemon_CP_1875_elements(140) & SoftwareRegisterAccessDaemon_CP_1875_elements(132) & SoftwareRegisterAccessDaemon_CP_1875_elements(128);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Sample/ra
      -- 
    ra_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1135_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	150 
    -- CP-element group 125: 	126 
    -- CP-element group 125: 	138 
    -- CP-element group 125: 	142 
    -- CP-element group 125: 	130 
    -- CP-element group 125: 	134 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	32 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	51 
    -- CP-element group 125: 	70 
    -- CP-element group 125:  members (29) 
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/RPIPE_AFB_NIC_REQUEST_1135_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_word_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_root_address_calculated
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_offset_calculated
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_resized_0
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_scaled_0
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_computed_0
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_resize_0/$entry
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_resize_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_resize_0/index_resize_req
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_resize_0/index_resize_ack
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_scale_0/$entry
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_scale_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_scale_0/scale_rename_req
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_index_scale_0/scale_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_final_index_sum_regn/$entry
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_final_index_sum_regn/$exit
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_final_index_sum_regn/req
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_final_index_sum_regn/ack
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_base_plus_offset/$entry
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_base_plus_offset/$exit
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_base_plus_offset/sum_rename_req
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_base_plus_offset/sum_rename_ack
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_word_addrgen/$entry
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_word_addrgen/$exit
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_word_addrgen/root_register_req
      -- CP-element group 125: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_word_addrgen/root_register_ack
      -- 
    ca_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1135_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	149 
    -- CP-element group 126: 	128 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (5) 
      -- CP-element group 126: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/word_access_start/$entry
      -- CP-element group 126: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/word_access_start/word_0/$entry
      -- CP-element group 126: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/word_access_start/word_0/rr
      -- 
    rr_2336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(126), ack => array_obj_ref_1188_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(125) & SoftwareRegisterAccessDaemon_CP_1875_elements(149) & SoftwareRegisterAccessDaemon_CP_1875_elements(128);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	148 
    -- CP-element group 127: 	155 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (5) 
      -- CP-element group 127: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_update_start_
      -- CP-element group 127: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/word_access_complete/$entry
      -- CP-element group 127: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/word_access_complete/word_0/$entry
      -- CP-element group 127: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/word_access_complete/word_0/cr
      -- 
    cr_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(127), ack => array_obj_ref_1188_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(148) & SoftwareRegisterAccessDaemon_CP_1875_elements(155);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	162 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: 	123 
    -- CP-element group 128:  members (5) 
      -- CP-element group 128: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/word_access_start/$exit
      -- CP-element group 128: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/word_access_start/word_0/$exit
      -- CP-element group 128: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Sample/word_access_start/word_0/ra
      -- 
    ra_2337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1188_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	146 
    -- CP-element group 129: 	154 
    -- CP-element group 129:  members (9) 
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/word_access_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/word_access_complete/word_0/$exit
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/word_access_complete/word_0/ca
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/array_obj_ref_1188_Merge/$entry
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/array_obj_ref_1188_Merge/$exit
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/array_obj_ref_1188_Merge/merge_req
      -- CP-element group 129: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_Update/array_obj_ref_1188_Merge/merge_ack
      -- 
    ca_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1188_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	125 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Sample/req
      -- 
    req_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(130), ack => W_rwbar_1166_delayed_5_0_1190_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(125) & SoftwareRegisterAccessDaemon_CP_1875_elements(132);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	148 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_update_start_
      -- CP-element group 131: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Update/req
      -- 
    req_2366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(131), ack => W_rwbar_1166_delayed_5_0_1190_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: 	123 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Sample/ack
      -- 
    ack_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1166_delayed_5_0_1190_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	146 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1192_Update/ack
      -- 
    ack_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1166_delayed_5_0_1190_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	125 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	136 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Sample/req
      -- 
    req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(134), ack => W_bmask_1167_delayed_5_0_1193_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(125) & SoftwareRegisterAccessDaemon_CP_1875_elements(136);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	148 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_update_start_
      -- CP-element group 135: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Update/req
      -- 
    req_2380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(135), ack => W_bmask_1167_delayed_5_0_1193_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: 	123 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Sample/ack
      -- 
    ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1167_delayed_5_0_1193_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	146 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1195_Update/ack
      -- 
    ack_2381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1167_delayed_5_0_1193_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(137)); -- 
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	125 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Sample/req
      -- 
    req_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(138), ack => W_wdata_1169_delayed_5_0_1196_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(125) & SoftwareRegisterAccessDaemon_CP_1875_elements(140);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	148 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_update_start_
      -- CP-element group 139: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Update/req
      -- 
    req_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(139), ack => W_wdata_1169_delayed_5_0_1196_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: 	123 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Sample/ack
      -- 
    ack_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1169_delayed_5_0_1196_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	146 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1198_Update/ack
      -- 
    ack_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1169_delayed_5_0_1196_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	125 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Sample/req
      -- 
    req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(142), ack => W_index_1170_delayed_5_0_1199_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(125) & SoftwareRegisterAccessDaemon_CP_1875_elements(144);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	148 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_update_start_
      -- CP-element group 143: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Update/req
      -- 
    req_2408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(143), ack => W_index_1170_delayed_5_0_1199_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: 	123 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Sample/ack
      -- 
    ack_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1170_delayed_5_0_1199_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1201_Update/ack
      -- 
    ack_2409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1170_delayed_5_0_1199_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: 	159 
    -- CP-element group 146: 	160 
    -- CP-element group 146: 	161 
    -- CP-element group 146: 	162 
    -- CP-element group 146: 	158 
    -- CP-element group 146: 	137 
    -- CP-element group 146: 	141 
    -- CP-element group 146: 	129 
    -- CP-element group 146: 	133 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Sample/crr
      -- 
    crr_2417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(146), ack => call_stmt_1208_call_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(145) & SoftwareRegisterAccessDaemon_CP_1875_elements(159) & SoftwareRegisterAccessDaemon_CP_1875_elements(160) & SoftwareRegisterAccessDaemon_CP_1875_elements(161) & SoftwareRegisterAccessDaemon_CP_1875_elements(162) & SoftwareRegisterAccessDaemon_CP_1875_elements(158) & SoftwareRegisterAccessDaemon_CP_1875_elements(137) & SoftwareRegisterAccessDaemon_CP_1875_elements(141) & SoftwareRegisterAccessDaemon_CP_1875_elements(129) & SoftwareRegisterAccessDaemon_CP_1875_elements(133) & SoftwareRegisterAccessDaemon_CP_1875_elements(148);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_update_start_
      -- CP-element group 147: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Update/ccr
      -- 
    ccr_2422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(147), ack => call_stmt_1208_call_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	143 
    -- CP-element group 148: 	146 
    -- CP-element group 148: 	127 
    -- CP-element group 148: 	135 
    -- CP-element group 148: 	139 
    -- CP-element group 148: 	131 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Sample/cra
      -- 
    cra_2418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1208_call_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	163 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	126 
    -- CP-element group 149: 	100 
    -- CP-element group 149: 	115 
    -- CP-element group 149: 	89 
    -- CP-element group 149: 	93 
    -- CP-element group 149:  members (4) 
      -- CP-element group 149: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/call_stmt_1208_Update/cca
      -- CP-element group 149: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/ring_reenable_memory_space_0
      -- 
    cca_2423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1208_call_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	125 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Sample/req
      -- 
    req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(150), ack => W_rwbar_1174_delayed_5_0_1209_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(125) & SoftwareRegisterAccessDaemon_CP_1875_elements(152);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	155 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Update/req
      -- 
    req_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(151), ack => W_rwbar_1174_delayed_5_0_1209_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1875_elements(155);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: 	123 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Sample/ack
      -- 
    ack_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1174_delayed_5_0_1209_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/assign_stmt_1211_Update/ack
      -- 
    ack_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1174_delayed_5_0_1209_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: 	129 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Sample/req
      -- 
    req_2445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(154), ack => WPIPE_AFB_NIC_RESPONSE_1225_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(153) & SoftwareRegisterAccessDaemon_CP_1875_elements(129) & SoftwareRegisterAccessDaemon_CP_1875_elements(156);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	127 
    -- CP-element group 155: 	151 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Sample/ack
      -- CP-element group 155: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Update/req
      -- 
    ack_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1225_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(155)); -- 
    req_2450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1875_elements(155), ack => WPIPE_AFB_NIC_RESPONSE_1225_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	163 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/WPIPE_AFB_NIC_RESPONSE_1225_Update/ack
      -- 
    ack_2451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1225_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(156)); -- 
    -- CP-element group 157:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	9 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	10 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(157) is a control-delay.
    cp_element_157_delay: control_delay_element  generic map(name => " 157_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(9), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(157), clk => clk, reset =>reset);
    -- CP-element group 158:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	91 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	146 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1080_call_stmt_1208_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(158) is a control-delay.
    cp_element_158_delay: control_delay_element  generic map(name => " 158_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(91), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(158), clk => clk, reset =>reset);
    -- CP-element group 159:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	95 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	146 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1111_call_stmt_1208_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(159) is a control-delay.
    cp_element_159_delay: control_delay_element  generic map(name => " 159_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(95), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(159), clk => clk, reset =>reset);
    -- CP-element group 160:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	102 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	146 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1116_call_stmt_1208_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(160) is a control-delay.
    cp_element_160_delay: control_delay_element  generic map(name => " 160_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(102), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(160), clk => clk, reset =>reset);
    -- CP-element group 161:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	117 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	146 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1132_call_stmt_1208_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(161) is a control-delay.
    cp_element_161_delay: control_delay_element  generic map(name => " 161_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(117), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(161), clk => clk, reset =>reset);
    -- CP-element group 162:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	128 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	146 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/array_obj_ref_1188_call_stmt_1208_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1875_elements(162) is a control-delay.
    cp_element_162_delay: control_delay_element  generic map(name => " 162_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1875_elements(128), ack => SoftwareRegisterAccessDaemon_CP_1875_elements(162), clk => clk, reset =>reset);
    -- CP-element group 163:  join  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	12 
    -- CP-element group 163: 	149 
    -- CP-element group 163: 	156 
    -- CP-element group 163: 	99 
    -- CP-element group 163: 	121 
    -- CP-element group 163: 	114 
    -- CP-element group 163: 	92 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	6 
    -- CP-element group 163:  members (1) 
      -- CP-element group 163: 	 branch_block_stmt_1052/do_while_stmt_1053/do_while_stmt_1053_loop_body/$exit
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31,6 => 31);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1875_elements(12) & SoftwareRegisterAccessDaemon_CP_1875_elements(149) & SoftwareRegisterAccessDaemon_CP_1875_elements(156) & SoftwareRegisterAccessDaemon_CP_1875_elements(99) & SoftwareRegisterAccessDaemon_CP_1875_elements(121) & SoftwareRegisterAccessDaemon_CP_1875_elements(114) & SoftwareRegisterAccessDaemon_CP_1875_elements(92);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	5 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_exit/$exit
      -- CP-element group 164: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_exit/ack
      -- 
    ack_2462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1053_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	5 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_taken/$exit
      -- CP-element group 165: 	 branch_block_stmt_1052/do_while_stmt_1053/loop_taken/ack
      -- 
    ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1053_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1875_elements(165)); -- 
    -- CP-element group 166:  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	3 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	1 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_1052/do_while_stmt_1053/$exit
      -- 
    SoftwareRegisterAccessDaemon_CP_1875_elements(166) <= SoftwareRegisterAccessDaemon_CP_1875_elements(3);
    SoftwareRegisterAccessDaemon_do_while_stmt_1053_terminator_2467: loop_terminator -- 
      generic map (name => " SoftwareRegisterAccessDaemon_do_while_stmt_1053_terminator_2467", max_iterations_in_flight =>31) 
      port map(loop_body_exit => SoftwareRegisterAccessDaemon_CP_1875_elements(6),loop_continue => SoftwareRegisterAccessDaemon_CP_1875_elements(165),loop_terminate => SoftwareRegisterAccessDaemon_CP_1875_elements(164),loop_back => SoftwareRegisterAccessDaemon_CP_1875_elements(4),loop_exit => SoftwareRegisterAccessDaemon_CP_1875_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1055_phi_seq_1938_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(21);
      SoftwareRegisterAccessDaemon_CP_1875_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(24);
      SoftwareRegisterAccessDaemon_CP_1875_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(26);
      SoftwareRegisterAccessDaemon_CP_1875_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(19);
      SoftwareRegisterAccessDaemon_CP_1875_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(28);
      SoftwareRegisterAccessDaemon_CP_1875_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(30);
      SoftwareRegisterAccessDaemon_CP_1875_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1055_phi_seq_1938 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1055_phi_seq_1938") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1875_elements(11), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(17), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1875_elements(13), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(18), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1061_phi_seq_1982_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(40);
      SoftwareRegisterAccessDaemon_CP_1875_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(43);
      SoftwareRegisterAccessDaemon_CP_1875_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(45);
      SoftwareRegisterAccessDaemon_CP_1875_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(38);
      SoftwareRegisterAccessDaemon_CP_1875_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(49);
      SoftwareRegisterAccessDaemon_CP_1875_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(50);
      SoftwareRegisterAccessDaemon_CP_1875_elements(39) <= phi_mux_reqs(1);
      phi_stmt_1061_phi_seq_1982 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1061_phi_seq_1982") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1875_elements(34), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(35), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1875_elements(36), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(37), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1066_phi_seq_2026_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(59);
      SoftwareRegisterAccessDaemon_CP_1875_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(62);
      SoftwareRegisterAccessDaemon_CP_1875_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(64);
      SoftwareRegisterAccessDaemon_CP_1875_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(57);
      SoftwareRegisterAccessDaemon_CP_1875_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(68);
      SoftwareRegisterAccessDaemon_CP_1875_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(69);
      SoftwareRegisterAccessDaemon_CP_1875_elements(58) <= phi_mux_reqs(1);
      phi_stmt_1066_phi_seq_2026 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1066_phi_seq_2026") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1875_elements(53), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(54), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1875_elements(55), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(56), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1071_phi_seq_2070_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(78);
      SoftwareRegisterAccessDaemon_CP_1875_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(81);
      SoftwareRegisterAccessDaemon_CP_1875_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(83);
      SoftwareRegisterAccessDaemon_CP_1875_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(76);
      SoftwareRegisterAccessDaemon_CP_1875_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(87);
      SoftwareRegisterAccessDaemon_CP_1875_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(88);
      SoftwareRegisterAccessDaemon_CP_1875_elements(77) <= phi_mux_reqs(1);
      phi_stmt_1071_phi_seq_2070 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1071_phi_seq_2070") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1875_elements(72), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(73), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1875_elements(74), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(75), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1875_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1900_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(7);
        preds(1)  <= SoftwareRegisterAccessDaemon_CP_1875_elements(8);
        entry_tmerge_1900 : transition_merge -- 
          generic map(name => " entry_tmerge_1900")
          port map (preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1875_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1089_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1097_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1105_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u32_u35_1126_wire : std_logic_vector(34 downto 0);
    signal EQ_u1_u1_1165_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1174_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1183_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1162_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1171_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1180_wire : std_logic_vector(0 downto 0);
    signal FREE_Q_32_1117 : std_logic_vector(31 downto 0);
    signal INIT_1055 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1086_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1094_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1102_wire : std_logic_vector(0 downto 0);
    signal R_index_1187_resized : std_logic_vector(5 downto 0);
    signal R_index_1187_scaled : std_logic_vector(5 downto 0);
    signal addr_1150 : std_logic_vector(35 downto 0);
    signal array_obj_ref_1080_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1080_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1111_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1111_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1111_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1116_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1116_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1132_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1132_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1132_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1188_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1188_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_1188_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1188_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1188_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1188_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1188_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_1146 : std_logic_vector(3 downto 0);
    signal bmask_1167_delayed_5_0_1195 : std_logic_vector(3 downto 0);
    signal check_control_regsiter_1167 : std_logic_vector(0 downto 0);
    signal check_control_regsiter_1167_1065_buffered : std_logic_vector(0 downto 0);
    signal check_free_q_1176 : std_logic_vector(0 downto 0);
    signal check_free_q_1176_1070_buffered : std_logic_vector(0 downto 0);
    signal check_num_server_1185 : std_logic_vector(0 downto 0);
    signal check_num_server_1185_1075_buffered : std_logic_vector(0 downto 0);
    signal control_data_1081 : std_logic_vector(31 downto 0);
    signal control_register_1061 : std_logic_vector(0 downto 0);
    signal free_q_1066 : std_logic_vector(0 downto 0);
    signal index_1158 : std_logic_vector(5 downto 0);
    signal index_1170_delayed_5_0_1201 : std_logic_vector(5 downto 0);
    signal konst_1161_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1164_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1170_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1173_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1179_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1182_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1229_wire_constant : std_logic_vector(0 downto 0);
    signal num_server_1071 : std_logic_vector(0 downto 0);
    signal rdata_1218 : std_logic_vector(31 downto 0);
    signal req_1136 : std_logic_vector(73 downto 0);
    signal resp_1224 : std_logic_vector(32 downto 0);
    signal rval_1189 : std_logic_vector(31 downto 0);
    signal rwbar_1142 : std_logic_vector(0 downto 0);
    signal rwbar_1166_delayed_5_0_1192 : std_logic_vector(0 downto 0);
    signal rwbar_1174_delayed_5_0_1211 : std_logic_vector(0 downto 0);
    signal type_cast_1058_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1060_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1064_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1069_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1074_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1125_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_1127_wire : std_logic_vector(35 downto 0);
    signal type_cast_1216_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1221_wire_constant : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_1091 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1093_delayed_5_0_1120 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1099 : std_logic_vector(0 downto 0);
    signal update_server_num_1107 : std_logic_vector(0 downto 0);
    signal wdata_1154 : std_logic_vector(31 downto 0);
    signal wdata_1169_delayed_5_0_1198 : std_logic_vector(31 downto 0);
    signal wval_1208 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1080_word_address_0 <= "000000";
    array_obj_ref_1111_word_address_0 <= "000000";
    array_obj_ref_1116_word_address_0 <= "010010";
    array_obj_ref_1132_word_address_0 <= "000001";
    array_obj_ref_1188_offset_scale_factor_0 <= "000001";
    array_obj_ref_1188_resized_base_address <= "000000";
    array_obj_ref_1188_word_offset_0 <= "000000";
    konst_1161_wire_constant <= "000000";
    konst_1164_wire_constant <= "0";
    konst_1170_wire_constant <= "010010";
    konst_1173_wire_constant <= "0";
    konst_1179_wire_constant <= "000001";
    konst_1182_wire_constant <= "0";
    konst_1229_wire_constant <= "1";
    type_cast_1058_wire_constant <= "0";
    type_cast_1060_wire_constant <= "1";
    type_cast_1064_wire_constant <= "0";
    type_cast_1069_wire_constant <= "0";
    type_cast_1074_wire_constant <= "0";
    type_cast_1125_wire_constant <= "000";
    type_cast_1216_wire_constant <= "00000000000000000000000000000000";
    type_cast_1221_wire_constant <= "0";
    phi_stmt_1055: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1058_wire_constant & type_cast_1060_wire_constant;
      req <= phi_stmt_1055_req_0 & phi_stmt_1055_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1055",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1055_ack_0,
          idata => idata,
          odata => INIT_1055,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1055
    phi_stmt_1061: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1064_wire_constant & check_control_regsiter_1167_1065_buffered;
      req <= phi_stmt_1061_req_0 & phi_stmt_1061_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1061",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1061_ack_0,
          idata => idata,
          odata => control_register_1061,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1061
    phi_stmt_1066: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1069_wire_constant & check_free_q_1176_1070_buffered;
      req <= phi_stmt_1066_req_0 & phi_stmt_1066_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1066",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1066_ack_0,
          idata => idata,
          odata => free_q_1066,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1066
    phi_stmt_1071: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1074_wire_constant & check_num_server_1185_1075_buffered;
      req <= phi_stmt_1071_req_0 & phi_stmt_1071_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1071",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1071_ack_0,
          idata => idata,
          odata => num_server_1071,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1071
    -- flow-through select operator MUX_1217_inst
    rdata_1218 <= rval_1189 when (rwbar_1174_delayed_5_0_1211(0) /=  '0') else type_cast_1216_wire_constant;
    -- flow-through slice operator slice_1141_inst
    rwbar_1142 <= req_1136(72 downto 72);
    -- flow-through slice operator slice_1145_inst
    bmask_1146 <= req_1136(71 downto 68);
    -- flow-through slice operator slice_1149_inst
    addr_1150 <= req_1136(67 downto 32);
    -- flow-through slice operator slice_1153_inst
    wdata_1154 <= req_1136(31 downto 0);
    -- flow-through slice operator slice_1157_inst
    index_1158 <= addr_1150(5 downto 0);
    W_bmask_1167_delayed_5_0_1193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_1167_delayed_5_0_1193_inst_req_0;
      W_bmask_1167_delayed_5_0_1193_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_1167_delayed_5_0_1193_inst_req_1;
      W_bmask_1167_delayed_5_0_1193_inst_ack_1<= rack(0);
      W_bmask_1167_delayed_5_0_1193_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_1167_delayed_5_0_1193_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_1146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_1167_delayed_5_0_1195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_1170_delayed_5_0_1199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_1170_delayed_5_0_1199_inst_req_0;
      W_index_1170_delayed_5_0_1199_inst_ack_0<= wack(0);
      rreq(0) <= W_index_1170_delayed_5_0_1199_inst_req_1;
      W_index_1170_delayed_5_0_1199_inst_ack_1<= rack(0);
      W_index_1170_delayed_5_0_1199_inst : InterlockBuffer generic map ( -- 
        name => "W_index_1170_delayed_5_0_1199_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_1158,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_1170_delayed_5_0_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1166_delayed_5_0_1190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1166_delayed_5_0_1190_inst_req_0;
      W_rwbar_1166_delayed_5_0_1190_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1166_delayed_5_0_1190_inst_req_1;
      W_rwbar_1166_delayed_5_0_1190_inst_ack_1<= rack(0);
      W_rwbar_1166_delayed_5_0_1190_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1166_delayed_5_0_1190_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1166_delayed_5_0_1192,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1174_delayed_5_0_1209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1174_delayed_5_0_1209_inst_req_0;
      W_rwbar_1174_delayed_5_0_1209_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1174_delayed_5_0_1209_inst_req_1;
      W_rwbar_1174_delayed_5_0_1209_inst_ack_1<= rack(0);
      W_rwbar_1174_delayed_5_0_1209_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1174_delayed_5_0_1209_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1142,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1174_delayed_5_0_1211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_update_free_q_pipe_1093_delayed_5_0_1118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_update_free_q_pipe_1093_delayed_5_0_1118_inst_req_0;
      W_update_free_q_pipe_1093_delayed_5_0_1118_inst_ack_0<= wack(0);
      rreq(0) <= W_update_free_q_pipe_1093_delayed_5_0_1118_inst_req_1;
      W_update_free_q_pipe_1093_delayed_5_0_1118_inst_ack_1<= rack(0);
      W_update_free_q_pipe_1093_delayed_5_0_1118_inst : InterlockBuffer generic map ( -- 
        name => "W_update_free_q_pipe_1093_delayed_5_0_1118_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => update_free_q_pipe_1099,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => update_free_q_pipe_1093_delayed_5_0_1120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_1169_delayed_5_0_1196_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_1169_delayed_5_0_1196_inst_req_0;
      W_wdata_1169_delayed_5_0_1196_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_1169_delayed_5_0_1196_inst_req_1;
      W_wdata_1169_delayed_5_0_1196_inst_ack_1<= rack(0);
      W_wdata_1169_delayed_5_0_1196_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_1169_delayed_5_0_1196_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_1154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_1169_delayed_5_0_1198,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_control_regsiter_1167_1065_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_control_regsiter_1167_1065_buf_req_0;
      check_control_regsiter_1167_1065_buf_ack_0<= wack(0);
      rreq(0) <= check_control_regsiter_1167_1065_buf_req_1;
      check_control_regsiter_1167_1065_buf_ack_1<= rack(0);
      check_control_regsiter_1167_1065_buf : InterlockBuffer generic map ( -- 
        name => "check_control_regsiter_1167_1065_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_control_regsiter_1167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_control_regsiter_1167_1065_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_free_q_1176_1070_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_free_q_1176_1070_buf_req_0;
      check_free_q_1176_1070_buf_ack_0<= wack(0);
      rreq(0) <= check_free_q_1176_1070_buf_req_1;
      check_free_q_1176_1070_buf_ack_1<= rack(0);
      check_free_q_1176_1070_buf : InterlockBuffer generic map ( -- 
        name => "check_free_q_1176_1070_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_free_q_1176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_free_q_1176_1070_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_num_server_1185_1075_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_num_server_1185_1075_buf_req_0;
      check_num_server_1185_1075_buf_ack_0<= wack(0);
      rreq(0) <= check_num_server_1185_1075_buf_req_1;
      check_num_server_1185_1075_buf_ack_1<= rack(0);
      check_num_server_1185_1075_buf : InterlockBuffer generic map ( -- 
        name => "check_num_server_1185_1075_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_num_server_1185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_num_server_1185_1075_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1127_inst_req_0;
      type_cast_1127_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1127_inst_req_1;
      type_cast_1127_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  update_free_q_pipe_1093_delayed_5_0_1120(0);
      type_cast_1127_inst_gI: SplitGuardInterface generic map(name => "type_cast_1127_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 35,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => CONCAT_u32_u35_1126_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1127_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1080_gather_scatter
    process(array_obj_ref_1080_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1080_data_0;
      ov(31 downto 0) := iv;
      control_data_1081 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1111_gather_scatter
    process(array_obj_ref_1111_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1111_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1111_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1116_gather_scatter
    process(array_obj_ref_1116_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1116_data_0;
      ov(31 downto 0) := iv;
      FREE_Q_32_1117 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1132_gather_scatter
    process(array_obj_ref_1132_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1132_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1132_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_addr_0
    process(array_obj_ref_1188_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1188_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_1188_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_gather_scatter
    process(array_obj_ref_1188_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1188_data_0;
      ov(31 downto 0) := iv;
      rval_1189 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_index_0_rename
    process(R_index_1187_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1187_resized;
      ov(5 downto 0) := iv;
      R_index_1187_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_index_0_resize
    process(index_1158) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_1158;
      ov(5 downto 0) := iv;
      R_index_1187_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_index_offset
    process(R_index_1187_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1187_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_1188_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1188_root_address_inst
    process(array_obj_ref_1188_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1188_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_1188_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_1053_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1229_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1053_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1053_branch_req_0,
          ack0 => do_while_stmt_1053_branch_ack_0,
          ack1 => do_while_stmt_1053_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1089_inst
    process(INIT_1055, control_register_1061) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1055, control_register_1061, tmp_var);
      AND_u1_u1_1089_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1097_inst
    process(INIT_1055, free_q_1066) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1055, free_q_1066, tmp_var);
      AND_u1_u1_1097_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1105_inst
    process(INIT_1055, num_server_1071) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1055, num_server_1071, tmp_var);
      AND_u1_u1_1105_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1166_inst
    process(EQ_u6_u1_1162_wire, EQ_u1_u1_1165_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1162_wire, EQ_u1_u1_1165_wire, tmp_var);
      check_control_regsiter_1167 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1175_inst
    process(EQ_u6_u1_1171_wire, EQ_u1_u1_1174_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1171_wire, EQ_u1_u1_1174_wire, tmp_var);
      check_free_q_1176 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1184_inst
    process(EQ_u6_u1_1180_wire, EQ_u1_u1_1183_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1180_wire, EQ_u1_u1_1183_wire, tmp_var);
      check_num_server_1185 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_1223_inst
    process(type_cast_1221_wire_constant, rdata_1218) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1221_wire_constant, rdata_1218, tmp_var);
      resp_1224 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u35_1126_inst
    process(FREE_Q_32_1117) -- 
      variable tmp_var : std_logic_vector(34 downto 0); -- 
    begin -- 
      ApConcat_proc(FREE_Q_32_1117, type_cast_1125_wire_constant, tmp_var);
      CONCAT_u32_u35_1126_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1165_inst
    process(rwbar_1142) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1142, konst_1164_wire_constant, tmp_var);
      EQ_u1_u1_1165_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1174_inst
    process(rwbar_1142) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1142, konst_1173_wire_constant, tmp_var);
      EQ_u1_u1_1174_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1183_inst
    process(rwbar_1142) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1142, konst_1182_wire_constant, tmp_var);
      EQ_u1_u1_1183_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1162_inst
    process(index_1158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1158, konst_1161_wire_constant, tmp_var);
      EQ_u6_u1_1162_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1171_inst
    process(index_1158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1158, konst_1170_wire_constant, tmp_var);
      EQ_u6_u1_1171_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1180_inst
    process(index_1158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1158, konst_1179_wire_constant, tmp_var);
      EQ_u6_u1_1180_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1086_inst
    process(INIT_1055) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1055, tmp_var);
      NOT_u1_u1_1086_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1094_inst
    process(INIT_1055) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1055, tmp_var);
      NOT_u1_u1_1094_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1102_inst
    process(INIT_1055) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1055, tmp_var);
      NOT_u1_u1_1102_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1090_inst
    process(NOT_u1_u1_1086_wire, AND_u1_u1_1089_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1086_wire, AND_u1_u1_1089_wire, tmp_var);
      update_control_register_pipe_1091 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1098_inst
    process(NOT_u1_u1_1094_wire, AND_u1_u1_1097_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1094_wire, AND_u1_u1_1097_wire, tmp_var);
      update_free_q_pipe_1099 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1106_inst
    process(NOT_u1_u1_1102_wire, AND_u1_u1_1105_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1102_wire, AND_u1_u1_1105_wire, tmp_var);
      update_server_num_1107 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_1132_load_0 array_obj_ref_1188_load_0 array_obj_ref_1116_load_0 array_obj_ref_1111_load_0 array_obj_ref_1080_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => true, 2 => true, 3 => false, 4 => true);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5, 4 => 5);
      -- 
    begin -- 
      reqL_unguarded(4) <= array_obj_ref_1132_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_1188_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1116_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1111_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1080_load_0_req_0;
      array_obj_ref_1132_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_1188_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1116_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1111_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1080_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= array_obj_ref_1132_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_1188_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1116_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1111_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1080_load_0_req_1;
      array_obj_ref_1132_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_1188_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1116_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1111_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1080_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= update_control_register_pipe_1091(0);
      guard_vector(2)  <= update_free_q_pipe_1099(0);
      guard_vector(3)  <=  '1';
      guard_vector(4)  <= update_server_num_1107(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1132_word_address_0 & array_obj_ref_1188_word_address_0 & array_obj_ref_1116_word_address_0 & array_obj_ref_1111_word_address_0 & array_obj_ref_1080_word_address_0;
      array_obj_ref_1132_data_0 <= data_out(159 downto 128);
      array_obj_ref_1188_data_0 <= data_out(127 downto 96);
      array_obj_ref_1116_data_0 <= data_out(95 downto 64);
      array_obj_ref_1111_data_0 <= data_out(63 downto 32);
      array_obj_ref_1080_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_AFB_NIC_REQUEST_1135_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(73 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1135_inst_req_0;
      RPIPE_AFB_NIC_REQUEST_1135_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1135_inst_req_1;
      RPIPE_AFB_NIC_REQUEST_1135_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_1136 <= data_out(73 downto 0);
      AFB_NIC_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST_read_0", data_width => 74,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_REQUEST_pipe_read_req(0),
          oack => AFB_NIC_REQUEST_pipe_read_ack(0),
          odata => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_AFB_NIC_RESPONSE_1225_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1225_inst_req_0;
      WPIPE_AFB_NIC_RESPONSE_1225_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1225_inst_req_1;
      WPIPE_AFB_NIC_RESPONSE_1225_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_1224;
      AFB_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_RESPONSE_pipe_write_req(0),
          oack => AFB_NIC_RESPONSE_pipe_write_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_CONTROL_REGISTER_1109_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1109_inst_req_0;
      WPIPE_CONTROL_REGISTER_1109_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1109_inst_req_1;
      WPIPE_CONTROL_REGISTER_1109_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_1091(0);
      data_in <= array_obj_ref_1111_wire;
      CONTROL_REGISTER_write_1_gI: SplitGuardInterface generic map(name => "CONTROL_REGISTER_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      CONTROL_REGISTER_write_1: OutputPortRevised -- 
        generic map ( name => "CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => CONTROL_REGISTER_pipe_write_req(0),
          oack => CONTROL_REGISTER_pipe_write_ack(0),
          odata => CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_FREE_Q_1122_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_FREE_Q_1122_inst_req_0;
      WPIPE_FREE_Q_1122_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_FREE_Q_1122_inst_req_1;
      WPIPE_FREE_Q_1122_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_free_q_pipe_1093_delayed_5_0_1120(0);
      data_in <= type_cast_1127_wire;
      FREE_Q_write_2_gI: SplitGuardInterface generic map(name => "FREE_Q_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      FREE_Q_write_2: OutputPortRevised -- 
        generic map ( name => "FREE_Q", data_width => 36, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => FREE_Q_pipe_write_req(0),
          oack => FREE_Q_pipe_write_ack(0),
          odata => FREE_Q_pipe_write_data(35 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_NUMBER_OF_SERVERS_1130_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1130_inst_req_0;
      WPIPE_NUMBER_OF_SERVERS_1130_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1130_inst_req_1;
      WPIPE_NUMBER_OF_SERVERS_1130_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_server_num_1107(0);
      data_in <= array_obj_ref_1132_wire;
      NUMBER_OF_SERVERS_write_3_gI: SplitGuardInterface generic map(name => "NUMBER_OF_SERVERS_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NUMBER_OF_SERVERS_write_3: OutputPortRevised -- 
        generic map ( name => "NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1208_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1208_call_req_0;
      call_stmt_1208_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1208_call_req_1;
      call_stmt_1208_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_1166_delayed_5_0_1192(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_1167_delayed_5_0_1195 & rval_1189 & wdata_1169_delayed_5_0_1198 & index_1170_delayed_5_0_1201;
      wval_1208 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end SoftwareRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity UpdateRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    bmask : in  std_logic_vector(3 downto 0);
    rval : in  std_logic_vector(31 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    index : in  std_logic_vector(5 downto 0);
    wval : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity UpdateRegister;
architecture UpdateRegister_arch of UpdateRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 74)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal rval_buffer :  std_logic_vector(31 downto 0);
  signal rval_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(5 downto 0);
  signal index_update_enable: Boolean;
  -- output port buffer signals
  signal wval_buffer :  std_logic_vector(31 downto 0);
  signal wval_update_enable: Boolean;
  signal UpdateRegister_CP_34_start: Boolean;
  signal UpdateRegister_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u16_u32_170_inst_req_0 : boolean;
  signal CONCAT_u16_u32_170_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_170_inst_req_1 : boolean;
  signal CONCAT_u16_u32_170_inst_ack_1 : boolean;
  signal array_obj_ref_173_store_0_req_0 : boolean;
  signal array_obj_ref_173_store_0_ack_0 : boolean;
  signal array_obj_ref_173_store_0_req_1 : boolean;
  signal array_obj_ref_173_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "UpdateRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 74) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(3 downto 0) <= bmask;
  bmask_buffer <= in_buffer_data_out(3 downto 0);
  in_buffer_data_in(35 downto 4) <= rval;
  rval_buffer <= in_buffer_data_out(35 downto 4);
  in_buffer_data_in(67 downto 36) <= wdata;
  wdata_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(73 downto 68) <= index;
  index_buffer <= in_buffer_data_out(73 downto 68);
  in_buffer_data_in(tag_length + 73 downto 74) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 73 downto 74);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  UpdateRegister_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "UpdateRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wval_buffer;
  wval <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  UpdateRegister_CP_34: Block -- control-path 
    signal UpdateRegister_CP_34_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    UpdateRegister_CP_34_elements(0) <= UpdateRegister_CP_34_start;
    UpdateRegister_CP_34_symbol <= UpdateRegister_CP_34_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	5 
    -- CP-element group 0:  members (39) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_sample_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_update_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/rr
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/cr
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_update_start_
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_offset_calculated
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resized_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_computed_0
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_word_addrgen/root_register_ack
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/cr
      -- 
    cr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => array_obj_ref_173_store_0_req_1); -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_170_inst_req_0); -- 
    cr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_170_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_sample_completed_
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Sample/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_170_inst_ack_0, ack => UpdateRegister_CP_34_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_update_completed_
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/$exit
      -- CP-element group 2: 	 assign_stmt_106_to_assign_stmt_175/CONCAT_u16_u32_170_Update/ca
      -- 
    ca_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_170_inst_ack_1, ack => UpdateRegister_CP_34_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_sample_start_
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/$exit
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/split_req
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/array_obj_ref_173_Split/split_ack
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/rr
      -- 
    rr_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(3), ack => array_obj_ref_173_store_0_req_0); -- 
    UpdateRegister_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "UpdateRegister_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= UpdateRegister_CP_34_elements(2) & UpdateRegister_CP_34_elements(0);
      gj_UpdateRegister_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => UpdateRegister_CP_34_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_sample_completed_
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Sample/word_access_start/word_0/ra
      -- 
    ra_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_store_0_ack_0, ack => UpdateRegister_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_update_completed_
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_106_to_assign_stmt_175/array_obj_ref_173_Update/word_access_complete/word_0/ca
      -- 
    ca_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_173_store_0_ack_1, ack => UpdateRegister_CP_34_elements(5)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_160_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_169_wire : std_logic_vector(15 downto 0);
    signal MUX_155_wire : std_logic_vector(7 downto 0);
    signal MUX_159_wire : std_logic_vector(7 downto 0);
    signal MUX_164_wire : std_logic_vector(7 downto 0);
    signal MUX_168_wire : std_logic_vector(7 downto 0);
    signal R_index_172_resized : std_logic_vector(5 downto 0);
    signal R_index_172_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_173_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_173_word_offset_0 : std_logic_vector(5 downto 0);
    signal b0_106 : std_logic_vector(0 downto 0);
    signal b1_110 : std_logic_vector(0 downto 0);
    signal b2_114 : std_logic_vector(0 downto 0);
    signal b3_118 : std_logic_vector(0 downto 0);
    signal r0_122 : std_logic_vector(7 downto 0);
    signal r1_126 : std_logic_vector(7 downto 0);
    signal r2_130 : std_logic_vector(7 downto 0);
    signal r3_134 : std_logic_vector(7 downto 0);
    signal w0_138 : std_logic_vector(7 downto 0);
    signal w1_142 : std_logic_vector(7 downto 0);
    signal w2_146 : std_logic_vector(7 downto 0);
    signal w3_150 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_173_offset_scale_factor_0 <= "000001";
    array_obj_ref_173_resized_base_address <= "000000";
    array_obj_ref_173_word_offset_0 <= "000000";
    -- flow-through select operator MUX_155_inst
    MUX_155_wire <= w0_138 when (b0_106(0) /=  '0') else r0_122;
    -- flow-through select operator MUX_159_inst
    MUX_159_wire <= w1_142 when (b1_110(0) /=  '0') else r1_126;
    -- flow-through select operator MUX_164_inst
    MUX_164_wire <= w2_146 when (b2_114(0) /=  '0') else r2_130;
    -- flow-through select operator MUX_168_inst
    MUX_168_wire <= w3_150 when (b3_118(0) /=  '0') else r3_134;
    -- flow-through slice operator slice_105_inst
    b0_106 <= bmask_buffer(3 downto 3);
    -- flow-through slice operator slice_109_inst
    b1_110 <= bmask_buffer(2 downto 2);
    -- flow-through slice operator slice_113_inst
    b2_114 <= bmask_buffer(1 downto 1);
    -- flow-through slice operator slice_117_inst
    b3_118 <= bmask_buffer(0 downto 0);
    -- flow-through slice operator slice_121_inst
    r0_122 <= rval_buffer(31 downto 24);
    -- flow-through slice operator slice_125_inst
    r1_126 <= rval_buffer(23 downto 16);
    -- flow-through slice operator slice_129_inst
    r2_130 <= rval_buffer(15 downto 8);
    -- flow-through slice operator slice_133_inst
    r3_134 <= rval_buffer(7 downto 0);
    -- flow-through slice operator slice_137_inst
    w0_138 <= wdata_buffer(31 downto 24);
    -- flow-through slice operator slice_141_inst
    w1_142 <= wdata_buffer(23 downto 16);
    -- flow-through slice operator slice_145_inst
    w2_146 <= wdata_buffer(15 downto 8);
    -- flow-through slice operator slice_149_inst
    w3_150 <= wdata_buffer(7 downto 0);
    -- equivalence array_obj_ref_173_addr_0
    process(array_obj_ref_173_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_173_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_173_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_gather_scatter
    process(wval_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := wval_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_173_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_0_rename
    process(R_index_172_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_172_resized;
      ov(5 downto 0) := iv;
      R_index_172_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(5 downto 0) := iv;
      R_index_172_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_index_offset
    process(R_index_172_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_172_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_173_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_173_root_address_inst
    process(array_obj_ref_173_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_173_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_173_root_address <= ov(5 downto 0);
      --
    end process;
    -- shared split operator group (0) : CONCAT_u16_u32_170_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_160_wire & CONCAT_u8_u16_169_wire;
      wval_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_170_inst_req_0;
      CONCAT_u16_u32_170_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_170_inst_req_1;
      CONCAT_u16_u32_170_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator CONCAT_u8_u16_160_inst
    process(MUX_155_wire, MUX_159_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_155_wire, MUX_159_wire, tmp_var);
      CONCAT_u8_u16_160_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_169_inst
    process(MUX_164_wire, MUX_168_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_164_wire, MUX_168_wire, tmp_var);
      CONCAT_u8_u16_169_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_173_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_173_store_0_req_0;
      array_obj_ref_173_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_173_store_0_req_1;
      array_obj_ref_173_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_173_word_address_0;
      data_in <= array_obj_ref_173_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(5 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end UpdateRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity accessMemory is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(7 downto 0);
    addr : in  std_logic_vector(35 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemory;
architecture accessMemory_arch of accessMemory is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 110)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(7 downto 0);
  signal bmask_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemory_CP_329_start: Boolean;
  signal accessMemory_CP_329_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemory_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 110) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(9 downto 2) <= bmask;
  bmask_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(45 downto 10) <= addr;
  addr_buffer <= in_buffer_data_out(45 downto 10);
  in_buffer_data_in(109 downto 46) <= wdata;
  wdata_buffer <= in_buffer_data_out(109 downto 46);
  in_buffer_data_in(tag_length + 109 downto 110) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 109 downto 110);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= lock_update_enable & rwbar_update_enable & bmask_update_enable & addr_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemory_CP_329_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemory_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_329_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemory_CP_329_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_329_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemory_CP_329: Block -- control-path 
    signal accessMemory_CP_329_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    accessMemory_CP_329_elements(0) <= accessMemory_CP_329_start;
    accessMemory_CP_329_symbol <= accessMemory_CP_329_elements(22);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	11 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_267_to_stmt_287/$entry
      -- 
    accessMemory_CP_329_elements(1) <= accessMemory_CP_329_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_267_to_stmt_287/lock_update_enable
      -- CP-element group 2: 	 assign_stmt_267_to_stmt_287/lock_update_enable_out
      -- 
    accessMemory_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	9 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_267_to_stmt_287/rwbar_update_enable
      -- CP-element group 3: 	 assign_stmt_267_to_stmt_287/rwbar_update_enable_out
      -- 
    accessMemory_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	9 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	18 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_267_to_stmt_287/bmask_update_enable
      -- CP-element group 4: 	 assign_stmt_267_to_stmt_287/bmask_update_enable_out
      -- 
    accessMemory_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	9 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_267_to_stmt_287/addr_update_enable
      -- CP-element group 5: 	 assign_stmt_267_to_stmt_287/addr_update_enable_out
      -- 
    accessMemory_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	20 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_267_to_stmt_287/wdata_update_enable
      -- CP-element group 6: 	 assign_stmt_267_to_stmt_287/wdata_update_enable_out
      -- 
    accessMemory_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_329_elements(9);
      gj_accessMemory_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	21 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_267_to_stmt_287/rdata_update_enable
      -- CP-element group 7: 	 assign_stmt_267_to_stmt_287/rdata_update_enable_in
      -- 
    accessMemory_CP_329_elements(7) <= accessMemory_CP_329_elements(21);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_sample_start_
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/req
      -- 
    req_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(8), ack => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0); -- 
    accessMemory_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(1) & accessMemory_CP_329_elements(10);
      gj_accessMemory_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: 	3 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	5 
    -- CP-element group 9: 	6 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_sample_completed_
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_update_start_
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Sample/ack
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/$entry
      -- CP-element group 9: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/req
      -- 
    ack_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0, ack => accessMemory_CP_329_elements(9)); -- 
    req_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(9), ack => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_update_completed_
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/$exit
      -- CP-element group 10: 	 assign_stmt_267_to_stmt_287/WPIPE_NIC_TO_MEMORY_REQUEST_268_Update/ack
      -- 
    ack_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1, ack => accessMemory_CP_329_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_sample_start_
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/rr
      -- 
    rr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(11), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0); -- 
    accessMemory_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(1) & accessMemory_CP_329_elements(14);
      gj_accessMemory_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	7 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_update_start_
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/$entry
      -- CP-element group 12: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/cr
      -- 
    cr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_329_elements(12), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1); -- 
    accessMemory_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(13) & accessMemory_CP_329_elements(7);
      gj_accessMemory_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	12 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_sample_completed_
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Sample/ra
      -- 
    ra_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0, ack => accessMemory_CP_329_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_update_completed_
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/$exit
      -- CP-element group 14: 	 assign_stmt_267_to_stmt_287/RPIPE_MEMORY_TO_NIC_RESPONSE_272_Update/ca
      -- 
    ca_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1, ack => accessMemory_CP_329_elements(14)); -- 
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 assign_stmt_267_to_stmt_287/$exit
      -- 
    accessMemory_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_329_elements(14) & accessMemory_CP_329_elements(10);
      gj_accessMemory_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_329_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 lock_update_enable
      -- 
    accessMemory_CP_329_elements(16) <= accessMemory_CP_329_elements(2);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 rwbar_update_enable
      -- 
    accessMemory_CP_329_elements(17) <= accessMemory_CP_329_elements(3);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	4 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 bmask_update_enable
      -- 
    accessMemory_CP_329_elements(18) <= accessMemory_CP_329_elements(4);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 addr_update_enable
      -- 
    accessMemory_CP_329_elements(19) <= accessMemory_CP_329_elements(5);
    -- CP-element group 20:  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 wdata_update_enable
      -- 
    accessMemory_CP_329_elements(20) <= accessMemory_CP_329_elements(6);
    -- CP-element group 21:  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	7 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 rdata_update_enable
      -- 
    -- CP-element group 22:  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 $exit
      -- 
    accessMemory_CP_329_elements(22) <= accessMemory_CP_329_elements(15);
    --  hookup: inputs to control-path 
    accessMemory_CP_329_elements(21) <= rdata_update_enable;
    -- hookup: output from control-path 
    lock_update_enable <= accessMemory_CP_329_elements(16);
    rwbar_update_enable <= accessMemory_CP_329_elements(17);
    bmask_update_enable <= accessMemory_CP_329_elements(18);
    addr_update_enable <= accessMemory_CP_329_elements(19);
    wdata_update_enable <= accessMemory_CP_329_elements(20);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_260_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_262_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_265_wire : std_logic_vector(99 downto 0);
    signal err_277 : std_logic_vector(0 downto 0);
    signal request_267 : std_logic_vector(109 downto 0);
    signal response_273 : std_logic_vector(64 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_276_inst
    err_277 <= response_273(64 downto 64);
    -- flow-through slice operator slice_280_inst
    rdata_buffer <= response_273(63 downto 0);
    -- binary operator CONCAT_u10_u110_266_inst
    process(CONCAT_u2_u10_262_wire, CONCAT_u36_u100_265_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_262_wire, CONCAT_u36_u100_265_wire, tmp_var);
      request_267 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_260_inst
    process(lock_buffer, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(lock_buffer, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_260_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u10_262_inst
    process(CONCAT_u1_u2_260_wire, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_260_wire, bmask_buffer, tmp_var);
      CONCAT_u2_u10_262_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_265_inst
    process(addr_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_buffer, wdata_buffer, tmp_var);
      CONCAT_u36_u100_265_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_0;
      RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_req_1;
      RPIPE_MEMORY_TO_NIC_RESPONSE_272_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_273 <= data_out(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE_read_0", data_width => 65,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_TO_MEMORY_REQUEST_268_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_0;
      WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_req_1;
      WPIPE_NIC_TO_MEMORY_REQUEST_268_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_267;
      NIC_TO_MEMORY_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_write_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemory_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity acquireMutex is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    m_ok : out  std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity acquireMutex;
architecture acquireMutex_arch of acquireMutex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal m_ok_buffer :  std_logic_vector(0 downto 0);
  signal acquireMutex_CP_381_start: Boolean;
  signal acquireMutex_CP_381_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal if_stmt_313_branch_ack_0 : boolean;
  signal call_stmt_308_call_req_1 : boolean;
  signal if_stmt_313_branch_ack_1 : boolean;
  signal call_stmt_336_call_req_1 : boolean;
  signal call_stmt_336_call_ack_1 : boolean;
  signal if_stmt_313_branch_req_0 : boolean;
  signal call_stmt_336_call_ack_0 : boolean;
  signal call_stmt_308_call_ack_0 : boolean;
  signal call_stmt_336_call_req_0 : boolean;
  signal call_stmt_308_call_req_0 : boolean;
  signal call_stmt_308_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "acquireMutex_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  acquireMutex_CP_381_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "acquireMutex_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  m_ok_buffer <= "1";
  out_buffer_data_in(0 downto 0) <= m_ok_buffer;
  m_ok <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireMutex_CP_381_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= acquireMutex_CP_381_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireMutex_CP_381_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  acquireMutex_CP_381: Block -- control-path 
    signal acquireMutex_CP_381_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    acquireMutex_CP_381_elements(0) <= acquireMutex_CP_381_start;
    acquireMutex_CP_381_symbol <= acquireMutex_CP_381_elements(6);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295/$exit
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296__entry__
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295__exit__
      -- CP-element group 0: 	 branch_block_stmt_292/assign_stmt_295__entry__
      -- CP-element group 0: 	 branch_block_stmt_292/branch_block_stmt_292__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_292/$entry
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_292/merge_stmt_296__entry___PhiReq/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	7 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_sample_completed_
      -- 
    cra_413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_308_call_ack_0, ack => acquireMutex_CP_381_elements(1)); -- 
    -- CP-element group 2:  branch  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (27) 
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_else_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312__exit__
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_if_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/EQ_u32_u1_316_place
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/EQ_u32_u1_316_inputs/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/branch_req
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/EQ_u32_u1_316_inputs/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/ca
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/$exit
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_eval_test/EQ_u32_u1_316/SplitProtocol/Update/cr
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313__entry__
      -- CP-element group 2: 	 branch_block_stmt_292/if_stmt_313_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/cca
      -- 
    cca_418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_308_call_ack_1, ack => acquireMutex_CP_381_elements(2)); -- 
    branch_req_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(2), ack => if_stmt_313_branch_req_0); -- 
    -- CP-element group 3:  transition  place  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	7 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_292/if_stmt_313_if_link/if_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_292/if_stmt_313_if_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_292/loopback_PhiReq/$exit
      -- CP-element group 3: 	 branch_block_stmt_292/loopback_PhiReq/$entry
      -- CP-element group 3: 	 branch_block_stmt_292/loopback
      -- 
    if_choice_transition_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_313_branch_ack_1, ack => acquireMutex_CP_381_elements(3)); -- 
    -- CP-element group 4:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (11) 
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_313_else_link/else_choice_transition
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_313_else_link/$exit
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Update/ccr
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Sample/crr
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_update_start_
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336__entry__
      -- CP-element group 4: 	 branch_block_stmt_292/if_stmt_313__exit__
      -- CP-element group 4: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/$entry
      -- 
    else_choice_transition_454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_313_branch_ack_0, ack => acquireMutex_CP_381_elements(4)); -- 
    ccr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(4), ack => call_stmt_336_call_req_1); -- 
    crr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(4), ack => call_stmt_336_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Sample/cra
      -- CP-element group 5: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_sample_completed_
      -- 
    cra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_336_call_ack_0, ack => acquireMutex_CP_381_elements(5)); -- 
    -- CP-element group 6:  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (10) 
      -- CP-element group 6: 	 $exit
      -- CP-element group 6: 	 assign_stmt_341/$exit
      -- CP-element group 6: 	 assign_stmt_341/$entry
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Update/cca
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/call_stmt_336_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_292/branch_block_stmt_292__exit__
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336__exit__
      -- CP-element group 6: 	 branch_block_stmt_292/assign_stmt_325_to_call_stmt_336/$exit
      -- CP-element group 6: 	 branch_block_stmt_292/$exit
      -- 
    cca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_336_call_ack_1, ack => acquireMutex_CP_381_elements(6)); -- 
    -- CP-element group 7:  merge  fork  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: 	3 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: 	2 
    -- CP-element group 7:  members (13) 
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/ccr
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312__entry__
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/$entry
      -- CP-element group 7: 	 branch_block_stmt_292/merge_stmt_296__exit__
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/crr
      -- CP-element group 7: 	 branch_block_stmt_292/merge_stmt_296_PhiAck/dummy
      -- CP-element group 7: 	 branch_block_stmt_292/merge_stmt_296_PhiAck/$exit
      -- CP-element group 7: 	 branch_block_stmt_292/merge_stmt_296_PhiAck/$entry
      -- CP-element group 7: 	 branch_block_stmt_292/merge_stmt_296_PhiReqMerge
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_update_start_
      -- CP-element group 7: 	 branch_block_stmt_292/call_stmt_308_to_assign_stmt_312/call_stmt_308_sample_start_
      -- 
    ccr_417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(7), ack => call_stmt_308_call_req_1); -- 
    crr_412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_381_elements(7), ack => call_stmt_308_call_req_0); -- 
    acquireMutex_CP_381_elements(7) <= OrReduce(acquireMutex_CP_381_elements(0) & acquireMutex_CP_381_elements(3));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u32_u1_316_wire : std_logic_vector(0 downto 0);
    signal NOT_u8_u8_303_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_332_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_336 : std_logic_vector(63 downto 0);
    signal konst_315_wire_constant : std_logic_vector(31 downto 0);
    signal mutex_address_295 : std_logic_vector(35 downto 0);
    signal mutex_plus_nentries_308 : std_logic_vector(63 downto 0);
    signal mutex_val_312 : std_logic_vector(31 downto 0);
    signal slice_323_wire : std_logic_vector(31 downto 0);
    signal type_cast_298_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_300_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_306_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_321_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_327_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_329_wire_constant : std_logic_vector(0 downto 0);
    signal wval_325 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_303_wire_constant <= "11111111";
    NOT_u8_u8_332_wire_constant <= "11111111";
    konst_315_wire_constant <= "00000000000000000000000000000001";
    type_cast_298_wire_constant <= "1";
    type_cast_300_wire_constant <= "1";
    type_cast_306_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_321_wire_constant <= "00000000000000000000000000000001";
    type_cast_327_wire_constant <= "0";
    type_cast_329_wire_constant <= "0";
    -- flow-through slice operator slice_311_inst
    mutex_val_312 <= mutex_plus_nentries_308(63 downto 32);
    -- flow-through slice operator slice_323_inst
    slice_323_wire <= mutex_plus_nentries_308(31 downto 0);
    -- interlock W_mutex_address_293_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 35 downto 0) := q_base_address_buffer(35 downto 0);
      mutex_address_295 <= tmp_var; -- 
    end process;
    if_stmt_313_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u32_u1_316_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_313_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_313_branch_req_0,
          ack0 => if_stmt_313_branch_ack_0,
          ack1 => if_stmt_313_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u32_u64_324_inst
    process(type_cast_321_wire_constant, slice_323_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_321_wire_constant, slice_323_wire, tmp_var);
      wval_325 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_316_inst
    process(mutex_val_312) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mutex_val_312, konst_315_wire_constant, tmp_var);
      EQ_u32_u1_316_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_336_call call_stmt_308_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_336_call_req_0;
      reqL_unguarded(0) <= call_stmt_308_call_req_0;
      call_stmt_336_call_ack_0 <= ackL_unguarded(1);
      call_stmt_308_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_336_call_req_1;
      reqR_unguarded(0) <= call_stmt_308_call_req_1;
      call_stmt_336_call_ack_1 <= ackR_unguarded(1);
      call_stmt_308_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_327_wire_constant & type_cast_329_wire_constant & NOT_u8_u8_332_wire_constant & mutex_address_295 & wval_325 & type_cast_298_wire_constant & type_cast_300_wire_constant & NOT_u8_u8_303_wire_constant & mutex_address_295 & type_cast_306_wire_constant;
      ignore_336 <= data_out(127 downto 64);
      mutex_plus_nentries_308 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end acquireMutex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity delay_time_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    T : in  std_logic_vector(31 downto 0);
    delay_done : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity delay_time_Operator;
architecture delay_time_Operator_arch of delay_time_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal T_buffer :  std_logic_vector(31 downto 0);
  signal T_update_enable: Boolean;
  signal T_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal delay_done_buffer :  std_logic_vector(0 downto 0);
  signal delay_time_CP_1212_start: Boolean;
  signal delay_time_CP_1212_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_845_branch_req_0 : boolean;
  signal phi_stmt_847_req_0 : boolean;
  signal phi_stmt_847_req_1 : boolean;
  signal phi_stmt_847_ack_0 : boolean;
  signal nR_856_849_buf_req_0 : boolean;
  signal nR_856_849_buf_ack_0 : boolean;
  signal nR_856_849_buf_req_1 : boolean;
  signal nR_856_849_buf_ack_1 : boolean;
  signal T_850_buf_req_0 : boolean;
  signal T_850_buf_ack_0 : boolean;
  signal T_850_buf_req_1 : boolean;
  signal T_850_buf_ack_1 : boolean;
  signal do_while_stmt_845_branch_ack_0 : boolean;
  signal do_while_stmt_845_branch_ack_1 : boolean;
  -- 
begin --  
  sample_ack <= delay_time_CP_1212_symbol;
  -- input handling ------------------------------------------------
  T_buffer <= T;
  delay_time_CP_1212_start <= sample_req;
  -- output handling  -------------------------------------------------------
  delay_done_buffer <= "1";
  delay_done <= delay_done_buffer;
  update_ack_symbol <= delay_time_CP_1212_symbol;
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  delay_time_CP_1212: Block -- control-path 
    signal delay_time_CP_1212_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    delay_time_CP_1212_elements(0) <= delay_time_CP_1212_start;
    delay_time_CP_1212_symbol <= delay_time_CP_1212_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_844/$entry
      -- CP-element group 0: 	 branch_block_stmt_844/branch_block_stmt_844__entry__
      -- CP-element group 0: 	 branch_block_stmt_844/do_while_stmt_845__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	32 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (8) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_844/$exit
      -- CP-element group 1: 	 branch_block_stmt_844/branch_block_stmt_844__exit__
      -- CP-element group 1: 	 branch_block_stmt_844/do_while_stmt_845__exit__
      -- CP-element group 1: 	 branch_block_stmt_844/assign_stmt_863__entry__
      -- CP-element group 1: 	 branch_block_stmt_844/assign_stmt_863__exit__
      -- CP-element group 1: 	 branch_block_stmt_844/assign_stmt_863/$entry
      -- CP-element group 1: 	 branch_block_stmt_844/assign_stmt_863/$exit
      -- 
    delay_time_CP_1212_elements(1) <= delay_time_CP_1212_elements(32);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_844/do_while_stmt_845/$entry
      -- CP-element group 2: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845__entry__
      -- 
    delay_time_CP_1212_elements(2) <= delay_time_CP_1212_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	32 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845__exit__
      -- 
    -- Element group delay_time_CP_1212_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_844/do_while_stmt_845/loop_back
      -- 
    -- Element group delay_time_CP_1212_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	31 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_844/do_while_stmt_845/condition_done
      -- CP-element group 5: 	 branch_block_stmt_844/do_while_stmt_845/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_844/do_while_stmt_845/loop_taken/$entry
      -- 
    delay_time_CP_1212_elements(5) <= delay_time_CP_1212_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	14 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_844/do_while_stmt_845/loop_body_done
      -- 
    delay_time_CP_1212_elements(6) <= delay_time_CP_1212_elements(14);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/back_edge_to_loop_body
      -- 
    delay_time_CP_1212_elements(7) <= delay_time_CP_1212_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/first_time_through_loop_body
      -- 
    delay_time_CP_1212_elements(8) <= delay_time_CP_1212_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	29 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/loop_body_start
      -- 
    -- Element group delay_time_CP_1212_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	29 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/condition_evaluated
      -- 
    condition_evaluated_1238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1212_elements(10), ack => do_while_stmt_845_branch_req_0); -- 
    delay_time_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1212_elements(29) & delay_time_CP_1212_elements(15);
      gj_delay_time_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1212_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_sample_start__ps
      -- 
    delay_time_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1212_elements(12) & delay_time_CP_1212_elements(15);
      gj_delay_time_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1212_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_sample_start_
      -- 
    delay_time_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1212_elements(9) & delay_time_CP_1212_elements(14);
      gj_delay_time_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1212_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_update_start_
      -- CP-element group 13: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_update_start__ps
      -- 
    delay_time_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1212_elements(9) & delay_time_CP_1212_elements(15);
      gj_delay_time_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1212_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/$exit
      -- CP-element group 14: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_sample_completed__ps
      -- 
    -- Element group delay_time_CP_1212_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_update_completed__ps
      -- 
    -- Element group delay_time_CP_1212_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_loopback_trigger
      -- 
    delay_time_CP_1212_elements(16) <= delay_time_CP_1212_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_loopback_sample_req_ps
      -- 
    phi_stmt_847_loopback_sample_req_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_847_loopback_sample_req_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1212_elements(17), ack => phi_stmt_847_req_0); -- 
    -- Element group delay_time_CP_1212_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_entry_trigger
      -- 
    delay_time_CP_1212_elements(18) <= delay_time_CP_1212_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_entry_sample_req_ps
      -- 
    phi_stmt_847_entry_sample_req_1256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_847_entry_sample_req_1256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1212_elements(19), ack => phi_stmt_847_req_1); -- 
    -- Element group delay_time_CP_1212_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/phi_stmt_847_phi_mux_ack_ps
      -- 
    phi_stmt_847_phi_mux_ack_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_847_ack_0, ack => delay_time_CP_1212_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Sample/req
      -- 
    req_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1212_elements(21), ack => nR_856_849_buf_req_0); -- 
    -- Element group delay_time_CP_1212_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_update_start_
      -- CP-element group 22: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Update/req
      -- 
    req_1277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1212_elements(22), ack => nR_856_849_buf_req_1); -- 
    -- Element group delay_time_CP_1212_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_sample_completed__ps
      -- CP-element group 23: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Sample/ack
      -- 
    ack_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_856_849_buf_ack_0, ack => delay_time_CP_1212_elements(23)); -- 
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_nR_849_Update/ack
      -- 
    ack_1278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_856_849_buf_ack_1, ack => delay_time_CP_1212_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Sample/req
      -- 
    req_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1212_elements(25), ack => T_850_buf_req_0); -- 
    -- Element group delay_time_CP_1212_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_update_start_
      -- CP-element group 26: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Update/req
      -- 
    req_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1212_elements(26), ack => T_850_buf_req_1); -- 
    -- Element group delay_time_CP_1212_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Sample/ack
      -- 
    ack_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_850_buf_ack_0, ack => delay_time_CP_1212_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/R_T_850_Update/ack
      -- 
    ack_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_850_buf_ack_1, ack => delay_time_CP_1212_elements(28)); -- 
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	9 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	10 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_844/do_while_stmt_845/do_while_stmt_845_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group delay_time_CP_1212_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => delay_time_CP_1212_elements(9), ack => delay_time_CP_1212_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_844/do_while_stmt_845/loop_exit/$exit
      -- CP-element group 30: 	 branch_block_stmt_844/do_while_stmt_845/loop_exit/ack
      -- 
    ack_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_845_branch_ack_0, ack => delay_time_CP_1212_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_844/do_while_stmt_845/loop_taken/$exit
      -- CP-element group 31: 	 branch_block_stmt_844/do_while_stmt_845/loop_taken/ack
      -- 
    ack_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_845_branch_ack_1, ack => delay_time_CP_1212_elements(31)); -- 
    -- CP-element group 32:  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	3 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	1 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_844/do_while_stmt_845/$exit
      -- 
    delay_time_CP_1212_elements(32) <= delay_time_CP_1212_elements(3);
    delay_time_do_while_stmt_845_terminator_1307: loop_terminator -- 
      generic map (name => " delay_time_do_while_stmt_845_terminator_1307", max_iterations_in_flight =>7) 
      port map(loop_body_exit => delay_time_CP_1212_elements(6),loop_continue => delay_time_CP_1212_elements(31),loop_terminate => delay_time_CP_1212_elements(30),loop_back => delay_time_CP_1212_elements(4),loop_exit => delay_time_CP_1212_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_847_phi_seq_1297_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= delay_time_CP_1212_elements(16);
      delay_time_CP_1212_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= delay_time_CP_1212_elements(23);
      delay_time_CP_1212_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= delay_time_CP_1212_elements(24);
      delay_time_CP_1212_elements(17) <= phi_mux_reqs(0);
      triggers(1)  <= delay_time_CP_1212_elements(18);
      delay_time_CP_1212_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= delay_time_CP_1212_elements(27);
      delay_time_CP_1212_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= delay_time_CP_1212_elements(28);
      delay_time_CP_1212_elements(19) <= phi_mux_reqs(1);
      phi_stmt_847_phi_seq_1297 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_847_phi_seq_1297") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => delay_time_CP_1212_elements(11), 
          phi_sample_ack => delay_time_CP_1212_elements(14), 
          phi_update_req => delay_time_CP_1212_elements(13), 
          phi_update_ack => delay_time_CP_1212_elements(15), 
          phi_mux_ack => delay_time_CP_1212_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1239_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= delay_time_CP_1212_elements(7);
        preds(1)  <= delay_time_CP_1212_elements(8);
        entry_tmerge_1239 : transition_merge -- 
          generic map(name => " entry_tmerge_1239")
          port map (preds => preds, symbol_out => delay_time_CP_1212_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_847 : std_logic_vector(31 downto 0);
    signal T_850_buffered : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_860_wire : std_logic_vector(0 downto 0);
    signal konst_854_wire_constant : std_logic_vector(31 downto 0);
    signal konst_859_wire_constant : std_logic_vector(31 downto 0);
    signal nR_856 : std_logic_vector(31 downto 0);
    signal nR_856_849_buffered : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_854_wire_constant <= "00000000000000000000000000000001";
    konst_859_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_847: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nR_856_849_buffered & T_850_buffered;
      req <= phi_stmt_847_req_0 & phi_stmt_847_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_847",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_847_ack_0,
          idata => idata,
          odata => R_847,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_847
    T_850_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= T_850_buf_req_0;
      T_850_buf_ack_0<= wack(0);
      rreq(0) <= T_850_buf_req_1;
      T_850_buf_ack_1<= rack(0);
      T_850_buf : InterlockBuffer generic map ( -- 
        name => "T_850_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_850_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nR_856_849_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_856_849_buf_req_0;
      nR_856_849_buf_ack_0<= wack(0);
      rreq(0) <= nR_856_849_buf_req_1;
      nR_856_849_buf_ack_1<= rack(0);
      nR_856_849_buf : InterlockBuffer generic map ( -- 
        name => "nR_856_849_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_856_849_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_845_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u32_u1_860_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_845_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_845_branch_req_0,
          ack0 => do_while_stmt_845_branch_ack_0,
          ack1 => do_while_stmt_845_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator SUB_u32_u32_855_inst
    process(R_847) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_847, konst_854_wire_constant, tmp_var);
      nR_856 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_860_inst
    process(R_847) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(R_847, konst_859_wire_constant, tmp_var);
      UGT_u32_u1_860_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end delay_time_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    read_pointer : in  std_logic_vector(31 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueElement;
architecture getQueueElement_arch of getQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal read_pointer_buffer :  std_logic_vector(31 downto 0);
  signal read_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal getQueueElement_CP_511_start: Boolean;
  signal getQueueElement_CP_511_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_408_call_ack_0 : boolean;
  signal MUX_423_inst_ack_1 : boolean;
  signal call_stmt_408_call_req_0 : boolean;
  signal MUX_423_inst_req_1 : boolean;
  signal call_stmt_408_call_ack_1 : boolean;
  signal call_stmt_408_call_req_1 : boolean;
  signal MUX_423_inst_req_0 : boolean;
  signal MUX_423_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= read_pointer;
  read_pointer_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueElement_CP_511_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_511_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueElement_CP_511_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_511_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueElement_CP_511: Block -- control-path 
    signal getQueueElement_CP_511_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueElement_CP_511_elements(0) <= getQueueElement_CP_511_start;
    getQueueElement_CP_511_symbol <= getQueueElement_CP_511_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Sample/crr
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_complete/req
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_update_start_
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_sample_start_
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_update_start_
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Update/ccr
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Update/$entry
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_complete/$entry
      -- 
    crr_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_511_elements(0), ack => call_stmt_408_call_req_0); -- 
    ccr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_511_elements(0), ack => call_stmt_408_call_req_1); -- 
    req_543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_511_elements(0), ack => MUX_423_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Sample/cra
      -- CP-element group 1: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_sample_completed_
      -- 
    cra_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_408_call_ack_0, ack => getQueueElement_CP_511_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_start/$entry
      -- CP-element group 2: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_update_completed_
      -- CP-element group 2: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Update/cca
      -- CP-element group 2: 	 assign_stmt_383_to_assign_stmt_424/call_stmt_408_Update/$exit
      -- CP-element group 2: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_sample_start_
      -- CP-element group 2: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_start/req
      -- 
    cca_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_408_call_ack_1, ack => getQueueElement_CP_511_elements(2)); -- 
    req_538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_511_elements(2), ack => MUX_423_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_sample_completed_
      -- CP-element group 3: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_start/$exit
      -- CP-element group 3: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_start/ack
      -- 
    ack_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_423_inst_ack_0, ack => getQueueElement_CP_511_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_complete/ack
      -- CP-element group 4: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_complete/$exit
      -- CP-element group 4: 	 assign_stmt_383_to_assign_stmt_424/$exit
      -- CP-element group 4: 	 assign_stmt_383_to_assign_stmt_424/MUX_423_update_completed_
      -- CP-element group 4: 	 $exit
      -- 
    ack_544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_423_inst_ack_1, ack => getQueueElement_CP_511_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_420_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_392_wire : std_logic_vector(33 downto 0);
    signal NOT_u8_u8_403_wire_constant : std_logic_vector(7 downto 0);
    signal buffer_address_383 : std_logic_vector(35 downto 0);
    signal e0_412 : std_logic_vector(31 downto 0);
    signal e1_416 : std_logic_vector(31 downto 0);
    signal element_pair_408 : std_logic_vector(63 downto 0);
    signal element_pair_address_396 : std_logic_vector(35 downto 0);
    signal konst_419_wire_constant : std_logic_vector(31 downto 0);
    signal slice_388_wire : std_logic_vector(30 downto 0);
    signal type_cast_381_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_391_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_394_wire : std_logic_vector(35 downto 0);
    signal type_cast_398_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_400_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_406_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_403_wire_constant <= "11111111";
    konst_419_wire_constant <= "00000000000000000000000000000000";
    type_cast_381_wire_constant <= "000000000000000000000000000000010000";
    type_cast_391_wire_constant <= "000";
    type_cast_398_wire_constant <= "0";
    type_cast_400_wire_constant <= "1";
    type_cast_406_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    MUX_423_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_423_inst_req_0;
      MUX_423_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_423_inst_req_1;
      MUX_423_inst_ack_1<= update_ack(0);
      MUX_423_inst: SelectSplitProtocol generic map(name => "MUX_423_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => e1_416, y => e0_412, sel => BITSEL_u32_u1_420_wire, z => q_r_data_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_388_inst
    slice_388_wire <= read_pointer_buffer(31 downto 1);
    -- flow-through slice operator slice_411_inst
    e0_412 <= element_pair_408(63 downto 32);
    -- flow-through slice operator slice_415_inst
    e1_416 <= element_pair_408(31 downto 0);
    -- interlock type_cast_394_inst
    process(CONCAT_u31_u34_392_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_392_wire(33 downto 0);
      type_cast_394_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_382_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_381_wire_constant, tmp_var);
      buffer_address_383 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_395_inst
    process(buffer_address_383, type_cast_394_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_383, type_cast_394_wire, tmp_var);
      element_pair_address_396 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_420_inst
    process(read_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(read_pointer_buffer, konst_419_wire_constant, tmp_var);
      BITSEL_u32_u1_420_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_392_inst
    process(slice_388_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_388_wire, type_cast_391_wire_constant, tmp_var);
      CONCAT_u31_u34_392_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_408_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_408_call_req_0;
      call_stmt_408_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_408_call_req_1;
      call_stmt_408_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_398_wire_constant & type_cast_400_wire_constant & NOT_u8_u8_403_wire_constant & element_pair_address_396 & type_cast_406_wire_constant;
      element_pair_408 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : out  std_logic_vector(31 downto 0);
    rp : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointers;
architecture getQueuePointers_arch of getQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  signal getQueuePointers_CP_491_start: Boolean;
  signal getQueuePointers_CP_491_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_360_call_req_1 : boolean;
  signal call_stmt_360_call_ack_0 : boolean;
  signal call_stmt_360_call_req_0 : boolean;
  signal call_stmt_360_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointers_CP_491_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wp_buffer;
  wp <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= rp_buffer;
  rp <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_491_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointers_CP_491_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_491_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointers_CP_491: Block -- control-path 
    signal getQueuePointers_CP_491_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    getQueuePointers_CP_491_elements(0) <= getQueuePointers_CP_491_start;
    getQueuePointers_CP_491_symbol <= getQueuePointers_CP_491_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Update/ccr
      -- CP-element group 0: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_sample_start_
      -- CP-element group 0: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Update/$entry
      -- CP-element group 0: 	 call_stmt_360_to_assign_stmt_368/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Sample/crr
      -- CP-element group 0: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Sample/$entry
      -- CP-element group 0: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_update_start_
      -- 
    crr_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_491_elements(0), ack => call_stmt_360_call_req_0); -- 
    ccr_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_491_elements(0), ack => call_stmt_360_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_sample_completed_
      -- CP-element group 1: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Sample/cra
      -- CP-element group 1: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Sample/$exit
      -- 
    cra_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_360_call_ack_0, ack => getQueuePointers_CP_491_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Update/$exit
      -- CP-element group 2: 	 call_stmt_360_to_assign_stmt_368/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_Update/cca
      -- CP-element group 2: 	 call_stmt_360_to_assign_stmt_368/call_stmt_360_update_completed_
      -- 
    cca_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_360_call_ack_1, ack => getQueuePointers_CP_491_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_356_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_353_wire_constant : std_logic_vector(7 downto 0);
    signal konst_355_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_348_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_358_wire_constant : std_logic_vector(63 downto 0);
    signal wp_rp_360 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_353_wire_constant <= "11111111";
    konst_355_wire_constant <= "000000000000000000000000000000001000";
    type_cast_348_wire_constant <= "0";
    type_cast_350_wire_constant <= "1";
    type_cast_358_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through slice operator slice_363_inst
    wp_buffer <= wp_rp_360(63 downto 32);
    -- flow-through slice operator slice_367_inst
    rp_buffer <= wp_rp_360(31 downto 0);
    -- binary operator ADD_u36_u36_356_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_355_wire_constant, tmp_var);
      ADD_u36_u36_356_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_360_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_360_call_req_0;
      call_stmt_360_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_360_call_req_1;
      call_stmt_360_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_348_wire_constant & type_cast_350_wire_constant & NOT_u8_u8_353_wire_constant & ADD_u36_u36_356_wire & type_cast_358_wire_constant;
      wp_rp_360 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity getTxPacketPointerFromServer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_index : in  std_logic_vector(5 downto 0);
    pkt_pointer : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTxPacketPointerFromServer;
architecture getTxPacketPointerFromServer_arch of getTxPacketPointerFromServer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 6)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_index_buffer :  std_logic_vector(5 downto 0);
  signal queue_index_update_enable: Boolean;
  -- output port buffer signals
  signal pkt_pointer_buffer :  std_logic_vector(31 downto 0);
  signal pkt_pointer_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal getTxPacketPointerFromServer_CP_2468_start: Boolean;
  signal getTxPacketPointerFromServer_CP_2468_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1263_call_req_1 : boolean;
  signal call_stmt_1263_call_ack_1 : boolean;
  signal call_stmt_1263_call_ack_0 : boolean;
  signal call_stmt_1263_call_req_0 : boolean;
  signal call_stmt_1251_call_ack_1 : boolean;
  signal call_stmt_1251_call_req_1 : boolean;
  signal call_stmt_1251_call_ack_0 : boolean;
  signal call_stmt_1251_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 6) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= queue_index;
  queue_index_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(tag_length + 5 downto 6) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 5 downto 6);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 7);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= queue_index_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTxPacketPointerFromServer_CP_2468_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= pkt_pointer_buffer;
  pkt_pointer <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2468_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  pkt_pointer_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "pkt_pointer_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_pkt_pointer_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => pkt_pointer_update_enable, clk => clk, reset => reset); --
  end block;
  status_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "status_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_status_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => status_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2468_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2468_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTxPacketPointerFromServer_CP_2468: Block -- control-path 
    signal getTxPacketPointerFromServer_CP_2468_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    getTxPacketPointerFromServer_CP_2468_elements(0) <= getTxPacketPointerFromServer_CP_2468_start;
    getTxPacketPointerFromServer_CP_2468_symbol <= getTxPacketPointerFromServer_CP_2468_elements(16);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_1241_to_stmt_1268/$entry
      -- 
    getTxPacketPointerFromServer_CP_2468_elements(1) <= getTxPacketPointerFromServer_CP_2468_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_1241_to_stmt_1268/queue_index_update_enable_out
      -- CP-element group 2: 	 assign_stmt_1241_to_stmt_1268/queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_2468_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2468_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	14 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_1241_to_stmt_1268/pkt_pointer_update_enable_in
      -- CP-element group 3: 	 assign_stmt_1241_to_stmt_1268/pkt_pointer_update_enable
      -- 
    getTxPacketPointerFromServer_CP_2468_elements(3) <= getTxPacketPointerFromServer_CP_2468_elements(14);
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_1241_to_stmt_1268/status_update_enable_in
      -- CP-element group 4: 	 assign_stmt_1241_to_stmt_1268/status_update_enable
      -- 
    getTxPacketPointerFromServer_CP_2468_elements(4) <= getTxPacketPointerFromServer_CP_2468_elements(15);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_sample_start_
      -- CP-element group 5: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Sample/crr
      -- CP-element group 5: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Sample/$entry
      -- 
    crr_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2468_elements(5), ack => call_stmt_1251_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2468_elements(1) & getTxPacketPointerFromServer_CP_2468_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2468_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_update_start_
      -- CP-element group 6: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Update/ccr
      -- CP-element group 6: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Update/$entry
      -- 
    ccr_2492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2468_elements(6), ack => call_stmt_1251_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2468_elements(8) & getTxPacketPointerFromServer_CP_2468_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2468_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_sample_completed_
      -- CP-element group 7: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Sample/cra
      -- CP-element group 7: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Sample/$exit
      -- 
    cra_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1251_call_ack_0, ack => getTxPacketPointerFromServer_CP_2468_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Update/cca
      -- CP-element group 8: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_Update/$exit
      -- CP-element group 8: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1251_update_completed_
      -- 
    cca_2493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1251_call_ack_1, ack => getTxPacketPointerFromServer_CP_2468_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_sample_start_
      -- CP-element group 9: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Sample/crr
      -- CP-element group 9: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Sample/$entry
      -- 
    crr_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2468_elements(9), ack => call_stmt_1263_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2468_elements(8) & getTxPacketPointerFromServer_CP_2468_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2468_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Update/ccr
      -- CP-element group 10: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Update/$entry
      -- CP-element group 10: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_update_start_
      -- 
    ccr_2506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2468_elements(10), ack => call_stmt_1263_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "getTxPacketPointerFromServer_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2468_elements(3) & getTxPacketPointerFromServer_CP_2468_elements(4) & getTxPacketPointerFromServer_CP_2468_elements(12);
      gj_getTxPacketPointerFromServer_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2468_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_sample_completed_
      -- CP-element group 11: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Sample/cra
      -- CP-element group 11: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Sample/$exit
      -- 
    cra_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1263_call_ack_0, ack => getTxPacketPointerFromServer_CP_2468_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Update/cca
      -- CP-element group 12: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_Update/$exit
      -- CP-element group 12: 	 assign_stmt_1241_to_stmt_1268/$exit
      -- CP-element group 12: 	 assign_stmt_1241_to_stmt_1268/call_stmt_1263_update_completed_
      -- 
    cca_2507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1263_call_ack_1, ack => getTxPacketPointerFromServer_CP_2468_elements(12)); -- 
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_CP_2468_elements(13) <= getTxPacketPointerFromServer_CP_2468_elements(2);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 pkt_pointer_update_enable
      -- 
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 status_update_enable
      -- 
    -- CP-element group 16:  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 $exit
      -- 
    getTxPacketPointerFromServer_CP_2468_elements(16) <= getTxPacketPointerFromServer_CP_2468_elements(12);
    --  hookup: inputs to control-path 
    getTxPacketPointerFromServer_CP_2468_elements(15) <= status_update_enable;
    getTxPacketPointerFromServer_CP_2468_elements(14) <= pkt_pointer_update_enable;
    -- hookup: output from control-path 
    queue_index_update_enable <= getTxPacketPointerFromServer_CP_2468_elements(13);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1239_wire : std_logic_vector(5 downto 0);
    signal NOT_u4_u4_1246_wire_constant : std_logic_vector(3 downto 0);
    signal R_TX_QUEUES_REG_START_OFFSET_1238_wire_constant : std_logic_vector(5 downto 0);
    signal register_index_1241 : std_logic_vector(5 downto 0);
    signal tx_queue_pointer_32_1251 : std_logic_vector(31 downto 0);
    signal tx_queue_pointer_36_1257 : std_logic_vector(35 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1249_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1255_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1259_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1246_wire_constant <= "1111";
    R_TX_QUEUES_REG_START_OFFSET_1238_wire_constant <= "001010";
    type_cast_1243_wire_constant <= "1";
    type_cast_1249_wire_constant <= "00000000000000000000000000000000";
    type_cast_1255_wire_constant <= "0000";
    type_cast_1259_wire_constant <= "0";
    -- interlock type_cast_1240_inst
    process(ADD_u6_u6_1239_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1239_wire(5 downto 0);
      register_index_1241 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u6_u6_1239_inst
    process(queue_index_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(queue_index_buffer, R_TX_QUEUES_REG_START_OFFSET_1238_wire_constant, tmp_var);
      ADD_u6_u6_1239_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u36_1256_inst
    process(tx_queue_pointer_32_1251) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(tx_queue_pointer_32_1251, type_cast_1255_wire_constant, tmp_var);
      tx_queue_pointer_36_1257 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1251_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1251_call_req_0;
      call_stmt_1251_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1251_call_req_1;
      call_stmt_1251_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1243_wire_constant & NOT_u4_u4_1246_wire_constant & register_index_1241 & type_cast_1249_wire_constant;
      tx_queue_pointer_32_1251 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1263_call 
    popFromQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1263_call_req_0;
      call_stmt_1263_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1263_call_req_1;
      call_stmt_1263_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_1_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1259_wire_constant & tx_queue_pointer_36_1257;
      pkt_pointer_buffer <= data_out(32 downto 1);
      status_buffer <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getTxPacketPointerFromServer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity loadBuffer is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
    writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
    writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
    writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadBuffer;
architecture loadBuffer_arch of loadBuffer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal loadBuffer_CP_1000_start: Boolean;
  signal loadBuffer_CP_1000_symbol: Boolean;
  -- volatile/operator module components. 
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_699_call_req_1 : boolean;
  signal W_rx_buffer_pointer_691_delayed_8_0_703_inst_req_1 : boolean;
  signal call_stmt_699_call_ack_1 : boolean;
  signal call_stmt_699_call_req_0 : boolean;
  signal call_stmt_699_call_ack_0 : boolean;
  signal call_stmt_690_call_req_1 : boolean;
  signal call_stmt_690_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_684_delayed_4_0_691_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_691_delayed_8_0_703_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_691_delayed_8_0_703_inst_req_0 : boolean;
  signal call_stmt_710_call_req_1 : boolean;
  signal call_stmt_710_call_ack_1 : boolean;
  signal W_bad_packet_identifier_690_delayed_8_0_700_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_684_delayed_4_0_691_inst_req_1 : boolean;
  signal call_stmt_690_call_ack_0 : boolean;
  signal call_stmt_690_call_req_0 : boolean;
  signal W_rx_buffer_pointer_684_delayed_4_0_691_inst_ack_0 : boolean;
  signal W_bad_packet_identifier_690_delayed_8_0_700_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_691_delayed_8_0_703_inst_ack_1 : boolean;
  signal call_stmt_710_call_req_0 : boolean;
  signal call_stmt_710_call_ack_0 : boolean;
  signal W_bad_packet_identifier_690_delayed_8_0_700_inst_req_0 : boolean;
  signal W_bad_packet_identifier_690_delayed_8_0_700_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_684_delayed_4_0_691_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadBuffer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 31);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_buffer_pointer_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadBuffer_CP_1000_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadBuffer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1000_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  bad_packet_identifier_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 40) := "bad_packet_identifier_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_bad_packet_identifier_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => bad_packet_identifier_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 31,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadBuffer_CP_1000_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1000_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadBuffer_CP_1000: Block -- control-path 
    signal loadBuffer_CP_1000_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    loadBuffer_CP_1000_elements(0) <= loadBuffer_CP_1000_start;
    loadBuffer_CP_1000_symbol <= loadBuffer_CP_1000_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	20 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_690_to_call_stmt_710/$entry
      -- 
    loadBuffer_CP_1000_elements(1) <= loadBuffer_CP_1000_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	22 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	28 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_690_to_call_stmt_710/rx_buffer_pointer_update_enable_out
      -- CP-element group 2: 	 call_stmt_690_to_call_stmt_710/rx_buffer_pointer_update_enable
      -- 
    loadBuffer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(6) & loadBuffer_CP_1000_elements(10) & loadBuffer_CP_1000_elements(22);
      gj_loadBuffer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	29 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_690_to_call_stmt_710/bad_packet_identifier_update_enable
      -- CP-element group 3: 	 call_stmt_690_to_call_stmt_710/bad_packet_identifier_update_enable_in
      -- 
    loadBuffer_CP_1000_elements(3) <= loadBuffer_CP_1000_elements(29);
    -- CP-element group 4:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	27 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_sample_start_
      -- CP-element group 4: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Sample/crr
      -- CP-element group 4: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Sample/$entry
      -- 
    crr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(4), ack => call_stmt_690_call_req_0); -- 
    loadBuffer_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(1) & loadBuffer_CP_1000_elements(6) & loadBuffer_CP_1000_elements(27);
      gj_loadBuffer_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	14 
    -- CP-element group 5: 	7 
    -- CP-element group 5: 	27 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Update/ccr
      -- CP-element group 5: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Update/$entry
      -- CP-element group 5: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_update_start_
      -- 
    ccr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(5), ack => call_stmt_690_call_req_1); -- 
    loadBuffer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(14) & loadBuffer_CP_1000_elements(7) & loadBuffer_CP_1000_elements(27);
      gj_loadBuffer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: marked-successors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: 	4 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_sample_completed_
      -- CP-element group 6: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Sample/cra
      -- CP-element group 6: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Sample/$exit
      -- 
    cra_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_690_call_ack_0, ack => loadBuffer_CP_1000_elements(6)); -- 
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Update/$exit
      -- CP-element group 7: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_Update/cca
      -- CP-element group 7: 	 call_stmt_690_to_call_stmt_710/call_stmt_690_update_completed_
      -- 
    cca_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_690_call_ack_1, ack => loadBuffer_CP_1000_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Sample/$entry
      -- CP-element group 8: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_sample_start_
      -- CP-element group 8: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Sample/req
      -- 
    req_1031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(8), ack => W_rx_buffer_pointer_684_delayed_4_0_691_inst_req_0); -- 
    loadBuffer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(1) & loadBuffer_CP_1000_elements(10);
      gj_loadBuffer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Update/$entry
      -- CP-element group 9: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_update_start_
      -- CP-element group 9: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Update/req
      -- 
    req_1036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(9), ack => W_rx_buffer_pointer_684_delayed_4_0_691_inst_req_1); -- 
    loadBuffer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(14) & loadBuffer_CP_1000_elements(11);
      gj_loadBuffer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: 	2 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_sample_completed_
      -- CP-element group 10: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Sample/ack
      -- CP-element group 10: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Sample/$exit
      -- 
    ack_1032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_684_delayed_4_0_691_inst_ack_0, ack => loadBuffer_CP_1000_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Update/$exit
      -- CP-element group 11: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_Update/ack
      -- CP-element group 11: 	 call_stmt_690_to_call_stmt_710/assign_stmt_693_update_completed_
      -- 
    ack_1037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_684_delayed_4_0_691_inst_ack_1, ack => loadBuffer_CP_1000_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Sample/crr
      -- CP-element group 12: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Sample/$entry
      -- CP-element group 12: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_sample_start_
      -- 
    crr_1045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(12), ack => call_stmt_699_call_req_0); -- 
    loadBuffer_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(7) & loadBuffer_CP_1000_elements(11) & loadBuffer_CP_1000_elements(14);
      gj_loadBuffer_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	26 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Update/ccr
      -- CP-element group 13: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_update_start_
      -- CP-element group 13: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Update/$entry
      -- 
    ccr_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(13), ack => call_stmt_699_call_req_1); -- 
    loadBuffer_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(3) & loadBuffer_CP_1000_elements(15) & loadBuffer_CP_1000_elements(18) & loadBuffer_CP_1000_elements(26);
      gj_loadBuffer_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	5 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Sample/$exit
      -- CP-element group 14: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Sample/cra
      -- CP-element group 14: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_sample_completed_
      -- 
    cra_1046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_699_call_ack_0, ack => loadBuffer_CP_1000_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	24 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Update/cca
      -- CP-element group 15: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_Update/$exit
      -- CP-element group 15: 	 call_stmt_690_to_call_stmt_710/call_stmt_699_update_completed_
      -- 
    cca_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_699_call_ack_1, ack => loadBuffer_CP_1000_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Sample/$entry
      -- CP-element group 16: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_sample_start_
      -- CP-element group 16: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Sample/req
      -- 
    req_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(16), ack => W_bad_packet_identifier_690_delayed_8_0_700_inst_req_0); -- 
    loadBuffer_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(15) & loadBuffer_CP_1000_elements(18);
      gj_loadBuffer_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	26 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_update_start_
      -- CP-element group 17: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Update/req
      -- CP-element group 17: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Update/$entry
      -- 
    req_1064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(17), ack => W_bad_packet_identifier_690_delayed_8_0_700_inst_req_1); -- 
    loadBuffer_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(19) & loadBuffer_CP_1000_elements(26);
      gj_loadBuffer_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	13 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Sample/$exit
      -- CP-element group 18: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_sample_completed_
      -- CP-element group 18: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Sample/ack
      -- 
    ack_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_690_delayed_8_0_700_inst_ack_0, ack => loadBuffer_CP_1000_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Update/ack
      -- CP-element group 19: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_update_completed_
      -- CP-element group 19: 	 call_stmt_690_to_call_stmt_710/assign_stmt_702_Update/$exit
      -- 
    ack_1065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_690_delayed_8_0_700_inst_ack_1, ack => loadBuffer_CP_1000_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	1 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Sample/$entry
      -- CP-element group 20: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Sample/req
      -- CP-element group 20: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_sample_start_
      -- 
    req_1073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(20), ack => W_rx_buffer_pointer_691_delayed_8_0_703_inst_req_0); -- 
    loadBuffer_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(1) & loadBuffer_CP_1000_elements(22);
      gj_loadBuffer_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	26 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Update/req
      -- CP-element group 21: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_update_start_
      -- CP-element group 21: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Update/$entry
      -- 
    req_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(21), ack => W_rx_buffer_pointer_691_delayed_8_0_703_inst_req_1); -- 
    loadBuffer_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(23) & loadBuffer_CP_1000_elements(26);
      gj_loadBuffer_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	2 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_sample_completed_
      -- CP-element group 22: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Sample/ack
      -- CP-element group 22: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Sample/$exit
      -- 
    ack_1074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_691_delayed_8_0_703_inst_ack_0, ack => loadBuffer_CP_1000_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Update/$exit
      -- CP-element group 23: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_update_completed_
      -- CP-element group 23: 	 call_stmt_690_to_call_stmt_710/assign_stmt_705_Update/ack
      -- 
    ack_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_691_delayed_8_0_703_inst_ack_1, ack => loadBuffer_CP_1000_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Sample/$entry
      -- CP-element group 24: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_sample_start_
      -- CP-element group 24: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Sample/crr
      -- 
    crr_1087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(24), ack => call_stmt_710_call_req_0); -- 
    loadBuffer_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1000_elements(15) & loadBuffer_CP_1000_elements(19) & loadBuffer_CP_1000_elements(23) & loadBuffer_CP_1000_elements(26);
      gj_loadBuffer_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_update_start_
      -- CP-element group 25: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Update/$entry
      -- CP-element group 25: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Update/ccr
      -- 
    ccr_1092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1000_elements(25), ack => call_stmt_710_call_req_1); -- 
    loadBuffer_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadBuffer_CP_1000_elements(27);
      gj_loadBuffer_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1000_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	17 
    -- CP-element group 26: 	21 
    -- CP-element group 26: 	13 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Sample/$exit
      -- CP-element group 26: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Sample/cra
      -- CP-element group 26: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_sample_completed_
      -- 
    cra_1088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_0, ack => loadBuffer_CP_1000_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: 	4 
    -- CP-element group 27: 	5 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Update/$exit
      -- CP-element group 27: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_Update/cca
      -- CP-element group 27: 	 call_stmt_690_to_call_stmt_710/$exit
      -- CP-element group 27: 	 call_stmt_690_to_call_stmt_710/call_stmt_710_update_completed_
      -- 
    cca_1093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_710_call_ack_1, ack => loadBuffer_CP_1000_elements(27)); -- 
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 rx_buffer_pointer_update_enable
      -- 
    loadBuffer_CP_1000_elements(28) <= loadBuffer_CP_1000_elements(2);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	3 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 bad_packet_identifier_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    loadBuffer_CP_1000_elements(30) <= loadBuffer_CP_1000_elements(27);
    --  hookup: inputs to control-path 
    loadBuffer_CP_1000_elements(29) <= bad_packet_identifier_update_enable;
    -- hookup: output from control-path 
    rx_buffer_pointer_update_enable <= loadBuffer_CP_1000_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal bad_packet_identifier_690_delayed_8_0_702 : std_logic_vector(0 downto 0);
    signal last_keep_699 : std_logic_vector(7 downto 0);
    signal new_buf_pointer_690 : std_logic_vector(35 downto 0);
    signal packet_size_699 : std_logic_vector(7 downto 0);
    signal rx_buffer_pointer_684_delayed_4_0_693 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_691_delayed_8_0_705 : std_logic_vector(35 downto 0);
    -- 
  begin -- 
    W_bad_packet_identifier_690_delayed_8_0_700_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bad_packet_identifier_690_delayed_8_0_700_inst_req_0;
      W_bad_packet_identifier_690_delayed_8_0_700_inst_ack_0<= wack(0);
      rreq(0) <= W_bad_packet_identifier_690_delayed_8_0_700_inst_req_1;
      W_bad_packet_identifier_690_delayed_8_0_700_inst_ack_1<= rack(0);
      W_bad_packet_identifier_690_delayed_8_0_700_inst : InterlockBuffer generic map ( -- 
        name => "W_bad_packet_identifier_690_delayed_8_0_700_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bad_packet_identifier_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bad_packet_identifier_690_delayed_8_0_702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_684_delayed_4_0_691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_684_delayed_4_0_691_inst_req_0;
      W_rx_buffer_pointer_684_delayed_4_0_691_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_684_delayed_4_0_691_inst_req_1;
      W_rx_buffer_pointer_684_delayed_4_0_691_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_684_delayed_4_0_691_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_684_delayed_4_0_691_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_684_delayed_4_0_693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_691_delayed_8_0_703_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_691_delayed_8_0_703_inst_req_0;
      W_rx_buffer_pointer_691_delayed_8_0_703_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_691_delayed_8_0_703_inst_req_1;
      W_rx_buffer_pointer_691_delayed_8_0_703_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_691_delayed_8_0_703_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_691_delayed_8_0_703_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_691_delayed_8_0_705,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared call operator group (0) : call_stmt_690_call 
    writeEthernetHeaderToMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_690_call_req_0;
      call_stmt_690_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_690_call_req_1;
      call_stmt_690_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeEthernetHeaderToMem_call_group_0_gI: SplitGuardInterface generic map(name => "writeEthernetHeaderToMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer;
      new_buf_pointer_690 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeEthernetHeaderToMem_call_reqs(0),
          ackR => writeEthernetHeaderToMem_call_acks(0),
          dataR => writeEthernetHeaderToMem_call_data(35 downto 0),
          tagR => writeEthernetHeaderToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeEthernetHeaderToMem_return_acks(0), -- cross-over
          ackL => writeEthernetHeaderToMem_return_reqs(0), -- cross-over
          dataL => writeEthernetHeaderToMem_return_data(35 downto 0),
          tagL => writeEthernetHeaderToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_699_call 
    writePayloadToMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(16 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_699_call_req_0;
      call_stmt_699_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_699_call_req_1;
      call_stmt_699_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writePayloadToMem_call_group_1_gI: SplitGuardInterface generic map(name => "writePayloadToMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_684_delayed_4_0_693 & new_buf_pointer_690;
      packet_size_699 <= data_out(16 downto 9);
      bad_packet_identifier_buffer <= data_out(8 downto 8);
      last_keep_699 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writePayloadToMem_call_reqs(0),
          ackR => writePayloadToMem_call_acks(0),
          dataR => writePayloadToMem_call_data(71 downto 0),
          tagR => writePayloadToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 17,
          owidth => 17,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writePayloadToMem_return_acks(0), -- cross-over
          ackL => writePayloadToMem_return_reqs(0), -- cross-over
          dataL => writePayloadToMem_return_data(16 downto 0),
          tagL => writePayloadToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_710_call 
    writeControlInformationToMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(51 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_710_call_req_0;
      call_stmt_710_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_710_call_req_1;
      call_stmt_710_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not bad_packet_identifier_690_delayed_8_0_702(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeControlInformationToMem_call_group_2_gI: SplitGuardInterface generic map(name => "writeControlInformationToMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_691_delayed_8_0_705 & packet_size_699 & last_keep_699;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 52,
        owidth => 52,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeControlInformationToMem_call_reqs(0),
          ackR => writeControlInformationToMem_call_acks(0),
          dataR => writeControlInformationToMem_call_data(51 downto 0),
          tagR => writeControlInformationToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeControlInformationToMem_return_acks(0), -- cross-over
          ackL => writeControlInformationToMem_return_reqs(0), -- cross-over
          tagL => writeControlInformationToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end loadBuffer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nextLSTATE_Volatile is -- 
  port ( -- 
    RX : in  std_logic_vector(72 downto 0);
    LSTATE : in  std_logic_vector(1 downto 0);
    nLSTATE : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity nextLSTATE_Volatile;
architecture nextLSTATE_Volatile_arch of nextLSTATE_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal RX_buffer :  std_logic_vector(72 downto 0);
  signal LSTATE_buffer :  std_logic_vector(1 downto 0);
  -- output port buffer signals
  signal nLSTATE_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  RX_buffer <= RX;
  LSTATE_buffer <= LSTATE;
  -- output handling  -------------------------------------------------------
  nLSTATE <= nLSTATE_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1305_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1313_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1289_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1295_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1302_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1311_wire : std_logic_vector(0 downto 0);
    signal MUX_1292_wire : std_logic_vector(1 downto 0);
    signal MUX_1298_wire : std_logic_vector(1 downto 0);
    signal MUX_1308_wire : std_logic_vector(1 downto 0);
    signal MUX_1316_wire : std_logic_vector(1 downto 0);
    signal NOT_u1_u1_1304_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_1299_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_1317_wire : std_logic_vector(1 downto 0);
    signal R_S0_1288_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1314_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1290_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1294_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1296_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1301_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1306_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1310_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1283_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1291_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1297_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1307_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1315_wire_constant : std_logic_vector(1 downto 0);
    signal last_word_1285 : std_logic_vector(0 downto 0);
    signal tlast_1280 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_S0_1288_wire_constant <= "00";
    R_S0_1314_wire_constant <= "00";
    R_S1_1290_wire_constant <= "01";
    R_S1_1294_wire_constant <= "01";
    R_S2_1296_wire_constant <= "10";
    R_S2_1301_wire_constant <= "10";
    R_S2_1306_wire_constant <= "10";
    R_S2_1310_wire_constant <= "10";
    konst_1283_wire_constant <= "1";
    konst_1291_wire_constant <= "00";
    konst_1297_wire_constant <= "00";
    konst_1307_wire_constant <= "00";
    konst_1315_wire_constant <= "00";
    -- flow-through select operator MUX_1292_inst
    MUX_1292_wire <= R_S1_1290_wire_constant when (EQ_u2_u1_1289_wire(0) /=  '0') else konst_1291_wire_constant;
    -- flow-through select operator MUX_1298_inst
    MUX_1298_wire <= R_S2_1296_wire_constant when (EQ_u2_u1_1295_wire(0) /=  '0') else konst_1297_wire_constant;
    -- flow-through select operator MUX_1308_inst
    MUX_1308_wire <= R_S2_1306_wire_constant when (AND_u1_u1_1305_wire(0) /=  '0') else konst_1307_wire_constant;
    -- flow-through select operator MUX_1316_inst
    MUX_1316_wire <= R_S0_1314_wire_constant when (AND_u1_u1_1313_wire(0) /=  '0') else konst_1315_wire_constant;
    -- flow-through slice operator slice_1279_inst
    tlast_1280 <= RX_buffer(72 downto 72);
    -- binary operator AND_u1_u1_1305_inst
    process(EQ_u2_u1_1302_wire, NOT_u1_u1_1304_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1302_wire, NOT_u1_u1_1304_wire, tmp_var);
      AND_u1_u1_1305_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1313_inst
    process(EQ_u2_u1_1311_wire, last_word_1285) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1311_wire, last_word_1285, tmp_var);
      AND_u1_u1_1313_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1284_inst
    process(tlast_1280) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tlast_1280, konst_1283_wire_constant, tmp_var);
      last_word_1285 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1289_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S0_1288_wire_constant, tmp_var);
      EQ_u2_u1_1289_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1295_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S1_1294_wire_constant, tmp_var);
      EQ_u2_u1_1295_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1302_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1301_wire_constant, tmp_var);
      EQ_u2_u1_1302_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1311_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1310_wire_constant, tmp_var);
      EQ_u2_u1_1311_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1304_inst
    process(last_word_1285) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_word_1285, tmp_var);
      NOT_u1_u1_1304_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u2_u2_1299_inst
    process(MUX_1292_wire, MUX_1298_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1292_wire, MUX_1298_wire, tmp_var);
      OR_u2_u2_1299_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1317_inst
    process(MUX_1308_wire, MUX_1316_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1308_wire, MUX_1316_wire, tmp_var);
      OR_u2_u2_1317_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_1318_inst
    process(OR_u2_u2_1299_wire, OR_u2_u2_1317_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_1299_wire, OR_u2_u2_1317_wire, tmp_var);
      nLSTATE_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end nextLSTATE_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity nicRxFromMacDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
    nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicRxFromMacDaemon;
architecture nicRxFromMacDaemon_arch of nicRxFromMacDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicRxFromMacDaemon_CP_2517_start: Boolean;
  signal nicRxFromMacDaemon_CP_2517_symbol: Boolean;
  -- volatile/operator module components. 
  component nextLSTATE_Volatile is -- 
    port ( -- 
      RX : in  std_logic_vector(72 downto 0);
      LSTATE : in  std_logic_vector(1 downto 0);
      nLSTATE : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal WPIPE_nic_rx_to_packet_1371_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1371_inst_ack_1 : boolean;
  signal do_while_stmt_1333_branch_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1371_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1371_inst_req_1 : boolean;
  signal do_while_stmt_1333_branch_ack_1 : boolean;
  signal if_stmt_1325_branch_req_0 : boolean;
  signal if_stmt_1325_branch_ack_1 : boolean;
  signal if_stmt_1325_branch_ack_0 : boolean;
  signal do_while_stmt_1333_branch_req_0 : boolean;
  signal phi_stmt_1335_req_0 : boolean;
  signal phi_stmt_1335_req_1 : boolean;
  signal phi_stmt_1335_ack_0 : boolean;
  signal nLSTATE_1349_1337_buf_req_0 : boolean;
  signal nLSTATE_1349_1337_buf_ack_0 : boolean;
  signal nLSTATE_1349_1337_buf_req_1 : boolean;
  signal nLSTATE_1349_1337_buf_ack_1 : boolean;
  signal RPIPE_mac_to_nic_data_1341_inst_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_1341_inst_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_1341_inst_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_1341_inst_ack_1 : boolean;
  signal MUX_1369_inst_req_0 : boolean;
  signal MUX_1369_inst_ack_0 : boolean;
  signal MUX_1369_inst_req_1 : boolean;
  signal MUX_1369_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_1360_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_header_1360_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_header_1360_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_header_1360_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicRxFromMacDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicRxFromMacDaemon_CP_2517_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicRxFromMacDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2517_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2517_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2517_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicRxFromMacDaemon_CP_2517: Block -- control-path 
    signal nicRxFromMacDaemon_CP_2517_elements: BooleanArray(55 downto 0);
    -- 
  begin -- 
    nicRxFromMacDaemon_CP_2517_elements(0) <= nicRxFromMacDaemon_CP_2517_start;
    nicRxFromMacDaemon_CP_2517_symbol <= nicRxFromMacDaemon_CP_2517_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	55 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_1322/merge_stmt_1324_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1322/merge_stmt_1324__entry___PhiReq/$exit
      -- CP-element group 0: 	 branch_block_stmt_1322/merge_stmt_1324__entry___PhiReq/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1322/$entry
      -- CP-element group 0: 	 branch_block_stmt_1322/branch_block_stmt_1322__entry__
      -- CP-element group 0: 	 branch_block_stmt_1322/merge_stmt_1324__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1322/$exit
      -- CP-element group 1: 	 branch_block_stmt_1322/branch_block_stmt_1322__exit__
      -- 
    nicRxFromMacDaemon_CP_2517_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	54 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	55 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_1322/disable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/disable_loopback_PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_1322/do_while_stmt_1333__exit__
      -- CP-element group 2: 	 branch_block_stmt_1322/disable_loopback
      -- 
    nicRxFromMacDaemon_CP_2517_elements(2) <= nicRxFromMacDaemon_CP_2517_elements(54);
    -- CP-element group 3:  transition  place  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	55 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	55 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1322/not_enabled_yet_loopback_PhiReq/$exit
      -- CP-element group 3: 	 branch_block_stmt_1322/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 3: 	 branch_block_stmt_1322/if_stmt_1325_if_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_1322/if_stmt_1325_if_link/if_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_1322/not_enabled_yet_loopback
      -- 
    if_choice_transition_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1325_branch_ack_1, ack => nicRxFromMacDaemon_CP_2517_elements(3)); -- 
    -- CP-element group 4:  merge  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	55 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1322/if_stmt_1325__exit__
      -- CP-element group 4: 	 branch_block_stmt_1322/do_while_stmt_1333__entry__
      -- CP-element group 4: 	 branch_block_stmt_1322/if_stmt_1325_else_link/$exit
      -- CP-element group 4: 	 branch_block_stmt_1322/if_stmt_1325_else_link/else_choice_transition
      -- 
    else_choice_transition_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1325_branch_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(4)); -- 
    -- CP-element group 5:  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	11 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_1322/do_while_stmt_1333/$entry
      -- CP-element group 5: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333__entry__
      -- 
    nicRxFromMacDaemon_CP_2517_elements(5) <= nicRxFromMacDaemon_CP_2517_elements(4);
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	54 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333__exit__
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(6) is bound as output of CP function.
    -- CP-element group 7:  merge  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_back
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(7) is bound as output of CP function.
    -- CP-element group 8:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	52 
    -- CP-element group 8: 	53 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_exit/$entry
      -- CP-element group 8: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_taken/$entry
      -- CP-element group 8: 	 branch_block_stmt_1322/do_while_stmt_1333/condition_done
      -- 
    nicRxFromMacDaemon_CP_2517_elements(8) <= nicRxFromMacDaemon_CP_2517_elements(13);
    -- CP-element group 9:  branch  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	51 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_body_done
      -- 
    nicRxFromMacDaemon_CP_2517_elements(9) <= nicRxFromMacDaemon_CP_2517_elements(51);
    -- CP-element group 10:  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	22 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/back_edge_to_loop_body
      -- 
    nicRxFromMacDaemon_CP_2517_elements(10) <= nicRxFromMacDaemon_CP_2517_elements(7);
    -- CP-element group 11:  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	24 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/first_time_through_loop_body
      -- 
    nicRxFromMacDaemon_CP_2517_elements(11) <= nicRxFromMacDaemon_CP_2517_elements(5);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	50 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/$entry
      -- CP-element group 12: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/loop_body_start
      -- CP-element group 12: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1339_sample_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(12) is bound as output of CP function.
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: 	50 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	8 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/condition_evaluated
      -- 
    condition_evaluated_2612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(13), ack => do_while_stmt_1333_branch_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(17) & nicRxFromMacDaemon_CP_2517_elements(50);
      gj_nicRxFromMacDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	18 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/aggregated_phi_sample_req
      -- CP-element group 14: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_sample_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(12) & nicRxFromMacDaemon_CP_2517_elements(18) & nicRxFromMacDaemon_CP_2517_elements(17);
      gj_nicRxFromMacDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	51 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/aggregated_phi_sample_ack
      -- CP-element group 15: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1339_sample_completed_
      -- 
    nicRxFromMacDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(38) & nicRxFromMacDaemon_CP_2517_elements(20);
      gj_nicRxFromMacDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	35 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	37 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/aggregated_phi_update_req
      -- CP-element group 16: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_update_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(35) & nicRxFromMacDaemon_CP_2517_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	39 
    -- CP-element group 17: 	21 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/aggregated_phi_update_ack
      -- 
    nicRxFromMacDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(39) & nicRxFromMacDaemon_CP_2517_elements(21);
      gj_nicRxFromMacDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	12 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(12) & nicRxFromMacDaemon_CP_2517_elements(15);
      gj_nicRxFromMacDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	12 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	45 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(12) & nicRxFromMacDaemon_CP_2517_elements(42) & nicRxFromMacDaemon_CP_2517_elements(45);
      gj_nicRxFromMacDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	44 
    -- CP-element group 21: 	40 
    -- CP-element group 21: 	17 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_update_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	10 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_2517_elements(22) <= nicRxFromMacDaemon_CP_2517_elements(10);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_loopback_sample_req
      -- CP-element group 23: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_loopback_sample_req_ps
      -- 
    phi_stmt_1335_loopback_sample_req_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1335_loopback_sample_req_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(23), ack => phi_stmt_1335_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	11 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_2517_elements(24) <= nicRxFromMacDaemon_CP_2517_elements(11);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_entry_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_entry_sample_req_ps
      -- 
    phi_stmt_1335_entry_sample_req_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1335_entry_sample_req_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(25), ack => phi_stmt_1335_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_phi_mux_ack
      -- CP-element group 26: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1335_phi_mux_ack_ps
      -- 
    phi_stmt_1335_phi_mux_ack_2633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1335_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_sample_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Sample/req
      -- 
    req_2646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(27), ack => nLSTATE_1349_1337_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_update_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Update/req
      -- 
    req_2651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(28), ack => nLSTATE_1349_1337_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Sample/ack
      -- 
    ack_2647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1349_1337_buf_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(29)); -- 
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_nLSTATE_1337_Update/ack
      -- 
    ack_2652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1349_1337_buf_ack_1, ack => nicRxFromMacDaemon_CP_2517_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_sample_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_update_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_2517_elements(33) <= nicRxFromMacDaemon_CP_2517_elements(34);
    -- CP-element group 34:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	33 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/R_S0_1338_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(34) is a control-delay.
    cp_element_34_delay: control_delay_element  generic map(name => " 34_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2517_elements(32), ack => nicRxFromMacDaemon_CP_2517_elements(34), clk => clk, reset =>reset);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	42 
    -- CP-element group 35: 	48 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	16 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1339_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(12) & nicRxFromMacDaemon_CP_2517_elements(42) & nicRxFromMacDaemon_CP_2517_elements(48);
      gj_nicRxFromMacDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	39 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Sample/rr
      -- 
    rr_2673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(36), ack => RPIPE_mac_to_nic_data_1341_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(14) & nicRxFromMacDaemon_CP_2517_elements(39);
      gj_nicRxFromMacDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	16 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Update/cr
      -- 
    cr_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(37), ack => RPIPE_mac_to_nic_data_1341_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(38) & nicRxFromMacDaemon_CP_2517_elements(16);
      gj_nicRxFromMacDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	15 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Sample/ra
      -- 
    ra_2674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1341_inst_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	47 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	17 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	36 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/phi_stmt_1339_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/RPIPE_mac_to_nic_data_1341_Update/ca
      -- 
    ca_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1341_inst_ack_1, ack => nicRxFromMacDaemon_CP_2517_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: 	21 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_start/$entry
      -- CP-element group 40: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_start/req
      -- 
    req_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(40), ack => MUX_1369_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(39) & nicRxFromMacDaemon_CP_2517_elements(21) & nicRxFromMacDaemon_CP_2517_elements(42);
      gj_nicRxFromMacDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	45 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_update_start_
      -- CP-element group 41: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_complete/$entry
      -- CP-element group 41: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_complete/req
      -- 
    req_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(41), ack => MUX_1369_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicRxFromMacDaemon_CP_2517_elements(45);
      gj_nicRxFromMacDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	35 
    -- CP-element group 42: 	40 
    -- CP-element group 42: 	19 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_start/ack
      -- 
    ack_2688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1369_inst_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/MUX_1369_complete/ack
      -- 
    ack_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1369_inst_ack_1, ack => nicRxFromMacDaemon_CP_2517_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	21 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Sample/req
      -- 
    req_2701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(44), ack => WPIPE_nic_rx_to_header_1360_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(43) & nicRxFromMacDaemon_CP_2517_elements(21) & nicRxFromMacDaemon_CP_2517_elements(46);
      gj_nicRxFromMacDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	41 
    -- CP-element group 45: 	19 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Update/req
      -- 
    ack_2702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1360_inst_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(45)); -- 
    req_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(45), ack => WPIPE_nic_rx_to_header_1360_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	51 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_header_1360_Update/ack
      -- 
    ack_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1360_inst_ack_1, ack => nicRxFromMacDaemon_CP_2517_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	39 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_sample_start_
      -- 
    req_2715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(47), ack => WPIPE_nic_rx_to_packet_1371_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(39) & nicRxFromMacDaemon_CP_2517_elements(49);
      gj_nicRxFromMacDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	35 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Update/req
      -- CP-element group 48: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_sample_completed_
      -- 
    ack_2716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1371_inst_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(48)); -- 
    req_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(48), ack => WPIPE_nic_rx_to_packet_1371_inst_req_1); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/WPIPE_nic_rx_to_packet_1371_Update/$exit
      -- 
    ack_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1371_inst_ack_1, ack => nicRxFromMacDaemon_CP_2517_elements(49)); -- 
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	12 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	13 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_2517_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2517_elements(12), ack => nicRxFromMacDaemon_CP_2517_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	46 
    -- CP-element group 51: 	15 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	9 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1322/do_while_stmt_1333/do_while_stmt_1333_loop_body/$exit
      -- 
    nicRxFromMacDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2517_elements(46) & nicRxFromMacDaemon_CP_2517_elements(15) & nicRxFromMacDaemon_CP_2517_elements(49);
      gj_nicRxFromMacDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	8 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (2) 
      -- CP-element group 52: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_exit/ack
      -- CP-element group 52: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_exit/$exit
      -- 
    ack_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1333_branch_ack_0, ack => nicRxFromMacDaemon_CP_2517_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	8 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_taken/$exit
      -- CP-element group 53: 	 branch_block_stmt_1322/do_while_stmt_1333/loop_taken/ack
      -- 
    ack_2730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1333_branch_ack_1, ack => nicRxFromMacDaemon_CP_2517_elements(53)); -- 
    -- CP-element group 54:  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	6 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	2 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1322/do_while_stmt_1333/$exit
      -- 
    nicRxFromMacDaemon_CP_2517_elements(54) <= nicRxFromMacDaemon_CP_2517_elements(6);
    -- CP-element group 55:  merge  branch  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	2 
    -- CP-element group 55: 	0 
    -- CP-element group 55: 	3 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	3 
    -- CP-element group 55: 	4 
    -- CP-element group 55:  members (49) 
      -- CP-element group 55: 	 branch_block_stmt_1322/merge_stmt_1324_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/merge_stmt_1324_PhiAck/dummy
      -- CP-element group 55: 	 branch_block_stmt_1322/merge_stmt_1324_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/merge_stmt_1324_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_1322/merge_stmt_1324__exit__
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325__entry__
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Sample/req
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Update/req
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/BITSEL_u32_u1_1328_inputs/RPIPE_CONTROL_REGISTER_1326/Update/ack
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/BITSEL_u32_u1_1328/SplitProtocol/Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/NOT_u1_u1_1329/SplitProtocol/Update/ca
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_1322/NOT_u1_u1_1329_place
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_1322/if_stmt_1325_else_link/$entry
      -- 
    branch_req_2587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2517_elements(55), ack => if_stmt_1325_branch_req_0); -- 
    nicRxFromMacDaemon_CP_2517_elements(55) <= OrReduce(nicRxFromMacDaemon_CP_2517_elements(2) & nicRxFromMacDaemon_CP_2517_elements(0) & nicRxFromMacDaemon_CP_2517_elements(3));
    nicRxFromMacDaemon_do_while_stmt_1333_terminator_2731: loop_terminator -- 
      generic map (name => " nicRxFromMacDaemon_do_while_stmt_1333_terminator_2731", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicRxFromMacDaemon_CP_2517_elements(9),loop_continue => nicRxFromMacDaemon_CP_2517_elements(53),loop_terminate => nicRxFromMacDaemon_CP_2517_elements(52),loop_back => nicRxFromMacDaemon_CP_2517_elements(7),loop_exit => nicRxFromMacDaemon_CP_2517_elements(6),clk => clk, reset => reset); -- 
    phi_stmt_1335_phi_seq_2661_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_2517_elements(22);
      nicRxFromMacDaemon_CP_2517_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_2517_elements(29);
      nicRxFromMacDaemon_CP_2517_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_2517_elements(30);
      nicRxFromMacDaemon_CP_2517_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_2517_elements(24);
      nicRxFromMacDaemon_CP_2517_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_2517_elements(31);
      nicRxFromMacDaemon_CP_2517_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_2517_elements(33);
      nicRxFromMacDaemon_CP_2517_elements(25) <= phi_mux_reqs(1);
      phi_stmt_1335_phi_seq_2661 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1335_phi_seq_2661") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_2517_elements(14), 
          phi_sample_ack => nicRxFromMacDaemon_CP_2517_elements(20), 
          phi_update_req => nicRxFromMacDaemon_CP_2517_elements(16), 
          phi_update_ack => nicRxFromMacDaemon_CP_2517_elements(21), 
          phi_mux_ack => nicRxFromMacDaemon_CP_2517_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2613_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicRxFromMacDaemon_CP_2517_elements(10);
        preds(1)  <= nicRxFromMacDaemon_CP_2517_elements(11);
        entry_tmerge_2613 : transition_merge -- 
          generic map(name => " entry_tmerge_2613")
          port map (preds => preds, symbol_out => nicRxFromMacDaemon_CP_2517_elements(12));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1328_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1380_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u65_u73_1367_wire : std_logic_vector(72 downto 0);
    signal EQ_u2_u1_1353_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1356_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1363_wire : std_logic_vector(0 downto 0);
    signal LSTATE_1335 : std_logic_vector(1 downto 0);
    signal MUX_1369_wire : std_logic_vector(72 downto 0);
    signal NOT_u1_u1_1329_wire : std_logic_vector(0 downto 0);
    signal RPIPE_CONTROL_REGISTER_1326_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1378_wire : std_logic_vector(31 downto 0);
    signal RPIPE_mac_to_nic_data_1341_wire : std_logic_vector(72 downto 0);
    signal RX_1339 : std_logic_vector(72 downto 0);
    signal R_HEADER_TKEEP_1366_wire_constant : std_logic_vector(7 downto 0);
    signal R_S0_1338_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1352_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1355_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1362_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1327_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1379_wire_constant : std_logic_vector(31 downto 0);
    signal nLSTATE_1349 : std_logic_vector(1 downto 0);
    signal nLSTATE_1349_1337_buffered : std_logic_vector(1 downto 0);
    signal slice_1365_wire : std_logic_vector(64 downto 0);
    signal write_to_header_1358 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_HEADER_TKEEP_1366_wire_constant <= "00111111";
    R_S0_1338_wire_constant <= "00";
    R_S0_1352_wire_constant <= "00";
    R_S1_1355_wire_constant <= "01";
    R_S1_1362_wire_constant <= "01";
    konst_1327_wire_constant <= "00000000000000000000000000000000";
    konst_1379_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_1335: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nLSTATE_1349_1337_buffered & R_S0_1338_wire_constant;
      req <= phi_stmt_1335_req_0 & phi_stmt_1335_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1335",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1335_ack_0,
          idata => idata,
          odata => LSTATE_1335,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1335
    MUX_1369_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= MUX_1369_inst_req_0;
      MUX_1369_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= MUX_1369_inst_req_1;
      MUX_1369_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  write_to_header_1358(0);
      MUX_1369_inst_gI: SplitGuardInterface generic map(name => "MUX_1369_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      MUX_1369_inst: SelectSplitProtocol generic map(name => "MUX_1369_inst", data_width => 73, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u65_u73_1367_wire, y => RX_1339, sel => EQ_u2_u1_1363_wire, z => MUX_1369_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_1365_inst
    slice_1365_wire <= RX_1339(72 downto 8);
    nLSTATE_1349_1337_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nLSTATE_1349_1337_buf_req_0;
      nLSTATE_1349_1337_buf_ack_0<= wack(0);
      rreq(0) <= nLSTATE_1349_1337_buf_req_1;
      nLSTATE_1349_1337_buf_ack_1<= rack(0);
      nLSTATE_1349_1337_buf : InterlockBuffer generic map ( -- 
        name => "nLSTATE_1349_1337_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nLSTATE_1349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nLSTATE_1349_1337_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1339
    process(RPIPE_mac_to_nic_data_1341_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_mac_to_nic_data_1341_wire(72 downto 0);
      RX_1339 <= tmp_var; -- 
    end process;
    do_while_stmt_1333_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1380_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1333_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1333_branch_req_0,
          ack0 => do_while_stmt_1333_branch_ack_0,
          ack1 => do_while_stmt_1333_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1325_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1329_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1325_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1325_branch_req_0,
          ack0 => if_stmt_1325_branch_ack_0,
          ack1 => if_stmt_1325_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator BITSEL_u32_u1_1328_inst
    process(RPIPE_CONTROL_REGISTER_1326_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1326_wire, konst_1327_wire_constant, tmp_var);
      BITSEL_u32_u1_1328_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1380_inst
    process(RPIPE_CONTROL_REGISTER_1378_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1378_wire, konst_1379_wire_constant, tmp_var);
      BITSEL_u32_u1_1380_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u65_u73_1367_inst
    process(slice_1365_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1365_wire, R_HEADER_TKEEP_1366_wire_constant, tmp_var);
      CONCAT_u65_u73_1367_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1353_inst
    process(LSTATE_1335) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1335, R_S0_1352_wire_constant, tmp_var);
      EQ_u2_u1_1353_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1356_inst
    process(LSTATE_1335) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1335, R_S1_1355_wire_constant, tmp_var);
      EQ_u2_u1_1356_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1363_inst
    process(LSTATE_1335) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1335, R_S1_1362_wire_constant, tmp_var);
      EQ_u2_u1_1363_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1329_inst
    process(BITSEL_u32_u1_1328_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1328_wire, tmp_var);
      NOT_u1_u1_1329_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1357_inst
    process(EQ_u2_u1_1353_wire, EQ_u2_u1_1356_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_1353_wire, EQ_u2_u1_1356_wire, tmp_var);
      write_to_header_1358 <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1326_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1378_wire <= CONTROL_REGISTER;
    -- shared inport operator group (2) : RPIPE_mac_to_nic_data_1341_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_1341_inst_req_0;
      RPIPE_mac_to_nic_data_1341_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_1341_inst_req_1;
      RPIPE_mac_to_nic_data_1341_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_1341_wire <= data_out(72 downto 0);
      mac_to_nic_data_read_2_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_read_2: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_read_2", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_pipe_read_req(0),
          oack => mac_to_nic_data_pipe_read_ack(0),
          odata => mac_to_nic_data_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_nic_rx_to_header_1360_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_header_1360_inst_req_0;
      WPIPE_nic_rx_to_header_1360_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_header_1360_inst_req_1;
      WPIPE_nic_rx_to_header_1360_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_to_header_1358(0);
      data_in <= MUX_1369_wire;
      nic_rx_to_header_write_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_write_0: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_header", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_header_pipe_write_req(0),
          oack => nic_rx_to_header_pipe_write_ack(0),
          odata => nic_rx_to_header_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_rx_to_packet_1371_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1371_inst_req_0;
      WPIPE_nic_rx_to_packet_1371_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1371_inst_req_1;
      WPIPE_nic_rx_to_packet_1371_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= RX_1339;
      nic_rx_to_packet_write_1_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_write_1: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_packet", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_packet_pipe_write_req(0),
          oack => nic_rx_to_packet_pipe_write_ack(0),
          odata => nic_rx_to_packet_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    volatile_operator_nextLSTATE_3791: nextLSTATE_Volatile port map(RX => RX_1339, LSTATE => LSTATE_1335, nLSTATE => nLSTATE_1349); 
    -- 
  end Block; -- data_path
  -- 
end nicRxFromMacDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity popFromQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_call_data : out  std_logic_vector(35 downto 0);
    releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_call_data : out  std_logic_vector(67 downto 0);
    getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_return_data : in   std_logic_vector(31 downto 0);
    getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_call_data : out  std_logic_vector(35 downto 0);
    acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_return_data : in   std_logic_vector(0 downto 0);
    acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity popFromQueue;
architecture popFromQueue_arch of popFromQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 37)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal popFromQueue_CP_585_start: Boolean;
  signal popFromQueue_CP_585_symbol: Boolean;
  -- volatile/operator module components. 
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_pointer : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_511_call_req_1 : boolean;
  signal call_stmt_511_call_ack_1 : boolean;
  signal call_stmt_486_call_req_1 : boolean;
  signal call_stmt_486_call_ack_1 : boolean;
  signal call_stmt_486_call_req_0 : boolean;
  signal call_stmt_486_call_ack_0 : boolean;
  signal call_stmt_481_call_req_1 : boolean;
  signal call_stmt_481_call_ack_1 : boolean;
  signal call_stmt_527_call_req_0 : boolean;
  signal call_stmt_527_call_ack_0 : boolean;
  signal call_stmt_527_call_req_1 : boolean;
  signal call_stmt_527_call_ack_1 : boolean;
  signal call_stmt_516_call_req_1 : boolean;
  signal call_stmt_481_call_ack_0 : boolean;
  signal call_stmt_481_call_req_0 : boolean;
  signal call_stmt_511_call_req_0 : boolean;
  signal call_stmt_511_call_ack_0 : boolean;
  signal W_status_528_inst_req_0 : boolean;
  signal W_status_528_inst_ack_0 : boolean;
  signal W_status_528_inst_req_1 : boolean;
  signal W_status_528_inst_ack_1 : boolean;
  signal call_stmt_516_call_req_0 : boolean;
  signal call_stmt_516_call_ack_0 : boolean;
  signal call_stmt_516_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "popFromQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 37) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(tag_length + 36 downto 37) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 36 downto 37);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  popFromQueue_CP_585_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "popFromQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_585_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= popFromQueue_CP_585_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_585_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  popFromQueue_CP_585: Block -- control-path 
    signal popFromQueue_CP_585_elements: BooleanArray(14 downto 0);
    -- 
  begin -- 
    popFromQueue_CP_585_elements(0) <= popFromQueue_CP_585_start;
    popFromQueue_CP_585_symbol <= popFromQueue_CP_585_elements(14);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_481/$entry
      -- CP-element group 0: 	 call_stmt_481/call_stmt_481_sample_start_
      -- CP-element group 0: 	 call_stmt_481/call_stmt_481_Update/ccr
      -- CP-element group 0: 	 call_stmt_481/call_stmt_481_Update/$entry
      -- CP-element group 0: 	 call_stmt_481/call_stmt_481_update_start_
      -- CP-element group 0: 	 call_stmt_481/call_stmt_481_Sample/$entry
      -- CP-element group 0: 	 call_stmt_481/call_stmt_481_Sample/crr
      -- CP-element group 0: 	 $entry
      -- 
    crr_598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(0), ack => call_stmt_481_call_req_0); -- 
    ccr_603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(0), ack => call_stmt_481_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_481/call_stmt_481_sample_completed_
      -- CP-element group 1: 	 call_stmt_481/call_stmt_481_Sample/cra
      -- CP-element group 1: 	 call_stmt_481/call_stmt_481_Sample/$exit
      -- 
    cra_599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_481_call_ack_0, ack => popFromQueue_CP_585_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (17) 
      -- CP-element group 2: 	 call_stmt_481/call_stmt_481_update_completed_
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Update/ccr
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Update/$entry
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Update/ccr
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Update/$entry
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Sample/crr
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Sample/$entry
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_update_start_
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_sample_start_
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/$entry
      -- CP-element group 2: 	 call_stmt_481/call_stmt_481_Update/cca
      -- CP-element group 2: 	 call_stmt_481/call_stmt_481_Update/$exit
      -- CP-element group 2: 	 call_stmt_481/$exit
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_update_start_
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Update/$entry
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Update/ccr
      -- CP-element group 2: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_update_start_
      -- 
    cca_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_481_call_ack_1, ack => popFromQueue_CP_585_elements(2)); -- 
    ccr_634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(2), ack => call_stmt_511_call_req_1); -- 
    ccr_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(2), ack => call_stmt_486_call_req_1); -- 
    crr_615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(2), ack => call_stmt_486_call_req_0); -- 
    ccr_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(2), ack => call_stmt_516_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Sample/cra
      -- CP-element group 3: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Sample/$exit
      -- CP-element group 3: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_sample_completed_
      -- 
    cra_616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_486_call_ack_0, ack => popFromQueue_CP_585_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Sample/$entry
      -- CP-element group 4: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Update/cca
      -- CP-element group 4: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_Update/$exit
      -- CP-element group 4: 	 call_stmt_486_to_call_stmt_516/call_stmt_486_update_completed_
      -- CP-element group 4: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_sample_start_
      -- CP-element group 4: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Sample/crr
      -- 
    cca_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_486_call_ack_1, ack => popFromQueue_CP_585_elements(4)); -- 
    crr_629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(4), ack => call_stmt_511_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Sample/$exit
      -- CP-element group 5: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_sample_completed_
      -- CP-element group 5: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Sample/cra
      -- 
    cra_630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_511_call_ack_0, ack => popFromQueue_CP_585_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Update/cca
      -- CP-element group 6: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_Update/$exit
      -- CP-element group 6: 	 call_stmt_486_to_call_stmt_516/call_stmt_511_update_completed_
      -- 
    cca_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_511_call_ack_1, ack => popFromQueue_CP_585_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Sample/crr
      -- CP-element group 7: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Sample/$entry
      -- CP-element group 7: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_sample_start_
      -- 
    crr_643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(7), ack => call_stmt_516_call_req_0); -- 
    popFromQueue_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "popFromQueue_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_585_elements(4) & popFromQueue_CP_585_elements(6);
      gj_popFromQueue_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_585_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Sample/cra
      -- CP-element group 8: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Sample/$exit
      -- CP-element group 8: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_sample_completed_
      -- 
    cra_644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_516_call_ack_0, ack => popFromQueue_CP_585_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (17) 
      -- CP-element group 9: 	 call_stmt_486_to_call_stmt_516/$exit
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Sample/$entry
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Sample/crr
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Update/$entry
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Update/ccr
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_sample_start_
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_update_start_
      -- CP-element group 9: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_update_completed_
      -- CP-element group 9: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Update/$exit
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/$entry
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Sample/$entry
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Sample/req
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Update/$entry
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Update/req
      -- CP-element group 9: 	 call_stmt_486_to_call_stmt_516/call_stmt_516_Update/cca
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_sample_start_
      -- CP-element group 9: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_update_start_
      -- 
    cca_649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_516_call_ack_1, ack => popFromQueue_CP_585_elements(9)); -- 
    ccr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(9), ack => call_stmt_527_call_req_1); -- 
    crr_660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(9), ack => call_stmt_527_call_req_0); -- 
    req_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(9), ack => W_status_528_inst_req_0); -- 
    req_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_585_elements(9), ack => W_status_528_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Sample/$exit
      -- CP-element group 10: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Sample/cra
      -- CP-element group 10: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_sample_completed_
      -- 
    cra_661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_527_call_ack_0, ack => popFromQueue_CP_585_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Update/$exit
      -- CP-element group 11: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_Update/cca
      -- CP-element group 11: 	 call_stmt_527_to_assign_stmt_530/call_stmt_527_update_completed_
      -- 
    cca_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_527_call_ack_1, ack => popFromQueue_CP_585_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_sample_completed_
      -- CP-element group 12: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Sample/$exit
      -- CP-element group 12: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Sample/ack
      -- 
    ack_675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_528_inst_ack_0, ack => popFromQueue_CP_585_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_update_completed_
      -- CP-element group 13: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Update/$exit
      -- CP-element group 13: 	 call_stmt_527_to_assign_stmt_530/assign_stmt_530_Update/ack
      -- 
    ack_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_528_inst_ack_1, ack => popFromQueue_CP_585_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 $exit
      -- CP-element group 14: 	 call_stmt_527_to_assign_stmt_530/$exit
      -- 
    popFromQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_585_elements(11) & popFromQueue_CP_585_elements(13);
      gj_popFromQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_585_elements(14), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_504_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_496_wire_constant : std_logic_vector(31 downto 0);
    signal konst_501_wire_constant : std_logic_vector(31 downto 0);
    signal konst_503_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_481 : std_logic_vector(0 downto 0);
    signal next_rp_506 : std_logic_vector(31 downto 0);
    signal q_empty_491 : std_logic_vector(0 downto 0);
    signal read_pointer_486 : std_logic_vector(31 downto 0);
    signal round_off_498 : std_logic_vector(0 downto 0);
    signal write_pointer_486 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    SUB_u32_u32_496_wire_constant <= "00000000000000000000000000000111";
    konst_501_wire_constant <= "00000000000000000000000000000000";
    konst_503_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_505_inst
    next_rp_506 <= konst_501_wire_constant when (round_off_498(0) /=  '0') else ADD_u32_u32_504_wire;
    W_status_528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_528_inst_req_0;
      W_status_528_inst_ack_0<= wack(0);
      rreq(0) <= W_status_528_inst_req_1;
      W_status_528_inst_ack_1<= rack(0);
      W_status_528_inst : InterlockBuffer generic map ( -- 
        name => "W_status_528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_empty_491,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator ADD_u32_u32_504_inst
    process(read_pointer_486) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(read_pointer_486, konst_503_wire_constant, tmp_var);
      ADD_u32_u32_504_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_490_inst
    process(write_pointer_486, read_pointer_486) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_pointer_486, read_pointer_486, tmp_var);
      q_empty_491 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_497_inst
    process(read_pointer_486) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(read_pointer_486, SUB_u32_u32_496_wire_constant, tmp_var);
      round_off_498 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_481_call 
    acquireMutex_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_481_call_req_0;
      call_stmt_481_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_481_call_req_1;
      call_stmt_481_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireMutex_call_group_0_gI: SplitGuardInterface generic map(name => "acquireMutex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_481 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireMutex_call_reqs(0),
          ackR => acquireMutex_call_acks(0),
          dataR => acquireMutex_call_data(35 downto 0),
          tagR => acquireMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireMutex_return_acks(0), -- cross-over
          ackL => acquireMutex_return_reqs(0), -- cross-over
          dataL => acquireMutex_return_data(0 downto 0),
          tagL => acquireMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_486_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_486_call_req_0;
      call_stmt_486_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_486_call_req_1;
      call_stmt_486_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_pointer_486 <= data_out(63 downto 32);
      read_pointer_486 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_511_call 
    getQueueElement_call_group_2: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_511_call_req_0;
      call_stmt_511_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_511_call_req_1;
      call_stmt_511_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_491(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueElement_call_group_2_gI: SplitGuardInterface generic map(name => "getQueueElement_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & read_pointer_486;
      q_r_data_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueElement_call_reqs(0),
          ackR => getQueueElement_call_acks(0),
          dataR => getQueueElement_call_data(67 downto 0),
          tagR => getQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueElement_return_acks(0), -- cross-over
          ackL => getQueueElement_return_reqs(0), -- cross-over
          dataL => getQueueElement_return_data(31 downto 0),
          tagL => getQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_516_call 
    setQueuePointers_call_group_3: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_516_call_req_0;
      call_stmt_516_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_516_call_req_1;
      call_stmt_516_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_491(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_3_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_pointer_486 & next_rp_506;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_527_call 
    releaseMutex_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_527_call_req_0;
      call_stmt_527_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_527_call_req_1;
      call_stmt_527_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseMutex_call_group_4_gI: SplitGuardInterface generic map(name => "releaseMutex_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseMutex_call_reqs(0),
          ackR => releaseMutex_call_acks(0),
          dataR => releaseMutex_call_data(35 downto 0),
          tagR => releaseMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseMutex_return_acks(0), -- cross-over
          ackL => releaseMutex_return_reqs(0), -- cross-over
          tagL => releaseMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end popFromQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity populateRxQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity populateRxQueue;
architecture populateRxQueue_arch of populateRxQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal populateRxQueue_CP_1311_start: Boolean;
  signal populateRxQueue_CP_1311_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component delay_time_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      T : in  std_logic_vector(31 downto 0);
      delay_done : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal if_stmt_940_branch_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_req_1 : boolean;
  signal if_stmt_940_branch_req_0 : boolean;
  signal AND_u6_u6_929_inst_ack_0 : boolean;
  signal n_q_index_930_882_buf_ack_0 : boolean;
  signal call_stmt_939_call_req_0 : boolean;
  signal call_stmt_903_call_req_0 : boolean;
  signal if_stmt_940_branch_ack_1 : boolean;
  signal if_stmt_934_branch_ack_0 : boolean;
  signal call_stmt_920_call_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_ack_0 : boolean;
  signal n_q_index_930_882_buf_req_1 : boolean;
  signal n_q_index_930_882_buf_ack_1 : boolean;
  signal AND_u6_u6_881_inst_req_0 : boolean;
  signal AND_u6_u6_881_inst_ack_0 : boolean;
  signal call_stmt_903_call_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_req_0 : boolean;
  signal call_stmt_903_call_req_1 : boolean;
  signal AND_u6_u6_929_inst_req_0 : boolean;
  signal AND_u6_u6_881_inst_req_1 : boolean;
  signal phi_stmt_872_ack_0 : boolean;
  signal AND_u6_u6_881_inst_ack_1 : boolean;
  signal phi_stmt_872_req_0 : boolean;
  signal call_stmt_939_call_ack_0 : boolean;
  signal n_q_index_930_882_buf_req_0 : boolean;
  signal call_stmt_903_call_ack_1 : boolean;
  signal if_stmt_934_branch_req_0 : boolean;
  signal if_stmt_934_branch_ack_1 : boolean;
  signal call_stmt_920_call_req_1 : boolean;
  signal phi_stmt_872_req_1 : boolean;
  signal AND_u6_u6_929_inst_ack_1 : boolean;
  signal AND_u6_u6_929_inst_req_1 : boolean;
  signal call_stmt_920_call_ack_0 : boolean;
  signal call_stmt_939_call_ack_1 : boolean;
  signal call_stmt_920_call_req_0 : boolean;
  signal call_stmt_939_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "populateRxQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  populateRxQueue_CP_1311_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "populateRxQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1311_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= populateRxQueue_CP_1311_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1311_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  populateRxQueue_CP_1311: Block -- control-path 
    signal populateRxQueue_CP_1311_elements: BooleanArray(25 downto 0);
    -- 
  begin -- 
    populateRxQueue_CP_1311_elements(0) <= populateRxQueue_CP_1311_start;
    populateRxQueue_CP_1311_symbol <= populateRxQueue_CP_1311_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	17 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 branch_block_stmt_870/merge_stmt_871_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_870/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_870/merge_stmt_871__entry__
      -- CP-element group 0: 	 branch_block_stmt_870/branch_block_stmt_870__entry__
      -- 
    -- CP-element group 1:  merge  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	16 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_870/if_stmt_934__exit__
      -- CP-element group 1: 	 branch_block_stmt_870/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_870/branch_block_stmt_870__exit__
      -- 
    populateRxQueue_CP_1311_elements(1) <= OrReduce(populateRxQueue_CP_1311_elements(14) & populateRxQueue_CP_1311_elements(16));
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	25 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Sample/cra
      -- CP-element group 2: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_sample_completed_
      -- 
    cra_1336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_903_call_ack_0, ack => populateRxQueue_CP_1311_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	25 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Sample/crr
      -- 
    cca_1341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_903_call_ack_1, ack => populateRxQueue_CP_1311_elements(3)); -- 
    crr_1349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(3), ack => call_stmt_920_call_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Sample/cra
      -- CP-element group 4: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Sample/$exit
      -- 
    cra_1350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_920_call_ack_0, ack => populateRxQueue_CP_1311_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Update/cca
      -- CP-element group 5: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Update/$exit
      -- 
    cca_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_920_call_ack_1, ack => populateRxQueue_CP_1311_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	25 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Sample/$exit
      -- 
    ra_1364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_929_inst_ack_0, ack => populateRxQueue_CP_1311_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	25 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Update/$exit
      -- 
    ca_1369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_929_inst_ack_1, ack => populateRxQueue_CP_1311_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (22) 
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_else_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/$exit
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/NOT_u1_u1_936_place
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/branch_req
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_eval_test/NOT_u1_u1_936/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/$exit
      -- CP-element group 8: 	 branch_block_stmt_870/if_stmt_934__entry__
      -- CP-element group 8: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930__exit__
      -- 
    branch_req_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(8), ack => if_stmt_934_branch_req_0); -- 
    populateRxQueue_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "populateRxQueue_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1311_elements(5) & populateRxQueue_CP_1311_elements(7);
      gj_populateRxQueue_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1311_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_870/if_stmt_934_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939__entry__
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_update_start_
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Sample/crr
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939/$entry
      -- CP-element group 9: 	 branch_block_stmt_870/if_stmt_934_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Update/ccr
      -- CP-element group 9: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Update/$entry
      -- 
    if_choice_transition_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_934_branch_ack_1, ack => populateRxQueue_CP_1311_elements(9)); -- 
    crr_1417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(9), ack => call_stmt_939_call_req_0); -- 
    ccr_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(9), ack => call_stmt_939_call_req_1); -- 
    -- CP-element group 10:  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_870/assign_stmt_949/$entry
      -- CP-element group 10: 	 branch_block_stmt_870/if_stmt_934_else_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_870/if_stmt_934_else_link/else_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Sample/req
      -- CP-element group 10: 	 branch_block_stmt_870/assign_stmt_949__entry__
      -- 
    else_choice_transition_1402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_934_branch_ack_0, ack => populateRxQueue_CP_1311_elements(10)); -- 
    req_1473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(10), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Sample/cra
      -- 
    cra_1418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_939_call_ack_0, ack => populateRxQueue_CP_1311_elements(11)); -- 
    -- CP-element group 12:  branch  transition  place  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (27) 
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/EQ_u1_u1_943_inputs/$exit
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/$exit
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/$exit
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940__entry__
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_else_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Update/cr
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/SplitProtocol/Update/ca
      -- CP-element group 12: 	 branch_block_stmt_870/EQ_u1_u1_943_place
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/EQ_u1_u1_943_inputs/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/if_stmt_940_eval_test/EQ_u1_u1_943/$entry
      -- CP-element group 12: 	 branch_block_stmt_870/call_stmt_939__exit__
      -- CP-element group 12: 	 branch_block_stmt_870/call_stmt_939/$exit
      -- CP-element group 12: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Update/cca
      -- CP-element group 12: 	 branch_block_stmt_870/call_stmt_939/call_stmt_939_Update/$exit
      -- 
    cca_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_939_call_ack_1, ack => populateRxQueue_CP_1311_elements(12)); -- 
    branch_req_1450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(12), ack => if_stmt_940_branch_req_0); -- 
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	21 
    -- CP-element group 13: 	22 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_870/if_stmt_940_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_870/if_stmt_940_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Update/req
      -- CP-element group 13: 	 branch_block_stmt_870/loopback
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Sample/req
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/$entry
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/$entry
      -- 
    if_choice_transition_1455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_940_branch_ack_1, ack => populateRxQueue_CP_1311_elements(13)); -- 
    req_1613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(13), ack => n_q_index_930_882_buf_req_1); -- 
    req_1608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(13), ack => n_q_index_930_882_buf_req_0); -- 
    -- CP-element group 14:  merge  transition  place  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	1 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_870/if_stmt_940_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_870/if_stmt_940__exit__
      -- CP-element group 14: 	 branch_block_stmt_870/if_stmt_940_else_link/$exit
      -- 
    else_choice_transition_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_940_branch_ack_0, ack => populateRxQueue_CP_1311_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Update/req
      -- CP-element group 15: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_update_start_
      -- CP-element group 15: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Sample/ack
      -- 
    ack_1474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_ack_0, ack => populateRxQueue_CP_1311_elements(15)); -- 
    req_1478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(15), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_req_1); -- 
    -- CP-element group 16:  transition  place  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	1 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Update/ack
      -- CP-element group 16: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_870/assign_stmt_949/$exit
      -- CP-element group 16: 	 branch_block_stmt_870/assign_stmt_949/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_870/assign_stmt_949__exit__
      -- 
    ack_1479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_ack_1, ack => populateRxQueue_CP_1311_elements(16)); -- 
    -- CP-element group 17:  join  fork  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (71) 
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Update/req
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/RPIPE_NUMBER_OF_SERVERS_877/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SUB_u32_u32_879_inputs/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Sample/req
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Update/ca
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Update/cr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/SplitProtocol/$entry
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Update/ack
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/type_cast_880/SUB_u32_u32_879/SplitProtocol/Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Update/req
      -- CP-element group 17: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/AND_u6_u6_881_inputs/ADD_u6_u6_876/ADD_u6_u6_876_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874/Update/$exit
      -- 
    cr_1590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(17), ack => AND_u6_u6_881_inst_req_1); -- 
    rr_1585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(17), ack => AND_u6_u6_881_inst_req_0); -- 
    populateRxQueue_CP_1311_elements(17) <= populateRxQueue_CP_1311_elements(0);
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Sample/ra
      -- 
    ra_1586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_881_inst_ack_0, ack => populateRxQueue_CP_1311_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/Update/ca
      -- 
    ca_1591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_881_inst_ack_1, ack => populateRxQueue_CP_1311_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	24 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/$exit
      -- CP-element group 20: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/$exit
      -- CP-element group 20: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/SplitProtocol/$exit
      -- CP-element group 20: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/$exit
      -- CP-element group 20: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_req
      -- CP-element group 20: 	 branch_block_stmt_870/merge_stmt_871__entry___PhiReq/phi_stmt_872/phi_stmt_872_sources/AND_u6_u6_881/$exit
      -- 
    phi_stmt_872_req_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_872_req_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(20), ack => phi_stmt_872_req_0); -- 
    populateRxQueue_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1311_elements(19) & populateRxQueue_CP_1311_elements(18);
      gj_populateRxQueue_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1311_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	13 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Sample/ack
      -- CP-element group 21: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Sample/$exit
      -- 
    ack_1609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_930_882_buf_ack_0, ack => populateRxQueue_CP_1311_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/Update/ack
      -- 
    ack_1614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_930_882_buf_ack_1, ack => populateRxQueue_CP_1311_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/Interlock/$exit
      -- CP-element group 23: 	 branch_block_stmt_870/loopback_PhiReq/$exit
      -- CP-element group 23: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/$exit
      -- CP-element group 23: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_req
      -- CP-element group 23: 	 branch_block_stmt_870/loopback_PhiReq/phi_stmt_872/phi_stmt_872_sources/$exit
      -- 
    phi_stmt_872_req_1615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_872_req_1615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(23), ack => phi_stmt_872_req_1); -- 
    populateRxQueue_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1311_elements(21) & populateRxQueue_CP_1311_elements(22);
      gj_populateRxQueue_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1311_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  merge  transition  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	20 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_870/merge_stmt_871_PhiReqMerge
      -- CP-element group 24: 	 branch_block_stmt_870/merge_stmt_871_PhiAck/$entry
      -- 
    populateRxQueue_CP_1311_elements(24) <= OrReduce(populateRxQueue_CP_1311_elements(20) & populateRxQueue_CP_1311_elements(23));
    -- CP-element group 25:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	5 
    -- CP-element group 25: 	6 
    -- CP-element group 25: 	7 
    -- CP-element group 25: 	3 
    -- CP-element group 25: 	2 
    -- CP-element group 25:  members (20) 
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_update_start_
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Sample/crr
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_update_start_
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Update/ccr
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_870/merge_stmt_871_PhiAck/phi_stmt_872_ack
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_update_start_
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_870/merge_stmt_871_PhiAck/$exit
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_920_Update/ccr
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/call_stmt_903_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/$entry
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930/AND_u6_u6_929_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_870/assign_stmt_891_to_assign_stmt_930__entry__
      -- CP-element group 25: 	 branch_block_stmt_870/merge_stmt_871__exit__
      -- 
    phi_stmt_872_ack_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_872_ack_0, ack => populateRxQueue_CP_1311_elements(25)); -- 
    crr_1335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(25), ack => call_stmt_903_call_req_0); -- 
    ccr_1340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(25), ack => call_stmt_903_call_req_1); -- 
    rr_1363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(25), ack => AND_u6_u6_929_inst_req_0); -- 
    ccr_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(25), ack => call_stmt_920_call_req_1); -- 
    cr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1311_elements(25), ack => AND_u6_u6_929_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_876_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_889_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_924_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_881_wire : std_logic_vector(5 downto 0);
    signal EQ_u1_u1_943_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_936_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_898_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_877_wire : std_logic_vector(31 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_925_wire : std_logic_vector(31 downto 0);
    signal R_RX_QUEUES_REG_START_OFFSET_888_wire_constant : std_logic_vector(5 downto 0);
    signal SUB_u32_u32_879_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_927_wire : std_logic_vector(31 downto 0);
    signal konst_875_wire_constant : std_logic_vector(5 downto 0);
    signal konst_878_wire_constant : std_logic_vector(31 downto 0);
    signal konst_923_wire_constant : std_logic_vector(5 downto 0);
    signal konst_926_wire_constant : std_logic_vector(31 downto 0);
    signal konst_937_wire_constant : std_logic_vector(31 downto 0);
    signal konst_942_wire_constant : std_logic_vector(0 downto 0);
    signal n_q_index_930 : std_logic_vector(5 downto 0);
    signal n_q_index_930_882_buffered : std_logic_vector(5 downto 0);
    signal push_status_920 : std_logic_vector(0 downto 0);
    signal q_index_872 : std_logic_vector(5 downto 0);
    signal register_index_891 : std_logic_vector(5 downto 0);
    signal rx_queue_pointer_32_903 : std_logic_vector(31 downto 0);
    signal rx_queue_pointer_36_909 : std_logic_vector(35 downto 0);
    signal slice_918_wire : std_logic_vector(31 downto 0);
    signal status_939 : std_logic_vector(0 downto 0);
    signal type_cast_880_wire : std_logic_vector(5 downto 0);
    signal type_cast_895_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_901_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_907_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_928_wire : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_898_wire_constant <= "1111";
    R_RX_QUEUES_REG_START_OFFSET_888_wire_constant <= "000010";
    konst_875_wire_constant <= "000001";
    konst_878_wire_constant <= "00000000000000000000000000000001";
    konst_923_wire_constant <= "000001";
    konst_926_wire_constant <= "00000000000000000000000000000001";
    konst_937_wire_constant <= "00000000000000000000000000100000";
    konst_942_wire_constant <= "0";
    type_cast_895_wire_constant <= "1";
    type_cast_901_wire_constant <= "00000000000000000000000000000000";
    type_cast_907_wire_constant <= "0000";
    type_cast_915_wire_constant <= "0";
    phi_stmt_872: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= AND_u6_u6_881_wire & n_q_index_930_882_buffered;
      req <= phi_stmt_872_req_0 & phi_stmt_872_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_872",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_872_ack_0,
          idata => idata,
          odata => q_index_872,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_872
    -- flow-through slice operator slice_918_inst
    slice_918_wire <= rx_buffer_pointer_buffer(35 downto 4);
    n_q_index_930_882_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_q_index_930_882_buf_req_0;
      n_q_index_930_882_buf_ack_0<= wack(0);
      rreq(0) <= n_q_index_930_882_buf_req_1;
      n_q_index_930_882_buf_ack_1<= rack(0);
      n_q_index_930_882_buf : InterlockBuffer generic map ( -- 
        name => "n_q_index_930_882_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_q_index_930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_q_index_930_882_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_880_inst
    process(SUB_u32_u32_879_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_879_wire(5 downto 0);
      type_cast_880_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_890_inst
    process(ADD_u6_u6_889_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_889_wire(5 downto 0);
      register_index_891 <= tmp_var; -- 
    end process;
    -- interlock type_cast_928_inst
    process(SUB_u32_u32_927_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_927_wire(5 downto 0);
      type_cast_928_wire <= tmp_var; -- 
    end process;
    if_stmt_934_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_936_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_934_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_934_branch_req_0,
          ack0 => if_stmt_934_branch_ack_0,
          ack1 => if_stmt_934_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_940_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_943_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_940_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_940_branch_req_0,
          ack0 => if_stmt_940_branch_ack_0,
          ack1 => if_stmt_940_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u6_u6_876_inst
    process(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874_wire, konst_875_wire_constant, tmp_var);
      ADD_u6_u6_876_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_889_inst
    process(q_index_872) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_872, R_RX_QUEUES_REG_START_OFFSET_888_wire_constant, tmp_var);
      ADD_u6_u6_889_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_924_inst
    process(q_index_872) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_872, konst_923_wire_constant, tmp_var);
      ADD_u6_u6_924_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_881_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_876_wire & type_cast_880_wire;
      AND_u6_u6_881_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_881_inst_req_0;
      AND_u6_u6_881_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_881_inst_req_1;
      AND_u6_u6_881_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : AND_u6_u6_929_inst 
    ApIntAnd_group_4: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_924_wire & type_cast_928_wire;
      n_q_index_930 <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_929_inst_req_0;
      AND_u6_u6_929_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_929_inst_req_1;
      AND_u6_u6_929_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator CONCAT_u32_u36_908_inst
    process(rx_queue_pointer_32_903) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(rx_queue_pointer_32_903, type_cast_907_wire_constant, tmp_var);
      rx_queue_pointer_36_909 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_943_inst
    process(status_939) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(status_939, konst_942_wire_constant, tmp_var);
      EQ_u1_u1_943_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_936_inst
    process(push_status_920) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", push_status_920, tmp_var);
      NOT_u1_u1_936_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u32_u32_879_inst
    process(RPIPE_NUMBER_OF_SERVERS_877_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_877_wire, konst_878_wire_constant, tmp_var);
      SUB_u32_u32_879_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_927_inst
    process(RPIPE_NUMBER_OF_SERVERS_925_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_925_wire, konst_926_wire_constant, tmp_var);
      SUB_u32_u32_927_wire <= tmp_var; --
    end process;
    -- read from input-signal LAST_WRITTEN_RX_QUEUE_INDEX
    RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_874_wire <= LAST_WRITTEN_RX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_925_wire <= NUMBER_OF_SERVERS;
    RPIPE_NUMBER_OF_SERVERS_877_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_947_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= q_index_872;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_903_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_903_call_req_0;
      call_stmt_903_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_903_call_req_1;
      call_stmt_903_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_895_wire_constant & NOT_u4_u4_898_wire_constant & register_index_891 & type_cast_901_wire_constant;
      rx_queue_pointer_32_903 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_920_call 
    pushIntoQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_920_call_req_0;
      call_stmt_920_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_920_call_req_1;
      call_stmt_920_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_1_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_915_wire_constant & rx_queue_pointer_36_909 & slice_918_wire;
      push_status_920 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    operator_delay_time_2296_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_939_call_req_0;
      call_stmt_939_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_939_call_req_1;
      call_stmt_939_call_ack_1<= update_ack(0);
      call_stmt_939_call: delay_time_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        T => konst_937_wire_constant,
        delay_done => status_939,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end populateRxQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity pushIntoQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_call_data : out  std_logic_vector(35 downto 0);
    releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_call_data : out  std_logic_vector(35 downto 0);
    acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_return_data : in   std_logic_vector(0 downto 0);
    acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
    setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_call_data : out  std_logic_vector(99 downto 0);
    setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity pushIntoQueue;
architecture pushIntoQueue_arch of pushIntoQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 69)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal pushIntoQueue_CP_1116_start: Boolean;
  signal pushIntoQueue_CP_1116_symbol: Boolean;
  -- volatile/operator module components. 
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_pointer : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_787_call_req_0 : boolean;
  signal call_stmt_787_call_ack_0 : boolean;
  signal call_stmt_787_call_req_1 : boolean;
  signal call_stmt_787_call_ack_1 : boolean;
  signal call_stmt_795_call_req_0 : boolean;
  signal call_stmt_795_call_ack_0 : boolean;
  signal call_stmt_795_call_req_1 : boolean;
  signal call_stmt_795_call_ack_1 : boolean;
  signal call_stmt_826_call_req_0 : boolean;
  signal call_stmt_826_call_ack_0 : boolean;
  signal call_stmt_826_call_req_1 : boolean;
  signal call_stmt_826_call_ack_1 : boolean;
  signal call_stmt_831_call_req_0 : boolean;
  signal call_stmt_831_call_ack_0 : boolean;
  signal call_stmt_831_call_req_1 : boolean;
  signal call_stmt_831_call_ack_1 : boolean;
  signal call_stmt_835_call_req_0 : boolean;
  signal call_stmt_835_call_ack_0 : boolean;
  signal call_stmt_835_call_req_1 : boolean;
  signal call_stmt_835_call_ack_1 : boolean;
  signal NOT_u1_u1_838_inst_req_0 : boolean;
  signal NOT_u1_u1_838_inst_ack_0 : boolean;
  signal NOT_u1_u1_838_inst_req_1 : boolean;
  signal NOT_u1_u1_838_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "pushIntoQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 69) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(68 downto 37) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(68 downto 37);
  in_buffer_data_in(tag_length + 68 downto 69) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 68 downto 69);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  pushIntoQueue_CP_1116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "pushIntoQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  pushIntoQueue_CP_1116: Block -- control-path 
    signal pushIntoQueue_CP_1116_elements: BooleanArray(14 downto 0);
    -- 
  begin -- 
    pushIntoQueue_CP_1116_elements(0) <= pushIntoQueue_CP_1116_start;
    pushIntoQueue_CP_1116_symbol <= pushIntoQueue_CP_1116_elements(14);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_787/$entry
      -- CP-element group 0: 	 call_stmt_787/call_stmt_787_sample_start_
      -- CP-element group 0: 	 call_stmt_787/call_stmt_787_update_start_
      -- CP-element group 0: 	 call_stmt_787/call_stmt_787_Sample/$entry
      -- CP-element group 0: 	 call_stmt_787/call_stmt_787_Sample/crr
      -- CP-element group 0: 	 call_stmt_787/call_stmt_787_Update/$entry
      -- CP-element group 0: 	 call_stmt_787/call_stmt_787_Update/ccr
      -- 
    crr_1129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(0), ack => call_stmt_787_call_req_0); -- 
    ccr_1134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(0), ack => call_stmt_787_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_787/call_stmt_787_sample_completed_
      -- CP-element group 1: 	 call_stmt_787/call_stmt_787_Sample/$exit
      -- CP-element group 1: 	 call_stmt_787/call_stmt_787_Sample/cra
      -- 
    cra_1130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_787_call_ack_0, ack => pushIntoQueue_CP_1116_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (17) 
      -- CP-element group 2: 	 call_stmt_787/$exit
      -- CP-element group 2: 	 call_stmt_787/call_stmt_787_update_completed_
      -- CP-element group 2: 	 call_stmt_787/call_stmt_787_Update/$exit
      -- CP-element group 2: 	 call_stmt_787/call_stmt_787_Update/cca
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/$entry
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_sample_start_
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_update_start_
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Sample/$entry
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Sample/crr
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Update/$entry
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Update/ccr
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_update_start_
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Update/$entry
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Update/ccr
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_update_start_
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Update/$entry
      -- CP-element group 2: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Update/ccr
      -- 
    cca_1135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_787_call_ack_1, ack => pushIntoQueue_CP_1116_elements(2)); -- 
    crr_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(2), ack => call_stmt_795_call_req_0); -- 
    ccr_1151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(2), ack => call_stmt_795_call_req_1); -- 
    ccr_1179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(2), ack => call_stmt_831_call_req_1); -- 
    ccr_1165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(2), ack => call_stmt_826_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_sample_completed_
      -- CP-element group 3: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Sample/$exit
      -- CP-element group 3: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Sample/cra
      -- 
    cra_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_795_call_ack_0, ack => pushIntoQueue_CP_1116_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_update_completed_
      -- CP-element group 4: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Update/$exit
      -- CP-element group 4: 	 call_stmt_795_to_call_stmt_831/call_stmt_795_Update/cca
      -- CP-element group 4: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_sample_start_
      -- CP-element group 4: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Sample/$entry
      -- CP-element group 4: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Sample/crr
      -- 
    cca_1152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_795_call_ack_1, ack => pushIntoQueue_CP_1116_elements(4)); -- 
    crr_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(4), ack => call_stmt_826_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_sample_completed_
      -- CP-element group 5: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Sample/$exit
      -- CP-element group 5: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Sample/cra
      -- 
    cra_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_826_call_ack_0, ack => pushIntoQueue_CP_1116_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_update_completed_
      -- CP-element group 6: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Update/$exit
      -- CP-element group 6: 	 call_stmt_795_to_call_stmt_831/call_stmt_826_Update/cca
      -- 
    cca_1166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_826_call_ack_1, ack => pushIntoQueue_CP_1116_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_sample_start_
      -- CP-element group 7: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Sample/$entry
      -- CP-element group 7: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Sample/crr
      -- 
    crr_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(7), ack => call_stmt_831_call_req_0); -- 
    pushIntoQueue_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "pushIntoQueue_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1116_elements(6) & pushIntoQueue_CP_1116_elements(4);
      gj_pushIntoQueue_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1116_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_sample_completed_
      -- CP-element group 8: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Sample/$exit
      -- CP-element group 8: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Sample/cra
      -- 
    cra_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_831_call_ack_0, ack => pushIntoQueue_CP_1116_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (17) 
      -- CP-element group 9: 	 call_stmt_795_to_call_stmt_831/$exit
      -- CP-element group 9: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_update_completed_
      -- CP-element group 9: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Update/$exit
      -- CP-element group 9: 	 call_stmt_795_to_call_stmt_831/call_stmt_831_Update/cca
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/$entry
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_sample_start_
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_update_start_
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Sample/$entry
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Sample/crr
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Update/$entry
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Update/ccr
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_sample_start_
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_update_start_
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Sample/$entry
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Sample/rr
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Update/$entry
      -- CP-element group 9: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Update/cr
      -- 
    cca_1180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_831_call_ack_1, ack => pushIntoQueue_CP_1116_elements(9)); -- 
    crr_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(9), ack => call_stmt_835_call_req_0); -- 
    ccr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(9), ack => call_stmt_835_call_req_1); -- 
    rr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(9), ack => NOT_u1_u1_838_inst_req_0); -- 
    cr_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1116_elements(9), ack => NOT_u1_u1_838_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_sample_completed_
      -- CP-element group 10: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Sample/$exit
      -- CP-element group 10: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Sample/cra
      -- 
    cra_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_835_call_ack_0, ack => pushIntoQueue_CP_1116_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_update_completed_
      -- CP-element group 11: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Update/$exit
      -- CP-element group 11: 	 call_stmt_835_to_assign_stmt_839/call_stmt_835_Update/cca
      -- 
    cca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_835_call_ack_1, ack => pushIntoQueue_CP_1116_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_sample_completed_
      -- CP-element group 12: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Sample/$exit
      -- CP-element group 12: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Sample/ra
      -- 
    ra_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_838_inst_ack_0, ack => pushIntoQueue_CP_1116_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_update_completed_
      -- CP-element group 13: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Update/$exit
      -- CP-element group 13: 	 call_stmt_835_to_assign_stmt_839/NOT_u1_u1_838_Update/ca
      -- 
    ca_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_838_inst_ack_1, ack => pushIntoQueue_CP_1116_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 $exit
      -- CP-element group 14: 	 call_stmt_835_to_assign_stmt_839/$exit
      -- 
    pushIntoQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1116_elements(11) & pushIntoQueue_CP_1116_elements(13);
      gj_pushIntoQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1116_elements(14), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_808_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_800_wire_constant : std_logic_vector(31 downto 0);
    signal konst_805_wire_constant : std_logic_vector(31 downto 0);
    signal konst_807_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_787 : std_logic_vector(0 downto 0);
    signal next_wp_810 : std_logic_vector(31 downto 0);
    signal q_full_815 : std_logic_vector(0 downto 0);
    signal read_pointer_795 : std_logic_vector(31 downto 0);
    signal round_off_802 : std_logic_vector(0 downto 0);
    signal write_pointer_795 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    SUB_u32_u32_800_wire_constant <= "00000000000000000000000000000111";
    konst_805_wire_constant <= "00000000000000000000000000000000";
    konst_807_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_809_inst
    next_wp_810 <= konst_805_wire_constant when (round_off_802(0) /=  '0') else ADD_u32_u32_808_wire;
    -- binary operator ADD_u32_u32_808_inst
    process(write_pointer_795) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(write_pointer_795, konst_807_wire_constant, tmp_var);
      ADD_u32_u32_808_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_801_inst
    process(write_pointer_795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_pointer_795, SUB_u32_u32_800_wire_constant, tmp_var);
      round_off_802 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_814_inst
    process(next_wp_810, read_pointer_795) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_wp_810, read_pointer_795, tmp_var);
      q_full_815 <= tmp_var; --
    end process;
    -- shared split operator group (3) : NOT_u1_u1_838_inst 
    ApIntNot_group_3: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= q_full_815;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_838_inst_req_0;
      NOT_u1_u1_838_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_838_inst_req_1;
      NOT_u1_u1_838_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_3_gI: SplitGuardInterface generic map(name => "ApIntNot_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared call operator group (0) : call_stmt_787_call 
    acquireMutex_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_787_call_req_0;
      call_stmt_787_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_787_call_req_1;
      call_stmt_787_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireMutex_call_group_0_gI: SplitGuardInterface generic map(name => "acquireMutex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_787 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireMutex_call_reqs(0),
          ackR => acquireMutex_call_acks(0),
          dataR => acquireMutex_call_data(35 downto 0),
          tagR => acquireMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireMutex_return_acks(0), -- cross-over
          ackL => acquireMutex_return_reqs(0), -- cross-over
          dataL => acquireMutex_return_data(0 downto 0),
          tagL => acquireMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_795_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_795_call_req_0;
      call_stmt_795_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_795_call_req_1;
      call_stmt_795_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_pointer_795 <= data_out(63 downto 32);
      read_pointer_795 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_826_call 
    setQueueElement_call_group_2: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_826_call_req_0;
      call_stmt_826_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_826_call_req_1;
      call_stmt_826_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_815(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueueElement_call_group_2_gI: SplitGuardInterface generic map(name => "setQueueElement_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_pointer_795 & q_w_data_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueueElement_call_reqs(0),
          ackR => setQueueElement_call_acks(0),
          dataR => setQueueElement_call_data(99 downto 0),
          tagR => setQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueueElement_return_acks(0), -- cross-over
          ackL => setQueueElement_return_reqs(0), -- cross-over
          tagL => setQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_831_call 
    setQueuePointers_call_group_3: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_831_call_req_0;
      call_stmt_831_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_831_call_req_1;
      call_stmt_831_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_815(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_3_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & next_wp_810 & read_pointer_795;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_835_call 
    releaseMutex_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_835_call_req_0;
      call_stmt_835_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_835_call_req_1;
      call_stmt_835_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseMutex_call_group_4_gI: SplitGuardInterface generic map(name => "releaseMutex_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseMutex_call_reqs(0),
          ackR => releaseMutex_call_acks(0),
          dataR => releaseMutex_call_data(35 downto 0),
          tagR => releaseMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseMutex_return_acks(0), -- cross-over
          ackL => releaseMutex_return_reqs(0), -- cross-over
          tagL => releaseMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end pushIntoQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity releaseMutex is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity releaseMutex;
architecture releaseMutex_arch of releaseMutex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal releaseMutex_CP_565_start: Boolean;
  signal releaseMutex_CP_565_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_471_call_ack_1 : boolean;
  signal call_stmt_471_call_req_1 : boolean;
  signal call_stmt_471_call_req_0 : boolean;
  signal call_stmt_471_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "releaseMutex_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  releaseMutex_CP_565_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "releaseMutex_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseMutex_CP_565_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= releaseMutex_CP_565_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseMutex_CP_565_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  releaseMutex_CP_565: Block -- control-path 
    signal releaseMutex_CP_565_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    releaseMutex_CP_565_elements(0) <= releaseMutex_CP_565_start;
    releaseMutex_CP_565_symbol <= releaseMutex_CP_565_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_471/call_stmt_471_Update/ccr
      -- CP-element group 0: 	 call_stmt_471/call_stmt_471_Update/$entry
      -- CP-element group 0: 	 call_stmt_471/call_stmt_471_Sample/crr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_471/$entry
      -- CP-element group 0: 	 call_stmt_471/call_stmt_471_Sample/$entry
      -- CP-element group 0: 	 call_stmt_471/call_stmt_471_update_start_
      -- CP-element group 0: 	 call_stmt_471/call_stmt_471_sample_start_
      -- 
    crr_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseMutex_CP_565_elements(0), ack => call_stmt_471_call_req_0); -- 
    ccr_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseMutex_CP_565_elements(0), ack => call_stmt_471_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_471/call_stmt_471_sample_completed_
      -- CP-element group 1: 	 call_stmt_471/call_stmt_471_Sample/cra
      -- CP-element group 1: 	 call_stmt_471/call_stmt_471_Sample/$exit
      -- 
    cra_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_471_call_ack_0, ack => releaseMutex_CP_565_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_471/call_stmt_471_Update/cca
      -- CP-element group 2: 	 call_stmt_471/call_stmt_471_Update/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_471/$exit
      -- CP-element group 2: 	 call_stmt_471/call_stmt_471_update_completed_
      -- 
    cca_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_471_call_ack_1, ack => releaseMutex_CP_565_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u4_u8_466_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_471 : std_logic_vector(63 downto 0);
    signal type_cast_458_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_460_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_469_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_466_wire_constant <= "11110000";
    type_cast_458_wire_constant <= "0";
    type_cast_460_wire_constant <= "0";
    type_cast_469_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- shared call operator group (0) : call_stmt_471_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_471_call_req_0;
      call_stmt_471_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_471_call_req_1;
      call_stmt_471_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_458_wire_constant & type_cast_460_wire_constant & CONCAT_u4_u8_466_wire_constant & q_base_address_buffer & type_cast_469_wire_constant;
      ignore_471 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end releaseMutex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    write_pointer : in  std_logic_vector(31 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueueElement;
architecture setQueueElement_arch of setQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal write_pointer_buffer :  std_logic_vector(31 downto 0);
  signal write_pointer_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal setQueueElement_CP_1096_start: Boolean;
  signal setQueueElement_CP_1096_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_777_call_req_0 : boolean;
  signal call_stmt_777_call_ack_0 : boolean;
  signal call_stmt_777_call_req_1 : boolean;
  signal call_stmt_777_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= write_pointer;
  write_pointer_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueueElement_CP_1096_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1096_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueueElement_CP_1096_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1096_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueueElement_CP_1096: Block -- control-path 
    signal setQueueElement_CP_1096_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueueElement_CP_1096_elements(0) <= setQueueElement_CP_1096_start;
    setQueueElement_CP_1096_symbol <= setQueueElement_CP_1096_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_721_to_call_stmt_777/$entry
      -- CP-element group 0: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_sample_start_
      -- CP-element group 0: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_update_start_
      -- CP-element group 0: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Sample/crr
      -- CP-element group 0: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Update/$entry
      -- CP-element group 0: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Update/ccr
      -- 
    crr_1109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1096_elements(0), ack => call_stmt_777_call_req_0); -- 
    ccr_1114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1096_elements(0), ack => call_stmt_777_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_sample_completed_
      -- CP-element group 1: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Sample/cra
      -- 
    cra_1110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_777_call_ack_0, ack => setQueueElement_CP_1096_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_721_to_call_stmt_777/$exit
      -- CP-element group 2: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_update_completed_
      -- CP-element group 2: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Update/$exit
      -- CP-element group 2: 	 assign_stmt_721_to_call_stmt_777/call_stmt_777_Update/cca
      -- 
    cca_1115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_777_call_ack_1, ack => setQueueElement_CP_1096_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_735_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_753_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_728_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u32_u64_757_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_761_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_741_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_747_wire_constant : std_logic_vector(7 downto 0);
    signal bmask_749 : std_logic_vector(7 downto 0);
    signal buffer_address_721 : std_logic_vector(35 downto 0);
    signal element_pair_address_731 : std_logic_vector(35 downto 0);
    signal ignore_777 : std_logic_vector(63 downto 0);
    signal konst_734_wire_constant : std_logic_vector(31 downto 0);
    signal konst_752_wire_constant : std_logic_vector(31 downto 0);
    signal slice_725_wire : std_logic_vector(30 downto 0);
    signal type_cast_719_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_727_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_729_wire : std_logic_vector(35 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_770_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_772_wire_constant : std_logic_vector(0 downto 0);
    signal wval_763 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_741_wire_constant <= "00001111";
    CONCAT_u4_u8_747_wire_constant <= "11110000";
    konst_734_wire_constant <= "00000000000000000000000000000000";
    konst_752_wire_constant <= "00000000000000000000000000000000";
    type_cast_719_wire_constant <= "000000000000000000000000000000010000";
    type_cast_727_wire_constant <= "000";
    type_cast_755_wire_constant <= "00000000000000000000000000000000";
    type_cast_760_wire_constant <= "00000000000000000000000000000000";
    type_cast_770_wire_constant <= "0";
    type_cast_772_wire_constant <= "0";
    -- flow-through select operator MUX_748_inst
    bmask_749 <= CONCAT_u4_u8_741_wire_constant when (BITSEL_u32_u1_735_wire(0) /=  '0') else CONCAT_u4_u8_747_wire_constant;
    -- flow-through select operator MUX_762_inst
    wval_763 <= CONCAT_u32_u64_757_wire when (BITSEL_u32_u1_753_wire(0) /=  '0') else CONCAT_u32_u64_761_wire;
    -- flow-through slice operator slice_725_inst
    slice_725_wire <= write_pointer_buffer(31 downto 1);
    -- interlock type_cast_729_inst
    process(CONCAT_u31_u34_728_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_728_wire(33 downto 0);
      type_cast_729_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_720_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_719_wire_constant, tmp_var);
      buffer_address_721 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_730_inst
    process(buffer_address_721, type_cast_729_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_721, type_cast_729_wire, tmp_var);
      element_pair_address_731 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_735_inst
    process(write_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_pointer_buffer, konst_734_wire_constant, tmp_var);
      BITSEL_u32_u1_735_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_753_inst
    process(write_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_pointer_buffer, konst_752_wire_constant, tmp_var);
      BITSEL_u32_u1_753_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_728_inst
    process(slice_725_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_725_wire, type_cast_727_wire_constant, tmp_var);
      CONCAT_u31_u34_728_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_757_inst
    process(type_cast_755_wire_constant, q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_755_wire_constant, q_w_data_buffer, tmp_var);
      CONCAT_u32_u64_757_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_761_inst
    process(q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(q_w_data_buffer, type_cast_760_wire_constant, tmp_var);
      CONCAT_u32_u64_761_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_777_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_777_call_req_0;
      call_stmt_777_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_777_call_req_1;
      call_stmt_777_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_770_wire_constant & type_cast_772_wire_constant & bmask_749 & element_pair_address_731 & wval_763;
      ignore_777 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity setQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : in  std_logic_vector(31 downto 0);
    rp : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueuePointers;
architecture setQueuePointers_arch of setQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  -- output port buffer signals
  signal setQueuePointers_CP_545_start: Boolean;
  signal setQueuePointers_CP_545_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_453_call_ack_1 : boolean;
  signal call_stmt_453_call_req_1 : boolean;
  signal call_stmt_453_call_ack_0 : boolean;
  signal call_stmt_453_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= wp;
  wp_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= rp;
  rp_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueuePointers_CP_545_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_545_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueuePointers_CP_545_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_545_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueuePointers_CP_545: Block -- control-path 
    signal setQueuePointers_CP_545_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueuePointers_CP_545_elements(0) <= setQueuePointers_CP_545_start;
    setQueuePointers_CP_545_symbol <= setQueuePointers_CP_545_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_453/call_stmt_453_sample_start_
      -- CP-element group 0: 	 call_stmt_453/call_stmt_453_Update/ccr
      -- CP-element group 0: 	 call_stmt_453/call_stmt_453_Sample/$entry
      -- CP-element group 0: 	 call_stmt_453/call_stmt_453_Update/$entry
      -- CP-element group 0: 	 call_stmt_453/call_stmt_453_Sample/crr
      -- CP-element group 0: 	 call_stmt_453/$entry
      -- CP-element group 0: 	 call_stmt_453/call_stmt_453_update_start_
      -- CP-element group 0: 	 $entry
      -- 
    crr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_545_elements(0), ack => call_stmt_453_call_req_0); -- 
    ccr_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_545_elements(0), ack => call_stmt_453_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_453/call_stmt_453_Sample/cra
      -- CP-element group 1: 	 call_stmt_453/call_stmt_453_Sample/$exit
      -- CP-element group 1: 	 call_stmt_453/call_stmt_453_sample_completed_
      -- 
    cra_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_453_call_ack_0, ack => setQueuePointers_CP_545_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_453/call_stmt_453_Update/cca
      -- CP-element group 2: 	 call_stmt_453/call_stmt_453_update_completed_
      -- CP-element group 2: 	 call_stmt_453/call_stmt_453_Update/$exit
      -- CP-element group 2: 	 call_stmt_453/$exit
      -- CP-element group 2: 	 $exit
      -- 
    cca_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_453_call_ack_1, ack => setQueuePointers_CP_545_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_448_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u32_u64_451_wire : std_logic_vector(63 downto 0);
    signal NOT_u8_u8_445_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_453 : std_logic_vector(63 downto 0);
    signal konst_447_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_440_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_442_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_445_wire_constant <= "11111111";
    konst_447_wire_constant <= "000000000000000000000000000000001000";
    type_cast_440_wire_constant <= "0";
    type_cast_442_wire_constant <= "0";
    -- binary operator ADD_u36_u36_448_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_447_wire_constant, tmp_var);
      ADD_u36_u36_448_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_451_inst
    process(wp_buffer, rp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(wp_buffer, rp_buffer, tmp_var);
      CONCAT_u32_u64_451_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_453_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_453_call_req_0;
      call_stmt_453_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_453_call_req_1;
      call_stmt_453_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_440_wire_constant & type_cast_442_wire_constant & NOT_u8_u8_445_wire_constant & ADD_u36_u36_448_wire & CONCAT_u32_u64_451_wire;
      ignore_453 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
    getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
    getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
    transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_call_data : out  std_logic_vector(31 downto 0);
    transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
    transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_return_data : in   std_logic_vector(0 downto 0);
    transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitEngineDaemon;
architecture transmitEngineDaemon_arch of transmitEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal transmitEngineDaemon_CP_3018_start: Boolean;
  signal transmitEngineDaemon_CP_3018_symbol: Boolean;
  -- volatile/operator module components. 
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_ack_1 : boolean;
  signal if_stmt_1514_branch_req_0 : boolean;
  signal if_stmt_1514_branch_ack_1 : boolean;
  signal if_stmt_1514_branch_ack_0 : boolean;
  signal do_while_stmt_1522_branch_req_0 : boolean;
  signal AND_u6_u6_1533_inst_req_0 : boolean;
  signal AND_u6_u6_1533_inst_ack_0 : boolean;
  signal AND_u6_u6_1533_inst_req_1 : boolean;
  signal AND_u6_u6_1533_inst_ack_1 : boolean;
  signal call_stmt_1540_call_req_0 : boolean;
  signal call_stmt_1540_call_ack_0 : boolean;
  signal call_stmt_1540_call_req_1 : boolean;
  signal call_stmt_1540_call_ack_1 : boolean;
  signal call_stmt_1544_call_req_0 : boolean;
  signal call_stmt_1544_call_ack_0 : boolean;
  signal call_stmt_1544_call_req_1 : boolean;
  signal call_stmt_1544_call_ack_1 : boolean;
  signal NOT_u1_u1_1554_inst_req_0 : boolean;
  signal NOT_u1_u1_1554_inst_ack_0 : boolean;
  signal NOT_u1_u1_1554_inst_req_1 : boolean;
  signal NOT_u1_u1_1554_inst_ack_1 : boolean;
  signal W_pkt_pointer_1539_delayed_4_0_1564_inst_req_0 : boolean;
  signal W_pkt_pointer_1539_delayed_4_0_1564_inst_ack_0 : boolean;
  signal W_pkt_pointer_1539_delayed_4_0_1564_inst_req_1 : boolean;
  signal W_pkt_pointer_1539_delayed_4_0_1564_inst_ack_1 : boolean;
  signal call_stmt_1573_call_req_0 : boolean;
  signal call_stmt_1573_call_ack_0 : boolean;
  signal call_stmt_1573_call_req_1 : boolean;
  signal call_stmt_1573_call_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_ack_1 : boolean;
  signal do_while_stmt_1522_branch_ack_0 : boolean;
  signal do_while_stmt_1522_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitEngineDaemon_CP_3018_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3018_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3018_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3018_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitEngineDaemon_CP_3018: Block -- control-path 
    signal transmitEngineDaemon_CP_3018_elements: BooleanArray(50 downto 0);
    -- 
  begin -- 
    transmitEngineDaemon_CP_3018_elements(0) <= transmitEngineDaemon_CP_3018_start;
    transmitEngineDaemon_CP_3018_symbol <= transmitEngineDaemon_CP_3018_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1511/$entry
      -- CP-element group 0: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_sample_start_
      -- CP-element group 0: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Sample/req
      -- 
    req_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(0), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_update_start_
      -- CP-element group 1: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Update/req
      -- 
    ack_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_ack_0, ack => transmitEngineDaemon_CP_3018_elements(1)); -- 
    req_3036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(1), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	50 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_1511/$exit
      -- CP-element group 2: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_update_completed_
      -- CP-element group 2: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1511/WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_1512/$entry
      -- CP-element group 2: 	 branch_block_stmt_1512/branch_block_stmt_1512__entry__
      -- CP-element group 2: 	 branch_block_stmt_1512/merge_stmt_1513__entry__
      -- CP-element group 2: 	 branch_block_stmt_1512/merge_stmt_1513_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1512/merge_stmt_1513__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1512/merge_stmt_1513__entry___PhiReq/$exit
      -- 
    ack_3037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_ack_1, ack => transmitEngineDaemon_CP_3018_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_1512/$exit
      -- CP-element group 3: 	 branch_block_stmt_1512/branch_block_stmt_1512__exit__
      -- 
    transmitEngineDaemon_CP_3018_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	49 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	50 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1512/do_while_stmt_1522__exit__
      -- CP-element group 4: 	 branch_block_stmt_1512/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_1512/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1512/disable_loopback_PhiReq/$exit
      -- 
    transmitEngineDaemon_CP_3018_elements(4) <= transmitEngineDaemon_CP_3018_elements(49);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	50 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1512/if_stmt_1514_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1512/if_stmt_1514_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1512/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1512/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1512/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_3110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1514_branch_ack_1, ack => transmitEngineDaemon_CP_3018_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	50 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_1512/if_stmt_1514__exit__
      -- CP-element group 6: 	 branch_block_stmt_1512/do_while_stmt_1522__entry__
      -- CP-element group 6: 	 branch_block_stmt_1512/if_stmt_1514_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1512/if_stmt_1514_else_link/else_choice_transition
      -- 
    else_choice_transition_3114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1514_branch_ack_0, ack => transmitEngineDaemon_CP_3018_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1512/do_while_stmt_1522/$entry
      -- CP-element group 7: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522__entry__
      -- 
    transmitEngineDaemon_CP_3018_elements(7) <= transmitEngineDaemon_CP_3018_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	49 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522__exit__
      -- 
    -- Element group transmitEngineDaemon_CP_3018_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_back
      -- 
    -- Element group transmitEngineDaemon_CP_3018_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	47 
    -- CP-element group 10: 	48 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1512/do_while_stmt_1522/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_taken/$entry
      -- 
    transmitEngineDaemon_CP_3018_elements(10) <= transmitEngineDaemon_CP_3018_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	46 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_body_done
      -- 
    transmitEngineDaemon_CP_3018_elements(11) <= transmitEngineDaemon_CP_3018_elements(46);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/back_edge_to_loop_body
      -- 
    transmitEngineDaemon_CP_3018_elements(12) <= transmitEngineDaemon_CP_3018_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/first_time_through_loop_body
      -- 
    transmitEngineDaemon_CP_3018_elements(13) <= transmitEngineDaemon_CP_3018_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	45 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/phi_stmt_1524_sample_start_
      -- 
    -- Element group transmitEngineDaemon_CP_3018_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	45 
    -- CP-element group 15: 	21 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/condition_evaluated
      -- 
    condition_evaluated_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(15), ack => do_while_stmt_1522_branch_req_0); -- 
    transmitEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(45) & transmitEngineDaemon_CP_3018_elements(21);
      gj_transmitEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/aggregated_phi_sample_req
      -- 
    transmitEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(14) & transmitEngineDaemon_CP_3018_elements(21);
      gj_transmitEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	43 
    -- CP-element group 17: 	24 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/aggregated_phi_update_req
      -- CP-element group 17: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/phi_stmt_1524_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(14) & transmitEngineDaemon_CP_3018_elements(43) & transmitEngineDaemon_CP_3018_elements(24);
      gj_transmitEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Sample/rr
      -- 
    rr_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(18), ack => AND_u6_u6_1533_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(16) & transmitEngineDaemon_CP_3018_elements(20);
      gj_transmitEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Update/cr
      -- 
    cr_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(19), ack => AND_u6_u6_1533_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(17) & transmitEngineDaemon_CP_3018_elements(21);
      gj_transmitEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	46 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/aggregated_phi_sample_ack
      -- CP-element group 20: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/phi_stmt_1524_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Sample/ra
      -- 
    ra_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1533_inst_ack_0, ack => transmitEngineDaemon_CP_3018_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: 	42 
    -- CP-element group 21: 	22 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/aggregated_phi_update_ack
      -- CP-element group 21: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/phi_stmt_1524_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/AND_u6_u6_1533_Update/ca
      -- 
    ca_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1533_inst_ack_1, ack => transmitEngineDaemon_CP_3018_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	41 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Sample/crr
      -- 
    crr_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(22), ack => call_stmt_1540_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(21) & transmitEngineDaemon_CP_3018_elements(41) & transmitEngineDaemon_CP_3018_elements(24);
      gj_transmitEngineDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	32 
    -- CP-element group 23: 	36 
    -- CP-element group 23: 	41 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Update/ccr
      -- 
    ccr_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(23), ack => call_stmt_1540_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(28) & transmitEngineDaemon_CP_3018_elements(32) & transmitEngineDaemon_CP_3018_elements(36) & transmitEngineDaemon_CP_3018_elements(41);
      gj_transmitEngineDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Sample/cra
      -- 
    cra_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1540_call_ack_0, ack => transmitEngineDaemon_CP_3018_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	30 
    -- CP-element group 25: 	34 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1540_Update/cca
      -- 
    cca_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1540_call_ack_1, ack => transmitEngineDaemon_CP_3018_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Sample/crr
      -- 
    crr_3175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(26), ack => call_stmt_1544_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(25) & transmitEngineDaemon_CP_3018_elements(28);
      gj_transmitEngineDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	40 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Update/ccr
      -- 
    ccr_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(27), ack => call_stmt_1544_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3018_elements(40);
      gj_transmitEngineDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Sample/cra
      -- 
    cra_3176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1544_call_ack_0, ack => transmitEngineDaemon_CP_3018_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	38 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1544_Update/cca
      -- 
    cca_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1544_call_ack_1, ack => transmitEngineDaemon_CP_3018_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	25 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Sample/rr
      -- 
    rr_3189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(30), ack => NOT_u1_u1_1554_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(25) & transmitEngineDaemon_CP_3018_elements(32);
      gj_transmitEngineDaemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	40 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Update/cr
      -- 
    cr_3194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(31), ack => NOT_u1_u1_1554_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3018_elements(40);
      gj_transmitEngineDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: 	23 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Sample/ra
      -- 
    ra_3190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1554_inst_ack_0, ack => transmitEngineDaemon_CP_3018_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	38 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/NOT_u1_u1_1554_Update/ca
      -- 
    ca_3195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1554_inst_ack_1, ack => transmitEngineDaemon_CP_3018_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	25 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Sample/req
      -- 
    req_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(34), ack => W_pkt_pointer_1539_delayed_4_0_1564_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(25) & transmitEngineDaemon_CP_3018_elements(36);
      gj_transmitEngineDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	40 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Update/req
      -- 
    req_3208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(35), ack => W_pkt_pointer_1539_delayed_4_0_1564_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3018_elements(40);
      gj_transmitEngineDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	23 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Sample/ack
      -- 
    ack_3204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_1539_delayed_4_0_1564_inst_ack_0, ack => transmitEngineDaemon_CP_3018_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/assign_stmt_1566_Update/ack
      -- 
    ack_3209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_1539_delayed_4_0_1564_inst_ack_1, ack => transmitEngineDaemon_CP_3018_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	29 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	37 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Sample/crr
      -- 
    crr_3217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(38), ack => call_stmt_1573_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(29) & transmitEngineDaemon_CP_3018_elements(33) & transmitEngineDaemon_CP_3018_elements(37) & transmitEngineDaemon_CP_3018_elements(40);
      gj_transmitEngineDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Update/ccr
      -- 
    ccr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(39), ack => call_stmt_1573_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3018_elements(41);
      gj_transmitEngineDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	31 
    -- CP-element group 40: 	35 
    -- CP-element group 40: 	38 
    -- CP-element group 40: 	27 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Sample/cra
      -- 
    cra_3218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1573_call_ack_0, ack => transmitEngineDaemon_CP_3018_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	46 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	22 
    -- CP-element group 41: 	23 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/call_stmt_1573_Update/cca
      -- 
    cca_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1573_call_ack_1, ack => transmitEngineDaemon_CP_3018_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	21 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Sample/req
      -- 
    req_3231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(42), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(21) & transmitEngineDaemon_CP_3018_elements(44);
      gj_transmitEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	17 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Update/req
      -- 
    ack_3232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_ack_0, ack => transmitEngineDaemon_CP_3018_elements(43)); -- 
    req_3236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(43), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_req_1); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_Update/ack
      -- 
    ack_3237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_ack_1, ack => transmitEngineDaemon_CP_3018_elements(44)); -- 
    -- CP-element group 45:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	14 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	15 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitEngineDaemon_CP_3018_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3018_elements(14), ack => transmitEngineDaemon_CP_3018_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	41 
    -- CP-element group 46: 	20 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	11 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1512/do_while_stmt_1522/do_while_stmt_1522_loop_body/$exit
      -- 
    transmitEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3018_elements(44) & transmitEngineDaemon_CP_3018_elements(41) & transmitEngineDaemon_CP_3018_elements(20);
      gj_transmitEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	10 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_exit/$exit
      -- CP-element group 47: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_exit/ack
      -- 
    ack_3242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1522_branch_ack_0, ack => transmitEngineDaemon_CP_3018_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	10 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_taken/$exit
      -- CP-element group 48: 	 branch_block_stmt_1512/do_while_stmt_1522/loop_taken/ack
      -- 
    ack_3246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1522_branch_ack_1, ack => transmitEngineDaemon_CP_3018_elements(48)); -- 
    -- CP-element group 49:  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	8 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	4 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1512/do_while_stmt_1522/$exit
      -- 
    transmitEngineDaemon_CP_3018_elements(49) <= transmitEngineDaemon_CP_3018_elements(8);
    -- CP-element group 50:  merge  branch  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	2 
    -- CP-element group 50: 	4 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	6 
    -- CP-element group 50: 	5 
    -- CP-element group 50:  members (49) 
      -- CP-element group 50: 	 branch_block_stmt_1512/merge_stmt_1513__exit__
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514__entry__
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Sample/req
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Update/req
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/BITSEL_u32_u1_1517_inputs/RPIPE_CONTROL_REGISTER_1515/Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Update/cr
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/BITSEL_u32_u1_1517/SplitProtocol/Update/ca
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Sample/ra
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Update/cr
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/NOT_u1_u1_1518/SplitProtocol/Update/ca
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_1512/NOT_u1_u1_1518_place
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/if_stmt_1514_else_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/merge_stmt_1513_PhiReqMerge
      -- CP-element group 50: 	 branch_block_stmt_1512/merge_stmt_1513_PhiAck/$entry
      -- CP-element group 50: 	 branch_block_stmt_1512/merge_stmt_1513_PhiAck/$exit
      -- CP-element group 50: 	 branch_block_stmt_1512/merge_stmt_1513_PhiAck/dummy
      -- 
    branch_req_3105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3018_elements(50), ack => if_stmt_1514_branch_req_0); -- 
    transmitEngineDaemon_CP_3018_elements(50) <= OrReduce(transmitEngineDaemon_CP_3018_elements(5) & transmitEngineDaemon_CP_3018_elements(2) & transmitEngineDaemon_CP_3018_elements(4));
    transmitEngineDaemon_do_while_stmt_1522_terminator_3247: loop_terminator -- 
      generic map (name => " transmitEngineDaemon_do_while_stmt_1522_terminator_3247", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitEngineDaemon_CP_3018_elements(11),loop_continue => transmitEngineDaemon_CP_3018_elements(48),loop_terminate => transmitEngineDaemon_CP_3018_elements(47),loop_back => transmitEngineDaemon_CP_3018_elements(9),loop_exit => transmitEngineDaemon_CP_3018_elements(8),clk => clk, reset => reset); -- 
    entry_tmerge_3131_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitEngineDaemon_CP_3018_elements(12);
        preds(1)  <= transmitEngineDaemon_CP_3018_elements(13);
        entry_tmerge_3131 : transition_merge -- 
          generic map(name => " entry_tmerge_3131")
          port map (preds => preds, symbol_out => transmitEngineDaemon_CP_3018_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1528_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_1533_wire : std_logic_vector(5 downto 0);
    signal BITSEL_u32_u1_1517_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1582_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1518_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1528_1528_delayed_4_0_1555 : std_logic_vector(0 downto 0);
    signal RPIPE_CONTROL_REGISTER_1515_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1580_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1570_wire : std_logic_vector(35 downto 0);
    signal RPIPE_LAST_READ_TX_QUEUE_INDEX_1526_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1529_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1531_wire : std_logic_vector(31 downto 0);
    signal konst_1510_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1516_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1527_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1530_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1581_wire_constant : std_logic_vector(31 downto 0);
    signal pkt_pointer_1539_delayed_4_0_1566 : std_logic_vector(31 downto 0);
    signal pkt_pointer_1540 : std_logic_vector(31 downto 0);
    signal push_pointer_back_to_free_Q_1560 : std_logic_vector(0 downto 0);
    signal push_status_1573 : std_logic_vector(0 downto 0);
    signal transmitted_flag_1544 : std_logic_vector(0 downto 0);
    signal tx_flag_1540 : std_logic_vector(0 downto 0);
    signal tx_q_index_1524 : std_logic_vector(5 downto 0);
    signal type_cast_1532_wire : std_logic_vector(5 downto 0);
    signal type_cast_1569_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1510_wire_constant <= "000000";
    konst_1516_wire_constant <= "00000000000000000000000000000000";
    konst_1527_wire_constant <= "000001";
    konst_1530_wire_constant <= "00000000000000000000000000000001";
    konst_1581_wire_constant <= "00000000000000000000000000000000";
    type_cast_1569_wire_constant <= "1";
    W_pkt_pointer_1539_delayed_4_0_1564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_pointer_1539_delayed_4_0_1564_inst_req_0;
      W_pkt_pointer_1539_delayed_4_0_1564_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_pointer_1539_delayed_4_0_1564_inst_req_1;
      W_pkt_pointer_1539_delayed_4_0_1564_inst_ack_1<= rack(0);
      W_pkt_pointer_1539_delayed_4_0_1564_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_pointer_1539_delayed_4_0_1564_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_pointer_1540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_pointer_1539_delayed_4_0_1566,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1524
    process(AND_u6_u6_1533_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := AND_u6_u6_1533_wire(5 downto 0);
      tx_q_index_1524 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1532_inst
    process(SUB_u32_u32_1531_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1531_wire(5 downto 0);
      type_cast_1532_wire <= tmp_var; -- 
    end process;
    do_while_stmt_1522_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1582_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1522_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1522_branch_req_0,
          ack0 => do_while_stmt_1522_branch_ack_0,
          ack1 => do_while_stmt_1522_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1514_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1518_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1514_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1514_branch_req_0,
          ack0 => if_stmt_1514_branch_ack_0,
          ack1 => if_stmt_1514_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u6_u6_1528_inst
    process(RPIPE_LAST_READ_TX_QUEUE_INDEX_1526_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_READ_TX_QUEUE_INDEX_1526_wire, konst_1527_wire_constant, tmp_var);
      ADD_u6_u6_1528_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1559_inst
    process(NOT_u1_u1_1528_1528_delayed_4_0_1555, transmitted_flag_1544) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1528_1528_delayed_4_0_1555, transmitted_flag_1544, tmp_var);
      push_pointer_back_to_free_Q_1560 <= tmp_var; --
    end process;
    -- shared split operator group (2) : AND_u6_u6_1533_inst 
    ApIntAnd_group_2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1528_wire & type_cast_1532_wire;
      AND_u6_u6_1533_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1533_inst_req_0;
      AND_u6_u6_1533_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1533_inst_req_1;
      AND_u6_u6_1533_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator BITSEL_u32_u1_1517_inst
    process(RPIPE_CONTROL_REGISTER_1515_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1515_wire, konst_1516_wire_constant, tmp_var);
      BITSEL_u32_u1_1517_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1582_inst
    process(RPIPE_CONTROL_REGISTER_1580_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1580_wire, konst_1581_wire_constant, tmp_var);
      BITSEL_u32_u1_1582_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1518_inst
    process(BITSEL_u32_u1_1517_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1517_wire, tmp_var);
      NOT_u1_u1_1518_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (6) : NOT_u1_u1_1554_inst 
    ApIntNot_group_6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tx_flag_1540;
      NOT_u1_u1_1528_1528_delayed_4_0_1555 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1554_inst_req_0;
      NOT_u1_u1_1554_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1554_inst_req_1;
      NOT_u1_u1_1554_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_6_gI: SplitGuardInterface generic map(name => "ApIntNot_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- binary operator SUB_u32_u32_1531_inst
    process(RPIPE_NUMBER_OF_SERVERS_1529_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1529_wire, konst_1530_wire_constant, tmp_var);
      SUB_u32_u32_1531_wire <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1515_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1580_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1570_wire <= FREE_Q;
    -- read from input-signal LAST_READ_TX_QUEUE_INDEX
    RPIPE_LAST_READ_TX_QUEUE_INDEX_1526_wire <= LAST_READ_TX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_1529_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1509_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_1510_wire_constant;
      LAST_READ_TX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 6),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1576_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= tx_q_index_1524;
      LAST_READ_TX_QUEUE_INDEX_write_1_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_1: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1540_call 
    getTxPacketPointerFromServer_call_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1540_call_req_0;
      call_stmt_1540_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1540_call_req_1;
      call_stmt_1540_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTxPacketPointerFromServer_call_group_0_gI: SplitGuardInterface generic map(name => "getTxPacketPointerFromServer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_q_index_1524;
      pkt_pointer_1540 <= data_out(32 downto 1);
      tx_flag_1540 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 6,
        owidth => 6,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTxPacketPointerFromServer_call_reqs(0),
          ackR => getTxPacketPointerFromServer_call_acks(0),
          dataR => getTxPacketPointerFromServer_call_data(5 downto 0),
          tagR => getTxPacketPointerFromServer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTxPacketPointerFromServer_return_acks(0), -- cross-over
          ackL => getTxPacketPointerFromServer_return_reqs(0), -- cross-over
          dataL => getTxPacketPointerFromServer_return_data(32 downto 0),
          tagL => getTxPacketPointerFromServer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1544_call 
    transmitPacket_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1544_call_req_0;
      call_stmt_1544_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1544_call_req_1;
      call_stmt_1544_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not tx_flag_1540(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      transmitPacket_call_group_1_gI: SplitGuardInterface generic map(name => "transmitPacket_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pkt_pointer_1540;
      transmitted_flag_1544 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => transmitPacket_call_reqs(0),
          ackR => transmitPacket_call_acks(0),
          dataR => transmitPacket_call_data(31 downto 0),
          tagR => transmitPacket_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => transmitPacket_return_acks(0), -- cross-over
          ackL => transmitPacket_return_reqs(0), -- cross-over
          dataL => transmitPacket_return_data(0 downto 0),
          tagL => transmitPacket_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1573_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1573_call_req_0;
      call_stmt_1573_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1573_call_req_1;
      call_stmt_1573_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_1560(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1569_wire_constant & RPIPE_FREE_Q_1570_wire & pkt_pointer_1539_delayed_4_0_1566;
      push_status_1573 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end transmitEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity transmitPacket is -- 
  generic (tag_length : integer); 
  port ( -- 
    packet_pointer : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_call_acks : in   std_logic_vector(1 downto 0);
    accessMemory_call_data : out  std_logic_vector(219 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_return_acks : in   std_logic_vector(1 downto 0);
    accessMemory_return_data : in   std_logic_vector(127 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitPacket;
architecture transmitPacket_arch of transmitPacket is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal packet_pointer_buffer :  std_logic_vector(31 downto 0);
  signal packet_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal transmitPacket_CP_2750_start: Boolean;
  signal transmitPacket_CP_2750_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ncount_down_1457_1427_buf_ack_1 : boolean;
  signal SUB_u8_u8_1426_inst_req_1 : boolean;
  signal ncount_down_1457_1427_buf_req_0 : boolean;
  signal phi_stmt_1422_req_0 : boolean;
  signal ADD_u36_u36_1432_inst_req_1 : boolean;
  signal CONCAT_u65_u73_1451_inst_req_0 : boolean;
  signal phi_stmt_1428_req_0 : boolean;
  signal nmem_addr_1462_1433_buf_ack_1 : boolean;
  signal phi_stmt_1428_req_1 : boolean;
  signal phi_stmt_1422_req_1 : boolean;
  signal SUB_u8_u8_1426_inst_req_0 : boolean;
  signal SUB_u8_u8_1426_inst_ack_1 : boolean;
  signal phi_stmt_1428_ack_0 : boolean;
  signal SUB_u8_u8_1426_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_1451_inst_req_1 : boolean;
  signal phi_stmt_1422_ack_0 : boolean;
  signal CONCAT_u65_u73_1451_inst_ack_1 : boolean;
  signal ncount_down_1457_1427_buf_ack_0 : boolean;
  signal do_while_stmt_1420_branch_ack_0 : boolean;
  signal nmem_addr_1462_1433_buf_ack_0 : boolean;
  signal ADD_u36_u36_1432_inst_ack_1 : boolean;
  signal call_stmt_1407_call_req_0 : boolean;
  signal call_stmt_1444_call_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1445_inst_req_1 : boolean;
  signal call_stmt_1407_call_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1445_inst_ack_1 : boolean;
  signal nmem_addr_1462_1433_buf_req_1 : boolean;
  signal call_stmt_1444_call_req_0 : boolean;
  signal ADD_u36_u36_1432_inst_req_0 : boolean;
  signal nmem_addr_1462_1433_buf_req_0 : boolean;
  signal do_while_stmt_1420_branch_req_0 : boolean;
  signal ADD_u36_u36_1432_inst_ack_0 : boolean;
  signal call_stmt_1444_call_ack_1 : boolean;
  signal ncount_down_1457_1427_buf_req_1 : boolean;
  signal CONCAT_u65_u73_1451_inst_ack_0 : boolean;
  signal call_stmt_1444_call_ack_0 : boolean;
  signal do_while_stmt_1420_branch_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1445_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1445_inst_req_0 : boolean;
  signal call_stmt_1407_call_ack_1 : boolean;
  signal call_stmt_1407_call_req_1 : boolean;
  signal call_stmt_1487_call_req_0 : boolean;
  signal call_stmt_1487_call_ack_0 : boolean;
  signal call_stmt_1487_call_req_1 : boolean;
  signal call_stmt_1487_call_ack_1 : boolean;
  signal CONCAT_u65_u73_1496_inst_req_0 : boolean;
  signal CONCAT_u65_u73_1496_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_1496_inst_req_1 : boolean;
  signal CONCAT_u65_u73_1496_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1490_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1490_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1490_inst_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1490_inst_ack_1 : boolean;
  signal EQ_u8_u1_1504_inst_req_0 : boolean;
  signal EQ_u8_u1_1504_inst_ack_0 : boolean;
  signal EQ_u8_u1_1504_inst_req_1 : boolean;
  signal EQ_u8_u1_1504_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitPacket_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= packet_pointer;
  packet_pointer_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitPacket_CP_2750_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitPacket_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_2750_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitPacket_CP_2750_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_2750_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitPacket_CP_2750: Block -- control-path 
    signal transmitPacket_CP_2750_elements: BooleanArray(81 downto 0);
    -- 
  begin -- 
    transmitPacket_CP_2750_elements(0) <= transmitPacket_CP_2750_start;
    transmitPacket_CP_2750_symbol <= transmitPacket_CP_2750_elements(81);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_update_start_
      -- CP-element group 0: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1394_to_assign_stmt_1415/$entry
      -- CP-element group 0: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Update/ccr
      -- 
    crr_2763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(0), ack => call_stmt_1407_call_req_0); -- 
    ccr_2768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(0), ack => call_stmt_1407_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Sample/cra
      -- CP-element group 1: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_sample_completed_
      -- 
    cra_2764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1407_call_ack_0, ack => transmitPacket_CP_2750_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_1394_to_assign_stmt_1415/$exit
      -- CP-element group 2: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1419/do_while_stmt_1420__entry__
      -- CP-element group 2: 	 branch_block_stmt_1419/branch_block_stmt_1419__entry__
      -- CP-element group 2: 	 branch_block_stmt_1419/$entry
      -- CP-element group 2: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Update/cca
      -- CP-element group 2: 	 assign_stmt_1394_to_assign_stmt_1415/call_stmt_1407_Update/$exit
      -- 
    cca_2769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1407_call_ack_1, ack => transmitPacket_CP_2750_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	72 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	73 
    -- CP-element group 3: 	74 
    -- CP-element group 3: 	79 
    -- CP-element group 3: 	76 
    -- CP-element group 3: 	80 
    -- CP-element group 3:  members (18) 
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505__entry__
      -- CP-element group 3: 	 branch_block_stmt_1419/do_while_stmt_1420__exit__
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/$entry
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Update/cr
      -- 
    crr_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(3), ack => call_stmt_1487_call_req_0); -- 
    ccr_2974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(3), ack => call_stmt_1487_call_req_1); -- 
    cr_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(3), ack => CONCAT_u65_u73_1496_inst_req_1); -- 
    rr_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(3), ack => EQ_u8_u1_1504_inst_req_0); -- 
    cr_3016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(3), ack => EQ_u8_u1_1504_inst_req_1); -- 
    transmitPacket_CP_2750_elements(3) <= transmitPacket_CP_2750_elements(72);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420__entry__
      -- CP-element group 4: 	 branch_block_stmt_1419/do_while_stmt_1420/$entry
      -- 
    transmitPacket_CP_2750_elements(4) <= transmitPacket_CP_2750_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	72 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420__exit__
      -- 
    -- Element group transmitPacket_CP_2750_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_back
      -- 
    -- Element group transmitPacket_CP_2750_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	70 
    -- CP-element group 7: 	71 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1419/do_while_stmt_1420/condition_done
      -- CP-element group 7: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_taken/$entry
      -- 
    transmitPacket_CP_2750_elements(7) <= transmitPacket_CP_2750_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	69 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_body_done
      -- 
    transmitPacket_CP_2750_elements(8) <= transmitPacket_CP_2750_elements(69);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	42 
    -- CP-element group 9: 	22 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/back_edge_to_loop_body
      -- 
    transmitPacket_CP_2750_elements(9) <= transmitPacket_CP_2750_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	44 
    -- CP-element group 10: 	24 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/first_time_through_loop_body
      -- 
    transmitPacket_CP_2750_elements(10) <= transmitPacket_CP_2750_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	68 
    -- CP-element group 11: 	38 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/$entry
      -- 
    -- Element group transmitPacket_CP_2750_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	68 
    -- CP-element group 12: 	21 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/condition_evaluated
      -- 
    condition_evaluated_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(12), ack => do_while_stmt_1420_branch_req_0); -- 
    transmitPacket_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(16) & transmitPacket_CP_2750_elements(68) & transmitPacket_CP_2750_elements(21);
      gj_transmitPacket_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	17 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	39 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_sample_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/aggregated_phi_sample_req
      -- 
    transmitPacket_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(37) & transmitPacket_CP_2750_elements(17) & transmitPacket_CP_2750_elements(16);
      gj_transmitPacket_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	40 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	69 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_sample_completed_
      -- 
    transmitPacket_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(19) & transmitPacket_CP_2750_elements(40);
      gj_transmitPacket_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	38 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/aggregated_phi_update_req
      -- CP-element group 15: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_update_start__ps
      -- 
    transmitPacket_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(18) & transmitPacket_CP_2750_elements(38);
      gj_transmitPacket_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	21 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/aggregated_phi_update_ack
      -- 
    transmitPacket_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(41) & transmitPacket_CP_2750_elements(21);
      gj_transmitPacket_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_sample_start_
      -- 
    transmitPacket_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(11) & transmitPacket_CP_2750_elements(14);
      gj_transmitPacket_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_update_start_
      -- 
    transmitPacket_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(11) & transmitPacket_CP_2750_elements(21);
      gj_transmitPacket_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_2750_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_update_start__ps
      -- 
    transmitPacket_CP_2750_elements(20) <= transmitPacket_CP_2750_elements(15);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	12 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_update_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_update_completed_
      -- 
    -- Element group transmitPacket_CP_2750_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	9 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_loopback_trigger
      -- 
    transmitPacket_CP_2750_elements(22) <= transmitPacket_CP_2750_elements(9);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_loopback_sample_req
      -- CP-element group 23: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_loopback_sample_req_ps
      -- 
    phi_stmt_1422_loopback_sample_req_2808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1422_loopback_sample_req_2808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(23), ack => phi_stmt_1422_req_1); -- 
    -- Element group transmitPacket_CP_2750_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	10 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_entry_trigger
      -- 
    transmitPacket_CP_2750_elements(24) <= transmitPacket_CP_2750_elements(10);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_entry_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_entry_sample_req_ps
      -- 
    phi_stmt_1422_entry_sample_req_2811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1422_entry_sample_req_2811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(25), ack => phi_stmt_1422_req_0); -- 
    -- Element group transmitPacket_CP_2750_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_phi_mux_ack
      -- CP-element group 26: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1422_phi_mux_ack_ps
      -- 
    phi_stmt_1422_phi_mux_ack_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1422_ack_0, ack => transmitPacket_CP_2750_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_2750_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_update_start__ps
      -- 
    -- Element group transmitPacket_CP_2750_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_sample_start_
      -- 
    rr_2827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(29), ack => SUB_u8_u8_1426_inst_req_0); -- 
    transmitPacket_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(27) & transmitPacket_CP_2750_elements(31);
      gj_transmitPacket_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Update/$entry
      -- 
    cr_2832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(30), ack => SUB_u8_u8_1426_inst_req_1); -- 
    transmitPacket_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(28) & transmitPacket_CP_2750_elements(32);
      gj_transmitPacket_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_sample_completed_
      -- 
    ra_2828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u8_u8_1426_inst_ack_0, ack => transmitPacket_CP_2750_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/SUB_u8_u8_1426_update_completed__ps
      -- 
    ca_2833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u8_u8_1426_inst_ack_1, ack => transmitPacket_CP_2750_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Sample/req
      -- CP-element group 33: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Sample/$entry
      -- 
    req_2845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(33), ack => ncount_down_1457_1427_buf_req_0); -- 
    -- Element group transmitPacket_CP_2750_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Update/req
      -- CP-element group 34: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Update/$entry
      -- 
    req_2850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(34), ack => ncount_down_1457_1427_buf_req_1); -- 
    -- Element group transmitPacket_CP_2750_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Sample/ack
      -- 
    ack_2846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1457_1427_buf_ack_0, ack => transmitPacket_CP_2750_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_ncount_down_1427_Update/$exit
      -- 
    ack_2851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1457_1427_buf_ack_1, ack => transmitPacket_CP_2750_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_sample_start_
      -- 
    transmitPacket_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(11) & transmitPacket_CP_2750_elements(14);
      gj_transmitPacket_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	59 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	15 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_update_start_
      -- 
    transmitPacket_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(11) & transmitPacket_CP_2750_elements(41) & transmitPacket_CP_2750_elements(59);
      gj_transmitPacket_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	13 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_sample_start__ps
      -- 
    transmitPacket_CP_2750_elements(39) <= transmitPacket_CP_2750_elements(13);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	14 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_2750_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	57 
    -- CP-element group 41: 	16 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	38 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_update_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_update_completed_
      -- 
    -- Element group transmitPacket_CP_2750_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	9 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_loopback_trigger
      -- 
    transmitPacket_CP_2750_elements(42) <= transmitPacket_CP_2750_elements(9);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_loopback_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_loopback_sample_req
      -- 
    phi_stmt_1428_loopback_sample_req_2862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1428_loopback_sample_req_2862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(43), ack => phi_stmt_1428_req_1); -- 
    -- Element group transmitPacket_CP_2750_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	10 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_entry_trigger
      -- 
    transmitPacket_CP_2750_elements(44) <= transmitPacket_CP_2750_elements(10);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_entry_sample_req_ps
      -- CP-element group 45: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_entry_sample_req
      -- 
    phi_stmt_1428_entry_sample_req_2865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1428_entry_sample_req_2865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(45), ack => phi_stmt_1428_req_0); -- 
    -- Element group transmitPacket_CP_2750_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/phi_stmt_1428_phi_mux_ack_ps
      -- 
    phi_stmt_1428_phi_mux_ack_2868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1428_ack_0, ack => transmitPacket_CP_2750_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_2750_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_update_start__ps
      -- 
    -- Element group transmitPacket_CP_2750_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Sample/rr
      -- 
    rr_2881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(49), ack => ADD_u36_u36_1432_inst_req_0); -- 
    transmitPacket_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(47) & transmitPacket_CP_2750_elements(51);
      gj_transmitPacket_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Update/cr
      -- CP-element group 50: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_update_start_
      -- 
    cr_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(50), ack => ADD_u36_u36_1432_inst_req_1); -- 
    transmitPacket_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(48) & transmitPacket_CP_2750_elements(52);
      gj_transmitPacket_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Sample/ra
      -- 
    ra_2882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1432_inst_ack_0, ack => transmitPacket_CP_2750_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/ADD_u36_u36_1432_update_completed_
      -- 
    ca_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1432_inst_ack_1, ack => transmitPacket_CP_2750_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Sample/req
      -- CP-element group 53: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_sample_start__ps
      -- 
    req_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(53), ack => nmem_addr_1462_1433_buf_req_0); -- 
    -- Element group transmitPacket_CP_2750_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Update/req
      -- CP-element group 54: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_update_start__ps
      -- 
    req_2904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(54), ack => nmem_addr_1462_1433_buf_req_1); -- 
    -- Element group transmitPacket_CP_2750_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Sample/$exit
      -- 
    ack_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1462_1433_buf_ack_0, ack => transmitPacket_CP_2750_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/R_nmem_addr_1433_update_completed_
      -- 
    ack_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1462_1433_buf_ack_1, ack => transmitPacket_CP_2750_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Sample/crr
      -- 
    crr_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(57), ack => call_stmt_1444_call_req_0); -- 
    transmitPacket_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(41) & transmitPacket_CP_2750_elements(59);
      gj_transmitPacket_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	63 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Update/ccr
      -- 
    ccr_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(58), ack => call_stmt_1444_call_req_1); -- 
    transmitPacket_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(60) & transmitPacket_CP_2750_elements(63);
      gj_transmitPacket_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: 	38 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Sample/cra
      -- 
    cra_2915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1444_call_ack_0, ack => transmitPacket_CP_2750_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/call_stmt_1444_Update/cca
      -- 
    cca_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1444_call_ack_1, ack => transmitPacket_CP_2750_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Sample/$entry
      -- 
    rr_2928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(61), ack => CONCAT_u65_u73_1451_inst_req_0); -- 
    transmitPacket_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(60) & transmitPacket_CP_2750_elements(63);
      gj_transmitPacket_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	66 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Update/$entry
      -- 
    cr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(62), ack => CONCAT_u65_u73_1451_inst_req_1); -- 
    transmitPacket_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(66) & transmitPacket_CP_2750_elements(64);
      gj_transmitPacket_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	58 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Sample/ra
      -- 
    ra_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1451_inst_ack_0, ack => transmitPacket_CP_2750_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/CONCAT_u65_u73_1451_update_completed_
      -- 
    ca_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1451_inst_ack_1, ack => transmitPacket_CP_2750_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_sample_start_
      -- 
    req_2942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(65), ack => WPIPE_nic_to_mac_transmit_pipe_1445_inst_req_0); -- 
    transmitPacket_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(64) & transmitPacket_CP_2750_elements(67);
      gj_transmitPacket_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	62 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Update/req
      -- CP-element group 66: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_update_start_
      -- CP-element group 66: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_sample_completed_
      -- 
    ack_2943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1445_inst_ack_0, ack => transmitPacket_CP_2750_elements(66)); -- 
    req_2947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(66), ack => WPIPE_nic_to_mac_transmit_pipe_1445_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/WPIPE_nic_to_mac_transmit_pipe_1445_update_completed_
      -- 
    ack_2948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1445_inst_ack_1, ack => transmitPacket_CP_2750_elements(67)); -- 
    -- CP-element group 68:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	11 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	12 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitPacket_CP_2750_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => transmitPacket_CP_2750_elements(11), ack => transmitPacket_CP_2750_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	14 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	8 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1419/do_while_stmt_1420/do_while_stmt_1420_loop_body/$exit
      -- 
    transmitPacket_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(67) & transmitPacket_CP_2750_elements(14);
      gj_transmitPacket_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	7 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_exit/ack
      -- CP-element group 70: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_exit/$exit
      -- 
    ack_2953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1420_branch_ack_0, ack => transmitPacket_CP_2750_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	7 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_taken/ack
      -- CP-element group 71: 	 branch_block_stmt_1419/do_while_stmt_1420/loop_taken/$exit
      -- 
    ack_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1420_branch_ack_1, ack => transmitPacket_CP_2750_elements(71)); -- 
    -- CP-element group 72:  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	5 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	3 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1419/do_while_stmt_1420/$exit
      -- 
    transmitPacket_CP_2750_elements(72) <= transmitPacket_CP_2750_elements(5);
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	3 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Sample/cra
      -- 
    cra_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1487_call_ack_0, ack => transmitPacket_CP_2750_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	3 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/call_stmt_1487_Update/cca
      -- CP-element group 74: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Sample/rr
      -- 
    cca_2975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1487_call_ack_1, ack => transmitPacket_CP_2750_elements(74)); -- 
    rr_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(74), ack => CONCAT_u65_u73_1496_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Sample/ra
      -- 
    ra_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1496_inst_ack_0, ack => transmitPacket_CP_2750_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	3 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/CONCAT_u65_u73_1496_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Sample/req
      -- 
    ca_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1496_inst_ack_1, ack => transmitPacket_CP_2750_elements(76)); -- 
    req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(76), ack => WPIPE_nic_to_mac_transmit_pipe_1490_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Update/req
      -- 
    ack_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1490_inst_ack_0, ack => transmitPacket_CP_2750_elements(77)); -- 
    req_3002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2750_elements(77), ack => WPIPE_nic_to_mac_transmit_pipe_1490_inst_req_1); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	81 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/WPIPE_nic_to_mac_transmit_pipe_1490_Update/ack
      -- 
    ack_3003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1490_inst_ack_1, ack => transmitPacket_CP_2750_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	3 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Sample/ra
      -- 
    ra_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_1504_inst_ack_0, ack => transmitPacket_CP_2750_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	3 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/EQ_u8_u1_1504_Update/ca
      -- 
    ca_3017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u8_u1_1504_inst_ack_1, ack => transmitPacket_CP_2750_elements(80)); -- 
    -- CP-element group 81:  join  transition  place  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	78 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1419/branch_block_stmt_1419__exit__
      -- CP-element group 81: 	 $exit
      -- CP-element group 81: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505__exit__
      -- CP-element group 81: 	 branch_block_stmt_1419/call_stmt_1487_to_assign_stmt_1505/$exit
      -- CP-element group 81: 	 branch_block_stmt_1419/$exit
      -- 
    transmitPacket_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2750_elements(78) & transmitPacket_CP_2750_elements(80);
      gj_transmitPacket_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2750_elements(81), clk => clk, reset => reset); --
    end block;
    transmitPacket_do_while_stmt_1420_terminator_2958: loop_terminator -- 
      generic map (name => " transmitPacket_do_while_stmt_1420_terminator_2958", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitPacket_CP_2750_elements(8),loop_continue => transmitPacket_CP_2750_elements(71),loop_terminate => transmitPacket_CP_2750_elements(70),loop_back => transmitPacket_CP_2750_elements(6),loop_exit => transmitPacket_CP_2750_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_1422_phi_seq_2852_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_2750_elements(24);
      transmitPacket_CP_2750_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_2750_elements(31);
      transmitPacket_CP_2750_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_2750_elements(32);
      transmitPacket_CP_2750_elements(25) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_2750_elements(22);
      transmitPacket_CP_2750_elements(33)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_2750_elements(35);
      transmitPacket_CP_2750_elements(34)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_2750_elements(36);
      transmitPacket_CP_2750_elements(23) <= phi_mux_reqs(1);
      phi_stmt_1422_phi_seq_2852 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1422_phi_seq_2852") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_2750_elements(13), 
          phi_sample_ack => transmitPacket_CP_2750_elements(19), 
          phi_update_req => transmitPacket_CP_2750_elements(20), 
          phi_update_ack => transmitPacket_CP_2750_elements(21), 
          phi_mux_ack => transmitPacket_CP_2750_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1428_phi_seq_2906_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_2750_elements(44);
      transmitPacket_CP_2750_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_2750_elements(51);
      transmitPacket_CP_2750_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_2750_elements(52);
      transmitPacket_CP_2750_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_2750_elements(42);
      transmitPacket_CP_2750_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_2750_elements(55);
      transmitPacket_CP_2750_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_2750_elements(56);
      transmitPacket_CP_2750_elements(43) <= phi_mux_reqs(1);
      phi_stmt_1428_phi_seq_2906 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1428_phi_seq_2906") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_2750_elements(39), 
          phi_sample_ack => transmitPacket_CP_2750_elements(40), 
          phi_update_req => transmitPacket_CP_2750_elements(15), 
          phi_update_ack => transmitPacket_CP_2750_elements(41), 
          phi_mux_ack => transmitPacket_CP_2750_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2794_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitPacket_CP_2750_elements(9);
        preds(1)  <= transmitPacket_CP_2750_elements(10);
        entry_tmerge_2794 : transition_merge -- 
          generic map(name => " entry_tmerge_2794")
          port map (preds => preds, symbol_out => transmitPacket_CP_2750_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1432_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u1_u65_1449_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u1_u65_1494_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u32_u36_1392_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u65_u73_1451_wire : std_logic_vector(72 downto 0);
    signal CONCAT_u65_u73_1496_wire : std_logic_vector(72 downto 0);
    signal R_FULL_BYTE_MASK_1402_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1439_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1450_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1482_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u36_u36_1502_wire : std_logic_vector(35 downto 0);
    signal SUB_u8_u8_1426_wire : std_logic_vector(7 downto 0);
    signal control_data_1407 : std_logic_vector(63 downto 0);
    signal control_data_addr_1394 : std_logic_vector(35 downto 0);
    signal count_down_1422 : std_logic_vector(7 downto 0);
    signal data_1444 : std_logic_vector(63 downto 0);
    signal konst_1425_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1431_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1455_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1460_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1471_wire_constant : std_logic_vector(7 downto 0);
    signal last_tkeep_1415 : std_logic_vector(7 downto 0);
    signal last_word_1487 : std_logic_vector(63 downto 0);
    signal mem_addr_1428 : std_logic_vector(35 downto 0);
    signal ncount_down_1457 : std_logic_vector(7 downto 0);
    signal ncount_down_1457_1427_buffered : std_logic_vector(7 downto 0);
    signal nmem_addr_1462 : std_logic_vector(35 downto 0);
    signal nmem_addr_1462_1433_buffered : std_logic_vector(35 downto 0);
    signal not_last_word_1473 : std_logic_vector(0 downto 0);
    signal packet_size_1411 : std_logic_vector(7 downto 0);
    signal slice_1389_wire : std_logic_vector(31 downto 0);
    signal type_cast_1391_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1399_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1401_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1405_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1436_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1442_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1447_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1479_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1481_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1485_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1492_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1503_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_1402_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1439_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1450_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1482_wire_constant <= "11111111";
    konst_1425_wire_constant <= "00010000";
    konst_1431_wire_constant <= "000000000000000000000000000000011000";
    konst_1455_wire_constant <= "00001000";
    konst_1460_wire_constant <= "000000000000000000000000000000001000";
    konst_1471_wire_constant <= "00001000";
    type_cast_1391_wire_constant <= "0000";
    type_cast_1399_wire_constant <= "0";
    type_cast_1401_wire_constant <= "1";
    type_cast_1405_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1436_wire_constant <= "0";
    type_cast_1438_wire_constant <= "1";
    type_cast_1442_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1447_wire_constant <= "0";
    type_cast_1479_wire_constant <= "0";
    type_cast_1481_wire_constant <= "1";
    type_cast_1485_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1492_wire_constant <= "1";
    phi_stmt_1422: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SUB_u8_u8_1426_wire & ncount_down_1457_1427_buffered;
      req <= phi_stmt_1422_req_0 & phi_stmt_1422_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1422",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1422_ack_0,
          idata => idata,
          odata => count_down_1422,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1422
    phi_stmt_1428: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_1432_wire & nmem_addr_1462_1433_buffered;
      req <= phi_stmt_1428_req_0 & phi_stmt_1428_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1428",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1428_ack_0,
          idata => idata,
          odata => mem_addr_1428,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1428
    -- flow-through slice operator slice_1389_inst
    slice_1389_wire <= packet_pointer_buffer(31 downto 0);
    -- flow-through slice operator slice_1410_inst
    packet_size_1411 <= control_data_1407(15 downto 8);
    -- flow-through slice operator slice_1414_inst
    last_tkeep_1415 <= control_data_1407(7 downto 0);
    ncount_down_1457_1427_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_down_1457_1427_buf_req_0;
      ncount_down_1457_1427_buf_ack_0<= wack(0);
      rreq(0) <= ncount_down_1457_1427_buf_req_1;
      ncount_down_1457_1427_buf_ack_1<= rack(0);
      ncount_down_1457_1427_buf : InterlockBuffer generic map ( -- 
        name => "ncount_down_1457_1427_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_down_1457,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_down_1457_1427_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmem_addr_1462_1433_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmem_addr_1462_1433_buf_req_0;
      nmem_addr_1462_1433_buf_ack_0<= wack(0);
      rreq(0) <= nmem_addr_1462_1433_buf_req_1;
      nmem_addr_1462_1433_buf_ack_1<= rack(0);
      nmem_addr_1462_1433_buf : InterlockBuffer generic map ( -- 
        name => "nmem_addr_1462_1433_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_1462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmem_addr_1462_1433_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1393_inst
    process(CONCAT_u32_u36_1392_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 35 downto 0) := CONCAT_u32_u36_1392_wire(35 downto 0);
      control_data_addr_1394 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1503_inst
    process(SUB_u36_u36_1502_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u36_u36_1502_wire(7 downto 0);
      type_cast_1503_wire <= tmp_var; -- 
    end process;
    do_while_stmt_1420_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= not_last_word_1473;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1420_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1420_branch_req_0,
          ack0 => do_while_stmt_1420_branch_ack_0,
          ack1 => do_while_stmt_1420_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1432_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= control_data_addr_1394;
      ADD_u36_u36_1432_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1432_inst_req_0;
      ADD_u36_u36_1432_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1432_inst_req_1;
      ADD_u36_u36_1432_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000011000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_1461_inst
    process(mem_addr_1428) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mem_addr_1428, konst_1460_wire_constant, tmp_var);
      nmem_addr_1462 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_1449_inst
    process(type_cast_1447_wire_constant, data_1444) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1447_wire_constant, data_1444, tmp_var);
      CONCAT_u1_u65_1449_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_1494_inst
    process(type_cast_1492_wire_constant, last_word_1487) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1492_wire_constant, last_word_1487, tmp_var);
      CONCAT_u1_u65_1494_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u36_1392_inst
    process(slice_1389_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1389_wire, type_cast_1391_wire_constant, tmp_var);
      CONCAT_u32_u36_1392_wire <= tmp_var; --
    end process;
    -- shared split operator group (5) : CONCAT_u65_u73_1451_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_1449_wire;
      CONCAT_u65_u73_1451_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_1451_inst_req_0;
      CONCAT_u65_u73_1451_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_1451_inst_req_1;
      CONCAT_u65_u73_1451_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : CONCAT_u65_u73_1496_inst 
    ApConcat_group_6: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_1494_wire & last_tkeep_1415;
      CONCAT_u65_u73_1496_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_1496_inst_req_0;
      CONCAT_u65_u73_1496_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_1496_inst_req_1;
      CONCAT_u65_u73_1496_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_6_gI: SplitGuardInterface generic map(name => "ApConcat_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : EQ_u8_u1_1504_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_1411 & type_cast_1503_wire;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u8_u1_1504_inst_req_0;
      EQ_u8_u1_1504_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u8_u1_1504_inst_req_1;
      EQ_u8_u1_1504_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u36_u36_1502_inst
    process(nmem_addr_1462, control_data_addr_1394) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(nmem_addr_1462, control_data_addr_1394, tmp_var);
      SUB_u36_u36_1502_wire <= tmp_var; --
    end process;
    -- shared split operator group (9) : SUB_u8_u8_1426_inst 
    ApIntSub_group_9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_1411;
      SUB_u8_u8_1426_wire <= data_out(7 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u8_u8_1426_inst_req_0;
      SUB_u8_u8_1426_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u8_u8_1426_inst_req_1;
      SUB_u8_u8_1426_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_9_gI: SplitGuardInterface generic map(name => "ApIntSub_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00010000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- binary operator SUB_u8_u8_1456_inst
    process(count_down_1422) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_1422, konst_1455_wire_constant, tmp_var);
      ncount_down_1457 <= tmp_var; --
    end process;
    -- binary operator UGT_u8_u1_1472_inst
    process(ncount_down_1457) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ncount_down_1457, konst_1471_wire_constant, tmp_var);
      not_last_word_1473 <= tmp_var; --
    end process;
    -- shared outport operator group (0) : WPIPE_nic_to_mac_transmit_pipe_1445_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1445_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_1445_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1445_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_1445_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_1451_wire;
      nic_to_mac_transmit_pipe_write_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(1),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(1),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 73),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_to_mac_transmit_pipe_1490_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1490_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_1490_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1490_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_1490_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_1496_wire;
      nic_to_mac_transmit_pipe_write_1_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1407_call call_stmt_1487_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1407_call_req_0;
      reqL_unguarded(0) <= call_stmt_1487_call_req_0;
      call_stmt_1407_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1487_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1407_call_req_1;
      reqR_unguarded(0) <= call_stmt_1487_call_req_1;
      call_stmt_1407_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1487_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1399_wire_constant & type_cast_1401_wire_constant & R_FULL_BYTE_MASK_1402_wire_constant & control_data_addr_1394 & type_cast_1405_wire_constant & type_cast_1479_wire_constant & type_cast_1481_wire_constant & R_FULL_BYTE_MASK_1482_wire_constant & nmem_addr_1462 & type_cast_1485_wire_constant;
      control_data_1407 <= data_out(127 downto 64);
      last_word_1487 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(1),
          ackR => accessMemory_call_acks(1),
          dataR => accessMemory_call_data(219 downto 110),
          tagR => accessMemory_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(1), -- cross-over
          ackL => accessMemory_return_reqs(1), -- cross-over
          dataL => accessMemory_return_data(127 downto 64),
          tagL => accessMemory_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1444_call 
    accessMemory_call_group_1: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1444_call_req_0;
      call_stmt_1444_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1444_call_req_1;
      call_stmt_1444_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1436_wire_constant & type_cast_1438_wire_constant & R_FULL_BYTE_MASK_1439_wire_constant & mem_addr_1428 & type_cast_1442_wire_constant;
      data_1444 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end transmitPacket_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeControlInformationToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buffer_pointer : in  std_logic_vector(35 downto 0);
    packet_size : in  std_logic_vector(7 downto 0);
    last_keep : in  std_logic_vector(7 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeControlInformationToMem;
architecture writeControlInformationToMem_arch of writeControlInformationToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 52)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buffer_pointer_update_enable: Boolean;
  signal packet_size_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  -- output port buffer signals
  signal writeControlInformationToMem_CP_980_start: Boolean;
  signal writeControlInformationToMem_CP_980_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_683_call_ack_1 : boolean;
  signal call_stmt_683_call_req_1 : boolean;
  signal call_stmt_683_call_ack_0 : boolean;
  signal call_stmt_683_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeControlInformationToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 52) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buffer_pointer;
  base_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(43 downto 36) <= packet_size;
  packet_size_buffer <= in_buffer_data_out(43 downto 36);
  in_buffer_data_in(51 downto 44) <= last_keep;
  last_keep_buffer <= in_buffer_data_out(51 downto 44);
  in_buffer_data_in(tag_length + 51 downto 52) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 51 downto 52);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeControlInformationToMem_CP_980_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeControlInformationToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_980_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_980_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_980_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeControlInformationToMem_CP_980: Block -- control-path 
    signal writeControlInformationToMem_CP_980_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeControlInformationToMem_CP_980_elements(0) <= writeControlInformationToMem_CP_980_start;
    writeControlInformationToMem_CP_980_symbol <= writeControlInformationToMem_CP_980_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_update_start_
      -- CP-element group 0: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Update/ccr
      -- CP-element group 0: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Update/$entry
      -- CP-element group 0: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_sample_start_
      -- CP-element group 0: 	 assign_stmt_674_to_call_stmt_683/$entry
      -- CP-element group 0: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Sample/crr
      -- CP-element group 0: 	 $entry
      -- 
    crr_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_980_elements(0), ack => call_stmt_683_call_req_0); -- 
    ccr_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_980_elements(0), ack => call_stmt_683_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_sample_completed_
      -- CP-element group 1: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Sample/cra
      -- CP-element group 1: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Sample/$exit
      -- 
    cra_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_683_call_ack_0, ack => writeControlInformationToMem_CP_980_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_update_completed_
      -- CP-element group 2: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Update/cca
      -- CP-element group 2: 	 assign_stmt_674_to_call_stmt_683/call_stmt_683_Update/$exit
      -- CP-element group 2: 	 assign_stmt_674_to_call_stmt_683/$exit
      -- CP-element group 2: 	 $exit
      -- 
    cca_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_683_call_ack_1, ack => writeControlInformationToMem_CP_980_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_672_wire : std_logic_vector(15 downto 0);
    signal R_FULL_BYTE_MASK_679_wire_constant : std_logic_vector(7 downto 0);
    signal control_data_674 : std_logic_vector(63 downto 0);
    signal ignore_return_683 : std_logic_vector(63 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_679_wire_constant <= "11111111";
    type_cast_676_wire_constant <= "0";
    type_cast_678_wire_constant <= "0";
    -- interlock type_cast_673_inst
    process(CONCAT_u8_u16_672_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := CONCAT_u8_u16_672_wire(15 downto 0);
      control_data_674 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u8_u16_672_inst
    process(packet_size_buffer, last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(packet_size_buffer, last_keep_buffer, tmp_var);
      CONCAT_u8_u16_672_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_683_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_683_call_req_0;
      call_stmt_683_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_683_call_req_1;
      call_stmt_683_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_676_wire_constant & type_cast_678_wire_constant & R_FULL_BYTE_MASK_679_wire_constant & base_buffer_pointer_buffer & control_data_674;
      ignore_return_683 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeControlInformationToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writeEthernetHeaderToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    buf_pointer : in  std_logic_vector(35 downto 0);
    buf_position : out  std_logic_vector(35 downto 0);
    nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeEthernetHeaderToMem;
architecture writeEthernetHeaderToMem_arch of writeEthernetHeaderToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal buf_position_buffer :  std_logic_vector(35 downto 0);
  signal buf_position_update_enable: Boolean;
  signal writeEthernetHeaderToMem_CP_681_start: Boolean;
  signal writeEthernetHeaderToMem_CP_681_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_536_branch_req_0 : boolean;
  signal phi_stmt_538_req_1 : boolean;
  signal phi_stmt_538_req_0 : boolean;
  signal phi_stmt_538_ack_0 : boolean;
  signal ADD_u36_u36_542_inst_req_0 : boolean;
  signal ADD_u36_u36_542_inst_ack_0 : boolean;
  signal ADD_u36_u36_542_inst_req_1 : boolean;
  signal ADD_u36_u36_542_inst_ack_1 : boolean;
  signal nbuf_position_582_543_buf_req_0 : boolean;
  signal nbuf_position_582_543_buf_ack_0 : boolean;
  signal nbuf_position_582_543_buf_req_1 : boolean;
  signal nbuf_position_582_543_buf_ack_1 : boolean;
  signal phi_stmt_544_req_1 : boolean;
  signal phi_stmt_544_req_0 : boolean;
  signal phi_stmt_544_ack_0 : boolean;
  signal nI_577_548_buf_req_0 : boolean;
  signal nI_577_548_buf_ack_0 : boolean;
  signal nI_577_548_buf_req_1 : boolean;
  signal nI_577_548_buf_ack_1 : boolean;
  signal RPIPE_nic_rx_to_header_551_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_header_551_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_551_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_header_551_inst_ack_1 : boolean;
  signal call_stmt_572_call_req_0 : boolean;
  signal call_stmt_572_call_ack_0 : boolean;
  signal call_stmt_572_call_req_1 : boolean;
  signal call_stmt_572_call_ack_1 : boolean;
  signal do_while_stmt_536_branch_ack_0 : boolean;
  signal do_while_stmt_536_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeEthernetHeaderToMem_CP_681_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(35 downto 0) <= buf_position_buffer;
  buf_position <= out_buffer_data_out(35 downto 0);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_681_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_681_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_681_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeEthernetHeaderToMem_CP_681: Block -- control-path 
    signal writeEthernetHeaderToMem_CP_681_elements: BooleanArray(66 downto 0);
    -- 
  begin -- 
    writeEthernetHeaderToMem_CP_681_elements(0) <= writeEthernetHeaderToMem_CP_681_start;
    writeEthernetHeaderToMem_CP_681_symbol <= writeEthernetHeaderToMem_CP_681_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_535/$entry
      -- CP-element group 0: 	 branch_block_stmt_535/branch_block_stmt_535__entry__
      -- CP-element group 0: 	 branch_block_stmt_535/do_while_stmt_536__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	66 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_535/$exit
      -- CP-element group 1: 	 branch_block_stmt_535/branch_block_stmt_535__exit__
      -- CP-element group 1: 	 branch_block_stmt_535/do_while_stmt_536__exit__
      -- 
    writeEthernetHeaderToMem_CP_681_elements(1) <= writeEthernetHeaderToMem_CP_681_elements(66);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_535/do_while_stmt_536/$entry
      -- CP-element group 2: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536__entry__
      -- 
    writeEthernetHeaderToMem_CP_681_elements(2) <= writeEthernetHeaderToMem_CP_681_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	66 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536__exit__
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_535/do_while_stmt_536/loop_back
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	64 
    -- CP-element group 5: 	65 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_535/do_while_stmt_536/condition_done
      -- CP-element group 5: 	 branch_block_stmt_535/do_while_stmt_536/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_535/do_while_stmt_536/loop_taken/$entry
      -- 
    writeEthernetHeaderToMem_CP_681_elements(5) <= writeEthernetHeaderToMem_CP_681_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	63 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_535/do_while_stmt_536/loop_body_done
      -- 
    writeEthernetHeaderToMem_CP_681_elements(6) <= writeEthernetHeaderToMem_CP_681_elements(63);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	40 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/back_edge_to_loop_body
      -- 
    writeEthernetHeaderToMem_CP_681_elements(7) <= writeEthernetHeaderToMem_CP_681_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	42 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/first_time_through_loop_body
      -- 
    writeEthernetHeaderToMem_CP_681_elements(8) <= writeEthernetHeaderToMem_CP_681_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	62 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_549_sample_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	62 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/condition_evaluated
      -- 
    condition_evaluated_705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(10), ack => do_while_stmt_536_branch_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(14) & writeEthernetHeaderToMem_CP_681_elements(62);
      gj_writeEthernetHeaderToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	54 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_sample_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(9) & writeEthernetHeaderToMem_CP_681_elements(15) & writeEthernetHeaderToMem_CP_681_elements(34) & writeEthernetHeaderToMem_CP_681_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	56 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	63 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_549_sample_completed_
      -- 
    writeEthernetHeaderToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(17) & writeEthernetHeaderToMem_CP_681_elements(37) & writeEthernetHeaderToMem_CP_681_elements(56);
      gj_writeEthernetHeaderToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	53 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	55 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_update_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(16) & writeEthernetHeaderToMem_CP_681_elements(35) & writeEthernetHeaderToMem_CP_681_elements(53);
      gj_writeEthernetHeaderToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	57 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/aggregated_phi_update_ack
      -- 
    writeEthernetHeaderToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(18) & writeEthernetHeaderToMem_CP_681_elements(39) & writeEthernetHeaderToMem_CP_681_elements(57);
      gj_writeEthernetHeaderToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(9) & writeEthernetHeaderToMem_CP_681_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(9) & writeEthernetHeaderToMem_CP_681_elements(18);
      gj_writeEthernetHeaderToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_681_elements(19) <= writeEthernetHeaderToMem_CP_681_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_loopback_sample_req_ps
      -- 
    phi_stmt_538_loopback_sample_req_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_538_loopback_sample_req_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(20), ack => phi_stmt_538_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_681_elements(21) <= writeEthernetHeaderToMem_CP_681_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_entry_sample_req_ps
      -- 
    phi_stmt_538_entry_sample_req_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_538_entry_sample_req_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(22), ack => phi_stmt_538_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_538_phi_mux_ack_ps
      -- 
    phi_stmt_538_phi_mux_ack_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_538_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Sample/rr
      -- 
    rr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(26), ack => ADD_u36_u36_542_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(24) & writeEthernetHeaderToMem_CP_681_elements(28);
      gj_writeEthernetHeaderToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_update_start_
      -- CP-element group 27: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Update/cr
      -- 
    cr_744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(27), ack => ADD_u36_u36_542_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(25) & writeEthernetHeaderToMem_CP_681_elements(29);
      gj_writeEthernetHeaderToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Sample/ra
      -- 
    ra_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_542_inst_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/ADD_u36_u36_542_Update/ca
      -- 
    ca_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_542_inst_ack_1, ack => writeEthernetHeaderToMem_CP_681_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Sample/req
      -- 
    req_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(30), ack => nbuf_position_582_543_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_update_start_
      -- CP-element group 31: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Update/req
      -- 
    req_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(31), ack => nbuf_position_582_543_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Sample/ack
      -- 
    ack_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_582_543_buf_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nbuf_position_543_Update/ack
      -- 
    ack_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_582_543_buf_ack_1, ack => writeEthernetHeaderToMem_CP_681_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(9) & writeEthernetHeaderToMem_CP_681_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	39 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(9) & writeEthernetHeaderToMem_CP_681_elements(39);
      gj_writeEthernetHeaderToMem_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_sample_start__ps
      -- 
    writeEthernetHeaderToMem_CP_681_elements(36) <= writeEthernetHeaderToMem_CP_681_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_update_start__ps
      -- 
    writeEthernetHeaderToMem_CP_681_elements(38) <= writeEthernetHeaderToMem_CP_681_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	35 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_681_elements(40) <= writeEthernetHeaderToMem_CP_681_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_loopback_sample_req_ps
      -- 
    phi_stmt_544_loopback_sample_req_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_544_loopback_sample_req_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(41), ack => phi_stmt_544_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_681_elements(42) <= writeEthernetHeaderToMem_CP_681_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_entry_sample_req_ps
      -- 
    phi_stmt_544_entry_sample_req_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_544_entry_sample_req_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(43), ack => phi_stmt_544_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_544_phi_mux_ack_ps
      -- 
    phi_stmt_544_phi_mux_ack_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_544_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_sample_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_update_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_681_elements(47) <= writeEthernetHeaderToMem_CP_681_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/type_cast_547_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_681_elements(46), ack => writeEthernetHeaderToMem_CP_681_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Sample/req
      -- 
    req_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(49), ack => nI_577_548_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_update_start_
      -- CP-element group 50: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Update/req
      -- 
    req_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(50), ack => nI_577_548_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Sample/ack
      -- 
    ack_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_577_548_buf_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/R_nI_548_Update/ack
      -- 
    ack_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_577_548_buf_ack_1, ack => writeEthernetHeaderToMem_CP_681_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	60 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	13 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_549_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(9) & writeEthernetHeaderToMem_CP_681_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Sample/rr
      -- 
    rr_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(54), ack => RPIPE_nic_rx_to_header_551_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(11) & writeEthernetHeaderToMem_CP_681_elements(57);
      gj_writeEthernetHeaderToMem_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: 	56 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_update_start_
      -- CP-element group 55: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Update/cr
      -- 
    cr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(55), ack => RPIPE_nic_rx_to_header_551_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(13) & writeEthernetHeaderToMem_CP_681_elements(56);
      gj_writeEthernetHeaderToMem_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56: 	55 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Sample/ra
      -- 
    ra_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_551_inst_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	14 
    -- CP-element group 57: 	58 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	54 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/phi_stmt_549_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/RPIPE_nic_rx_to_header_551_Update/ca
      -- 
    ca_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_551_inst_ack_1, ack => writeEthernetHeaderToMem_CP_681_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Sample/crr
      -- 
    crr_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(58), ack => call_stmt_572_call_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(57) & writeEthernetHeaderToMem_CP_681_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_update_start_
      -- CP-element group 59: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Update/ccr
      -- 
    ccr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_681_elements(59), ack => call_stmt_572_call_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_681_elements(61);
      gj_writeEthernetHeaderToMem_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	53 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Sample/cra
      -- 
    cra_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_572_call_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/call_stmt_572_Update/cca
      -- 
    cca_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_572_call_ack_1, ack => writeEthernetHeaderToMem_CP_681_elements(61)); -- 
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	9 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	10 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writeEthernetHeaderToMem_CP_681_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_681_elements(9), ack => writeEthernetHeaderToMem_CP_681_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	12 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	6 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_535/do_while_stmt_536/do_while_stmt_536_loop_body/$exit
      -- 
    writeEthernetHeaderToMem_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_681_elements(12) & writeEthernetHeaderToMem_CP_681_elements(61);
      gj_writeEthernetHeaderToMem_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	5 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_535/do_while_stmt_536/loop_exit/$exit
      -- CP-element group 64: 	 branch_block_stmt_535/do_while_stmt_536/loop_exit/ack
      -- 
    ack_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_536_branch_ack_0, ack => writeEthernetHeaderToMem_CP_681_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	5 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_535/do_while_stmt_536/loop_taken/$exit
      -- CP-element group 65: 	 branch_block_stmt_535/do_while_stmt_536/loop_taken/ack
      -- 
    ack_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_536_branch_ack_1, ack => writeEthernetHeaderToMem_CP_681_elements(65)); -- 
    -- CP-element group 66:  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	3 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	1 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_535/do_while_stmt_536/$exit
      -- 
    writeEthernetHeaderToMem_CP_681_elements(66) <= writeEthernetHeaderToMem_CP_681_elements(3);
    writeEthernetHeaderToMem_do_while_stmt_536_terminator_850: loop_terminator -- 
      generic map (name => " writeEthernetHeaderToMem_do_while_stmt_536_terminator_850", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeEthernetHeaderToMem_CP_681_elements(6),loop_continue => writeEthernetHeaderToMem_CP_681_elements(65),loop_terminate => writeEthernetHeaderToMem_CP_681_elements(64),loop_back => writeEthernetHeaderToMem_CP_681_elements(4),loop_exit => writeEthernetHeaderToMem_CP_681_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_538_phi_seq_764_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_681_elements(21);
      writeEthernetHeaderToMem_CP_681_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_681_elements(28);
      writeEthernetHeaderToMem_CP_681_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_681_elements(29);
      writeEthernetHeaderToMem_CP_681_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_681_elements(19);
      writeEthernetHeaderToMem_CP_681_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_681_elements(32);
      writeEthernetHeaderToMem_CP_681_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_681_elements(33);
      writeEthernetHeaderToMem_CP_681_elements(20) <= phi_mux_reqs(1);
      phi_stmt_538_phi_seq_764 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_538_phi_seq_764") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_681_elements(11), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_681_elements(17), 
          phi_update_req => writeEthernetHeaderToMem_CP_681_elements(13), 
          phi_update_ack => writeEthernetHeaderToMem_CP_681_elements(18), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_681_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_544_phi_seq_808_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_681_elements(42);
      writeEthernetHeaderToMem_CP_681_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_681_elements(45);
      writeEthernetHeaderToMem_CP_681_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_681_elements(47);
      writeEthernetHeaderToMem_CP_681_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_681_elements(40);
      writeEthernetHeaderToMem_CP_681_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_681_elements(51);
      writeEthernetHeaderToMem_CP_681_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_681_elements(52);
      writeEthernetHeaderToMem_CP_681_elements(41) <= phi_mux_reqs(1);
      phi_stmt_544_phi_seq_808 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_544_phi_seq_808") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_681_elements(36), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_681_elements(37), 
          phi_update_req => writeEthernetHeaderToMem_CP_681_elements(38), 
          phi_update_ack => writeEthernetHeaderToMem_CP_681_elements(39), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_681_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_706_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeEthernetHeaderToMem_CP_681_elements(7);
        preds(1)  <= writeEthernetHeaderToMem_CP_681_elements(8);
        entry_tmerge_706 : transition_merge -- 
          generic map(name => " entry_tmerge_706")
          port map (preds => preds, symbol_out => writeEthernetHeaderToMem_CP_681_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_542_wire : std_logic_vector(35 downto 0);
    signal I_544 : std_logic_vector(3 downto 0);
    signal RPIPE_nic_rx_to_header_551_wire : std_logic_vector(72 downto 0);
    signal ULE_u4_u1_586_wire : std_logic_vector(0 downto 0);
    signal ethernet_header_549 : std_logic_vector(72 downto 0);
    signal ignore_return_572 : std_logic_vector(63 downto 0);
    signal konst_541_wire_constant : std_logic_vector(35 downto 0);
    signal konst_575_wire_constant : std_logic_vector(3 downto 0);
    signal konst_580_wire_constant : std_logic_vector(35 downto 0);
    signal konst_585_wire_constant : std_logic_vector(3 downto 0);
    signal nI_577 : std_logic_vector(3 downto 0);
    signal nI_577_548_buffered : std_logic_vector(3 downto 0);
    signal nbuf_position_582 : std_logic_vector(35 downto 0);
    signal nbuf_position_582_543_buffered : std_logic_vector(35 downto 0);
    signal type_cast_547_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_565_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_559 : std_logic_vector(63 downto 0);
    signal wkeep_563 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_541_wire_constant <= "000000000000000000000000000000001000";
    konst_575_wire_constant <= "0001";
    konst_580_wire_constant <= "000000000000000000000000000000001000";
    konst_585_wire_constant <= "0001";
    type_cast_547_wire_constant <= "0000";
    type_cast_565_wire_constant <= "0";
    type_cast_567_wire_constant <= "0";
    phi_stmt_538: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_542_wire & nbuf_position_582_543_buffered;
      req <= phi_stmt_538_req_0 & phi_stmt_538_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_538",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_538_ack_0,
          idata => idata,
          odata => buf_position_buffer,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_538
    phi_stmt_544: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_547_wire_constant & nI_577_548_buffered;
      req <= phi_stmt_544_req_0 & phi_stmt_544_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_544",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_544_ack_0,
          idata => idata,
          odata => I_544,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_544
    -- flow-through slice operator slice_558_inst
    wdata_559 <= ethernet_header_549(71 downto 8);
    -- flow-through slice operator slice_562_inst
    wkeep_563 <= ethernet_header_549(7 downto 0);
    nI_577_548_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_577_548_buf_req_0;
      nI_577_548_buf_ack_0<= wack(0);
      rreq(0) <= nI_577_548_buf_req_1;
      nI_577_548_buf_ack_1<= rack(0);
      nI_577_548_buf : InterlockBuffer generic map ( -- 
        name => "nI_577_548_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_577_548_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nbuf_position_582_543_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nbuf_position_582_543_buf_req_0;
      nbuf_position_582_543_buf_ack_0<= wack(0);
      rreq(0) <= nbuf_position_582_543_buf_req_1;
      nbuf_position_582_543_buf_ack_1<= rack(0);
      nbuf_position_582_543_buf : InterlockBuffer generic map ( -- 
        name => "nbuf_position_582_543_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nbuf_position_582,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nbuf_position_582_543_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_549
    process(RPIPE_nic_rx_to_header_551_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_header_551_wire(72 downto 0);
      ethernet_header_549 <= tmp_var; -- 
    end process;
    do_while_stmt_536_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULE_u4_u1_586_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_536_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_536_branch_req_0,
          ack0 => do_while_stmt_536_branch_ack_0,
          ack1 => do_while_stmt_536_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_542_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_542_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_542_inst_req_0;
      ADD_u36_u36_542_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_542_inst_req_1;
      ADD_u36_u36_542_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_581_inst
    process(buf_position_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buf_position_buffer, konst_580_wire_constant, tmp_var);
      nbuf_position_582 <= tmp_var; --
    end process;
    -- binary operator ADD_u4_u4_576_inst
    process(I_544) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_544, konst_575_wire_constant, tmp_var);
      nI_577 <= tmp_var; --
    end process;
    -- binary operator ULE_u4_u1_586_inst
    process(nI_577) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(nI_577, konst_585_wire_constant, tmp_var);
      ULE_u4_u1_586_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_header_551_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_header_551_inst_req_0;
      RPIPE_nic_rx_to_header_551_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_header_551_inst_req_1;
      RPIPE_nic_rx_to_header_551_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_header_551_wire <= data_out(72 downto 0);
      nic_rx_to_header_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_header_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_header_pipe_read_req(0),
          oack => nic_rx_to_header_pipe_read_ack(0),
          odata => nic_rx_to_header_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_572_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_572_call_req_0;
      call_stmt_572_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_572_call_req_1;
      call_stmt_572_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_565_wire_constant & type_cast_567_wire_constant & wkeep_563 & buf_position_buffer & wdata_559;
      ignore_return_572 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeEthernetHeaderToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity writePayloadToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buf_pointer : in  std_logic_vector(35 downto 0);
    buf_pointer : in  std_logic_vector(35 downto 0);
    packet_size_32 : out  std_logic_vector(7 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    last_keep : out  std_logic_vector(7 downto 0);
    nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writePayloadToMem;
architecture writePayloadToMem_arch of writePayloadToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 17)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buf_pointer_update_enable: Boolean;
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal packet_size_32_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_32_update_enable: Boolean;
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  signal writePayloadToMem_CP_851_start: Boolean;
  signal writePayloadToMem_CP_851_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_596_branch_ack_1 : boolean;
  signal ADD_u36_u36_602_inst_req_1 : boolean;
  signal phi_stmt_598_req_0 : boolean;
  signal ADD_u36_u36_602_inst_ack_0 : boolean;
  signal do_while_stmt_596_branch_req_0 : boolean;
  signal ADD_u36_u36_602_inst_ack_1 : boolean;
  signal do_while_stmt_596_branch_ack_0 : boolean;
  signal call_stmt_635_call_req_0 : boolean;
  signal ADD_u36_u36_605_inst_ack_1 : boolean;
  signal call_stmt_635_call_ack_0 : boolean;
  signal ADD_u36_u36_605_inst_req_1 : boolean;
  signal ADD_u36_u36_602_inst_req_0 : boolean;
  signal phi_stmt_598_req_1 : boolean;
  signal ADD_u36_u36_605_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_608_inst_ack_1 : boolean;
  signal RPIPE_nic_rx_to_packet_608_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_packet_608_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_608_inst_req_0 : boolean;
  signal ADD_u36_u36_605_inst_req_0 : boolean;
  signal phi_stmt_598_ack_0 : boolean;
  signal call_stmt_635_call_ack_1 : boolean;
  signal call_stmt_635_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writePayloadToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buf_pointer;
  base_buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(71 downto 36) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(71 downto 36);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writePayloadToMem_CP_851_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writePayloadToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 17) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= packet_size_32_buffer;
  packet_size_32 <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(8 downto 8) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(8 downto 8);
  out_buffer_data_in(16 downto 9) <= last_keep_buffer;
  last_keep <= out_buffer_data_out(16 downto 9);
  out_buffer_data_in(tag_length + 16 downto 17) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 16 downto 17);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_851_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writePayloadToMem_CP_851_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_851_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writePayloadToMem_CP_851: Block -- control-path 
    signal writePayloadToMem_CP_851_elements: BooleanArray(49 downto 0);
    -- 
  begin -- 
    writePayloadToMem_CP_851_elements(0) <= writePayloadToMem_CP_851_start;
    writePayloadToMem_CP_851_symbol <= writePayloadToMem_CP_851_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_595/do_while_stmt_596__entry__
      -- CP-element group 0: 	 branch_block_stmt_595/branch_block_stmt_595__entry__
      -- CP-element group 0: 	 branch_block_stmt_595/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	49 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_595/do_while_stmt_596__exit__
      -- CP-element group 1: 	 assign_stmt_648_to_assign_stmt_663/$exit
      -- CP-element group 1: 	 assign_stmt_648_to_assign_stmt_663/$entry
      -- CP-element group 1: 	 branch_block_stmt_595/$exit
      -- CP-element group 1: 	 branch_block_stmt_595/branch_block_stmt_595__exit__
      -- CP-element group 1: 	 $exit
      -- 
    writePayloadToMem_CP_851_elements(1) <= writePayloadToMem_CP_851_elements(49);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_595/do_while_stmt_596/$entry
      -- CP-element group 2: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596__entry__
      -- 
    writePayloadToMem_CP_851_elements(2) <= writePayloadToMem_CP_851_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	49 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596__exit__
      -- 
    -- Element group writePayloadToMem_CP_851_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_595/do_while_stmt_596/loop_back
      -- 
    -- Element group writePayloadToMem_CP_851_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	47 
    -- CP-element group 5: 	48 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_595/do_while_stmt_596/condition_done
      -- CP-element group 5: 	 branch_block_stmt_595/do_while_stmt_596/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_595/do_while_stmt_596/loop_exit/$entry
      -- 
    writePayloadToMem_CP_851_elements(5) <= writePayloadToMem_CP_851_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	46 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_595/do_while_stmt_596/loop_body_done
      -- 
    writePayloadToMem_CP_851_elements(6) <= writePayloadToMem_CP_851_elements(46);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/back_edge_to_loop_body
      -- 
    writePayloadToMem_CP_851_elements(7) <= writePayloadToMem_CP_851_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/first_time_through_loop_body
      -- 
    writePayloadToMem_CP_851_elements(8) <= writePayloadToMem_CP_851_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	45 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_606_sample_start_
      -- 
    -- Element group writePayloadToMem_CP_851_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	45 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/condition_evaluated
      -- 
    condition_evaluated_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(10), ack => do_while_stmt_596_branch_req_0); -- 
    writePayloadToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(14) & writePayloadToMem_CP_851_elements(45);
      gj_writePayloadToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	37 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/aggregated_phi_sample_req
      -- 
    writePayloadToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(9) & writePayloadToMem_CP_851_elements(15) & writePayloadToMem_CP_851_elements(14);
      gj_writePayloadToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	39 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	46 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_606_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_sample_completed_
      -- 
    writePayloadToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(17) & writePayloadToMem_CP_851_elements(39);
      gj_writePayloadToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	36 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_update_start__ps
      -- 
    writePayloadToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(16) & writePayloadToMem_CP_851_elements(36);
      gj_writePayloadToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	40 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/aggregated_phi_update_ack
      -- 
    writePayloadToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(18) & writePayloadToMem_CP_851_elements(40);
      gj_writePayloadToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_sample_start_
      -- 
    writePayloadToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(9) & writePayloadToMem_CP_851_elements(12);
      gj_writePayloadToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	43 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_update_start_
      -- 
    writePayloadToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(9) & writePayloadToMem_CP_851_elements(43);
      gj_writePayloadToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_sample_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_851_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	41 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_update_completed_
      -- 
    -- Element group writePayloadToMem_CP_851_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_loopback_trigger
      -- 
    writePayloadToMem_CP_851_elements(19) <= writePayloadToMem_CP_851_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_loopback_sample_req
      -- 
    phi_stmt_598_loopback_sample_req_890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_598_loopback_sample_req_890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(20), ack => phi_stmt_598_req_1); -- 
    -- Element group writePayloadToMem_CP_851_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_entry_trigger
      -- 
    writePayloadToMem_CP_851_elements(21) <= writePayloadToMem_CP_851_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_entry_sample_req_ps
      -- 
    phi_stmt_598_entry_sample_req_893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_598_entry_sample_req_893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(22), ack => phi_stmt_598_req_0); -- 
    -- Element group writePayloadToMem_CP_851_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_598_phi_mux_ack
      -- 
    phi_stmt_598_phi_mux_ack_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_598_ack_0, ack => writePayloadToMem_CP_851_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_851_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_851_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_sample_start_
      -- 
    rr_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(26), ack => ADD_u36_u36_602_inst_req_0); -- 
    writePayloadToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(24) & writePayloadToMem_CP_851_elements(28);
      gj_writePayloadToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_update_start_
      -- CP-element group 27: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Update/cr
      -- 
    cr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(27), ack => ADD_u36_u36_602_inst_req_1); -- 
    writePayloadToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(25) & writePayloadToMem_CP_851_elements(29);
      gj_writePayloadToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_sample_completed__ps
      -- 
    ra_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_602_inst_ack_0, ack => writePayloadToMem_CP_851_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_602_update_completed__ps
      -- 
    ca_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_602_inst_ack_1, ack => writePayloadToMem_CP_851_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_851_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_851_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Sample/rr
      -- 
    rr_927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(32), ack => ADD_u36_u36_605_inst_req_0); -- 
    writePayloadToMem_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(30) & writePayloadToMem_CP_851_elements(34);
      gj_writePayloadToMem_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_update_start_
      -- CP-element group 33: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Update/$entry
      -- 
    cr_932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(33), ack => ADD_u36_u36_605_inst_req_1); -- 
    writePayloadToMem_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(31) & writePayloadToMem_CP_851_elements(35);
      gj_writePayloadToMem_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Sample/$exit
      -- 
    ra_928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_605_inst_ack_0, ack => writePayloadToMem_CP_851_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/ADD_u36_u36_605_Update/ca
      -- 
    ca_933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_605_inst_ack_1, ack => writePayloadToMem_CP_851_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	43 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	13 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_606_update_start_
      -- 
    writePayloadToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(9) & writePayloadToMem_CP_851_elements(43);
      gj_writePayloadToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	40 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Sample/rr
      -- CP-element group 37: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_sample_start_
      -- 
    rr_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(37), ack => RPIPE_nic_rx_to_packet_608_inst_req_0); -- 
    writePayloadToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(11) & writePayloadToMem_CP_851_elements(40);
      gj_writePayloadToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: 	39 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Update/cr
      -- CP-element group 38: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_update_start_
      -- 
    cr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(38), ack => RPIPE_nic_rx_to_packet_608_inst_req_1); -- 
    writePayloadToMem_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(13) & writePayloadToMem_CP_851_elements(39);
      gj_writePayloadToMem_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	12 
    -- CP-element group 39: 	38 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_sample_completed_
      -- 
    ra_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_608_inst_ack_0, ack => writePayloadToMem_CP_851_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	14 
    -- CP-element group 40: 	41 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	37 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/RPIPE_nic_rx_to_packet_608_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/phi_stmt_606_update_completed_
      -- 
    ca_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_608_inst_ack_1, ack => writePayloadToMem_CP_851_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: 	40 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Sample/crr
      -- 
    crr_960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(41), ack => call_stmt_635_call_req_0); -- 
    writePayloadToMem_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(18) & writePayloadToMem_CP_851_elements(40) & writePayloadToMem_CP_851_elements(43);
      gj_writePayloadToMem_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_update_start_
      -- CP-element group 42: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Update/ccr
      -- 
    ccr_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_851_elements(42), ack => call_stmt_635_call_req_1); -- 
    writePayloadToMem_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writePayloadToMem_CP_851_elements(44);
      gj_writePayloadToMem_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	16 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Sample/cra
      -- 
    cra_961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_635_call_ack_0, ack => writePayloadToMem_CP_851_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/call_stmt_635_Update/cca
      -- 
    cca_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_635_call_ack_1, ack => writePayloadToMem_CP_851_elements(44)); -- 
    -- CP-element group 45:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	9 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	10 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writePayloadToMem_CP_851_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_851_elements(9), ack => writePayloadToMem_CP_851_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	12 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	6 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_595/do_while_stmt_596/do_while_stmt_596_loop_body/$exit
      -- 
    writePayloadToMem_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_851_elements(12) & writePayloadToMem_CP_851_elements(44);
      gj_writePayloadToMem_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_851_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	5 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_595/do_while_stmt_596/loop_exit/$exit
      -- CP-element group 47: 	 branch_block_stmt_595/do_while_stmt_596/loop_exit/ack
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_596_branch_ack_0, ack => writePayloadToMem_CP_851_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	5 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_595/do_while_stmt_596/loop_taken/ack
      -- CP-element group 48: 	 branch_block_stmt_595/do_while_stmt_596/loop_taken/$exit
      -- 
    ack_975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_596_branch_ack_1, ack => writePayloadToMem_CP_851_elements(48)); -- 
    -- CP-element group 49:  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	3 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	1 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_595/do_while_stmt_596/$exit
      -- 
    writePayloadToMem_CP_851_elements(49) <= writePayloadToMem_CP_851_elements(3);
    writePayloadToMem_do_while_stmt_596_terminator_976: loop_terminator -- 
      generic map (name => " writePayloadToMem_do_while_stmt_596_terminator_976", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writePayloadToMem_CP_851_elements(6),loop_continue => writePayloadToMem_CP_851_elements(48),loop_terminate => writePayloadToMem_CP_851_elements(47),loop_back => writePayloadToMem_CP_851_elements(4),loop_exit => writePayloadToMem_CP_851_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_598_phi_seq_934_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writePayloadToMem_CP_851_elements(21);
      writePayloadToMem_CP_851_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writePayloadToMem_CP_851_elements(28);
      writePayloadToMem_CP_851_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writePayloadToMem_CP_851_elements(29);
      writePayloadToMem_CP_851_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writePayloadToMem_CP_851_elements(19);
      writePayloadToMem_CP_851_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writePayloadToMem_CP_851_elements(34);
      writePayloadToMem_CP_851_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writePayloadToMem_CP_851_elements(35);
      writePayloadToMem_CP_851_elements(20) <= phi_mux_reqs(1);
      phi_stmt_598_phi_seq_934 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_598_phi_seq_934") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writePayloadToMem_CP_851_elements(11), 
          phi_sample_ack => writePayloadToMem_CP_851_elements(17), 
          phi_update_req => writePayloadToMem_CP_851_elements(13), 
          phi_update_ack => writePayloadToMem_CP_851_elements(18), 
          phi_mux_ack => writePayloadToMem_CP_851_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_876_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writePayloadToMem_CP_851_elements(7);
        preds(1)  <= writePayloadToMem_CP_851_elements(8);
        entry_tmerge_876 : transition_merge -- 
          generic map(name => " entry_tmerge_876")
          port map (preds => preds, symbol_out => writePayloadToMem_CP_851_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_602_wire : std_logic_vector(35 downto 0);
    signal ADD_u36_u36_605_wire : std_logic_vector(35 downto 0);
    signal EQ_u64_u1_643_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_646_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_638_wire : std_logic_vector(0 downto 0);
    signal RPIPE_nic_rx_to_packet_608_wire : std_logic_vector(72 downto 0);
    signal R_BAD_PACKET_DATA_642_wire_constant : std_logic_vector(63 downto 0);
    signal SUB_u36_u36_652_wire : std_logic_vector(35 downto 0);
    signal buf_position_598 : std_logic_vector(35 downto 0);
    signal ignore_return_635 : std_logic_vector(63 downto 0);
    signal konst_601_wire_constant : std_logic_vector(35 downto 0);
    signal konst_604_wire_constant : std_logic_vector(35 downto 0);
    signal konst_645_wire_constant : std_logic_vector(7 downto 0);
    signal last_bit_613 : std_logic_vector(0 downto 0);
    signal packet_size_8_654 : std_logic_vector(7 downto 0);
    signal payload_data_606 : std_logic_vector(72 downto 0);
    signal type_cast_628_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_630_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_617 : std_logic_vector(63 downto 0);
    signal wkeep_621 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_BAD_PACKET_DATA_642_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    konst_601_wire_constant <= "000000000000000000000000000000001000";
    konst_604_wire_constant <= "000000000000000000000000000000001000";
    konst_645_wire_constant <= "00000000";
    type_cast_628_wire_constant <= "0";
    type_cast_630_wire_constant <= "0";
    phi_stmt_598: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_602_wire & ADD_u36_u36_605_wire;
      req <= phi_stmt_598_req_0 & phi_stmt_598_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_598",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_598_ack_0,
          idata => idata,
          odata => buf_position_598,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_598
    -- flow-through slice operator slice_612_inst
    last_bit_613 <= payload_data_606(72 downto 72);
    -- flow-through slice operator slice_616_inst
    wdata_617 <= payload_data_606(71 downto 8);
    -- flow-through slice operator slice_620_inst
    wkeep_621 <= payload_data_606(7 downto 0);
    -- interlock W_last_keep_661_inst
    process(wkeep_621) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := wkeep_621(7 downto 0);
      last_keep_buffer <= tmp_var; -- 
    end process;
    -- interlock W_packet_size_32_655_inst
    process(packet_size_8_654) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := packet_size_8_654(7 downto 0);
      packet_size_32_buffer <= tmp_var; -- 
    end process;
    -- interlock ssrc_phi_stmt_606
    process(RPIPE_nic_rx_to_packet_608_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_packet_608_wire(72 downto 0);
      payload_data_606 <= tmp_var; -- 
    end process;
    -- interlock type_cast_653_inst
    process(SUB_u36_u36_652_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := SUB_u36_u36_652_wire(7 downto 0);
      packet_size_8_654 <= tmp_var; -- 
    end process;
    do_while_stmt_596_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_638_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_596_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_596_branch_req_0,
          ack0 => do_while_stmt_596_branch_ack_0,
          ack1 => do_while_stmt_596_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_602_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_602_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_602_inst_req_0;
      ADD_u36_u36_602_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_602_inst_req_1;
      ADD_u36_u36_602_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : ADD_u36_u36_605_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_position_598;
      ADD_u36_u36_605_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_605_inst_req_0;
      ADD_u36_u36_605_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_605_inst_req_1;
      ADD_u36_u36_605_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- binary operator AND_u1_u1_647_inst
    process(EQ_u64_u1_643_wire, EQ_u8_u1_646_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u64_u1_643_wire, EQ_u8_u1_646_wire, tmp_var);
      bad_packet_identifier_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_643_inst
    process(wdata_617) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wdata_617, R_BAD_PACKET_DATA_642_wire_constant, tmp_var);
      EQ_u64_u1_643_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_646_inst
    process(wkeep_621) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wkeep_621, konst_645_wire_constant, tmp_var);
      EQ_u8_u1_646_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_638_inst
    process(last_bit_613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_613, tmp_var);
      NOT_u1_u1_638_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u36_u36_652_inst
    process(buf_position_598, base_buf_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(buf_position_598, base_buf_pointer_buffer, tmp_var);
      SUB_u36_u36_652_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_packet_608_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_packet_608_inst_req_0;
      RPIPE_nic_rx_to_packet_608_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_packet_608_inst_req_1;
      RPIPE_nic_rx_to_packet_608_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_packet_608_wire <= data_out(72 downto 0);
      nic_rx_to_packet_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_packet_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_packet_pipe_read_req(0),
          oack => nic_rx_to_packet_pipe_read_ack(0),
          odata => nic_rx_to_packet_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_635_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 3);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_635_call_req_0;
      call_stmt_635_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_635_call_req_1;
      call_stmt_635_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_628_wire_constant & type_cast_630_wire_constant & wkeep_621 & buf_position_598 & wdata_617;
      ignore_return_635 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writePayloadToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library ahir_system_global_packagelib;
use ahir_system_global_packagelib.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    AFB_NIC_REQUEST_pipe_write_data: in std_logic_vector(73 downto 0);
    AFB_NIC_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
    AFB_NIC_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_data: in std_logic_vector(72 downto 0);
    mac_to_nic_data_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_data: out std_logic_vector(72 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(11 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(5 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module AccessRegister
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module AccessRegister
  signal AccessRegister_rwbar :  std_logic_vector(0 downto 0);
  signal AccessRegister_bmask :  std_logic_vector(3 downto 0);
  signal AccessRegister_register_index :  std_logic_vector(5 downto 0);
  signal AccessRegister_wdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_rdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_in_args    : std_logic_vector(42 downto 0);
  signal AccessRegister_out_args   : std_logic_vector(31 downto 0);
  signal AccessRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal AccessRegister_tag_out   : std_logic_vector(2 downto 0);
  signal AccessRegister_start_req : std_logic;
  signal AccessRegister_start_ack : std_logic;
  signal AccessRegister_fin_req   : std_logic;
  signal AccessRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module AccessRegister
  signal AccessRegister_call_reqs: std_logic_vector(1 downto 0);
  signal AccessRegister_call_acks: std_logic_vector(1 downto 0);
  signal AccessRegister_return_reqs: std_logic_vector(1 downto 0);
  signal AccessRegister_return_acks: std_logic_vector(1 downto 0);
  signal AccessRegister_call_data: std_logic_vector(85 downto 0);
  signal AccessRegister_call_tag: std_logic_vector(1 downto 0);
  signal AccessRegister_return_data: std_logic_vector(63 downto 0);
  signal AccessRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module NicRegisterAccessDaemon
  component NicRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module NicRegisterAccessDaemon
  signal NicRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal NicRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal NicRegisterAccessDaemon_start_req : std_logic;
  signal NicRegisterAccessDaemon_start_ack : std_logic;
  signal NicRegisterAccessDaemon_fin_req   : std_logic;
  signal NicRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module ReceiveEngineDaemon
  component ReceiveEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      FREE_Q : in std_logic_vector(35 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_call_data : out  std_logic_vector(35 downto 0);
      loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
      loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_return_data : in   std_logic_vector(0 downto 0);
      loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
      populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
      populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ReceiveEngineDaemon
  signal ReceiveEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ReceiveEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal ReceiveEngineDaemon_start_req : std_logic;
  signal ReceiveEngineDaemon_start_ack : std_logic;
  signal ReceiveEngineDaemon_fin_req   : std_logic;
  signal ReceiveEngineDaemon_fin_ack : std_logic;
  -- declarations related to module SoftwareRegisterAccessDaemon
  component SoftwareRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
      FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
      AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
      CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module SoftwareRegisterAccessDaemon
  signal SoftwareRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal SoftwareRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal SoftwareRegisterAccessDaemon_start_req : std_logic;
  signal SoftwareRegisterAccessDaemon_start_ack : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_req   : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module UpdateRegister
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module UpdateRegister
  signal UpdateRegister_bmask :  std_logic_vector(3 downto 0);
  signal UpdateRegister_rval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_wdata :  std_logic_vector(31 downto 0);
  signal UpdateRegister_index :  std_logic_vector(5 downto 0);
  signal UpdateRegister_wval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_in_args    : std_logic_vector(73 downto 0);
  signal UpdateRegister_out_args   : std_logic_vector(31 downto 0);
  signal UpdateRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal UpdateRegister_tag_out   : std_logic_vector(2 downto 0);
  signal UpdateRegister_start_req : std_logic;
  signal UpdateRegister_start_ack : std_logic;
  signal UpdateRegister_fin_req   : std_logic;
  signal UpdateRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module UpdateRegister
  signal UpdateRegister_call_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_data: std_logic_vector(147 downto 0);
  signal UpdateRegister_call_tag: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_data: std_logic_vector(63 downto 0);
  signal UpdateRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMemory
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemory
  signal accessMemory_lock :  std_logic_vector(0 downto 0);
  signal accessMemory_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemory_bmask :  std_logic_vector(7 downto 0);
  signal accessMemory_addr :  std_logic_vector(35 downto 0);
  signal accessMemory_wdata :  std_logic_vector(63 downto 0);
  signal accessMemory_rdata :  std_logic_vector(63 downto 0);
  signal accessMemory_in_args    : std_logic_vector(109 downto 0);
  signal accessMemory_out_args   : std_logic_vector(63 downto 0);
  signal accessMemory_tag_in    : std_logic_vector(5 downto 0) := (others => '0');
  signal accessMemory_tag_out   : std_logic_vector(5 downto 0);
  signal accessMemory_start_req : std_logic;
  signal accessMemory_start_ack : std_logic;
  signal accessMemory_fin_req   : std_logic;
  signal accessMemory_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemory
  signal accessMemory_call_reqs: std_logic_vector(10 downto 0);
  signal accessMemory_call_acks: std_logic_vector(10 downto 0);
  signal accessMemory_return_reqs: std_logic_vector(10 downto 0);
  signal accessMemory_return_acks: std_logic_vector(10 downto 0);
  signal accessMemory_call_data: std_logic_vector(1209 downto 0);
  signal accessMemory_call_tag: std_logic_vector(21 downto 0);
  signal accessMemory_return_data: std_logic_vector(703 downto 0);
  signal accessMemory_return_tag: std_logic_vector(21 downto 0);
  -- declarations related to module acquireMutex
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module acquireMutex
  signal acquireMutex_q_base_address :  std_logic_vector(35 downto 0);
  signal acquireMutex_m_ok :  std_logic_vector(0 downto 0);
  signal acquireMutex_in_args    : std_logic_vector(35 downto 0);
  signal acquireMutex_out_args   : std_logic_vector(0 downto 0);
  signal acquireMutex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal acquireMutex_tag_out   : std_logic_vector(2 downto 0);
  signal acquireMutex_start_req : std_logic;
  signal acquireMutex_start_ack : std_logic;
  signal acquireMutex_fin_req   : std_logic;
  signal acquireMutex_fin_ack : std_logic;
  -- caller side aggregated signals for module acquireMutex
  signal acquireMutex_call_reqs: std_logic_vector(1 downto 0);
  signal acquireMutex_call_acks: std_logic_vector(1 downto 0);
  signal acquireMutex_return_reqs: std_logic_vector(1 downto 0);
  signal acquireMutex_return_acks: std_logic_vector(1 downto 0);
  signal acquireMutex_call_data: std_logic_vector(71 downto 0);
  signal acquireMutex_call_tag: std_logic_vector(1 downto 0);
  signal acquireMutex_return_data: std_logic_vector(1 downto 0);
  signal acquireMutex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module delay_time
  -- declarations related to module getQueueElement
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_pointer : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueElement
  signal getQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueElement_read_pointer :  std_logic_vector(31 downto 0);
  signal getQueueElement_q_r_data :  std_logic_vector(31 downto 0);
  signal getQueueElement_in_args    : std_logic_vector(67 downto 0);
  signal getQueueElement_out_args   : std_logic_vector(31 downto 0);
  signal getQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal getQueueElement_start_req : std_logic;
  signal getQueueElement_start_ack : std_logic;
  signal getQueueElement_fin_req   : std_logic;
  signal getQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueElement
  signal getQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_call_data: std_logic_vector(67 downto 0);
  signal getQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal getQueueElement_return_data: std_logic_vector(31 downto 0);
  signal getQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module getQueuePointers
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointers
  signal getQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_in_args    : std_logic_vector(35 downto 0);
  signal getQueuePointers_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointers_start_req : std_logic;
  signal getQueuePointers_start_ack : std_logic;
  signal getQueuePointers_fin_req   : std_logic;
  signal getQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointers
  signal getQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_data: std_logic_vector(71 downto 0);
  signal getQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTxPacketPointerFromServer
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_queue_index :  std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_pkt_pointer :  std_logic_vector(31 downto 0);
  signal getTxPacketPointerFromServer_status :  std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_in_args    : std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_out_args   : std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getTxPacketPointerFromServer_tag_out   : std_logic_vector(1 downto 0);
  signal getTxPacketPointerFromServer_start_req : std_logic;
  signal getTxPacketPointerFromServer_start_ack : std_logic;
  signal getTxPacketPointerFromServer_fin_req   : std_logic;
  signal getTxPacketPointerFromServer_fin_ack : std_logic;
  -- caller side aggregated signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_call_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_data: std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_call_tag: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_data: std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module loadBuffer
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadBuffer
  signal loadBuffer_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal loadBuffer_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal loadBuffer_in_args    : std_logic_vector(35 downto 0);
  signal loadBuffer_out_args   : std_logic_vector(0 downto 0);
  signal loadBuffer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadBuffer_tag_out   : std_logic_vector(1 downto 0);
  signal loadBuffer_start_req : std_logic;
  signal loadBuffer_start_ack : std_logic;
  signal loadBuffer_fin_req   : std_logic;
  signal loadBuffer_fin_ack : std_logic;
  -- caller side aggregated signals for module loadBuffer
  signal loadBuffer_call_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_call_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_return_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_return_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_call_data: std_logic_vector(35 downto 0);
  signal loadBuffer_call_tag: std_logic_vector(0 downto 0);
  signal loadBuffer_return_data: std_logic_vector(0 downto 0);
  signal loadBuffer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module nextLSTATE
  -- declarations related to module nicRxFromMacDaemon
  component nicRxFromMacDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
      nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicRxFromMacDaemon
  signal nicRxFromMacDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicRxFromMacDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal nicRxFromMacDaemon_start_req : std_logic;
  signal nicRxFromMacDaemon_start_ack : std_logic;
  signal nicRxFromMacDaemon_fin_req   : std_logic;
  signal nicRxFromMacDaemon_fin_ack : std_logic;
  -- declarations related to module popFromQueue
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module popFromQueue
  signal popFromQueue_lock :  std_logic_vector(0 downto 0);
  signal popFromQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal popFromQueue_q_r_data :  std_logic_vector(31 downto 0);
  signal popFromQueue_status :  std_logic_vector(0 downto 0);
  signal popFromQueue_in_args    : std_logic_vector(36 downto 0);
  signal popFromQueue_out_args   : std_logic_vector(32 downto 0);
  signal popFromQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal popFromQueue_tag_out   : std_logic_vector(2 downto 0);
  signal popFromQueue_start_req : std_logic;
  signal popFromQueue_start_ack : std_logic;
  signal popFromQueue_fin_req   : std_logic;
  signal popFromQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module popFromQueue
  signal popFromQueue_call_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_call_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_return_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_return_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_call_data: std_logic_vector(73 downto 0);
  signal popFromQueue_call_tag: std_logic_vector(1 downto 0);
  signal popFromQueue_return_data: std_logic_vector(65 downto 0);
  signal popFromQueue_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module populateRxQueue
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module populateRxQueue
  signal populateRxQueue_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal populateRxQueue_in_args    : std_logic_vector(35 downto 0);
  signal populateRxQueue_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal populateRxQueue_tag_out   : std_logic_vector(1 downto 0);
  signal populateRxQueue_start_req : std_logic;
  signal populateRxQueue_start_ack : std_logic;
  signal populateRxQueue_fin_req   : std_logic;
  signal populateRxQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module populateRxQueue
  signal populateRxQueue_call_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_data: std_logic_vector(35 downto 0);
  signal populateRxQueue_call_tag: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module pushIntoQueue
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module pushIntoQueue
  signal pushIntoQueue_lock :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal pushIntoQueue_q_w_data :  std_logic_vector(31 downto 0);
  signal pushIntoQueue_status :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_in_args    : std_logic_vector(68 downto 0);
  signal pushIntoQueue_out_args   : std_logic_vector(0 downto 0);
  signal pushIntoQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal pushIntoQueue_tag_out   : std_logic_vector(2 downto 0);
  signal pushIntoQueue_start_req : std_logic;
  signal pushIntoQueue_start_ack : std_logic;
  signal pushIntoQueue_fin_req   : std_logic;
  signal pushIntoQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module pushIntoQueue
  signal pushIntoQueue_call_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_data: std_logic_vector(206 downto 0);
  signal pushIntoQueue_call_tag: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_data: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module releaseMutex
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module releaseMutex
  signal releaseMutex_q_base_address :  std_logic_vector(35 downto 0);
  signal releaseMutex_in_args    : std_logic_vector(35 downto 0);
  signal releaseMutex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal releaseMutex_tag_out   : std_logic_vector(2 downto 0);
  signal releaseMutex_start_req : std_logic;
  signal releaseMutex_start_ack : std_logic;
  signal releaseMutex_fin_req   : std_logic;
  signal releaseMutex_fin_ack : std_logic;
  -- caller side aggregated signals for module releaseMutex
  signal releaseMutex_call_reqs: std_logic_vector(1 downto 0);
  signal releaseMutex_call_acks: std_logic_vector(1 downto 0);
  signal releaseMutex_return_reqs: std_logic_vector(1 downto 0);
  signal releaseMutex_return_acks: std_logic_vector(1 downto 0);
  signal releaseMutex_call_data: std_logic_vector(71 downto 0);
  signal releaseMutex_call_tag: std_logic_vector(1 downto 0);
  signal releaseMutex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setQueueElement
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_pointer : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueueElement
  signal setQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueueElement_write_pointer :  std_logic_vector(31 downto 0);
  signal setQueueElement_q_w_data :  std_logic_vector(31 downto 0);
  signal setQueueElement_in_args    : std_logic_vector(99 downto 0);
  signal setQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal setQueueElement_start_req : std_logic;
  signal setQueueElement_start_ack : std_logic;
  signal setQueueElement_fin_req   : std_logic;
  signal setQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueueElement
  signal setQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_call_data: std_logic_vector(99 downto 0);
  signal setQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal setQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueuePointers
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueuePointers
  signal setQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_in_args    : std_logic_vector(99 downto 0);
  signal setQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal setQueuePointers_start_req : std_logic;
  signal setQueuePointers_start_ack : std_logic;
  signal setQueuePointers_fin_req   : std_logic;
  signal setQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueuePointers
  signal setQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_data: std_logic_vector(199 downto 0);
  signal setQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module transmitEngineDaemon
  component transmitEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
      getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
      getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
      transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_call_data : out  std_logic_vector(31 downto 0);
      transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
      transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_return_data : in   std_logic_vector(0 downto 0);
      transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitEngineDaemon
  signal transmitEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal transmitEngineDaemon_start_req : std_logic;
  signal transmitEngineDaemon_start_ack : std_logic;
  signal transmitEngineDaemon_fin_req   : std_logic;
  signal transmitEngineDaemon_fin_ack : std_logic;
  -- declarations related to module transmitPacket
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitPacket
  signal transmitPacket_packet_pointer :  std_logic_vector(31 downto 0);
  signal transmitPacket_status :  std_logic_vector(0 downto 0);
  signal transmitPacket_in_args    : std_logic_vector(31 downto 0);
  signal transmitPacket_out_args   : std_logic_vector(0 downto 0);
  signal transmitPacket_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitPacket_tag_out   : std_logic_vector(1 downto 0);
  signal transmitPacket_start_req : std_logic;
  signal transmitPacket_start_ack : std_logic;
  signal transmitPacket_fin_req   : std_logic;
  signal transmitPacket_fin_ack : std_logic;
  -- caller side aggregated signals for module transmitPacket
  signal transmitPacket_call_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_call_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_return_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_return_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_call_data: std_logic_vector(31 downto 0);
  signal transmitPacket_call_tag: std_logic_vector(0 downto 0);
  signal transmitPacket_return_data: std_logic_vector(0 downto 0);
  signal transmitPacket_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeControlInformationToMem
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeControlInformationToMem
  signal writeControlInformationToMem_base_buffer_pointer :  std_logic_vector(35 downto 0);
  signal writeControlInformationToMem_packet_size :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_in_args    : std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeControlInformationToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeControlInformationToMem_start_req : std_logic;
  signal writeControlInformationToMem_start_ack : std_logic;
  signal writeControlInformationToMem_fin_req   : std_logic;
  signal writeControlInformationToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeControlInformationToMem
  signal writeControlInformationToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_data: std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeEthernetHeaderToMem
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_buf_position :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_in_args    : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_out_args   : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeEthernetHeaderToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeEthernetHeaderToMem_start_req : std_logic;
  signal writeEthernetHeaderToMem_start_ack : std_logic;
  signal writeEthernetHeaderToMem_fin_req   : std_logic;
  signal writeEthernetHeaderToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writePayloadToMem
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writePayloadToMem
  signal writePayloadToMem_base_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_packet_size_32 :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal writePayloadToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_in_args    : std_logic_vector(71 downto 0);
  signal writePayloadToMem_out_args   : std_logic_vector(16 downto 0);
  signal writePayloadToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writePayloadToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writePayloadToMem_start_req : std_logic;
  signal writePayloadToMem_start_ack : std_logic;
  signal writePayloadToMem_fin_req   : std_logic;
  signal writePayloadToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writePayloadToMem
  signal writePayloadToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_data: std_logic_vector(71 downto 0);
  signal writePayloadToMem_call_tag: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_data: std_logic_vector(16 downto 0);
  signal writePayloadToMem_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_read_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_write_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe CONTROL_REGISTER
  signal CONTROL_REGISTER_pipe_write_data: std_logic_vector(31 downto 0);
  signal CONTROL_REGISTER_pipe_write_req: std_logic_vector(0 downto 0);
  signal CONTROL_REGISTER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe CONTROL_REGISTER
  signal CONTROL_REGISTER: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe FREE_Q
  signal FREE_Q_pipe_write_data: std_logic_vector(35 downto 0);
  signal FREE_Q_pipe_write_req: std_logic_vector(0 downto 0);
  signal FREE_Q_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe FREE_Q
  signal FREE_Q: std_logic_vector(35 downto 0);
  -- aggregate signals for write to pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for read from pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS_pipe_write_data: std_logic_vector(31 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_req: std_logic_vector(0 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS: std_logic_vector(31 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_read_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_write_data: std_logic_vector(145 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module AccessRegister
  AccessRegister_rwbar <= AccessRegister_in_args(42 downto 42);
  AccessRegister_bmask <= AccessRegister_in_args(41 downto 38);
  AccessRegister_register_index <= AccessRegister_in_args(37 downto 32);
  AccessRegister_wdata <= AccessRegister_in_args(31 downto 0);
  AccessRegister_out_args <= AccessRegister_rdata ;
  -- call arbiter for module AccessRegister
  AccessRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 43,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => AccessRegister_call_reqs,
      call_acks => AccessRegister_call_acks,
      return_reqs => AccessRegister_return_reqs,
      return_acks => AccessRegister_return_acks,
      call_data  => AccessRegister_call_data,
      call_tag  => AccessRegister_call_tag,
      return_tag  => AccessRegister_return_tag,
      call_mtag => AccessRegister_tag_in,
      return_mtag => AccessRegister_tag_out,
      return_data =>AccessRegister_return_data,
      call_mreq => AccessRegister_start_req,
      call_mack => AccessRegister_start_ack,
      return_mreq => AccessRegister_fin_req,
      return_mack => AccessRegister_fin_ack,
      call_mdata => AccessRegister_in_args,
      return_mdata => AccessRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  AccessRegister_instance:AccessRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      rwbar => AccessRegister_rwbar,
      bmask => AccessRegister_bmask,
      register_index => AccessRegister_register_index,
      wdata => AccessRegister_wdata,
      rdata => AccessRegister_rdata,
      start_req => AccessRegister_start_req,
      start_ack => AccessRegister_start_ack,
      fin_req => AccessRegister_fin_req,
      fin_ack => AccessRegister_fin_ack,
      clk => clk,
      reset => reset,
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
      tag_in => AccessRegister_tag_in,
      tag_out => AccessRegister_tag_out-- 
    ); -- 
  -- module NicRegisterAccessDaemon
  NicRegisterAccessDaemon_instance:NicRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => NicRegisterAccessDaemon_start_req,
      start_ack => NicRegisterAccessDaemon_start_ack,
      fin_req => NicRegisterAccessDaemon_fin_req,
      fin_ack => NicRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(11 downto 6),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(1 downto 1),
      UpdateRegister_call_acks => UpdateRegister_call_acks(1 downto 1),
      UpdateRegister_call_data => UpdateRegister_call_data(147 downto 74),
      UpdateRegister_call_tag => UpdateRegister_call_tag(1 downto 1),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(1 downto 1),
      UpdateRegister_return_acks => UpdateRegister_return_acks(1 downto 1),
      UpdateRegister_return_data => UpdateRegister_return_data(63 downto 32),
      UpdateRegister_return_tag => UpdateRegister_return_tag(1 downto 1),
      tag_in => NicRegisterAccessDaemon_tag_in,
      tag_out => NicRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  NicRegisterAccessDaemon_tag_in <= (others => '0');
  NicRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => NicRegisterAccessDaemon_start_req, start_ack => NicRegisterAccessDaemon_start_ack,  fin_req => NicRegisterAccessDaemon_fin_req,  fin_ack => NicRegisterAccessDaemon_fin_ack);
  -- module ReceiveEngineDaemon
  ReceiveEngineDaemon_instance:ReceiveEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ReceiveEngineDaemon_start_req,
      start_ack => ReceiveEngineDaemon_start_ack,
      fin_req => ReceiveEngineDaemon_fin_req,
      fin_ack => ReceiveEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      FREE_Q => FREE_Q,
      CONTROL_REGISTER => CONTROL_REGISTER,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
      popFromQueue_call_reqs => popFromQueue_call_reqs(1 downto 1),
      popFromQueue_call_acks => popFromQueue_call_acks(1 downto 1),
      popFromQueue_call_data => popFromQueue_call_data(73 downto 37),
      popFromQueue_call_tag => popFromQueue_call_tag(1 downto 1),
      popFromQueue_return_reqs => popFromQueue_return_reqs(1 downto 1),
      popFromQueue_return_acks => popFromQueue_return_acks(1 downto 1),
      popFromQueue_return_data => popFromQueue_return_data(65 downto 33),
      popFromQueue_return_tag => popFromQueue_return_tag(1 downto 1),
      loadBuffer_call_reqs => loadBuffer_call_reqs(0 downto 0),
      loadBuffer_call_acks => loadBuffer_call_acks(0 downto 0),
      loadBuffer_call_data => loadBuffer_call_data(35 downto 0),
      loadBuffer_call_tag => loadBuffer_call_tag(0 downto 0),
      loadBuffer_return_reqs => loadBuffer_return_reqs(0 downto 0),
      loadBuffer_return_acks => loadBuffer_return_acks(0 downto 0),
      loadBuffer_return_data => loadBuffer_return_data(0 downto 0),
      loadBuffer_return_tag => loadBuffer_return_tag(0 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(1 downto 1),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(1 downto 1),
      pushIntoQueue_call_data => pushIntoQueue_call_data(137 downto 69),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(1 downto 1),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(1 downto 1),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(1 downto 1),
      pushIntoQueue_return_data => pushIntoQueue_return_data(1 downto 1),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(1 downto 1),
      populateRxQueue_call_reqs => populateRxQueue_call_reqs(0 downto 0),
      populateRxQueue_call_acks => populateRxQueue_call_acks(0 downto 0),
      populateRxQueue_call_data => populateRxQueue_call_data(35 downto 0),
      populateRxQueue_call_tag => populateRxQueue_call_tag(0 downto 0),
      populateRxQueue_return_reqs => populateRxQueue_return_reqs(0 downto 0),
      populateRxQueue_return_acks => populateRxQueue_return_acks(0 downto 0),
      populateRxQueue_return_tag => populateRxQueue_return_tag(0 downto 0),
      tag_in => ReceiveEngineDaemon_tag_in,
      tag_out => ReceiveEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  ReceiveEngineDaemon_tag_in <= (others => '0');
  ReceiveEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ReceiveEngineDaemon_start_req, start_ack => ReceiveEngineDaemon_start_ack,  fin_req => ReceiveEngineDaemon_fin_req,  fin_ack => ReceiveEngineDaemon_fin_ack);
  -- module SoftwareRegisterAccessDaemon
  SoftwareRegisterAccessDaemon_instance:SoftwareRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => SoftwareRegisterAccessDaemon_start_req,
      start_ack => SoftwareRegisterAccessDaemon_start_ack,
      fin_req => SoftwareRegisterAccessDaemon_fin_req,
      fin_ack => SoftwareRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(5 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      AFB_NIC_REQUEST_pipe_read_req => AFB_NIC_REQUEST_pipe_read_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_ack => AFB_NIC_REQUEST_pipe_read_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_data => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
      FREE_Q_pipe_write_req => FREE_Q_pipe_write_req(0 downto 0),
      FREE_Q_pipe_write_ack => FREE_Q_pipe_write_ack(0 downto 0),
      FREE_Q_pipe_write_data => FREE_Q_pipe_write_data(35 downto 0),
      AFB_NIC_RESPONSE_pipe_write_req => AFB_NIC_RESPONSE_pipe_write_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_ack => AFB_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_data => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
      CONTROL_REGISTER_pipe_write_req => CONTROL_REGISTER_pipe_write_req(0 downto 0),
      CONTROL_REGISTER_pipe_write_ack => CONTROL_REGISTER_pipe_write_ack(0 downto 0),
      CONTROL_REGISTER_pipe_write_data => CONTROL_REGISTER_pipe_write_data(31 downto 0),
      NUMBER_OF_SERVERS_pipe_write_req => NUMBER_OF_SERVERS_pipe_write_req(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_ack => NUMBER_OF_SERVERS_pipe_write_ack(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_data => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(0 downto 0),
      UpdateRegister_call_acks => UpdateRegister_call_acks(0 downto 0),
      UpdateRegister_call_data => UpdateRegister_call_data(73 downto 0),
      UpdateRegister_call_tag => UpdateRegister_call_tag(0 downto 0),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(0 downto 0),
      UpdateRegister_return_acks => UpdateRegister_return_acks(0 downto 0),
      UpdateRegister_return_data => UpdateRegister_return_data(31 downto 0),
      UpdateRegister_return_tag => UpdateRegister_return_tag(0 downto 0),
      tag_in => SoftwareRegisterAccessDaemon_tag_in,
      tag_out => SoftwareRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  SoftwareRegisterAccessDaemon_tag_in <= (others => '0');
  SoftwareRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => SoftwareRegisterAccessDaemon_start_req, start_ack => SoftwareRegisterAccessDaemon_start_ack,  fin_req => SoftwareRegisterAccessDaemon_fin_req,  fin_ack => SoftwareRegisterAccessDaemon_fin_ack);
  -- module UpdateRegister
  UpdateRegister_bmask <= UpdateRegister_in_args(73 downto 70);
  UpdateRegister_rval <= UpdateRegister_in_args(69 downto 38);
  UpdateRegister_wdata <= UpdateRegister_in_args(37 downto 6);
  UpdateRegister_index <= UpdateRegister_in_args(5 downto 0);
  UpdateRegister_out_args <= UpdateRegister_wval ;
  -- call arbiter for module UpdateRegister
  UpdateRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 74,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => UpdateRegister_call_reqs,
      call_acks => UpdateRegister_call_acks,
      return_reqs => UpdateRegister_return_reqs,
      return_acks => UpdateRegister_return_acks,
      call_data  => UpdateRegister_call_data,
      call_tag  => UpdateRegister_call_tag,
      return_tag  => UpdateRegister_return_tag,
      call_mtag => UpdateRegister_tag_in,
      return_mtag => UpdateRegister_tag_out,
      return_data =>UpdateRegister_return_data,
      call_mreq => UpdateRegister_start_req,
      call_mack => UpdateRegister_start_ack,
      return_mreq => UpdateRegister_fin_req,
      return_mack => UpdateRegister_fin_ack,
      call_mdata => UpdateRegister_in_args,
      return_mdata => UpdateRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  UpdateRegister_instance:UpdateRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      bmask => UpdateRegister_bmask,
      rval => UpdateRegister_rval,
      wdata => UpdateRegister_wdata,
      index => UpdateRegister_index,
      wval => UpdateRegister_wval,
      start_req => UpdateRegister_start_req,
      start_ack => UpdateRegister_start_ack,
      fin_req => UpdateRegister_fin_req,
      fin_ack => UpdateRegister_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(5 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => UpdateRegister_tag_in,
      tag_out => UpdateRegister_tag_out-- 
    ); -- 
  -- module accessMemory
  accessMemory_lock <= accessMemory_in_args(109 downto 109);
  accessMemory_rwbar <= accessMemory_in_args(108 downto 108);
  accessMemory_bmask <= accessMemory_in_args(107 downto 100);
  accessMemory_addr <= accessMemory_in_args(99 downto 64);
  accessMemory_wdata <= accessMemory_in_args(63 downto 0);
  accessMemory_out_args <= accessMemory_rdata ;
  -- call arbiter for module accessMemory
  accessMemory_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 11,
      call_data_width => 110,
      return_data_width => 64,
      callee_tag_length => 4,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessMemory_call_reqs,
      call_acks => accessMemory_call_acks,
      return_reqs => accessMemory_return_reqs,
      return_acks => accessMemory_return_acks,
      call_data  => accessMemory_call_data,
      call_tag  => accessMemory_call_tag,
      return_tag  => accessMemory_return_tag,
      call_mtag => accessMemory_tag_in,
      return_mtag => accessMemory_tag_out,
      return_data =>accessMemory_return_data,
      call_mreq => accessMemory_start_req,
      call_mack => accessMemory_start_ack,
      return_mreq => accessMemory_fin_req,
      return_mack => accessMemory_fin_ack,
      call_mdata => accessMemory_in_args,
      return_mdata => accessMemory_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemory_instance:accessMemory-- 
    generic map(tag_length => 6)
    port map(-- 
      lock => accessMemory_lock,
      rwbar => accessMemory_rwbar,
      bmask => accessMemory_bmask,
      addr => accessMemory_addr,
      wdata => accessMemory_wdata,
      rdata => accessMemory_rdata,
      start_req => accessMemory_start_req,
      start_ack => accessMemory_start_ack,
      fin_req => accessMemory_fin_req,
      fin_ack => accessMemory_fin_ack,
      clk => clk,
      reset => reset,
      MEMORY_TO_NIC_RESPONSE_pipe_read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessMemory_tag_in,
      tag_out => accessMemory_tag_out-- 
    ); -- 
  -- module acquireMutex
  acquireMutex_q_base_address <= acquireMutex_in_args(35 downto 0);
  acquireMutex_out_args <= acquireMutex_m_ok ;
  -- call arbiter for module acquireMutex
  acquireMutex_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => acquireMutex_call_reqs,
      call_acks => acquireMutex_call_acks,
      return_reqs => acquireMutex_return_reqs,
      return_acks => acquireMutex_return_acks,
      call_data  => acquireMutex_call_data,
      call_tag  => acquireMutex_call_tag,
      return_tag  => acquireMutex_return_tag,
      call_mtag => acquireMutex_tag_in,
      return_mtag => acquireMutex_tag_out,
      return_data =>acquireMutex_return_data,
      call_mreq => acquireMutex_start_req,
      call_mack => acquireMutex_start_ack,
      return_mreq => acquireMutex_fin_req,
      return_mack => acquireMutex_fin_ack,
      call_mdata => acquireMutex_in_args,
      return_mdata => acquireMutex_out_args,
      clk => clk, 
      reset => reset --
    ); --
  acquireMutex_instance:acquireMutex-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => acquireMutex_q_base_address,
      m_ok => acquireMutex_m_ok,
      start_req => acquireMutex_start_req,
      start_ack => acquireMutex_start_ack,
      fin_req => acquireMutex_fin_req,
      fin_ack => acquireMutex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(6 downto 6),
      accessMemory_call_acks => accessMemory_call_acks(6 downto 6),
      accessMemory_call_data => accessMemory_call_data(769 downto 660),
      accessMemory_call_tag => accessMemory_call_tag(13 downto 12),
      accessMemory_return_reqs => accessMemory_return_reqs(6 downto 6),
      accessMemory_return_acks => accessMemory_return_acks(6 downto 6),
      accessMemory_return_data => accessMemory_return_data(447 downto 384),
      accessMemory_return_tag => accessMemory_return_tag(13 downto 12),
      tag_in => acquireMutex_tag_in,
      tag_out => acquireMutex_tag_out-- 
    ); -- 
  -- module getQueueElement
  getQueueElement_q_base_address <= getQueueElement_in_args(67 downto 32);
  getQueueElement_read_pointer <= getQueueElement_in_args(31 downto 0);
  getQueueElement_out_args <= getQueueElement_q_r_data ;
  -- call arbiter for module getQueueElement
  getQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 68,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueElement_call_reqs,
      call_acks => getQueueElement_call_acks,
      return_reqs => getQueueElement_return_reqs,
      return_acks => getQueueElement_return_acks,
      call_data  => getQueueElement_call_data,
      call_tag  => getQueueElement_call_tag,
      return_tag  => getQueueElement_return_tag,
      call_mtag => getQueueElement_tag_in,
      return_mtag => getQueueElement_tag_out,
      return_data =>getQueueElement_return_data,
      call_mreq => getQueueElement_start_req,
      call_mack => getQueueElement_start_ack,
      return_mreq => getQueueElement_fin_req,
      return_mack => getQueueElement_fin_ack,
      call_mdata => getQueueElement_in_args,
      return_mdata => getQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueElement_instance:getQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => getQueueElement_q_base_address,
      read_pointer => getQueueElement_read_pointer,
      q_r_data => getQueueElement_q_r_data,
      start_req => getQueueElement_start_req,
      start_ack => getQueueElement_start_ack,
      fin_req => getQueueElement_fin_req,
      fin_ack => getQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(8 downto 8),
      accessMemory_call_acks => accessMemory_call_acks(8 downto 8),
      accessMemory_call_data => accessMemory_call_data(989 downto 880),
      accessMemory_call_tag => accessMemory_call_tag(17 downto 16),
      accessMemory_return_reqs => accessMemory_return_reqs(8 downto 8),
      accessMemory_return_acks => accessMemory_return_acks(8 downto 8),
      accessMemory_return_data => accessMemory_return_data(575 downto 512),
      accessMemory_return_tag => accessMemory_return_tag(17 downto 16),
      tag_in => getQueueElement_tag_in,
      tag_out => getQueueElement_tag_out-- 
    ); -- 
  -- module getQueuePointers
  getQueuePointers_q_base_address <= getQueuePointers_in_args(35 downto 0);
  getQueuePointers_out_args <= getQueuePointers_wp & getQueuePointers_rp ;
  -- call arbiter for module getQueuePointers
  getQueuePointers_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointers_call_reqs,
      call_acks => getQueuePointers_call_acks,
      return_reqs => getQueuePointers_return_reqs,
      return_acks => getQueuePointers_return_acks,
      call_data  => getQueuePointers_call_data,
      call_tag  => getQueuePointers_call_tag,
      return_tag  => getQueuePointers_return_tag,
      call_mtag => getQueuePointers_tag_in,
      return_mtag => getQueuePointers_tag_out,
      return_data =>getQueuePointers_return_data,
      call_mreq => getQueuePointers_start_req,
      call_mack => getQueuePointers_start_ack,
      return_mreq => getQueuePointers_fin_req,
      return_mack => getQueuePointers_fin_ack,
      call_mdata => getQueuePointers_in_args,
      return_mdata => getQueuePointers_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointers_instance:getQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueuePointers_q_base_address,
      wp => getQueuePointers_wp,
      rp => getQueuePointers_rp,
      start_req => getQueuePointers_start_req,
      start_ack => getQueuePointers_start_ack,
      fin_req => getQueuePointers_fin_req,
      fin_ack => getQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(7 downto 7),
      accessMemory_call_acks => accessMemory_call_acks(7 downto 7),
      accessMemory_call_data => accessMemory_call_data(879 downto 770),
      accessMemory_call_tag => accessMemory_call_tag(15 downto 14),
      accessMemory_return_reqs => accessMemory_return_reqs(7 downto 7),
      accessMemory_return_acks => accessMemory_return_acks(7 downto 7),
      accessMemory_return_data => accessMemory_return_data(511 downto 448),
      accessMemory_return_tag => accessMemory_return_tag(15 downto 14),
      tag_in => getQueuePointers_tag_in,
      tag_out => getQueuePointers_tag_out-- 
    ); -- 
  -- module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_queue_index <= getTxPacketPointerFromServer_in_args(5 downto 0);
  getTxPacketPointerFromServer_out_args <= getTxPacketPointerFromServer_pkt_pointer & getTxPacketPointerFromServer_status ;
  -- call arbiter for module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 6,
      return_data_width => 33,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTxPacketPointerFromServer_call_reqs,
      call_acks => getTxPacketPointerFromServer_call_acks,
      return_reqs => getTxPacketPointerFromServer_return_reqs,
      return_acks => getTxPacketPointerFromServer_return_acks,
      call_data  => getTxPacketPointerFromServer_call_data,
      call_tag  => getTxPacketPointerFromServer_call_tag,
      return_tag  => getTxPacketPointerFromServer_return_tag,
      call_mtag => getTxPacketPointerFromServer_tag_in,
      return_mtag => getTxPacketPointerFromServer_tag_out,
      return_data =>getTxPacketPointerFromServer_return_data,
      call_mreq => getTxPacketPointerFromServer_start_req,
      call_mack => getTxPacketPointerFromServer_start_ack,
      return_mreq => getTxPacketPointerFromServer_fin_req,
      return_mack => getTxPacketPointerFromServer_fin_ack,
      call_mdata => getTxPacketPointerFromServer_in_args,
      return_mdata => getTxPacketPointerFromServer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTxPacketPointerFromServer_instance:getTxPacketPointerFromServer-- 
    generic map(tag_length => 2)
    port map(-- 
      queue_index => getTxPacketPointerFromServer_queue_index,
      pkt_pointer => getTxPacketPointerFromServer_pkt_pointer,
      status => getTxPacketPointerFromServer_status,
      start_req => getTxPacketPointerFromServer_start_req,
      start_ack => getTxPacketPointerFromServer_start_ack,
      fin_req => getTxPacketPointerFromServer_fin_req,
      fin_ack => getTxPacketPointerFromServer_fin_ack,
      clk => clk,
      reset => reset,
      AccessRegister_call_reqs => AccessRegister_call_reqs(0 downto 0),
      AccessRegister_call_acks => AccessRegister_call_acks(0 downto 0),
      AccessRegister_call_data => AccessRegister_call_data(42 downto 0),
      AccessRegister_call_tag => AccessRegister_call_tag(0 downto 0),
      AccessRegister_return_reqs => AccessRegister_return_reqs(0 downto 0),
      AccessRegister_return_acks => AccessRegister_return_acks(0 downto 0),
      AccessRegister_return_data => AccessRegister_return_data(31 downto 0),
      AccessRegister_return_tag => AccessRegister_return_tag(0 downto 0),
      popFromQueue_call_reqs => popFromQueue_call_reqs(0 downto 0),
      popFromQueue_call_acks => popFromQueue_call_acks(0 downto 0),
      popFromQueue_call_data => popFromQueue_call_data(36 downto 0),
      popFromQueue_call_tag => popFromQueue_call_tag(0 downto 0),
      popFromQueue_return_reqs => popFromQueue_return_reqs(0 downto 0),
      popFromQueue_return_acks => popFromQueue_return_acks(0 downto 0),
      popFromQueue_return_data => popFromQueue_return_data(32 downto 0),
      popFromQueue_return_tag => popFromQueue_return_tag(0 downto 0),
      tag_in => getTxPacketPointerFromServer_tag_in,
      tag_out => getTxPacketPointerFromServer_tag_out-- 
    ); -- 
  -- module loadBuffer
  loadBuffer_rx_buffer_pointer <= loadBuffer_in_args(35 downto 0);
  loadBuffer_out_args <= loadBuffer_bad_packet_identifier ;
  -- call arbiter for module loadBuffer
  loadBuffer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadBuffer_call_reqs,
      call_acks => loadBuffer_call_acks,
      return_reqs => loadBuffer_return_reqs,
      return_acks => loadBuffer_return_acks,
      call_data  => loadBuffer_call_data,
      call_tag  => loadBuffer_call_tag,
      return_tag  => loadBuffer_return_tag,
      call_mtag => loadBuffer_tag_in,
      return_mtag => loadBuffer_tag_out,
      return_data =>loadBuffer_return_data,
      call_mreq => loadBuffer_start_req,
      call_mack => loadBuffer_start_ack,
      return_mreq => loadBuffer_fin_req,
      return_mack => loadBuffer_fin_ack,
      call_mdata => loadBuffer_in_args,
      return_mdata => loadBuffer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  loadBuffer_instance:loadBuffer-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => loadBuffer_rx_buffer_pointer,
      bad_packet_identifier => loadBuffer_bad_packet_identifier,
      start_req => loadBuffer_start_req,
      start_ack => loadBuffer_start_ack,
      fin_req => loadBuffer_fin_req,
      fin_ack => loadBuffer_fin_ack,
      clk => clk,
      reset => reset,
      writeEthernetHeaderToMem_call_reqs => writeEthernetHeaderToMem_call_reqs(0 downto 0),
      writeEthernetHeaderToMem_call_acks => writeEthernetHeaderToMem_call_acks(0 downto 0),
      writeEthernetHeaderToMem_call_data => writeEthernetHeaderToMem_call_data(35 downto 0),
      writeEthernetHeaderToMem_call_tag => writeEthernetHeaderToMem_call_tag(0 downto 0),
      writeEthernetHeaderToMem_return_reqs => writeEthernetHeaderToMem_return_reqs(0 downto 0),
      writeEthernetHeaderToMem_return_acks => writeEthernetHeaderToMem_return_acks(0 downto 0),
      writeEthernetHeaderToMem_return_data => writeEthernetHeaderToMem_return_data(35 downto 0),
      writeEthernetHeaderToMem_return_tag => writeEthernetHeaderToMem_return_tag(0 downto 0),
      writePayloadToMem_call_reqs => writePayloadToMem_call_reqs(0 downto 0),
      writePayloadToMem_call_acks => writePayloadToMem_call_acks(0 downto 0),
      writePayloadToMem_call_data => writePayloadToMem_call_data(71 downto 0),
      writePayloadToMem_call_tag => writePayloadToMem_call_tag(0 downto 0),
      writePayloadToMem_return_reqs => writePayloadToMem_return_reqs(0 downto 0),
      writePayloadToMem_return_acks => writePayloadToMem_return_acks(0 downto 0),
      writePayloadToMem_return_data => writePayloadToMem_return_data(16 downto 0),
      writePayloadToMem_return_tag => writePayloadToMem_return_tag(0 downto 0),
      writeControlInformationToMem_call_reqs => writeControlInformationToMem_call_reqs(0 downto 0),
      writeControlInformationToMem_call_acks => writeControlInformationToMem_call_acks(0 downto 0),
      writeControlInformationToMem_call_data => writeControlInformationToMem_call_data(51 downto 0),
      writeControlInformationToMem_call_tag => writeControlInformationToMem_call_tag(0 downto 0),
      writeControlInformationToMem_return_reqs => writeControlInformationToMem_return_reqs(0 downto 0),
      writeControlInformationToMem_return_acks => writeControlInformationToMem_return_acks(0 downto 0),
      writeControlInformationToMem_return_tag => writeControlInformationToMem_return_tag(0 downto 0),
      tag_in => loadBuffer_tag_in,
      tag_out => loadBuffer_tag_out-- 
    ); -- 
  -- module nicRxFromMacDaemon
  nicRxFromMacDaemon_instance:nicRxFromMacDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicRxFromMacDaemon_start_req,
      start_ack => nicRxFromMacDaemon_start_ack,
      fin_req => nicRxFromMacDaemon_fin_req,
      fin_ack => nicRxFromMacDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      mac_to_nic_data_pipe_read_req => mac_to_nic_data_pipe_read_req(0 downto 0),
      mac_to_nic_data_pipe_read_ack => mac_to_nic_data_pipe_read_ack(0 downto 0),
      mac_to_nic_data_pipe_read_data => mac_to_nic_data_pipe_read_data(72 downto 0),
      nic_rx_to_packet_pipe_write_req => nic_rx_to_packet_pipe_write_req(0 downto 0),
      nic_rx_to_packet_pipe_write_ack => nic_rx_to_packet_pipe_write_ack(0 downto 0),
      nic_rx_to_packet_pipe_write_data => nic_rx_to_packet_pipe_write_data(72 downto 0),
      nic_rx_to_header_pipe_write_req => nic_rx_to_header_pipe_write_req(0 downto 0),
      nic_rx_to_header_pipe_write_ack => nic_rx_to_header_pipe_write_ack(0 downto 0),
      nic_rx_to_header_pipe_write_data => nic_rx_to_header_pipe_write_data(72 downto 0),
      tag_in => nicRxFromMacDaemon_tag_in,
      tag_out => nicRxFromMacDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicRxFromMacDaemon_tag_in <= (others => '0');
  nicRxFromMacDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicRxFromMacDaemon_start_req, start_ack => nicRxFromMacDaemon_start_ack,  fin_req => nicRxFromMacDaemon_fin_req,  fin_ack => nicRxFromMacDaemon_fin_ack);
  -- module popFromQueue
  popFromQueue_lock <= popFromQueue_in_args(36 downto 36);
  popFromQueue_q_base_address <= popFromQueue_in_args(35 downto 0);
  popFromQueue_out_args <= popFromQueue_q_r_data & popFromQueue_status ;
  -- call arbiter for module popFromQueue
  popFromQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 37,
      return_data_width => 33,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => popFromQueue_call_reqs,
      call_acks => popFromQueue_call_acks,
      return_reqs => popFromQueue_return_reqs,
      return_acks => popFromQueue_return_acks,
      call_data  => popFromQueue_call_data,
      call_tag  => popFromQueue_call_tag,
      return_tag  => popFromQueue_return_tag,
      call_mtag => popFromQueue_tag_in,
      return_mtag => popFromQueue_tag_out,
      return_data =>popFromQueue_return_data,
      call_mreq => popFromQueue_start_req,
      call_mack => popFromQueue_start_ack,
      return_mreq => popFromQueue_fin_req,
      return_mack => popFromQueue_fin_ack,
      call_mdata => popFromQueue_in_args,
      return_mdata => popFromQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  popFromQueue_instance:popFromQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => popFromQueue_lock,
      q_base_address => popFromQueue_q_base_address,
      q_r_data => popFromQueue_q_r_data,
      status => popFromQueue_status,
      start_req => popFromQueue_start_req,
      start_ack => popFromQueue_start_ack,
      fin_req => popFromQueue_fin_req,
      fin_ack => popFromQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireMutex_call_reqs => acquireMutex_call_reqs(1 downto 1),
      acquireMutex_call_acks => acquireMutex_call_acks(1 downto 1),
      acquireMutex_call_data => acquireMutex_call_data(71 downto 36),
      acquireMutex_call_tag => acquireMutex_call_tag(1 downto 1),
      acquireMutex_return_reqs => acquireMutex_return_reqs(1 downto 1),
      acquireMutex_return_acks => acquireMutex_return_acks(1 downto 1),
      acquireMutex_return_data => acquireMutex_return_data(1 downto 1),
      acquireMutex_return_tag => acquireMutex_return_tag(1 downto 1),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(1 downto 1),
      getQueuePointers_call_acks => getQueuePointers_call_acks(1 downto 1),
      getQueuePointers_call_data => getQueuePointers_call_data(71 downto 36),
      getQueuePointers_call_tag => getQueuePointers_call_tag(1 downto 1),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(1 downto 1),
      getQueuePointers_return_acks => getQueuePointers_return_acks(1 downto 1),
      getQueuePointers_return_data => getQueuePointers_return_data(127 downto 64),
      getQueuePointers_return_tag => getQueuePointers_return_tag(1 downto 1),
      getQueueElement_call_reqs => getQueueElement_call_reqs(0 downto 0),
      getQueueElement_call_acks => getQueueElement_call_acks(0 downto 0),
      getQueueElement_call_data => getQueueElement_call_data(67 downto 0),
      getQueueElement_call_tag => getQueueElement_call_tag(0 downto 0),
      getQueueElement_return_reqs => getQueueElement_return_reqs(0 downto 0),
      getQueueElement_return_acks => getQueueElement_return_acks(0 downto 0),
      getQueueElement_return_data => getQueueElement_return_data(31 downto 0),
      getQueueElement_return_tag => getQueueElement_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(1 downto 1),
      setQueuePointers_call_acks => setQueuePointers_call_acks(1 downto 1),
      setQueuePointers_call_data => setQueuePointers_call_data(199 downto 100),
      setQueuePointers_call_tag => setQueuePointers_call_tag(1 downto 1),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(1 downto 1),
      setQueuePointers_return_acks => setQueuePointers_return_acks(1 downto 1),
      setQueuePointers_return_tag => setQueuePointers_return_tag(1 downto 1),
      releaseMutex_call_reqs => releaseMutex_call_reqs(1 downto 1),
      releaseMutex_call_acks => releaseMutex_call_acks(1 downto 1),
      releaseMutex_call_data => releaseMutex_call_data(71 downto 36),
      releaseMutex_call_tag => releaseMutex_call_tag(1 downto 1),
      releaseMutex_return_reqs => releaseMutex_return_reqs(1 downto 1),
      releaseMutex_return_acks => releaseMutex_return_acks(1 downto 1),
      releaseMutex_return_tag => releaseMutex_return_tag(1 downto 1),
      tag_in => popFromQueue_tag_in,
      tag_out => popFromQueue_tag_out-- 
    ); -- 
  -- module populateRxQueue
  populateRxQueue_rx_buffer_pointer <= populateRxQueue_in_args(35 downto 0);
  -- call arbiter for module populateRxQueue
  populateRxQueue_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => populateRxQueue_call_reqs,
      call_acks => populateRxQueue_call_acks,
      return_reqs => populateRxQueue_return_reqs,
      return_acks => populateRxQueue_return_acks,
      call_data  => populateRxQueue_call_data,
      call_tag  => populateRxQueue_call_tag,
      return_tag  => populateRxQueue_return_tag,
      call_mtag => populateRxQueue_tag_in,
      return_mtag => populateRxQueue_tag_out,
      call_mreq => populateRxQueue_start_req,
      call_mack => populateRxQueue_start_ack,
      return_mreq => populateRxQueue_fin_req,
      return_mack => populateRxQueue_fin_ack,
      call_mdata => populateRxQueue_in_args,
      clk => clk, 
      reset => reset --
    ); --
  populateRxQueue_instance:populateRxQueue-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => populateRxQueue_rx_buffer_pointer,
      start_req => populateRxQueue_start_req,
      start_ack => populateRxQueue_start_ack,
      fin_req => populateRxQueue_fin_req,
      fin_ack => populateRxQueue_fin_ack,
      clk => clk,
      reset => reset,
      LAST_WRITTEN_RX_QUEUE_INDEX => LAST_WRITTEN_RX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(11 downto 6),
      AccessRegister_call_reqs => AccessRegister_call_reqs(1 downto 1),
      AccessRegister_call_acks => AccessRegister_call_acks(1 downto 1),
      AccessRegister_call_data => AccessRegister_call_data(85 downto 43),
      AccessRegister_call_tag => AccessRegister_call_tag(1 downto 1),
      AccessRegister_return_reqs => AccessRegister_return_reqs(1 downto 1),
      AccessRegister_return_acks => AccessRegister_return_acks(1 downto 1),
      AccessRegister_return_data => AccessRegister_return_data(63 downto 32),
      AccessRegister_return_tag => AccessRegister_return_tag(1 downto 1),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(2 downto 2),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(2 downto 2),
      pushIntoQueue_call_data => pushIntoQueue_call_data(206 downto 138),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(2 downto 2),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(2 downto 2),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(2 downto 2),
      pushIntoQueue_return_data => pushIntoQueue_return_data(2 downto 2),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(2 downto 2),
      tag_in => populateRxQueue_tag_in,
      tag_out => populateRxQueue_tag_out-- 
    ); -- 
  -- module pushIntoQueue
  pushIntoQueue_lock <= pushIntoQueue_in_args(68 downto 68);
  pushIntoQueue_q_base_address <= pushIntoQueue_in_args(67 downto 32);
  pushIntoQueue_q_w_data <= pushIntoQueue_in_args(31 downto 0);
  pushIntoQueue_out_args <= pushIntoQueue_status ;
  -- call arbiter for module pushIntoQueue
  pushIntoQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 69,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => pushIntoQueue_call_reqs,
      call_acks => pushIntoQueue_call_acks,
      return_reqs => pushIntoQueue_return_reqs,
      return_acks => pushIntoQueue_return_acks,
      call_data  => pushIntoQueue_call_data,
      call_tag  => pushIntoQueue_call_tag,
      return_tag  => pushIntoQueue_return_tag,
      call_mtag => pushIntoQueue_tag_in,
      return_mtag => pushIntoQueue_tag_out,
      return_data =>pushIntoQueue_return_data,
      call_mreq => pushIntoQueue_start_req,
      call_mack => pushIntoQueue_start_ack,
      return_mreq => pushIntoQueue_fin_req,
      return_mack => pushIntoQueue_fin_ack,
      call_mdata => pushIntoQueue_in_args,
      return_mdata => pushIntoQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  pushIntoQueue_instance:pushIntoQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => pushIntoQueue_lock,
      q_base_address => pushIntoQueue_q_base_address,
      q_w_data => pushIntoQueue_q_w_data,
      status => pushIntoQueue_status,
      start_req => pushIntoQueue_start_req,
      start_ack => pushIntoQueue_start_ack,
      fin_req => pushIntoQueue_fin_req,
      fin_ack => pushIntoQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireMutex_call_reqs => acquireMutex_call_reqs(0 downto 0),
      acquireMutex_call_acks => acquireMutex_call_acks(0 downto 0),
      acquireMutex_call_data => acquireMutex_call_data(35 downto 0),
      acquireMutex_call_tag => acquireMutex_call_tag(0 downto 0),
      acquireMutex_return_reqs => acquireMutex_return_reqs(0 downto 0),
      acquireMutex_return_acks => acquireMutex_return_acks(0 downto 0),
      acquireMutex_return_data => acquireMutex_return_data(0 downto 0),
      acquireMutex_return_tag => acquireMutex_return_tag(0 downto 0),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(0 downto 0),
      getQueuePointers_call_acks => getQueuePointers_call_acks(0 downto 0),
      getQueuePointers_call_data => getQueuePointers_call_data(35 downto 0),
      getQueuePointers_call_tag => getQueuePointers_call_tag(0 downto 0),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(0 downto 0),
      getQueuePointers_return_acks => getQueuePointers_return_acks(0 downto 0),
      getQueuePointers_return_data => getQueuePointers_return_data(63 downto 0),
      getQueuePointers_return_tag => getQueuePointers_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(0 downto 0),
      setQueuePointers_call_acks => setQueuePointers_call_acks(0 downto 0),
      setQueuePointers_call_data => setQueuePointers_call_data(99 downto 0),
      setQueuePointers_call_tag => setQueuePointers_call_tag(0 downto 0),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(0 downto 0),
      setQueuePointers_return_acks => setQueuePointers_return_acks(0 downto 0),
      setQueuePointers_return_tag => setQueuePointers_return_tag(0 downto 0),
      releaseMutex_call_reqs => releaseMutex_call_reqs(0 downto 0),
      releaseMutex_call_acks => releaseMutex_call_acks(0 downto 0),
      releaseMutex_call_data => releaseMutex_call_data(35 downto 0),
      releaseMutex_call_tag => releaseMutex_call_tag(0 downto 0),
      releaseMutex_return_reqs => releaseMutex_return_reqs(0 downto 0),
      releaseMutex_return_acks => releaseMutex_return_acks(0 downto 0),
      releaseMutex_return_tag => releaseMutex_return_tag(0 downto 0),
      setQueueElement_call_reqs => setQueueElement_call_reqs(0 downto 0),
      setQueueElement_call_acks => setQueueElement_call_acks(0 downto 0),
      setQueueElement_call_data => setQueueElement_call_data(99 downto 0),
      setQueueElement_call_tag => setQueueElement_call_tag(0 downto 0),
      setQueueElement_return_reqs => setQueueElement_return_reqs(0 downto 0),
      setQueueElement_return_acks => setQueueElement_return_acks(0 downto 0),
      setQueueElement_return_tag => setQueueElement_return_tag(0 downto 0),
      tag_in => pushIntoQueue_tag_in,
      tag_out => pushIntoQueue_tag_out-- 
    ); -- 
  -- module releaseMutex
  releaseMutex_q_base_address <= releaseMutex_in_args(35 downto 0);
  -- call arbiter for module releaseMutex
  releaseMutex_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 36,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => releaseMutex_call_reqs,
      call_acks => releaseMutex_call_acks,
      return_reqs => releaseMutex_return_reqs,
      return_acks => releaseMutex_return_acks,
      call_data  => releaseMutex_call_data,
      call_tag  => releaseMutex_call_tag,
      return_tag  => releaseMutex_return_tag,
      call_mtag => releaseMutex_tag_in,
      return_mtag => releaseMutex_tag_out,
      call_mreq => releaseMutex_start_req,
      call_mack => releaseMutex_start_ack,
      return_mreq => releaseMutex_fin_req,
      return_mack => releaseMutex_fin_ack,
      call_mdata => releaseMutex_in_args,
      clk => clk, 
      reset => reset --
    ); --
  releaseMutex_instance:releaseMutex-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => releaseMutex_q_base_address,
      start_req => releaseMutex_start_req,
      start_ack => releaseMutex_start_ack,
      fin_req => releaseMutex_fin_req,
      fin_ack => releaseMutex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(10 downto 10),
      accessMemory_call_acks => accessMemory_call_acks(10 downto 10),
      accessMemory_call_data => accessMemory_call_data(1209 downto 1100),
      accessMemory_call_tag => accessMemory_call_tag(21 downto 20),
      accessMemory_return_reqs => accessMemory_return_reqs(10 downto 10),
      accessMemory_return_acks => accessMemory_return_acks(10 downto 10),
      accessMemory_return_data => accessMemory_return_data(703 downto 640),
      accessMemory_return_tag => accessMemory_return_tag(21 downto 20),
      tag_in => releaseMutex_tag_in,
      tag_out => releaseMutex_tag_out-- 
    ); -- 
  -- module setQueueElement
  setQueueElement_q_base_address <= setQueueElement_in_args(99 downto 64);
  setQueueElement_write_pointer <= setQueueElement_in_args(63 downto 32);
  setQueueElement_q_w_data <= setQueueElement_in_args(31 downto 0);
  -- call arbiter for module setQueueElement
  setQueueElement_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 100,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueueElement_call_reqs,
      call_acks => setQueueElement_call_acks,
      return_reqs => setQueueElement_return_reqs,
      return_acks => setQueueElement_return_acks,
      call_data  => setQueueElement_call_data,
      call_tag  => setQueueElement_call_tag,
      return_tag  => setQueueElement_return_tag,
      call_mtag => setQueueElement_tag_in,
      return_mtag => setQueueElement_tag_out,
      call_mreq => setQueueElement_start_req,
      call_mack => setQueueElement_start_ack,
      return_mreq => setQueueElement_fin_req,
      return_mack => setQueueElement_fin_ack,
      call_mdata => setQueueElement_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueueElement_instance:setQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => setQueueElement_q_base_address,
      write_pointer => setQueueElement_write_pointer,
      q_w_data => setQueueElement_q_w_data,
      start_req => setQueueElement_start_req,
      start_ack => setQueueElement_start_ack,
      fin_req => setQueueElement_fin_req,
      fin_ack => setQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(2 downto 2),
      accessMemory_call_acks => accessMemory_call_acks(2 downto 2),
      accessMemory_call_data => accessMemory_call_data(329 downto 220),
      accessMemory_call_tag => accessMemory_call_tag(5 downto 4),
      accessMemory_return_reqs => accessMemory_return_reqs(2 downto 2),
      accessMemory_return_acks => accessMemory_return_acks(2 downto 2),
      accessMemory_return_data => accessMemory_return_data(191 downto 128),
      accessMemory_return_tag => accessMemory_return_tag(5 downto 4),
      tag_in => setQueueElement_tag_in,
      tag_out => setQueueElement_tag_out-- 
    ); -- 
  -- module setQueuePointers
  setQueuePointers_q_base_address <= setQueuePointers_in_args(99 downto 64);
  setQueuePointers_wp <= setQueuePointers_in_args(63 downto 32);
  setQueuePointers_rp <= setQueuePointers_in_args(31 downto 0);
  -- call arbiter for module setQueuePointers
  setQueuePointers_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 100,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueuePointers_call_reqs,
      call_acks => setQueuePointers_call_acks,
      return_reqs => setQueuePointers_return_reqs,
      return_acks => setQueuePointers_return_acks,
      call_data  => setQueuePointers_call_data,
      call_tag  => setQueuePointers_call_tag,
      return_tag  => setQueuePointers_return_tag,
      call_mtag => setQueuePointers_tag_in,
      return_mtag => setQueuePointers_tag_out,
      call_mreq => setQueuePointers_start_req,
      call_mack => setQueuePointers_start_ack,
      return_mreq => setQueuePointers_fin_req,
      return_mack => setQueuePointers_fin_ack,
      call_mdata => setQueuePointers_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueuePointers_instance:setQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => setQueuePointers_q_base_address,
      wp => setQueuePointers_wp,
      rp => setQueuePointers_rp,
      start_req => setQueuePointers_start_req,
      start_ack => setQueuePointers_start_ack,
      fin_req => setQueuePointers_fin_req,
      fin_ack => setQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(9 downto 9),
      accessMemory_call_acks => accessMemory_call_acks(9 downto 9),
      accessMemory_call_data => accessMemory_call_data(1099 downto 990),
      accessMemory_call_tag => accessMemory_call_tag(19 downto 18),
      accessMemory_return_reqs => accessMemory_return_reqs(9 downto 9),
      accessMemory_return_acks => accessMemory_return_acks(9 downto 9),
      accessMemory_return_data => accessMemory_return_data(639 downto 576),
      accessMemory_return_tag => accessMemory_return_tag(19 downto 18),
      tag_in => setQueuePointers_tag_in,
      tag_out => setQueuePointers_tag_out-- 
    ); -- 
  -- module transmitEngineDaemon
  transmitEngineDaemon_instance:transmitEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => transmitEngineDaemon_start_req,
      start_ack => transmitEngineDaemon_start_ack,
      fin_req => transmitEngineDaemon_fin_req,
      fin_ack => transmitEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      FREE_Q => FREE_Q,
      LAST_READ_TX_QUEUE_INDEX => LAST_READ_TX_QUEUE_INDEX,
      CONTROL_REGISTER => CONTROL_REGISTER,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(0 downto 0),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(0 downto 0),
      pushIntoQueue_call_data => pushIntoQueue_call_data(68 downto 0),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(0 downto 0),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(0 downto 0),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(0 downto 0),
      pushIntoQueue_return_data => pushIntoQueue_return_data(0 downto 0),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(0 downto 0),
      getTxPacketPointerFromServer_call_reqs => getTxPacketPointerFromServer_call_reqs(0 downto 0),
      getTxPacketPointerFromServer_call_acks => getTxPacketPointerFromServer_call_acks(0 downto 0),
      getTxPacketPointerFromServer_call_data => getTxPacketPointerFromServer_call_data(5 downto 0),
      getTxPacketPointerFromServer_call_tag => getTxPacketPointerFromServer_call_tag(0 downto 0),
      getTxPacketPointerFromServer_return_reqs => getTxPacketPointerFromServer_return_reqs(0 downto 0),
      getTxPacketPointerFromServer_return_acks => getTxPacketPointerFromServer_return_acks(0 downto 0),
      getTxPacketPointerFromServer_return_data => getTxPacketPointerFromServer_return_data(32 downto 0),
      getTxPacketPointerFromServer_return_tag => getTxPacketPointerFromServer_return_tag(0 downto 0),
      transmitPacket_call_reqs => transmitPacket_call_reqs(0 downto 0),
      transmitPacket_call_acks => transmitPacket_call_acks(0 downto 0),
      transmitPacket_call_data => transmitPacket_call_data(31 downto 0),
      transmitPacket_call_tag => transmitPacket_call_tag(0 downto 0),
      transmitPacket_return_reqs => transmitPacket_return_reqs(0 downto 0),
      transmitPacket_return_acks => transmitPacket_return_acks(0 downto 0),
      transmitPacket_return_data => transmitPacket_return_data(0 downto 0),
      transmitPacket_return_tag => transmitPacket_return_tag(0 downto 0),
      tag_in => transmitEngineDaemon_tag_in,
      tag_out => transmitEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  transmitEngineDaemon_tag_in <= (others => '0');
  transmitEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => transmitEngineDaemon_start_req, start_ack => transmitEngineDaemon_start_ack,  fin_req => transmitEngineDaemon_fin_req,  fin_ack => transmitEngineDaemon_fin_ack);
  -- module transmitPacket
  transmitPacket_packet_pointer <= transmitPacket_in_args(31 downto 0);
  transmitPacket_out_args <= transmitPacket_status ;
  -- call arbiter for module transmitPacket
  transmitPacket_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => transmitPacket_call_reqs,
      call_acks => transmitPacket_call_acks,
      return_reqs => transmitPacket_return_reqs,
      return_acks => transmitPacket_return_acks,
      call_data  => transmitPacket_call_data,
      call_tag  => transmitPacket_call_tag,
      return_tag  => transmitPacket_return_tag,
      call_mtag => transmitPacket_tag_in,
      return_mtag => transmitPacket_tag_out,
      return_data =>transmitPacket_return_data,
      call_mreq => transmitPacket_start_req,
      call_mack => transmitPacket_start_ack,
      return_mreq => transmitPacket_fin_req,
      return_mack => transmitPacket_fin_ack,
      call_mdata => transmitPacket_in_args,
      return_mdata => transmitPacket_out_args,
      clk => clk, 
      reset => reset --
    ); --
  transmitPacket_instance:transmitPacket-- 
    generic map(tag_length => 2)
    port map(-- 
      packet_pointer => transmitPacket_packet_pointer,
      status => transmitPacket_status,
      start_req => transmitPacket_start_req,
      start_ack => transmitPacket_start_ack,
      fin_req => transmitPacket_fin_req,
      fin_ack => transmitPacket_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_write_req => nic_to_mac_transmit_pipe_pipe_write_req(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_ack => nic_to_mac_transmit_pipe_pipe_write_ack(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_data => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(1 downto 0),
      accessMemory_call_acks => accessMemory_call_acks(1 downto 0),
      accessMemory_call_data => accessMemory_call_data(219 downto 0),
      accessMemory_call_tag => accessMemory_call_tag(3 downto 0),
      accessMemory_return_reqs => accessMemory_return_reqs(1 downto 0),
      accessMemory_return_acks => accessMemory_return_acks(1 downto 0),
      accessMemory_return_data => accessMemory_return_data(127 downto 0),
      accessMemory_return_tag => accessMemory_return_tag(3 downto 0),
      tag_in => transmitPacket_tag_in,
      tag_out => transmitPacket_tag_out-- 
    ); -- 
  -- module writeControlInformationToMem
  writeControlInformationToMem_base_buffer_pointer <= writeControlInformationToMem_in_args(51 downto 16);
  writeControlInformationToMem_packet_size <= writeControlInformationToMem_in_args(15 downto 8);
  writeControlInformationToMem_last_keep <= writeControlInformationToMem_in_args(7 downto 0);
  -- call arbiter for module writeControlInformationToMem
  writeControlInformationToMem_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 52,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeControlInformationToMem_call_reqs,
      call_acks => writeControlInformationToMem_call_acks,
      return_reqs => writeControlInformationToMem_return_reqs,
      return_acks => writeControlInformationToMem_return_acks,
      call_data  => writeControlInformationToMem_call_data,
      call_tag  => writeControlInformationToMem_call_tag,
      return_tag  => writeControlInformationToMem_return_tag,
      call_mtag => writeControlInformationToMem_tag_in,
      return_mtag => writeControlInformationToMem_tag_out,
      call_mreq => writeControlInformationToMem_start_req,
      call_mack => writeControlInformationToMem_start_ack,
      return_mreq => writeControlInformationToMem_fin_req,
      return_mack => writeControlInformationToMem_fin_ack,
      call_mdata => writeControlInformationToMem_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeControlInformationToMem_instance:writeControlInformationToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buffer_pointer => writeControlInformationToMem_base_buffer_pointer,
      packet_size => writeControlInformationToMem_packet_size,
      last_keep => writeControlInformationToMem_last_keep,
      start_req => writeControlInformationToMem_start_req,
      start_ack => writeControlInformationToMem_start_ack,
      fin_req => writeControlInformationToMem_fin_req,
      fin_ack => writeControlInformationToMem_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(5 downto 5),
      accessMemory_call_acks => accessMemory_call_acks(5 downto 5),
      accessMemory_call_data => accessMemory_call_data(659 downto 550),
      accessMemory_call_tag => accessMemory_call_tag(11 downto 10),
      accessMemory_return_reqs => accessMemory_return_reqs(5 downto 5),
      accessMemory_return_acks => accessMemory_return_acks(5 downto 5),
      accessMemory_return_data => accessMemory_return_data(383 downto 320),
      accessMemory_return_tag => accessMemory_return_tag(11 downto 10),
      tag_in => writeControlInformationToMem_tag_in,
      tag_out => writeControlInformationToMem_tag_out-- 
    ); -- 
  -- module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_buf_pointer <= writeEthernetHeaderToMem_in_args(35 downto 0);
  writeEthernetHeaderToMem_out_args <= writeEthernetHeaderToMem_buf_position ;
  -- call arbiter for module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeEthernetHeaderToMem_call_reqs,
      call_acks => writeEthernetHeaderToMem_call_acks,
      return_reqs => writeEthernetHeaderToMem_return_reqs,
      return_acks => writeEthernetHeaderToMem_return_acks,
      call_data  => writeEthernetHeaderToMem_call_data,
      call_tag  => writeEthernetHeaderToMem_call_tag,
      return_tag  => writeEthernetHeaderToMem_return_tag,
      call_mtag => writeEthernetHeaderToMem_tag_in,
      return_mtag => writeEthernetHeaderToMem_tag_out,
      return_data =>writeEthernetHeaderToMem_return_data,
      call_mreq => writeEthernetHeaderToMem_start_req,
      call_mack => writeEthernetHeaderToMem_start_ack,
      return_mreq => writeEthernetHeaderToMem_fin_req,
      return_mack => writeEthernetHeaderToMem_fin_ack,
      call_mdata => writeEthernetHeaderToMem_in_args,
      return_mdata => writeEthernetHeaderToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeEthernetHeaderToMem_instance:writeEthernetHeaderToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      buf_pointer => writeEthernetHeaderToMem_buf_pointer,
      buf_position => writeEthernetHeaderToMem_buf_position,
      start_req => writeEthernetHeaderToMem_start_req,
      start_ack => writeEthernetHeaderToMem_start_ack,
      fin_req => writeEthernetHeaderToMem_fin_req,
      fin_ack => writeEthernetHeaderToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_header_pipe_read_req => nic_rx_to_header_pipe_read_req(0 downto 0),
      nic_rx_to_header_pipe_read_ack => nic_rx_to_header_pipe_read_ack(0 downto 0),
      nic_rx_to_header_pipe_read_data => nic_rx_to_header_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(4 downto 4),
      accessMemory_call_acks => accessMemory_call_acks(4 downto 4),
      accessMemory_call_data => accessMemory_call_data(549 downto 440),
      accessMemory_call_tag => accessMemory_call_tag(9 downto 8),
      accessMemory_return_reqs => accessMemory_return_reqs(4 downto 4),
      accessMemory_return_acks => accessMemory_return_acks(4 downto 4),
      accessMemory_return_data => accessMemory_return_data(319 downto 256),
      accessMemory_return_tag => accessMemory_return_tag(9 downto 8),
      tag_in => writeEthernetHeaderToMem_tag_in,
      tag_out => writeEthernetHeaderToMem_tag_out-- 
    ); -- 
  -- module writePayloadToMem
  writePayloadToMem_base_buf_pointer <= writePayloadToMem_in_args(71 downto 36);
  writePayloadToMem_buf_pointer <= writePayloadToMem_in_args(35 downto 0);
  writePayloadToMem_out_args <= writePayloadToMem_packet_size_32 & writePayloadToMem_bad_packet_identifier & writePayloadToMem_last_keep ;
  -- call arbiter for module writePayloadToMem
  writePayloadToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 17,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writePayloadToMem_call_reqs,
      call_acks => writePayloadToMem_call_acks,
      return_reqs => writePayloadToMem_return_reqs,
      return_acks => writePayloadToMem_return_acks,
      call_data  => writePayloadToMem_call_data,
      call_tag  => writePayloadToMem_call_tag,
      return_tag  => writePayloadToMem_return_tag,
      call_mtag => writePayloadToMem_tag_in,
      return_mtag => writePayloadToMem_tag_out,
      return_data =>writePayloadToMem_return_data,
      call_mreq => writePayloadToMem_start_req,
      call_mack => writePayloadToMem_start_ack,
      return_mreq => writePayloadToMem_fin_req,
      return_mack => writePayloadToMem_fin_ack,
      call_mdata => writePayloadToMem_in_args,
      return_mdata => writePayloadToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writePayloadToMem_instance:writePayloadToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buf_pointer => writePayloadToMem_base_buf_pointer,
      buf_pointer => writePayloadToMem_buf_pointer,
      packet_size_32 => writePayloadToMem_packet_size_32,
      bad_packet_identifier => writePayloadToMem_bad_packet_identifier,
      last_keep => writePayloadToMem_last_keep,
      start_req => writePayloadToMem_start_req,
      start_ack => writePayloadToMem_start_ack,
      fin_req => writePayloadToMem_fin_req,
      fin_ack => writePayloadToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_packet_pipe_read_req => nic_rx_to_packet_pipe_read_req(0 downto 0),
      nic_rx_to_packet_pipe_read_ack => nic_rx_to_packet_pipe_read_ack(0 downto 0),
      nic_rx_to_packet_pipe_read_data => nic_rx_to_packet_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(3 downto 3),
      accessMemory_call_acks => accessMemory_call_acks(3 downto 3),
      accessMemory_call_data => accessMemory_call_data(439 downto 330),
      accessMemory_call_tag => accessMemory_call_tag(7 downto 6),
      accessMemory_return_reqs => accessMemory_return_reqs(3 downto 3),
      accessMemory_return_acks => accessMemory_return_acks(3 downto 3),
      accessMemory_return_data => accessMemory_return_data(255 downto 192),
      accessMemory_return_tag => accessMemory_return_tag(7 downto 6),
      tag_in => writePayloadToMem_tag_in,
      tag_out => writePayloadToMem_tag_out-- 
    ); -- 
  AFB_NIC_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 74,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_REQUEST_pipe_read_req,
      read_ack => AFB_NIC_REQUEST_pipe_read_ack,
      read_data => AFB_NIC_REQUEST_pipe_read_data,
      write_req => AFB_NIC_REQUEST_pipe_write_req,
      write_ack => AFB_NIC_REQUEST_pipe_write_ack,
      write_data => AFB_NIC_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  AFB_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => AFB_NIC_RESPONSE_pipe_read_req,
      read_ack => AFB_NIC_RESPONSE_pipe_read_ack,
      read_data => AFB_NIC_RESPONSE_pipe_read_data,
      write_req => AFB_NIC_RESPONSE_pipe_write_req,
      write_ack => AFB_NIC_RESPONSE_pipe_write_ack,
      write_data => AFB_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  CONTROL_REGISTER_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe CONTROL_REGISTER",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => CONTROL_REGISTER,
      write_req => CONTROL_REGISTER_pipe_write_req,
      write_ack => CONTROL_REGISTER_pipe_write_ack,
      write_data => CONTROL_REGISTER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  FREE_Q_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe FREE_Q",
      volatile_flag => false,
      num_writes => 1,
      data_width => 36 --
    ) 
    port map( -- 
      read_data => FREE_Q,
      write_req => FREE_Q_pipe_write_req,
      write_ack => FREE_Q_pipe_write_ack,
      write_data => FREE_Q_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_READ_TX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_READ_TX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_READ_TX_QUEUE_INDEX,
      write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_WRITTEN_RX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_WRITTEN_RX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_WRITTEN_RX_QUEUE_INDEX,
      write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEMORY_TO_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEMORY_TO_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req,
      read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack,
      read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data,
      write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req,
      write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack,
      write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_REQUEST_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_REQUEST_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 43,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_RESPONSE_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_TO_MEMORY_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_TO_MEMORY_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req,
      read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack,
      read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data,
      write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req,
      write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack,
      write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NUMBER_OF_SERVERS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NUMBER_OF_SERVERS",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => NUMBER_OF_SERVERS,
      write_req => NUMBER_OF_SERVERS_pipe_write_req,
      write_ack => NUMBER_OF_SERVERS_pipe_write_ack,
      write_data => NUMBER_OF_SERVERS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => mac_to_nic_data_pipe_read_req,
      read_ack => mac_to_nic_data_pipe_read_ack,
      read_data => mac_to_nic_data_pipe_read_data,
      write_req => mac_to_nic_data_pipe_write_req,
      write_ack => mac_to_nic_data_pipe_write_ack,
      write_data => mac_to_nic_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_header_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_header",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 16 --
    )
    port map( -- 
      read_req => nic_rx_to_header_pipe_read_req,
      read_ack => nic_rx_to_header_pipe_read_ack,
      read_data => nic_rx_to_header_pipe_read_data,
      write_req => nic_rx_to_header_pipe_write_req,
      write_ack => nic_rx_to_header_pipe_write_ack,
      write_data => nic_rx_to_header_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_packet_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_packet",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 16 --
    )
    port map( -- 
      read_req => nic_rx_to_packet_pipe_read_req,
      read_ack => nic_rx_to_packet_pipe_read_ack,
      read_data => nic_rx_to_packet_pipe_read_data,
      write_req => nic_rx_to_packet_pipe_write_req,
      write_ack => nic_rx_to_packet_pipe_write_ack,
      write_data => nic_rx_to_packet_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_to_mac_transmit_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_to_mac_transmit_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => nic_to_mac_transmit_pipe_pipe_read_req,
      read_ack => nic_to_mac_transmit_pipe_pipe_read_ack,
      read_data => nic_to_mac_transmit_pipe_pipe_read_data,
      write_req => nic_to_mac_transmit_pipe_pipe_write_req,
      write_ack => nic_to_mac_transmit_pipe_pipe_write_ack,
      write_data => nic_to_mac_transmit_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 6,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 6,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
