-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package tx_deconcat_system_global_package is -- 
  -- 
end package tx_deconcat_system_global_package;
