-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity AccessRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(3 downto 0);
    register_index : in  std_logic_vector(5 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity AccessRegister;
architecture AccessRegister_arch of AccessRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 43)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal register_index_buffer :  std_logic_vector(5 downto 0);
  signal register_index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal AccessRegister_CP_0_start: Boolean;
  signal AccessRegister_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_1 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "AccessRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 43) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(4 downto 1) <= bmask;
  bmask_buffer <= in_buffer_data_out(4 downto 1);
  in_buffer_data_in(10 downto 5) <= register_index;
  register_index_buffer <= in_buffer_data_out(10 downto 5);
  in_buffer_data_in(42 downto 11) <= wdata;
  wdata_buffer <= in_buffer_data_out(42 downto 11);
  in_buffer_data_in(tag_length + 42 downto 43) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 42 downto 43);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  AccessRegister_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "AccessRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,AccessRegister_CP_0_start,"AccessRegister cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,AccessRegister_CP_0_symbol, "AccessRegister cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  AccessRegister_CP_0: Block -- control-path 
    signal AccessRegister_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    AccessRegister_CP_0_elements(0) <= AccessRegister_CP_0_start;
    AccessRegister_CP_0_symbol <= AccessRegister_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_92_to_assign_stmt_106/$entry
      -- CP-element group 0: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_sample_start_
      -- CP-element group 0: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Sample/req
      -- CP-element group 0: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_sample_start_
      -- CP-element group 0: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Sample/$entry
      -- 
    -- logger for CP element group AccessRegister_CP_0_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and AccessRegister_CP_0_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:AccessRegister_CP_0_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_0); -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_sample_completed_
      -- CP-element group 1: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_update_start_
      -- CP-element group 1: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Sample/ack
      -- CP-element group 1: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Update/$entry
      -- CP-element group 1: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Update/req
      -- 
    -- logger for CP element group AccessRegister_CP_0_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and AccessRegister_CP_0_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:AccessRegister_CP_0_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_0, ack => AccessRegister_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(1), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_update_completed_
      -- CP-element group 2: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Update/$exit
      -- CP-element group 2: 	 assign_stmt_92_to_assign_stmt_106/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_Update/ack
      -- 
    -- logger for CP element group AccessRegister_CP_0_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and AccessRegister_CP_0_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:AccessRegister_CP_0_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_1, ack => AccessRegister_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Sample/ra
      -- CP-element group 3: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Update/$entry
      -- CP-element group 3: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_sample_completed_
      -- CP-element group 3: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_update_start_
      -- CP-element group 3: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Update/cr
      -- 
    -- logger for CP element group AccessRegister_CP_0_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and AccessRegister_CP_0_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:AccessRegister_CP_0_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_0, ack => AccessRegister_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(3), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Update/$exit
      -- CP-element group 4: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_update_completed_
      -- CP-element group 4: 	 assign_stmt_92_to_assign_stmt_106/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_Update/ca
      -- 
    -- logger for CP element group AccessRegister_CP_0_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and AccessRegister_CP_0_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:AccessRegister_CP_0_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_1, ack => AccessRegister_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_92_to_assign_stmt_106/$exit
      -- 
    -- logger for CP element group AccessRegister_CP_0_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and AccessRegister_CP_0_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:AccessRegister:CP:AccessRegister_CP_0_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    AccessRegister_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "AccessRegister_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= AccessRegister_CP_0_elements(2) & AccessRegister_CP_0_elements(4);
      gj_AccessRegister_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => AccessRegister_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u5_87_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u6_u38_90_wire : std_logic_vector(37 downto 0);
    signal request_92 : std_logic_vector(42 downto 0);
    signal response_98 : std_logic_vector(32 downto 0);
    signal status_102 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- logger for split-operator slice_101_inst flow-through 
    process(status_102) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:slice_101_inst:flowthrough inputs: " & " response_98 = "& Convert_SLV_To_Hex_String(response_98) & " outputs:" & " status_102= "  & Convert_SLV_To_Hex_String(status_102));
      --
    end process; 
    -- flow-through slice operator slice_101_inst
    status_102 <= response_98(32 downto 32);
    -- logger for split-operator slice_105_inst flow-through 
    process(rdata_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:slice_105_inst:flowthrough inputs: " & " response_98 = "& Convert_SLV_To_Hex_String(response_98) & " outputs:" & " rdata_buffer= "  & Convert_SLV_To_Hex_String(rdata_buffer));
      --
    end process; 
    -- flow-through slice operator slice_105_inst
    rdata_buffer <= response_98(31 downto 0);
    -- logger for split-operator CONCAT_u1_u5_87_inst flow-through 
    process(CONCAT_u1_u5_87_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:CONCAT_u1_u5_87_inst:flowthrough inputs: " & " rwbar_buffer = "& Convert_SLV_To_Hex_String(rwbar_buffer) & " bmask_buffer = "& Convert_SLV_To_Hex_String(bmask_buffer) & " outputs:" & " CONCAT_u1_u5_87_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u5_87_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u5_87_inst
    process(rwbar_buffer, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(rwbar_buffer, bmask_buffer, tmp_var);
      CONCAT_u1_u5_87_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u5_u43_91_inst flow-through 
    process(request_92) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:CONCAT_u5_u43_91_inst:flowthrough inputs: " & " CONCAT_u1_u5_87_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u5_87_wire) & " CONCAT_u6_u38_90_wire = "& Convert_SLV_To_Hex_String(CONCAT_u6_u38_90_wire) & " outputs:" & " request_92= "  & Convert_SLV_To_Hex_String(request_92));
      --
    end process; 
    -- binary operator CONCAT_u5_u43_91_inst
    process(CONCAT_u1_u5_87_wire, CONCAT_u6_u38_90_wire) -- 
      variable tmp_var : std_logic_vector(42 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_87_wire, CONCAT_u6_u38_90_wire, tmp_var);
      request_92 <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u6_u38_90_inst flow-through 
    process(CONCAT_u6_u38_90_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:CONCAT_u6_u38_90_inst:flowthrough inputs: " & " register_index_buffer = "& Convert_SLV_To_Hex_String(register_index_buffer) & " wdata_buffer = "& Convert_SLV_To_Hex_String(wdata_buffer) & " outputs:" & " CONCAT_u6_u38_90_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u6_u38_90_wire));
      --
    end process; 
    -- binary operator CONCAT_u6_u38_90_inst
    process(register_index_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(37 downto 0); -- 
    begin -- 
      ApConcat_proc(register_index_buffer, wdata_buffer, tmp_var);
      CONCAT_u6_u38_90_wire <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst:started:   PipeRead from NIC_RESPONSE_REGISTER_ACCESS_PIPE inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst:finished:  outputs: " & " response_98= "  & Convert_SLV_To_Hex_String(response_98));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_0;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_req_1;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_97_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_98 <= data_out(32 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst:started:   PipeWrite to NIC_REQUEST_REGISTER_ACCESS_PIPE inputs: " & " request_92 = "& Convert_SLV_To_Hex_String(request_92));
          --
        end if; 
        if WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:AccessRegister:DP:WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_0;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_req_1;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_93_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_92;
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE", data_width => 43, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end AccessRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity NicRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity NicRegisterAccessDaemon;
architecture NicRegisterAccessDaemon_arch of NicRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal NicRegisterAccessDaemon_CP_116_start: Boolean;
  signal NicRegisterAccessDaemon_CP_116_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_1 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_1 : boolean;
  signal do_while_stmt_190_branch_req_0 : boolean;
  signal array_obj_ref_213_load_0_req_0 : boolean;
  signal array_obj_ref_213_load_0_ack_0 : boolean;
  signal array_obj_ref_213_load_0_req_1 : boolean;
  signal array_obj_ref_213_load_0_ack_1 : boolean;
  signal call_stmt_221_call_req_0 : boolean;
  signal call_stmt_221_call_ack_0 : boolean;
  signal call_stmt_221_call_req_1 : boolean;
  signal call_stmt_221_call_ack_1 : boolean;
  signal W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_0 : boolean;
  signal W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_0 : boolean;
  signal W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_1 : boolean;
  signal W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_1 : boolean;
  signal do_while_stmt_190_branch_ack_0 : boolean;
  signal do_while_stmt_190_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  NicRegisterAccessDaemon_CP_116_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_116_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,NicRegisterAccessDaemon_CP_116_start,"NicRegisterAccessDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,NicRegisterAccessDaemon_CP_116_symbol, "NicRegisterAccessDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  NicRegisterAccessDaemon_CP_116: Block -- control-path 
    signal NicRegisterAccessDaemon_CP_116_elements: BooleanArray(31 downto 0);
    -- 
  begin -- 
    NicRegisterAccessDaemon_CP_116_elements(0) <= NicRegisterAccessDaemon_CP_116_start;
    NicRegisterAccessDaemon_CP_116_symbol <= NicRegisterAccessDaemon_CP_116_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_189/$entry
      -- CP-element group 0: 	 branch_block_stmt_189/branch_block_stmt_189__entry__
      -- CP-element group 0: 	 branch_block_stmt_189/do_while_stmt_190__entry__
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	31 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_189/$exit
      -- CP-element group 1: 	 branch_block_stmt_189/branch_block_stmt_189__exit__
      -- CP-element group 1: 	 branch_block_stmt_189/do_while_stmt_190__exit__
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_CP_116_elements(1) <= NicRegisterAccessDaemon_CP_116_elements(31);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_189/do_while_stmt_190/$entry
      -- CP-element group 2: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190__entry__
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_CP_116_elements(2) <= NicRegisterAccessDaemon_CP_116_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	31 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190__exit__
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_189/do_while_stmt_190/loop_back
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	26 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	29 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_189/do_while_stmt_190/condition_done
      -- CP-element group 5: 	 branch_block_stmt_189/do_while_stmt_190/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_189/do_while_stmt_190/loop_taken/$entry
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_CP_116_elements(5) <= NicRegisterAccessDaemon_CP_116_elements(26);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	28 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_189/do_while_stmt_190/loop_body_done
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_CP_116_elements(6) <= NicRegisterAccessDaemon_CP_116_elements(28);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_CP_116_elements(7) <= NicRegisterAccessDaemon_CP_116_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_CP_116_elements(8) <= NicRegisterAccessDaemon_CP_116_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	26 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/loop_body_start
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Sample/rr
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(10), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(9) & NicRegisterAccessDaemon_CP_116_elements(13);
      gj_NicRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	20 
    -- CP-element group 11: 	24 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_update_start_
      -- CP-element group 11: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Update/cr
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(11), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(12) & NicRegisterAccessDaemon_CP_116_elements(20) & NicRegisterAccessDaemon_CP_116_elements(24);
      gj_NicRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Sample/ra
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: 	22 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (29) 
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_resized_0
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_scaled_0
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_computed_0
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_resize_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_resize_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_resize_0/index_resize_req
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_resize_0/index_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_scale_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_scale_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_scale_0/scale_rename_req
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_index_scale_0/scale_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_final_index_sum_regn/$entry
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_final_index_sum_regn/$exit
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_final_index_sum_regn/req
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_final_index_sum_regn/ack
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_word_addrgen/root_register_ack
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/word_access_start/$entry
      -- CP-element group 14: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/word_access_start/word_0/$entry
      -- CP-element group 14: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:array_obj_ref_213_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(14), ack => array_obj_ref_213_load_0_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(21) & NicRegisterAccessDaemon_CP_116_elements(16);
      gj_NicRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	24 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_update_start_
      -- CP-element group 15: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:array_obj_ref_213_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(15), ack => array_obj_ref_213_load_0_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(20) & NicRegisterAccessDaemon_CP_116_elements(24);
      gj_NicRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	27 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:array_obj_ref_213_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_load_0_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (9) 
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/array_obj_ref_213_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/array_obj_ref_213_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/array_obj_ref_213_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_Update/array_obj_ref_213_Merge/merge_ack
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:array_obj_ref_213_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_load_0_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	27 
    -- CP-element group 18: 	17 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Sample/crr
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:call_stmt_221_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(18), ack => call_stmt_221_call_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(27) & NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(20);
      gj_NicRegisterAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_update_start_
      -- CP-element group 19: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Update/ccr
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:call_stmt_221_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(19), ack => call_stmt_221_call_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(21);
      gj_NicRegisterAccessDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	11 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	15 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Sample/cra
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:call_stmt_221_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_221_call_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	28 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/call_stmt_221_Update/cca
      -- CP-element group 21: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/ring_reenable_memory_space_0
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:call_stmt_221_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_221_call_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: 	17 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Sample/req
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(22), ack => W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(13) & NicRegisterAccessDaemon_CP_116_elements(17) & NicRegisterAccessDaemon_CP_116_elements(24);
      gj_NicRegisterAccessDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_update_start_
      -- CP-element group 23: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Update/req
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(23), ack => W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_116_elements(25);
      gj_NicRegisterAccessDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	11 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	15 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Sample/ack
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/assign_stmt_237_Update/ack
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(25)); -- 
    -- CP-element group 26:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	9 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	5 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/condition_evaluated
      -- CP-element group 26: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:do_while_stmt_190_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_116_elements(26), ack => do_while_stmt_190_branch_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(26) is a control-delay.
    cp_element_26_delay: control_delay_element  generic map(name => " 26_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(9), ack => NicRegisterAccessDaemon_CP_116_elements(26), clk => clk, reset =>reset);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	16 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	18 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/array_obj_ref_213_call_stmt_221_delay
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group NicRegisterAccessDaemon_CP_116_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_116_elements(16), ack => NicRegisterAccessDaemon_CP_116_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	21 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	6 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_189/do_while_stmt_190/do_while_stmt_190_loop_body/$exit
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_116_elements(21) & NicRegisterAccessDaemon_CP_116_elements(25);
      gj_NicRegisterAccessDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	5 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_189/do_while_stmt_190/loop_exit/$exit
      -- CP-element group 29: 	 branch_block_stmt_189/do_while_stmt_190/loop_exit/ack
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:do_while_stmt_190_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_190_branch_ack_0, ack => NicRegisterAccessDaemon_CP_116_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_189/do_while_stmt_190/loop_taken/$exit
      -- CP-element group 30: 	 branch_block_stmt_189/do_while_stmt_190/loop_taken/ack
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:do_while_stmt_190_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_190_branch_ack_1, ack => NicRegisterAccessDaemon_CP_116_elements(30)); -- 
    -- CP-element group 31:  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	3 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	1 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_189/do_while_stmt_190/$exit
      -- 
    -- logger for CP element group NicRegisterAccessDaemon_CP_116_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and NicRegisterAccessDaemon_CP_116_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:NicRegisterAccessDaemon:CP:NicRegisterAccessDaemon_CP_116_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    NicRegisterAccessDaemon_CP_116_elements(31) <= NicRegisterAccessDaemon_CP_116_elements(3);
    NicRegisterAccessDaemon_do_while_stmt_190_terminator_258: loop_terminator -- 
      generic map (name => " NicRegisterAccessDaemon_do_while_stmt_190_terminator_258", max_iterations_in_flight =>31) 
      port map(loop_body_exit => NicRegisterAccessDaemon_CP_116_elements(6),loop_continue => NicRegisterAccessDaemon_CP_116_elements(30),loop_terminate => NicRegisterAccessDaemon_CP_116_elements(29),loop_back => NicRegisterAccessDaemon_CP_116_elements(4),loop_exit => NicRegisterAccessDaemon_CP_116_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_141_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= NicRegisterAccessDaemon_CP_116_elements(7);
        preds(1)  <= NicRegisterAccessDaemon_CP_116_elements(8);
        entry_tmerge_141 : transition_merge -- 
          generic map(name => " entry_tmerge_141")
          port map (preds => preds, symbol_out => NicRegisterAccessDaemon_CP_116_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NIC_RESPONE_REGISTER_ACCESS_PIPE_237 : std_logic_vector(32 downto 0);
    signal R_index_212_resized : std_logic_vector(5 downto 0);
    signal R_index_212_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_213_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_213_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_213_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_213_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_213_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_213_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_213_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_202 : std_logic_vector(3 downto 0);
    signal index_206 : std_logic_vector(5 downto 0);
    signal konst_239_wire_constant : std_logic_vector(0 downto 0);
    signal rdata_228 : std_logic_vector(31 downto 0);
    signal req_194 : std_logic_vector(42 downto 0);
    signal resp_234 : std_logic_vector(32 downto 0);
    signal rval_214 : std_logic_vector(31 downto 0);
    signal rwbar_198 : std_logic_vector(0 downto 0);
    signal type_cast_226_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_231_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_210 : std_logic_vector(31 downto 0);
    signal wval_221 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_213_offset_scale_factor_0 <= "000001";
    array_obj_ref_213_resized_base_address <= "000000";
    array_obj_ref_213_word_offset_0 <= "000000";
    konst_239_wire_constant <= "1";
    type_cast_226_wire_constant <= "00000000000000000000000000000000";
    type_cast_231_wire_constant <= "0";
    -- logger for split-operator MUX_227_inst flow-through 
    process(rdata_228) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:MUX_227_inst:flowthrough inputs: " & " rwbar_198 = "& Convert_SLV_To_Hex_String(rwbar_198) & " rval_214 = "& Convert_SLV_To_Hex_String(rval_214) & " type_cast_226_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_226_wire_constant) & " outputs:" & " rdata_228= "  & Convert_SLV_To_Hex_String(rdata_228));
      --
    end process; 
    -- flow-through select operator MUX_227_inst
    rdata_228 <= rval_214 when (rwbar_198(0) /=  '0') else type_cast_226_wire_constant;
    -- logger for split-operator slice_197_inst flow-through 
    process(rwbar_198) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:slice_197_inst:flowthrough inputs: " & " req_194 = "& Convert_SLV_To_Hex_String(req_194) & " outputs:" & " rwbar_198= "  & Convert_SLV_To_Hex_String(rwbar_198));
      --
    end process; 
    -- flow-through slice operator slice_197_inst
    rwbar_198 <= req_194(42 downto 42);
    -- logger for split-operator slice_201_inst flow-through 
    process(bmask_202) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:slice_201_inst:flowthrough inputs: " & " req_194 = "& Convert_SLV_To_Hex_String(req_194) & " outputs:" & " bmask_202= "  & Convert_SLV_To_Hex_String(bmask_202));
      --
    end process; 
    -- flow-through slice operator slice_201_inst
    bmask_202 <= req_194(41 downto 38);
    -- logger for split-operator slice_205_inst flow-through 
    process(index_206) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:slice_205_inst:flowthrough inputs: " & " req_194 = "& Convert_SLV_To_Hex_String(req_194) & " outputs:" & " index_206= "  & Convert_SLV_To_Hex_String(index_206));
      --
    end process; 
    -- flow-through slice operator slice_205_inst
    index_206 <= req_194(37 downto 32);
    -- logger for split-operator slice_209_inst flow-through 
    process(wdata_210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:slice_209_inst:flowthrough inputs: " & " req_194 = "& Convert_SLV_To_Hex_String(req_194) & " outputs:" & " wdata_210= "  & Convert_SLV_To_Hex_String(wdata_210));
      --
    end process; 
    -- flow-through slice operator slice_209_inst
    wdata_210 <= req_194(31 downto 0);
    -- logger for split-operator W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst:started:   inputs: " & " resp_234 = "& Convert_SLV_To_Hex_String(resp_234));
          --
        end if; 
        if W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst:finished:  outputs: " & " NIC_RESPONE_REGISTER_ACCESS_PIPE_237= "  & Convert_SLV_To_Hex_String(NIC_RESPONE_REGISTER_ACCESS_PIPE_237));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_0;
      W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_0<= wack(0);
      rreq(0) <= W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_req_1;
      W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst_ack_1<= rack(0);
      W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst : InterlockBuffer generic map ( -- 
        name => "W_NIC_RESPONE_REGISTER_ACCESS_PIPE_235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 33,
        out_data_width => 33,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => resp_234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => NIC_RESPONE_REGISTER_ACCESS_PIPE_237,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_213_addr_0 flow-through 
    process(array_obj_ref_213_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_addr_0:flowthrough  inputs: " & " array_obj_ref_213_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_213_root_address) & "outputs: " & " array_obj_ref_213_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_213_addr_0
    process(array_obj_ref_213_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_213_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_213_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_gather_scatter flow-through 
    process(rval_214) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_gather_scatter:flowthrough  inputs: " & " array_obj_ref_213_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_213_data_0) & "outputs: " & " rval_214= "  & Convert_SLV_To_Hex_String(rval_214));
      --
    end process; 
    -- equivalence array_obj_ref_213_gather_scatter
    process(array_obj_ref_213_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_213_data_0;
      ov(31 downto 0) := iv;
      rval_214 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_index_0_rename flow-through 
    process(R_index_212_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_index_0_rename:flowthrough  inputs: " & " R_index_212_resized = "& Convert_SLV_To_Hex_String(R_index_212_resized) & "outputs: " & " R_index_212_scaled= "  & Convert_SLV_To_Hex_String(R_index_212_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_213_index_0_rename
    process(R_index_212_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_212_resized;
      ov(5 downto 0) := iv;
      R_index_212_scaled <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_index_0_resize flow-through 
    process(R_index_212_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_index_0_resize:flowthrough  inputs: " & " index_206 = "& Convert_SLV_To_Hex_String(index_206) & "outputs: " & " R_index_212_resized= "  & Convert_SLV_To_Hex_String(R_index_212_resized));
      --
    end process; 
    -- equivalence array_obj_ref_213_index_0_resize
    process(index_206) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_206;
      ov(5 downto 0) := iv;
      R_index_212_resized <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_index_offset flow-through 
    process(array_obj_ref_213_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_index_offset:flowthrough  inputs: " & " R_index_212_scaled = "& Convert_SLV_To_Hex_String(R_index_212_scaled) & "outputs: " & " array_obj_ref_213_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_213_index_offset
    process(R_index_212_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_212_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_213_final_offset <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_213_root_address_inst flow-through 
    process(array_obj_ref_213_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_root_address_inst:flowthrough  inputs: " & " array_obj_ref_213_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_213_final_offset) & "outputs: " & " array_obj_ref_213_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_213_root_address_inst
    process(array_obj_ref_213_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_213_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_213_root_address <= ov(5 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_190_branch_req_0," req0 do_while_stmt_190_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_190_branch_ack_0," ack0 do_while_stmt_190_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_190_branch_ack_1," ack1 do_while_stmt_190_branch");
    do_while_stmt_190_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_239_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_190_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_190_branch_req_0,
          ack0 => do_while_stmt_190_branch_ack_0,
          ack1 => do_while_stmt_190_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator CONCAT_u1_u33_233_inst flow-through 
    process(resp_234) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:CONCAT_u1_u33_233_inst:flowthrough inputs: " & " type_cast_231_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_231_wire_constant) & " rdata_228 = "& Convert_SLV_To_Hex_String(rdata_228) & " outputs:" & " resp_234= "  & Convert_SLV_To_Hex_String(resp_234));
      --
    end process; 
    -- binary operator CONCAT_u1_u33_233_inst
    process(type_cast_231_wire_constant, rdata_228) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_231_wire_constant, rdata_228, tmp_var);
      resp_234 <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_213_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_213_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_load_0:started:   inputs: " & " array_obj_ref_213_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_213_word_address_0));
          --
        end if; 
        if array_obj_ref_213_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:array_obj_ref_213_load_0:finished:  outputs: " & " array_obj_ref_213_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_213_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_213_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_213_load_0_req_0,
        array_obj_ref_213_load_0_ack_0,
        array_obj_ref_213_load_0_req_1,
        array_obj_ref_213_load_0_ack_1,
        "array_obj_ref_213_load_0",
        "memory_space_0" ,
        array_obj_ref_213_data_0,
        array_obj_ref_213_word_address_0,
        "array_obj_ref_213_data_0",
        "array_obj_ref_213_word_address_0" -- 
      );
      reqL_unguarded(0) <= array_obj_ref_213_load_0_req_0;
      array_obj_ref_213_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_213_load_0_req_1;
      array_obj_ref_213_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_213_word_address_0;
      array_obj_ref_213_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst:started:   PipeRead from NIC_REQUEST_REGISTER_ACCESS_PIPE inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst:finished:  outputs: " & " req_194= "  & Convert_SLV_To_Hex_String(req_194));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(42 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_0;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_req_1;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_193_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_194 <= data_out(42 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0", data_width => 43,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator call_stmt_221_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_221_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:call_stmt_221_call:started:  Call to module UpdateRegister inputs: " & " rwbar_198 (guard complement )= " & Convert_SLV_To_String(rwbar_198) & " bmask_202 = "& Convert_SLV_To_Hex_String(bmask_202) & " rval_214 = "& Convert_SLV_To_Hex_String(rval_214) & " wdata_210 = "& Convert_SLV_To_Hex_String(wdata_210) & " index_206 = "& Convert_SLV_To_Hex_String(index_206));
          --
        end if; 
        if call_stmt_221_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:NicRegisterAccessDaemon:DP:call_stmt_221_call:finished:  outputs: " & " wval_221= "  & Convert_SLV_To_Hex_String(wval_221));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_221_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_221_call_req_0;
      call_stmt_221_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_221_call_req_1;
      call_stmt_221_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_198(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_202 & rval_214 & wdata_210 & index_206;
      wval_221 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end NicRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ReceiveEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_call_data : out  std_logic_vector(35 downto 0);
    loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
    loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_return_data : in   std_logic_vector(0 downto 0);
    loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
    populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ReceiveEngineDaemon;
architecture ReceiveEngineDaemon_arch of ReceiveEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ReceiveEngineDaemon_CP_1451_start: Boolean;
  signal ReceiveEngineDaemon_CP_1451_symbol: Boolean;
  -- volatile/operator module components. 
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_899_call_ack_0 : boolean;
  signal call_stmt_927_call_req_1 : boolean;
  signal call_stmt_911_call_req_0 : boolean;
  signal if_stmt_884_branch_ack_0 : boolean;
  signal call_stmt_911_call_ack_0 : boolean;
  signal call_stmt_899_call_req_1 : boolean;
  signal call_stmt_927_call_ack_1 : boolean;
  signal call_stmt_899_call_ack_1 : boolean;
  signal if_stmt_884_branch_req_0 : boolean;
  signal call_stmt_911_call_req_1 : boolean;
  signal call_stmt_911_call_ack_1 : boolean;
  signal if_stmt_884_branch_ack_1 : boolean;
  signal call_stmt_899_call_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_1 : boolean;
  signal call_stmt_937_call_ack_1 : boolean;
  signal call_stmt_937_call_ack_0 : boolean;
  signal do_while_stmt_891_branch_ack_0 : boolean;
  signal call_stmt_937_call_req_0 : boolean;
  signal do_while_stmt_891_branch_ack_1 : boolean;
  signal call_stmt_927_call_ack_0 : boolean;
  signal do_while_stmt_891_branch_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_0 : boolean;
  signal call_stmt_927_call_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_0 : boolean;
  signal call_stmt_937_call_req_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ReceiveEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ReceiveEngineDaemon_CP_1451_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ReceiveEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1451_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1451_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_1451_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,ReceiveEngineDaemon_CP_1451_start,"ReceiveEngineDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,ReceiveEngineDaemon_CP_1451_symbol, "ReceiveEngineDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ReceiveEngineDaemon_CP_1451: Block -- control-path 
    signal ReceiveEngineDaemon_CP_1451_elements: BooleanArray(35 downto 0);
    -- 
  begin -- 
    ReceiveEngineDaemon_CP_1451_elements(0) <= ReceiveEngineDaemon_CP_1451_start;
    ReceiveEngineDaemon_CP_1451_symbol <= ReceiveEngineDaemon_CP_1451_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_880/$entry
      -- CP-element group 0: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Sample/req
      -- CP-element group 0: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_sample_start_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(0), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Update/req
      -- CP-element group 1: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Update/$entry
      -- CP-element group 1: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Sample/ack
      -- CP-element group 1: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_update_start_
      -- CP-element group 1: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_sample_completed_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_0, ack => ReceiveEngineDaemon_CP_1451_elements(1)); -- 
    req_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(1), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	35 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 branch_block_stmt_881/branch_block_stmt_881__entry__
      -- CP-element group 2: 	 branch_block_stmt_881/merge_stmt_882__entry__
      -- CP-element group 2: 	 assign_stmt_880/$exit
      -- CP-element group 2: 	 branch_block_stmt_881/$entry
      -- CP-element group 2: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Update/ack
      -- CP-element group 2: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_881/merge_stmt_882_dead_link/$entry
      -- CP-element group 2: 	 assign_stmt_880/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_881/merge_stmt_882__entry___PhiReq/$exit
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_1, ack => ReceiveEngineDaemon_CP_1451_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_881/branch_block_stmt_881__exit__
      -- CP-element group 3: 	 branch_block_stmt_881/$exit
      -- CP-element group 3: 	 $exit
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	34 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	35 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_881/do_while_stmt_891__exit__
      -- CP-element group 4: 	 branch_block_stmt_881/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_881/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_881/disable_loopback_PhiReq/$exit
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(4) <= ReceiveEngineDaemon_CP_1451_elements(34);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	35 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	35 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_881/if_stmt_884_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_881/if_stmt_884_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_881/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_881/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_881/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:if_stmt_884_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_884_branch_ack_1, ack => ReceiveEngineDaemon_CP_1451_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	35 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_881/if_stmt_884__exit__
      -- CP-element group 6: 	 branch_block_stmt_881/if_stmt_884_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_881/do_while_stmt_891__entry__
      -- CP-element group 6: 	 branch_block_stmt_881/if_stmt_884_else_link/$exit
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:if_stmt_884_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_884_branch_ack_0, ack => ReceiveEngineDaemon_CP_1451_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891__entry__
      -- CP-element group 7: 	 branch_block_stmt_881/do_while_stmt_891/$entry
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(7) <= ReceiveEngineDaemon_CP_1451_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	34 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891__exit__
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group ReceiveEngineDaemon_CP_1451_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_881/do_while_stmt_891/loop_back
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group ReceiveEngineDaemon_CP_1451_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	31 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	32 
    -- CP-element group 10: 	33 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_881/do_while_stmt_891/condition_done
      -- CP-element group 10: 	 branch_block_stmt_881/do_while_stmt_891/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_881/do_while_stmt_891/loop_taken/$entry
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(10) <= ReceiveEngineDaemon_CP_1451_elements(31);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	30 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_881/do_while_stmt_891/loop_body_done
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(11) <= ReceiveEngineDaemon_CP_1451_elements(30);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(12) <= ReceiveEngineDaemon_CP_1451_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(13) <= ReceiveEngineDaemon_CP_1451_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/loop_body_start
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group ReceiveEngineDaemon_CP_1451_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	30 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Sample/crr
      -- CP-element group 15: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_sample_start_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_899_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(15), ack => call_stmt_899_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1451_elements(14) & ReceiveEngineDaemon_CP_1451_elements(17) & ReceiveEngineDaemon_CP_1451_elements(30);
      gj_ReceiveEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	25 
    -- CP-element group 16: 	29 
    -- CP-element group 16: 	30 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Update/ccr
      -- CP-element group 16: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_update_start_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_899_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(16), ack => call_stmt_899_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1451_elements(21) & ReceiveEngineDaemon_CP_1451_elements(25) & ReceiveEngineDaemon_CP_1451_elements(29) & ReceiveEngineDaemon_CP_1451_elements(30);
      gj_ReceiveEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Sample/cra
      -- CP-element group 17: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_sample_completed_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_899_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_899_call_ack_0, ack => ReceiveEngineDaemon_CP_1451_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	23 
    -- CP-element group 18: 	27 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Update/cca
      -- CP-element group 18: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_899_update_completed_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_899_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_899_call_ack_1, ack => ReceiveEngineDaemon_CP_1451_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Sample/crr
      -- CP-element group 19: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_sample_start_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_911_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(19), ack => call_stmt_911_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1451_elements(18) & ReceiveEngineDaemon_CP_1451_elements(21);
      gj_ReceiveEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	25 
    -- CP-element group 20: 	29 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Update/ccr
      -- CP-element group 20: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_update_start_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_911_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(20), ack => call_stmt_911_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1451_elements(25) & ReceiveEngineDaemon_CP_1451_elements(29);
      gj_ReceiveEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Sample/cra
      -- CP-element group 21: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_sample_completed_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_911_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_911_call_ack_0, ack => ReceiveEngineDaemon_CP_1451_elements(21)); -- 
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_Update/cca
      -- CP-element group 22: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_911_update_completed_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_911_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_911_call_ack_1, ack => ReceiveEngineDaemon_CP_1451_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	18 
    -- CP-element group 23: 	22 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Sample/crr
      -- CP-element group 23: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Sample/$entry
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_927_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(23), ack => call_stmt_927_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1451_elements(18) & ReceiveEngineDaemon_CP_1451_elements(22) & ReceiveEngineDaemon_CP_1451_elements(25);
      gj_ReceiveEngineDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_update_start_
      -- CP-element group 24: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Update/ccr
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_927_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(24), ack => call_stmt_927_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1451_elements(26);
      gj_ReceiveEngineDaemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	16 
    -- CP-element group 25: 	20 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Sample/cra
      -- CP-element group 25: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Sample/$exit
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_927_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_927_call_ack_0, ack => ReceiveEngineDaemon_CP_1451_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_927_Update/cca
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_927_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_927_call_ack_1, ack => ReceiveEngineDaemon_CP_1451_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	18 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	26 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Sample/crr
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_937_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(27), ack => call_stmt_937_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_1451_elements(18) & ReceiveEngineDaemon_CP_1451_elements(22) & ReceiveEngineDaemon_CP_1451_elements(26) & ReceiveEngineDaemon_CP_1451_elements(29);
      gj_ReceiveEngineDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_update_start_
      -- CP-element group 28: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Update/ccr
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_937_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_1603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(28), ack => call_stmt_937_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_1451_elements(30);
      gj_ReceiveEngineDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Sample/cra
      -- CP-element group 29: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_sample_completed_
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_937_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_937_call_ack_0, ack => ReceiveEngineDaemon_CP_1451_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	11 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: 	16 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/$exit
      -- CP-element group 30: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/call_stmt_937_Update/cca
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:call_stmt_937_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_937_call_ack_1, ack => ReceiveEngineDaemon_CP_1451_elements(30)); -- 
    -- CP-element group 31:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	14 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	10 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/loop_body_delay_to_condition_start
      -- CP-element group 31: 	 branch_block_stmt_881/do_while_stmt_891/do_while_stmt_891_loop_body/condition_evaluated
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:do_while_stmt_891_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_1547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(31), ack => do_while_stmt_891_branch_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_1451_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_1451_elements(14), ack => ReceiveEngineDaemon_CP_1451_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	10 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_881/do_while_stmt_891/loop_exit/$exit
      -- CP-element group 32: 	 branch_block_stmt_881/do_while_stmt_891/loop_exit/ack
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:do_while_stmt_891_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_891_branch_ack_0, ack => ReceiveEngineDaemon_CP_1451_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	10 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_881/do_while_stmt_891/loop_taken/$exit
      -- CP-element group 33: 	 branch_block_stmt_881/do_while_stmt_891/loop_taken/ack
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:do_while_stmt_891_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_891_branch_ack_1, ack => ReceiveEngineDaemon_CP_1451_elements(33)); -- 
    -- CP-element group 34:  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	8 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	4 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_881/do_while_stmt_891/$exit
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    ReceiveEngineDaemon_CP_1451_elements(34) <= ReceiveEngineDaemon_CP_1451_elements(8);
    -- CP-element group 35:  merge  branch  transition  place  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	5 
    -- CP-element group 35: 	4 
    -- CP-element group 35: 	2 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	5 
    -- CP-element group 35: 	6 
    -- CP-element group 35:  members (37) 
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Update/ack
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884__entry__
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/BITSEL_u32_u1_887_place
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/merge_stmt_882__exit__
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_if_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/branch_req
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_else_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_dead_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Update/cr
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/SplitProtocol/Update/ca
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Update/req
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Sample/req
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/if_stmt_884_eval_test/BITSEL_u32_u1_887/BITSEL_u32_u1_887_inputs/RPIPE_CONTROL_REGISTER_885/Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/merge_stmt_882_PhiReqMerge
      -- CP-element group 35: 	 branch_block_stmt_881/merge_stmt_882_PhiAck/$entry
      -- CP-element group 35: 	 branch_block_stmt_881/merge_stmt_882_PhiAck/$exit
      -- CP-element group 35: 	 branch_block_stmt_881/merge_stmt_882_PhiAck/dummy
      -- 
    -- logger for CP element group ReceiveEngineDaemon_CP_1451_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and ReceiveEngineDaemon_CP_1451_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:ReceiveEngineDaemon_CP_1451_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:ReceiveEngineDaemon:CP:if_stmt_884_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_1451_elements(35), ack => if_stmt_884_branch_req_0); -- 
    ReceiveEngineDaemon_CP_1451_elements(35) <= OrReduce(ReceiveEngineDaemon_CP_1451_elements(5) & ReceiveEngineDaemon_CP_1451_elements(4) & ReceiveEngineDaemon_CP_1451_elements(2));
    ReceiveEngineDaemon_do_while_stmt_891_terminator_1614: loop_terminator -- 
      generic map (name => " ReceiveEngineDaemon_do_while_stmt_891_terminator_1614", max_iterations_in_flight =>31) 
      port map(loop_body_exit => ReceiveEngineDaemon_CP_1451_elements(11),loop_continue => ReceiveEngineDaemon_CP_1451_elements(33),loop_terminate => ReceiveEngineDaemon_CP_1451_elements(32),loop_back => ReceiveEngineDaemon_CP_1451_elements(9),loop_exit => ReceiveEngineDaemon_CP_1451_elements(8),clk => clk, reset => reset); -- 
    entry_tmerge_1548_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ReceiveEngineDaemon_CP_1451_elements(12);
        preds(1)  <= ReceiveEngineDaemon_CP_1451_elements(13);
        entry_tmerge_1548 : transition_merge -- 
          generic map(name => " entry_tmerge_1548")
          port map (preds => preds, symbol_out => ReceiveEngineDaemon_CP_1451_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_887_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_942_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_915_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_943_wire : std_logic_vector(0 downto 0);
    signal RPIPE_CONTROL_REGISTER_885_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_940_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_896_wire : std_logic_vector(35 downto 0);
    signal RPIPE_FREE_Q_933_wire : std_logic_vector(35 downto 0);
    signal bad_packet_identifier_911 : std_logic_vector(0 downto 0);
    signal free_flag_922 : std_logic_vector(0 downto 0);
    signal konst_879_wire_constant : std_logic_vector(5 downto 0);
    signal konst_886_wire_constant : std_logic_vector(31 downto 0);
    signal konst_941_wire_constant : std_logic_vector(31 downto 0);
    signal ok_flag_917 : std_logic_vector(0 downto 0);
    signal push_status_937 : std_logic_vector(0 downto 0);
    signal rx_buffer_pointer_32_899 : std_logic_vector(31 downto 0);
    signal rx_buffer_pointer_36_905 : std_logic_vector(35 downto 0);
    signal slice_935_wire : std_logic_vector(31 downto 0);
    signal status_899 : std_logic_vector(0 downto 0);
    signal type_cast_895_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_903_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_932_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_879_wire_constant <= "000000";
    konst_886_wire_constant <= "00000000000000000000000000000000";
    konst_941_wire_constant <= "00000000000000000000000000000000";
    type_cast_895_wire_constant <= "1";
    type_cast_903_wire_constant <= "0000";
    type_cast_932_wire_constant <= "1";
    -- logger for split-operator slice_935_inst flow-through 
    process(slice_935_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:slice_935_inst:flowthrough inputs: " & " free_flag_922 (guard)= " & Convert_SLV_To_String(free_flag_922) & " rx_buffer_pointer_36_905 = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_36_905) & " outputs:" & " slice_935_wire= "  & Convert_SLV_To_Hex_String(slice_935_wire));
      --
    end process; 
    -- flow-through slice operator slice_935_inst
    slice_935_wire <= rx_buffer_pointer_36_905(35 downto 4);
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_891_branch_req_0," req0 do_while_stmt_891_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_891_branch_ack_0," ack0 do_while_stmt_891_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_891_branch_ack_1," ack1 do_while_stmt_891_branch");
    do_while_stmt_891_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_943_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_891_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_891_branch_req_0,
          ack0 => do_while_stmt_891_branch_ack_0,
          ack1 => do_while_stmt_891_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_884_branch_req_0," req0 if_stmt_884_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_884_branch_ack_0," ack0 if_stmt_884_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_884_branch_ack_1," ack1 if_stmt_884_branch");
    if_stmt_884_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_887_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_884_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_884_branch_req_0,
          ack0 => if_stmt_884_branch_ack_0,
          ack1 => if_stmt_884_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator AND_u1_u1_916_inst flow-through 
    process(ok_flag_917) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:AND_u1_u1_916_inst:flowthrough inputs: " & " status_899 = "& Convert_SLV_To_Hex_String(status_899) & " NOT_u1_u1_915_wire = "& Convert_SLV_To_Hex_String(NOT_u1_u1_915_wire) & " outputs:" & " ok_flag_917= "  & Convert_SLV_To_Hex_String(ok_flag_917));
      --
    end process; 
    -- binary operator AND_u1_u1_916_inst
    process(status_899, NOT_u1_u1_915_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(status_899, NOT_u1_u1_915_wire, tmp_var);
      ok_flag_917 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_921_inst flow-through 
    process(free_flag_922) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:AND_u1_u1_921_inst:flowthrough inputs: " & " status_899 = "& Convert_SLV_To_Hex_String(status_899) & " bad_packet_identifier_911 = "& Convert_SLV_To_Hex_String(bad_packet_identifier_911) & " outputs:" & " free_flag_922= "  & Convert_SLV_To_Hex_String(free_flag_922));
      --
    end process; 
    -- binary operator AND_u1_u1_921_inst
    process(status_899, bad_packet_identifier_911) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(status_899, bad_packet_identifier_911, tmp_var);
      free_flag_922 <= tmp_var; --
    end process;
    -- logger for split-operator BITSEL_u32_u1_887_inst flow-through 
    process(BITSEL_u32_u1_887_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:BITSEL_u32_u1_887_inst:flowthrough inputs: " & " RPIPE_CONTROL_REGISTER_885_wire = "& Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_885_wire) & " konst_886_wire_constant = "& Convert_SLV_To_Hex_String(konst_886_wire_constant) & " outputs:" & " BITSEL_u32_u1_887_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u32_u1_887_wire));
      --
    end process; 
    -- binary operator BITSEL_u32_u1_887_inst
    process(RPIPE_CONTROL_REGISTER_885_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_885_wire, konst_886_wire_constant, tmp_var);
      BITSEL_u32_u1_887_wire <= tmp_var; --
    end process;
    -- logger for split-operator BITSEL_u32_u1_942_inst flow-through 
    process(BITSEL_u32_u1_942_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:BITSEL_u32_u1_942_inst:flowthrough inputs: " & " RPIPE_CONTROL_REGISTER_940_wire = "& Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_940_wire) & " konst_941_wire_constant = "& Convert_SLV_To_Hex_String(konst_941_wire_constant) & " outputs:" & " BITSEL_u32_u1_942_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u32_u1_942_wire));
      --
    end process; 
    -- binary operator BITSEL_u32_u1_942_inst
    process(RPIPE_CONTROL_REGISTER_940_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_940_wire, konst_941_wire_constant, tmp_var);
      BITSEL_u32_u1_942_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u36_904_inst flow-through 
    process(rx_buffer_pointer_36_905) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:CONCAT_u32_u36_904_inst:flowthrough inputs: " & " rx_buffer_pointer_32_899 = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_32_899) & " type_cast_903_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_903_wire_constant) & " outputs:" & " rx_buffer_pointer_36_905= "  & Convert_SLV_To_Hex_String(rx_buffer_pointer_36_905));
      --
    end process; 
    -- binary operator CONCAT_u32_u36_904_inst
    process(rx_buffer_pointer_32_899) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(rx_buffer_pointer_32_899, type_cast_903_wire_constant, tmp_var);
      rx_buffer_pointer_36_905 <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_915_inst flow-through 
    process(NOT_u1_u1_915_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:NOT_u1_u1_915_inst:flowthrough inputs: " & " bad_packet_identifier_911 = "& Convert_SLV_To_Hex_String(bad_packet_identifier_911) & " outputs:" & " NOT_u1_u1_915_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_915_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_915_inst
    process(bad_packet_identifier_911) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", bad_packet_identifier_911, tmp_var);
      NOT_u1_u1_915_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator NOT_u1_u1_943_inst flow-through 
    process(NOT_u1_u1_943_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:NOT_u1_u1_943_inst:flowthrough inputs: " & " BITSEL_u32_u1_942_wire = "& Convert_SLV_To_Hex_String(BITSEL_u32_u1_942_wire) & " outputs:" & " NOT_u1_u1_943_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_943_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_943_inst
    process(BITSEL_u32_u1_942_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_942_wire, tmp_var);
      NOT_u1_u1_943_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator RPIPE_CONTROL_REGISTER_885_inst flow-through 
    process(RPIPE_CONTROL_REGISTER_885_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:RPIPE_CONTROL_REGISTER_885_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_CONTROL_REGISTER_885_wire= "  & Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_885_wire));
      --
    end process; 
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_885_wire <= CONTROL_REGISTER;
    -- logger for split-operator RPIPE_CONTROL_REGISTER_940_inst flow-through 
    process(RPIPE_CONTROL_REGISTER_940_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:RPIPE_CONTROL_REGISTER_940_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_CONTROL_REGISTER_940_wire= "  & Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_940_wire));
      --
    end process; 
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_940_wire <= CONTROL_REGISTER;
    -- logger for split-operator RPIPE_FREE_Q_896_inst flow-through 
    process(RPIPE_FREE_Q_896_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:RPIPE_FREE_Q_896_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_FREE_Q_896_wire= "  & Convert_SLV_To_Hex_String(RPIPE_FREE_Q_896_wire));
      --
    end process; 
    -- logger for split-operator RPIPE_FREE_Q_933_inst flow-through 
    process(RPIPE_FREE_Q_933_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:RPIPE_FREE_Q_933_inst:flowthrough inputs: " & " free_flag_922 (guard)= " & Convert_SLV_To_String(free_flag_922) & " outputs:" & " RPIPE_FREE_Q_933_wire= "  & Convert_SLV_To_Hex_String(RPIPE_FREE_Q_933_wire));
      --
    end process; 
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_896_wire <= FREE_Q;
    RPIPE_FREE_Q_933_wire <= FREE_Q;
    -- logger for split-operator WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst:started:   PipeWrite to LAST_WRITTEN_RX_QUEUE_INDEX inputs: " & " konst_879_wire_constant = "& Convert_SLV_To_Hex_String(konst_879_wire_constant));
          --
        end if; 
        if WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_878_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_879_wire_constant;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_899_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_899_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_899_call:started:  Call to module popFromQueue inputs: " & " type_cast_895_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_895_wire_constant) & " RPIPE_FREE_Q_896_wire = "& Convert_SLV_To_Hex_String(RPIPE_FREE_Q_896_wire));
          --
        end if; 
        if call_stmt_899_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_899_call:finished:  outputs: " & " rx_buffer_pointer_32_899= "  & Convert_SLV_To_Hex_String(rx_buffer_pointer_32_899) & " status_899= "  & Convert_SLV_To_Hex_String(status_899));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_899_call 
    popFromQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_899_call_req_0;
      call_stmt_899_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_899_call_req_1;
      call_stmt_899_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_0_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_895_wire_constant & RPIPE_FREE_Q_896_wire;
      rx_buffer_pointer_32_899 <= data_out(32 downto 1);
      status_899 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_911_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_911_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_911_call:started:  Call to module loadBuffer inputs: " & " status_899 (guard)= " & Convert_SLV_To_String(status_899) & " rx_buffer_pointer_36_905 = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_36_905));
          --
        end if; 
        if call_stmt_911_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_911_call:finished:  outputs: " & " bad_packet_identifier_911= "  & Convert_SLV_To_Hex_String(bad_packet_identifier_911));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_911_call 
    loadBuffer_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_911_call_req_0;
      call_stmt_911_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_911_call_req_1;
      call_stmt_911_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= status_899(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadBuffer_call_group_1_gI: SplitGuardInterface generic map(name => "loadBuffer_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_905;
      bad_packet_identifier_911 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadBuffer_call_reqs(0),
          ackR => loadBuffer_call_acks(0),
          dataR => loadBuffer_call_data(35 downto 0),
          tagR => loadBuffer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => loadBuffer_return_acks(0), -- cross-over
          ackL => loadBuffer_return_reqs(0), -- cross-over
          dataL => loadBuffer_return_data(0 downto 0),
          tagL => loadBuffer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_927_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_927_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_927_call:started:  Call to module populateRxQueue inputs: " & " ok_flag_917 (guard)= " & Convert_SLV_To_String(ok_flag_917) & " rx_buffer_pointer_36_905 = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_36_905));
          --
        end if; 
        if call_stmt_927_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_927_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_927_call 
    populateRxQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_927_call_req_0;
      call_stmt_927_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_927_call_req_1;
      call_stmt_927_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_917(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      populateRxQueue_call_group_2_gI: SplitGuardInterface generic map(name => "populateRxQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_905;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => populateRxQueue_call_reqs(0),
          ackR => populateRxQueue_call_acks(0),
          dataR => populateRxQueue_call_data(35 downto 0),
          tagR => populateRxQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => populateRxQueue_return_acks(0), -- cross-over
          ackL => populateRxQueue_return_reqs(0), -- cross-over
          tagL => populateRxQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- logger for split-operator call_stmt_937_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_937_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_937_call:started:  Call to module pushIntoQueue inputs: " & " free_flag_922 (guard)= " & Convert_SLV_To_String(free_flag_922) & " type_cast_932_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_932_wire_constant) & " RPIPE_FREE_Q_933_wire = "& Convert_SLV_To_Hex_String(RPIPE_FREE_Q_933_wire) & " slice_935_wire = "& Convert_SLV_To_Hex_String(slice_935_wire));
          --
        end if; 
        if call_stmt_937_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:ReceiveEngineDaemon:DP:call_stmt_937_call:finished:  outputs: " & " push_status_937= "  & Convert_SLV_To_Hex_String(push_status_937));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (3) : call_stmt_937_call 
    pushIntoQueue_call_group_3: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_937_call_req_0;
      call_stmt_937_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_937_call_req_1;
      call_stmt_937_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= free_flag_922(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_3_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_932_wire_constant & RPIPE_FREE_Q_933_wire & slice_935_wire;
      push_status_937 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end ReceiveEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity SoftwareRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
    CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
    AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
    NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity SoftwareRegisterAccessDaemon;
architecture SoftwareRegisterAccessDaemon_arch of SoftwareRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal SoftwareRegisterAccessDaemon_CP_1633_start: Boolean;
  signal SoftwareRegisterAccessDaemon_CP_1633_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal check_num_server_1076_972_buf_ack_0 : boolean;
  signal array_obj_ref_1007_load_0_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1101_inst_req_1 : boolean;
  signal array_obj_ref_1007_load_0_req_0 : boolean;
  signal check_num_server_1076_972_buf_req_1 : boolean;
  signal type_cast_1015_inst_ack_1 : boolean;
  signal type_cast_1015_inst_req_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1023_inst_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_1 : boolean;
  signal check_num_server_1076_972_buf_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1023_inst_req_1 : boolean;
  signal do_while_stmt_950_branch_ack_0 : boolean;
  signal type_cast_1015_inst_ack_0 : boolean;
  signal WPIPE_FREE_Q_1010_inst_ack_1 : boolean;
  signal type_cast_1015_inst_req_0 : boolean;
  signal WPIPE_FREE_Q_1010_inst_req_1 : boolean;
  signal array_obj_ref_1007_load_0_req_1 : boolean;
  signal check_num_server_1076_972_buf_ack_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1018_inst_req_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1018_inst_req_1 : boolean;
  signal do_while_stmt_950_branch_ack_1 : boolean;
  signal array_obj_ref_1007_load_0_ack_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_1 : boolean;
  signal array_obj_ref_1079_load_0_req_1 : boolean;
  signal array_obj_ref_1002_load_0_req_0 : boolean;
  signal array_obj_ref_1079_load_0_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_0 : boolean;
  signal array_obj_ref_1079_load_0_ack_0 : boolean;
  signal array_obj_ref_1079_load_0_req_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_1101_inst_req_0 : boolean;
  signal array_obj_ref_1020_load_0_ack_1 : boolean;
  signal array_obj_ref_1020_load_0_req_1 : boolean;
  signal do_while_stmt_950_branch_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1023_inst_ack_0 : boolean;
  signal phi_stmt_952_req_1 : boolean;
  signal phi_stmt_952_req_0 : boolean;
  signal phi_stmt_952_ack_0 : boolean;
  signal array_obj_ref_1020_load_0_ack_0 : boolean;
  signal array_obj_ref_1020_load_0_req_0 : boolean;
  signal call_stmt_1087_call_ack_1 : boolean;
  signal call_stmt_1087_call_req_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1000_inst_ack_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1000_inst_req_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1000_inst_ack_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1000_inst_req_0 : boolean;
  signal phi_stmt_958_req_1 : boolean;
  signal call_stmt_1087_call_ack_0 : boolean;
  signal phi_stmt_958_req_0 : boolean;
  signal call_stmt_1087_call_req_0 : boolean;
  signal phi_stmt_958_ack_0 : boolean;
  signal array_obj_ref_1002_load_0_ack_1 : boolean;
  signal array_obj_ref_1002_load_0_req_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1023_inst_req_0 : boolean;
  signal check_control_regsiter_1058_962_buf_req_0 : boolean;
  signal WPIPE_FREE_Q_1010_inst_ack_0 : boolean;
  signal check_control_regsiter_1058_962_buf_ack_0 : boolean;
  signal check_control_regsiter_1058_962_buf_req_1 : boolean;
  signal WPIPE_FREE_Q_1010_inst_req_0 : boolean;
  signal check_control_regsiter_1058_962_buf_ack_1 : boolean;
  signal array_obj_ref_1002_load_0_ack_0 : boolean;
  signal phi_stmt_963_req_1 : boolean;
  signal phi_stmt_963_req_0 : boolean;
  signal phi_stmt_963_ack_0 : boolean;
  signal check_free_q_1067_967_buf_req_0 : boolean;
  signal check_free_q_1067_967_buf_ack_0 : boolean;
  signal check_free_q_1067_967_buf_req_1 : boolean;
  signal check_free_q_1067_967_buf_ack_1 : boolean;
  signal phi_stmt_968_req_1 : boolean;
  signal phi_stmt_968_req_0 : boolean;
  signal phi_stmt_968_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  SoftwareRegisterAccessDaemon_CP_1633_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1633_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1633_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_1633_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,SoftwareRegisterAccessDaemon_CP_1633_start,"SoftwareRegisterAccessDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,SoftwareRegisterAccessDaemon_CP_1633_symbol, "SoftwareRegisterAccessDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  SoftwareRegisterAccessDaemon_CP_1633: Block -- control-path 
    signal SoftwareRegisterAccessDaemon_CP_1633_elements: BooleanArray(137 downto 0);
    -- 
  begin -- 
    SoftwareRegisterAccessDaemon_CP_1633_elements(0) <= SoftwareRegisterAccessDaemon_CP_1633_start;
    SoftwareRegisterAccessDaemon_CP_1633_symbol <= SoftwareRegisterAccessDaemon_CP_1633_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_949/$entry
      -- CP-element group 0: 	 branch_block_stmt_949/branch_block_stmt_949__entry__
      -- CP-element group 0: 	 branch_block_stmt_949/do_while_stmt_950__entry__
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	137 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_949/$exit
      -- CP-element group 1: 	 branch_block_stmt_949/branch_block_stmt_949__exit__
      -- CP-element group 1: 	 branch_block_stmt_949/do_while_stmt_950__exit__
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(1) <= SoftwareRegisterAccessDaemon_CP_1633_elements(137);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_949/do_while_stmt_950/$entry
      -- CP-element group 2: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950__entry__
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(2) <= SoftwareRegisterAccessDaemon_CP_1633_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	137 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950__exit__
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_949/do_while_stmt_950/loop_back
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	135 
    -- CP-element group 5: 	136 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_949/do_while_stmt_950/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_949/do_while_stmt_950/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_949/do_while_stmt_950/condition_done
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(5) <= SoftwareRegisterAccessDaemon_CP_1633_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	134 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_949/do_while_stmt_950/loop_body_done
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(6) <= SoftwareRegisterAccessDaemon_CP_1633_elements(134);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(7) <= SoftwareRegisterAccessDaemon_CP_1633_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	78 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	59 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(8) <= SoftwareRegisterAccessDaemon_CP_1633_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	71 
    -- CP-element group 9: 	114 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	89 
    -- CP-element group 9: 	107 
    -- CP-element group 9: 	96 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	52 
    -- CP-element group 9:  members (8) 
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_root_address_calculated
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	129 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/condition_evaluated
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:do_while_stmt_950_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_1657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(10), ack => do_while_stmt_950_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(14) & SoftwareRegisterAccessDaemon_CP_1633_elements(129);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	70 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_sample_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(15) & SoftwareRegisterAccessDaemon_CP_1633_elements(70) & SoftwareRegisterAccessDaemon_CP_1633_elements(32) & SoftwareRegisterAccessDaemon_CP_1633_elements(51) & SoftwareRegisterAccessDaemon_CP_1633_elements(14);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	54 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	134 
    -- CP-element group 12: 	115 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	70 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(17) & SoftwareRegisterAccessDaemon_CP_1633_elements(73) & SoftwareRegisterAccessDaemon_CP_1633_elements(35) & SoftwareRegisterAccessDaemon_CP_1633_elements(54);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	71 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	74 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_update_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(16) & SoftwareRegisterAccessDaemon_CP_1633_elements(71) & SoftwareRegisterAccessDaemon_CP_1633_elements(33) & SoftwareRegisterAccessDaemon_CP_1633_elements(52);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(75) & SoftwareRegisterAccessDaemon_CP_1633_elements(37) & SoftwareRegisterAccessDaemon_CP_1633_elements(56);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(12);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	112 
    -- CP-element group 16: 	91 
    -- CP-element group 16: 	105 
    -- CP-element group 16: 	109 
    -- CP-element group 16: 	102 
    -- CP-element group 16: 	94 
    -- CP-element group 16: 	98 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(112) & SoftwareRegisterAccessDaemon_CP_1633_elements(91) & SoftwareRegisterAccessDaemon_CP_1633_elements(105) & SoftwareRegisterAccessDaemon_CP_1633_elements(109) & SoftwareRegisterAccessDaemon_CP_1633_elements(102) & SoftwareRegisterAccessDaemon_CP_1633_elements(94) & SoftwareRegisterAccessDaemon_CP_1633_elements(98);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_sample_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	111 
    -- CP-element group 18: 	89 
    -- CP-element group 18: 	107 
    -- CP-element group 18: 	100 
    -- CP-element group 18: 	104 
    -- CP-element group 18: 	93 
    -- CP-element group 18: 	96 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_loopback_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(19) <= SoftwareRegisterAccessDaemon_CP_1633_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_loopback_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_952_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_952_loopback_sample_req_1672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_952_loopback_sample_req_1672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(20), ack => phi_stmt_952_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_entry_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(21) <= SoftwareRegisterAccessDaemon_CP_1633_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_entry_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_952_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_952_entry_sample_req_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_952_entry_sample_req_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(22), ack => phi_stmt_952_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_952_phi_mux_ack_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_952_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_952_phi_mux_ack_1678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_952_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(26) <= SoftwareRegisterAccessDaemon_CP_1633_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_955_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(25), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(30) <= SoftwareRegisterAccessDaemon_CP_1633_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_957_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(29), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: 	117 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(12) & SoftwareRegisterAccessDaemon_CP_1633_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	91 
    -- CP-element group 33: 	94 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(33) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(91) & SoftwareRegisterAccessDaemon_CP_1633_elements(94);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_sample_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(34) <= SoftwareRegisterAccessDaemon_CP_1633_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_sample_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_update_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(36) <= SoftwareRegisterAccessDaemon_CP_1633_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	89 
    -- CP-element group 37: 	93 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_loopback_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(38) <= SoftwareRegisterAccessDaemon_CP_1633_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_loopback_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_958_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_958_loopback_sample_req_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_958_loopback_sample_req_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(39), ack => phi_stmt_958_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_entry_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(40) <= SoftwareRegisterAccessDaemon_CP_1633_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_entry_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_958_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_958_entry_sample_req_1709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_958_entry_sample_req_1709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(41), ack => phi_stmt_958_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_958_phi_mux_ack_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_958_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_958_phi_mux_ack_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_958_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(43) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(45) <= SoftwareRegisterAccessDaemon_CP_1633_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_961_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(44), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Sample/req
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_control_regsiter_1058_962_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(47), ack => check_control_regsiter_1058_962_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_update_start_
      -- CP-element group 48: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Update/req
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_control_regsiter_1058_962_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(48), ack => check_control_regsiter_1058_962_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Sample/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_control_regsiter_1058_962_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1058_962_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_control_regsiter_962_Update/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_control_regsiter_1058_962_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1058_962_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: 	117 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(12) & SoftwareRegisterAccessDaemon_CP_1633_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	105 
    -- CP-element group 52: 	102 
    -- CP-element group 52: 	98 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(52) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(105) & SoftwareRegisterAccessDaemon_CP_1633_elements(102) & SoftwareRegisterAccessDaemon_CP_1633_elements(98);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_sample_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(53) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(53) <= SoftwareRegisterAccessDaemon_CP_1633_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_sample_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(54) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_update_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(55) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(55) <= SoftwareRegisterAccessDaemon_CP_1633_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: 	100 
    -- CP-element group 56: 	104 
    -- CP-element group 56: 	96 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(56) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_loopback_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(57) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(57) <= SoftwareRegisterAccessDaemon_CP_1633_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_loopback_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_963_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_963_loopback_sample_req_1750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_963_loopback_sample_req_1750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(58), ack => phi_stmt_963_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_entry_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(59) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(59) <= SoftwareRegisterAccessDaemon_CP_1633_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_entry_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_963_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_963_entry_sample_req_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_963_entry_sample_req_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(60), ack => phi_stmt_963_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_963_phi_mux_ack_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_963_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_963_phi_mux_ack_1756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_963_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(62) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(63) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(64) <= SoftwareRegisterAccessDaemon_CP_1633_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_966_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(65) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(63), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Sample/req
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_free_q_1067_967_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(66), ack => check_free_q_1067_967_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_update_start_
      -- CP-element group 67: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Update/req
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_free_q_1067_967_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(67), ack => check_free_q_1067_967_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Sample/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_free_q_1067_967_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1067_967_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_free_q_967_Update/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_free_q_1067_967_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_1067_967_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: 	117 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(12) & SoftwareRegisterAccessDaemon_CP_1633_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	112 
    -- CP-element group 71: 	109 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(71) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(112) & SoftwareRegisterAccessDaemon_CP_1633_elements(109);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_sample_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(72) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(72) <= SoftwareRegisterAccessDaemon_CP_1633_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_sample_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(73) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_update_start__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(74) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(74) <= SoftwareRegisterAccessDaemon_CP_1633_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	111 
    -- CP-element group 75: 	107 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(75) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_loopback_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(76) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(76) <= SoftwareRegisterAccessDaemon_CP_1633_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_loopback_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(77) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_968_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_968_loopback_sample_req_1794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_968_loopback_sample_req_1794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(77), ack => phi_stmt_968_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_entry_trigger
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(78)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(78)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(78) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(78) <= SoftwareRegisterAccessDaemon_CP_1633_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_entry_sample_req_ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(79)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(79)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(79) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_968_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_968_entry_sample_req_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_968_entry_sample_req_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(79), ack => phi_stmt_968_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_phi_mux_ack_ps
      -- CP-element group 80: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/phi_stmt_968_phi_mux_ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(80)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(80)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(80) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:phi_stmt_968_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_968_phi_mux_ack_1800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_968_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_sample_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(81)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(81)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(81) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(82)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(82)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(82) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(83)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(83)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(83) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(83) <= SoftwareRegisterAccessDaemon_CP_1633_elements(84);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	83 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_971_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(84)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(84)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(84) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(82), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(85)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(85)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(85) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_num_server_1076_972_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(85), ack => check_num_server_1076_972_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Update/req
      -- CP-element group 86: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(86)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(86)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(86) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_num_server_1076_972_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(86), ack => check_num_server_1076_972_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(87)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(87)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(87) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_num_server_1076_972_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1076_972_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/R_check_num_server_972_update_completed__ps
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(88)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(88)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(88) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:check_num_server_1076_972_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_1076_972_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	9 
    -- CP-element group 89: 	18 
    -- CP-element group 89: 	37 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	125 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/word_access_start/word_0/$entry
      -- CP-element group 89: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/word_access_start/$entry
      -- CP-element group 89: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/word_access_start/word_0/rr
      -- CP-element group 89: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/$entry
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(89)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(89)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(89) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1002_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(89), ack => array_obj_ref_1002_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(37) & SoftwareRegisterAccessDaemon_CP_1633_elements(125) & SoftwareRegisterAccessDaemon_CP_1633_elements(91);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	94 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_update_start_
      -- CP-element group 90: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/word_access_complete/word_0/cr
      -- CP-element group 90: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/word_access_complete/word_0/$entry
      -- CP-element group 90: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/word_access_complete/$entry
      -- CP-element group 90: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/$entry
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(90)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(90)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(90) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1002_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(90), ack => array_obj_ref_1002_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1633_elements(94);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	130 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	16 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	33 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/word_access_start/$exit
      -- CP-element group 91: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/word_access_start/word_0/$exit
      -- CP-element group 91: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(91)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(91)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(91) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1002_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1002_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/array_obj_ref_1002_Merge/merge_ack
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/array_obj_ref_1002_Merge/merge_req
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/array_obj_ref_1002_Merge/$exit
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/array_obj_ref_1002_Merge/$entry
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/word_access_complete/word_0/ca
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/word_access_complete/word_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/word_access_complete/$exit
      -- CP-element group 92: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_Update/$exit
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(92)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(92)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(92) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1002_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1002_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	18 
    -- CP-element group 93: 	92 
    -- CP-element group 93: 	37 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Sample/req
      -- CP-element group 93: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(93)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(93)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(93) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_CONTROL_REGISTER_1000_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(93), ack => WPIPE_CONTROL_REGISTER_1000_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(92) & SoftwareRegisterAccessDaemon_CP_1633_elements(37) & SoftwareRegisterAccessDaemon_CP_1633_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	16 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	33 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Update/req
      -- CP-element group 94: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Sample/ack
      -- CP-element group 94: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_update_start_
      -- CP-element group 94: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(94)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(94)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(94) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_CONTROL_REGISTER_1000_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_CONTROL_REGISTER_1000_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1000_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(94)); -- 
    req_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(94), ack => WPIPE_CONTROL_REGISTER_1000_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	134 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Update/ack
      -- CP-element group 95: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_CONTROL_REGISTER_1000_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(95)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(95)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(95) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_CONTROL_REGISTER_1000_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1000_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	9 
    -- CP-element group 96: 	18 
    -- CP-element group 96: 	56 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	125 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/word_access_start/word_0/rr
      -- CP-element group 96: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/word_access_start/$entry
      -- CP-element group 96: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/word_access_start/word_0/$entry
      -- CP-element group 96: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(96)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(96)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(96) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1007_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(96), ack => array_obj_ref_1007_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(56) & SoftwareRegisterAccessDaemon_CP_1633_elements(125) & SoftwareRegisterAccessDaemon_CP_1633_elements(98);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	102 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/word_access_complete/word_0/$entry
      -- CP-element group 97: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/word_access_complete/word_0/cr
      -- CP-element group 97: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/word_access_complete/$entry
      -- CP-element group 97: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(97)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(97)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(97) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1007_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(97), ack => array_obj_ref_1007_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1633_elements(102);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	131 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	16 
    -- CP-element group 98: 	96 
    -- CP-element group 98: 	52 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/word_access_start/word_0/ra
      -- CP-element group 98: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/word_access_start/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/word_access_start/$exit
      -- CP-element group 98: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(98)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(98)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(98) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1007_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1007_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/word_access_complete/$exit
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/word_access_complete/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/word_access_complete/word_0/ca
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/array_obj_ref_1007_Merge/$entry
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/array_obj_ref_1007_Merge/$exit
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/array_obj_ref_1007_Merge/merge_req
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_Update/array_obj_ref_1007_Merge/merge_ack
      -- CP-element group 99: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(99)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(99)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(99) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1007_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1007_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	18 
    -- CP-element group 100: 	99 
    -- CP-element group 100: 	56 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(100)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(100)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(100) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:type_cast_1015_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(100), ack => type_cast_1015_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(99) & SoftwareRegisterAccessDaemon_CP_1633_elements(56) & SoftwareRegisterAccessDaemon_CP_1633_elements(102);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	105 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Update/cr
      -- CP-element group 101: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(101)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(101)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(101) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:type_cast_1015_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(101), ack => type_cast_1015_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1633_elements(105);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	16 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	97 
    -- CP-element group 102: 	52 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(102)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(102)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(102) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:type_cast_1015_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/type_cast_1015_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(103)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(103)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(103) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:type_cast_1015_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	18 
    -- CP-element group 104: 	103 
    -- CP-element group 104: 	56 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Sample/req
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(104)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(104)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(104) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_FREE_Q_1010_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(104), ack => WPIPE_FREE_Q_1010_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(103) & SoftwareRegisterAccessDaemon_CP_1633_elements(56) & SoftwareRegisterAccessDaemon_CP_1633_elements(106);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: marked-successors 
    -- CP-element group 105: 	16 
    -- CP-element group 105: 	101 
    -- CP-element group 105: 	52 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_update_start_
      -- CP-element group 105: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Update/req
      -- CP-element group 105: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Sample/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(105)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(105)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(105) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_FREE_Q_1010_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_FREE_Q_1010_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1010_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(105)); -- 
    req_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(105), ack => WPIPE_FREE_Q_1010_inst_req_1); -- 
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	134 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Update/ack
      -- CP-element group 106: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_FREE_Q_1010_Update/$exit
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(106)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(106)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(106) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_FREE_Q_1010_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1010_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	9 
    -- CP-element group 107: 	18 
    -- CP-element group 107: 	75 
    -- CP-element group 107: marked-predecessors 
    -- CP-element group 107: 	125 
    -- CP-element group 107: 	109 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/word_access_start/word_0/rr
      -- CP-element group 107: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/word_access_start/word_0/$entry
      -- CP-element group 107: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/word_access_start/$entry
      -- CP-element group 107: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/$entry
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(107)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(107)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(107) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1020_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(107), ack => array_obj_ref_1020_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(75) & SoftwareRegisterAccessDaemon_CP_1633_elements(125) & SoftwareRegisterAccessDaemon_CP_1633_elements(109);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	112 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_update_start_
      -- CP-element group 108: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/word_access_complete/word_0/cr
      -- CP-element group 108: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/word_access_complete/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/word_access_complete/$entry
      -- CP-element group 108: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/$entry
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(108)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(108)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(108) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1020_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(108), ack => array_obj_ref_1020_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1633_elements(112);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	132 
    -- CP-element group 109: marked-successors 
    -- CP-element group 109: 	16 
    -- CP-element group 109: 	71 
    -- CP-element group 109: 	107 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/word_access_start/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/word_access_start/$exit
      -- CP-element group 109: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Sample/$exit
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(109)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(109)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(109) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1020_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1020_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/array_obj_ref_1020_Merge/merge_ack
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/array_obj_ref_1020_Merge/merge_req
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/array_obj_ref_1020_Merge/$exit
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/array_obj_ref_1020_Merge/$entry
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_Update/$exit
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(110)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(110)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(110) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1020_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1020_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	18 
    -- CP-element group 111: 	110 
    -- CP-element group 111: 	75 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Sample/req
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(111)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(111)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(111) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_NUMBER_OF_SERVERS_1018_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(111), ack => WPIPE_NUMBER_OF_SERVERS_1018_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(18) & SoftwareRegisterAccessDaemon_CP_1633_elements(110) & SoftwareRegisterAccessDaemon_CP_1633_elements(75) & SoftwareRegisterAccessDaemon_CP_1633_elements(113);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	16 
    -- CP-element group 112: 	71 
    -- CP-element group 112: 	108 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Sample/ack
      -- CP-element group 112: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_update_start_
      -- CP-element group 112: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Update/req
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(112)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(112)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(112) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_NUMBER_OF_SERVERS_1018_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(112)); -- 
    req_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(112), ack => WPIPE_NUMBER_OF_SERVERS_1018_inst_req_1); -- 
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	134 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_NUMBER_OF_SERVERS_1018_Update/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(113)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(113)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(113) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	9 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	117 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(114)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(114)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(114) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:RPIPE_AFB_NIC_REQUEST_1023_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(114), ack => RPIPE_AFB_NIC_REQUEST_1023_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(9) & SoftwareRegisterAccessDaemon_CP_1633_elements(117);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	12 
    -- CP-element group 115: 	116 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	127 
    -- CP-element group 115: 	124 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(115)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(115)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(115) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:RPIPE_AFB_NIC_REQUEST_1023_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(115), ack => RPIPE_AFB_NIC_REQUEST_1023_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(12) & SoftwareRegisterAccessDaemon_CP_1633_elements(116) & SoftwareRegisterAccessDaemon_CP_1633_elements(127) & SoftwareRegisterAccessDaemon_CP_1633_elements(124);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	115 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(116)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(116)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(116) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:RPIPE_AFB_NIC_REQUEST_1023_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1023_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(116)); -- 
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	126 
    -- CP-element group 117: 	118 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	114 
    -- CP-element group 117: 	70 
    -- CP-element group 117: 	32 
    -- CP-element group 117: 	51 
    -- CP-element group 117:  members (29) 
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_scale_0/$entry
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_resize_0/index_resize_ack
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_scale_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_scale_0/scale_rename_req
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_resize_0/index_resize_req
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_resize_0/$exit
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_resize_0/$entry
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_computed_0
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_scaled_0
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_word_addrgen/root_register_ack
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_word_addrgen/root_register_req
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_word_addrgen/$exit
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_word_addrgen/$entry
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_base_plus_offset/sum_rename_ack
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_base_plus_offset/sum_rename_req
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_base_plus_offset/$exit
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_base_plus_offset/$entry
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_resized_0
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_final_index_sum_regn/ack
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_final_index_sum_regn/req
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_final_index_sum_regn/$exit
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_final_index_sum_regn/$entry
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_index_scale_0/scale_rename_ack
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_offset_calculated
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_root_address_calculated
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_word_address_calculated
      -- CP-element group 117: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/RPIPE_AFB_NIC_REQUEST_1023_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(117)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(117)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(117) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:RPIPE_AFB_NIC_REQUEST_1023_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1023_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: 	125 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/word_access_start/word_0/rr
      -- CP-element group 118: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/word_access_start/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/word_access_start/$entry
      -- CP-element group 118: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/$entry
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(118)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(118)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(118) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1079_load_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(118), ack => array_obj_ref_1079_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(117) & SoftwareRegisterAccessDaemon_CP_1633_elements(120) & SoftwareRegisterAccessDaemon_CP_1633_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	127 
    -- CP-element group 119: 	124 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/word_access_complete/word_0/$entry
      -- CP-element group 119: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/word_access_complete/$entry
      -- CP-element group 119: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/word_access_complete/word_0/cr
      -- CP-element group 119: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(119)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(119)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(119) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1079_load_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(119), ack => array_obj_ref_1079_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(127) & SoftwareRegisterAccessDaemon_CP_1633_elements(124);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	133 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/word_access_start/word_0/ra
      -- CP-element group 120: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/word_access_start/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/word_access_start/$exit
      -- CP-element group 120: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(120)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(120)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(120) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1079_load_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(120)); -- 
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	126 
    -- CP-element group 121:  members (9) 
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/array_obj_ref_1079_Merge/merge_req
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/word_access_complete/$exit
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/array_obj_ref_1079_Merge/merge_ack
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/word_access_complete/word_0/$exit
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/word_access_complete/word_0/ca
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/array_obj_ref_1079_Merge/$entry
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_Update/array_obj_ref_1079_Merge/$exit
      -- CP-element group 121: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(121)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(121)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(121) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:array_obj_ref_1079_load_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	130 
    -- CP-element group 122: 	131 
    -- CP-element group 122: 	132 
    -- CP-element group 122: 	133 
    -- CP-element group 122: 	121 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Sample/crr
      -- CP-element group 122: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Sample/$entry
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(122)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(122)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(122) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:call_stmt_1087_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_2071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(122), ack => call_stmt_1087_call_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(130) & SoftwareRegisterAccessDaemon_CP_1633_elements(131) & SoftwareRegisterAccessDaemon_CP_1633_elements(132) & SoftwareRegisterAccessDaemon_CP_1633_elements(133) & SoftwareRegisterAccessDaemon_CP_1633_elements(121) & SoftwareRegisterAccessDaemon_CP_1633_elements(124);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Update/ccr
      -- CP-element group 123: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_update_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(123)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(123)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(123) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:call_stmt_1087_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_2076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(123), ack => call_stmt_1087_call_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_1633_elements(125);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: 	115 
    -- CP-element group 124: 	119 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Sample/cra
      -- CP-element group 124: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(124)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(124)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(124) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:call_stmt_1087_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1087_call_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	134 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	118 
    -- CP-element group 125: 	89 
    -- CP-element group 125: 	107 
    -- CP-element group 125: 	96 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/ring_reenable_memory_space_0
      -- CP-element group 125: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Update/cca
      -- CP-element group 125: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/call_stmt_1087_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(125)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(125)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(125) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:call_stmt_1087_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1087_call_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	121 
    -- CP-element group 126: 	117 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	128 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Sample/req
      -- CP-element group 126: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_sample_start_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(126)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(126)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(126) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_AFB_NIC_RESPONSE_1101_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(126), ack => WPIPE_AFB_NIC_RESPONSE_1101_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(121) & SoftwareRegisterAccessDaemon_CP_1633_elements(117) & SoftwareRegisterAccessDaemon_CP_1633_elements(128);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	115 
    -- CP-element group 127: 	119 
    -- CP-element group 127:  members (6) 
      -- CP-element group 127: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Update/req
      -- CP-element group 127: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Sample/ack
      -- CP-element group 127: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_update_start_
      -- CP-element group 127: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_sample_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(127)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(127)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(127) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_AFB_NIC_RESPONSE_1101_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(127)); -- 
    req_2090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_1633_elements(127), ack => WPIPE_AFB_NIC_RESPONSE_1101_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	134 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	126 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Update/ack
      -- CP-element group 128: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/WPIPE_AFB_NIC_RESPONSE_1101_update_completed_
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(128)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(128)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(128) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(128)); -- 
    -- CP-element group 129:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	10 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(129)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(129)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(129) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(129) is a control-delay.
    cp_element_129_delay: control_delay_element  generic map(name => " 129_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(9), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(129), clk => clk, reset =>reset);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	91 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	122 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1002_call_stmt_1087_delay
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(130)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(130)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(130) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(91), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	98 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	122 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1007_call_stmt_1087_delay
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(131)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(131)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(131) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(131) is a control-delay.
    cp_element_131_delay: control_delay_element  generic map(name => " 131_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(98), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(131), clk => clk, reset =>reset);
    -- CP-element group 132:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	109 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	122 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1020_call_stmt_1087_delay
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(132)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(132)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(132) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(132) is a control-delay.
    cp_element_132_delay: control_delay_element  generic map(name => " 132_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(109), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(132), clk => clk, reset =>reset);
    -- CP-element group 133:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	120 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	122 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/array_obj_ref_1079_call_stmt_1087_delay
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(133)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(133)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(133) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group SoftwareRegisterAccessDaemon_CP_1633_elements(133) is a control-delay.
    cp_element_133_delay: control_delay_element  generic map(name => " 133_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_1633_elements(120), ack => SoftwareRegisterAccessDaemon_CP_1633_elements(133), clk => clk, reset =>reset);
    -- CP-element group 134:  join  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	12 
    -- CP-element group 134: 	113 
    -- CP-element group 134: 	128 
    -- CP-element group 134: 	125 
    -- CP-element group 134: 	106 
    -- CP-element group 134: 	95 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	6 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_949/do_while_stmt_950/do_while_stmt_950_loop_body/$exit
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(134)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(134)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(134) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_1633_elements(12) & SoftwareRegisterAccessDaemon_CP_1633_elements(113) & SoftwareRegisterAccessDaemon_CP_1633_elements(128) & SoftwareRegisterAccessDaemon_CP_1633_elements(125) & SoftwareRegisterAccessDaemon_CP_1633_elements(106) & SoftwareRegisterAccessDaemon_CP_1633_elements(95);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	5 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (2) 
      -- CP-element group 135: 	 branch_block_stmt_949/do_while_stmt_950/loop_exit/$exit
      -- CP-element group 135: 	 branch_block_stmt_949/do_while_stmt_950/loop_exit/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(135)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(135)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(135) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:do_while_stmt_950_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_950_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	5 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_949/do_while_stmt_950/loop_taken/$exit
      -- CP-element group 136: 	 branch_block_stmt_949/do_while_stmt_950/loop_taken/ack
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(136)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(136)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(136) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:do_while_stmt_950_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_950_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_1633_elements(136)); -- 
    -- CP-element group 137:  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	3 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	1 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_949/do_while_stmt_950/$exit
      -- 
    -- logger for CP element group SoftwareRegisterAccessDaemon_CP_1633_elements(137)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and SoftwareRegisterAccessDaemon_CP_1633_elements(137)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:SoftwareRegisterAccessDaemon:CP:SoftwareRegisterAccessDaemon_CP_1633_elements(137) fired."); 
        -- 
      end if; --
    end process; 
    SoftwareRegisterAccessDaemon_CP_1633_elements(137) <= SoftwareRegisterAccessDaemon_CP_1633_elements(3);
    SoftwareRegisterAccessDaemon_do_while_stmt_950_terminator_2106: loop_terminator -- 
      generic map (name => " SoftwareRegisterAccessDaemon_do_while_stmt_950_terminator_2106", max_iterations_in_flight =>31) 
      port map(loop_body_exit => SoftwareRegisterAccessDaemon_CP_1633_elements(6),loop_continue => SoftwareRegisterAccessDaemon_CP_1633_elements(136),loop_terminate => SoftwareRegisterAccessDaemon_CP_1633_elements(135),loop_back => SoftwareRegisterAccessDaemon_CP_1633_elements(4),loop_exit => SoftwareRegisterAccessDaemon_CP_1633_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_952_phi_seq_1696_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(21);
      SoftwareRegisterAccessDaemon_CP_1633_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(24);
      SoftwareRegisterAccessDaemon_CP_1633_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(26);
      SoftwareRegisterAccessDaemon_CP_1633_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(19);
      SoftwareRegisterAccessDaemon_CP_1633_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(28);
      SoftwareRegisterAccessDaemon_CP_1633_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(30);
      SoftwareRegisterAccessDaemon_CP_1633_elements(20) <= phi_mux_reqs(1);
      phi_stmt_952_phi_seq_1696 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_952_phi_seq_1696") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1633_elements(11), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(17), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1633_elements(13), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(18), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_958_phi_seq_1740_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(40);
      SoftwareRegisterAccessDaemon_CP_1633_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(43);
      SoftwareRegisterAccessDaemon_CP_1633_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(45);
      SoftwareRegisterAccessDaemon_CP_1633_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(38);
      SoftwareRegisterAccessDaemon_CP_1633_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(49);
      SoftwareRegisterAccessDaemon_CP_1633_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(50);
      SoftwareRegisterAccessDaemon_CP_1633_elements(39) <= phi_mux_reqs(1);
      phi_stmt_958_phi_seq_1740 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_958_phi_seq_1740") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1633_elements(34), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(35), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1633_elements(36), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(37), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_963_phi_seq_1784_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(59);
      SoftwareRegisterAccessDaemon_CP_1633_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(62);
      SoftwareRegisterAccessDaemon_CP_1633_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(64);
      SoftwareRegisterAccessDaemon_CP_1633_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(57);
      SoftwareRegisterAccessDaemon_CP_1633_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(68);
      SoftwareRegisterAccessDaemon_CP_1633_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(69);
      SoftwareRegisterAccessDaemon_CP_1633_elements(58) <= phi_mux_reqs(1);
      phi_stmt_963_phi_seq_1784 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_963_phi_seq_1784") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1633_elements(53), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(54), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1633_elements(55), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(56), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_968_phi_seq_1828_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(78);
      SoftwareRegisterAccessDaemon_CP_1633_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(81);
      SoftwareRegisterAccessDaemon_CP_1633_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(83);
      SoftwareRegisterAccessDaemon_CP_1633_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(76);
      SoftwareRegisterAccessDaemon_CP_1633_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(87);
      SoftwareRegisterAccessDaemon_CP_1633_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(88);
      SoftwareRegisterAccessDaemon_CP_1633_elements(77) <= phi_mux_reqs(1);
      phi_stmt_968_phi_seq_1828 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_968_phi_seq_1828") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_1633_elements(72), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(73), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_1633_elements(74), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(75), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_1633_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1658_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(7);
        preds(1)  <= SoftwareRegisterAccessDaemon_CP_1633_elements(8);
        entry_tmerge_1658 : transition_merge -- 
          generic map(name => " entry_tmerge_1658")
          port map (preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_1633_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_980_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_988_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_996_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u32_u35_1014_wire : std_logic_vector(34 downto 0);
    signal EQ_u1_u1_1056_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1065_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1074_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1053_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1062_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1071_wire : std_logic_vector(0 downto 0);
    signal FREE_Q_32_1008 : std_logic_vector(31 downto 0);
    signal INIT_952 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_977_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_985_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_993_wire : std_logic_vector(0 downto 0);
    signal R_index_1078_resized : std_logic_vector(5 downto 0);
    signal R_index_1078_scaled : std_logic_vector(5 downto 0);
    signal addr_1041 : std_logic_vector(35 downto 0);
    signal array_obj_ref_1002_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1002_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1002_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1007_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1007_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1020_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1020_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1020_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1079_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1079_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_1079_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1079_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1079_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_1079_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1079_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_1037 : std_logic_vector(3 downto 0);
    signal check_control_regsiter_1058 : std_logic_vector(0 downto 0);
    signal check_control_regsiter_1058_962_buffered : std_logic_vector(0 downto 0);
    signal check_free_q_1067 : std_logic_vector(0 downto 0);
    signal check_free_q_1067_967_buffered : std_logic_vector(0 downto 0);
    signal check_num_server_1076 : std_logic_vector(0 downto 0);
    signal check_num_server_1076_972_buffered : std_logic_vector(0 downto 0);
    signal control_register_958 : std_logic_vector(0 downto 0);
    signal free_q_963 : std_logic_vector(0 downto 0);
    signal index_1049 : std_logic_vector(5 downto 0);
    signal konst_1052_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1055_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1061_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1064_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1070_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1073_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1105_wire_constant : std_logic_vector(0 downto 0);
    signal lock_1029 : std_logic_vector(0 downto 0);
    signal num_server_968 : std_logic_vector(0 downto 0);
    signal rdata_1094 : std_logic_vector(31 downto 0);
    signal req_1024 : std_logic_vector(73 downto 0);
    signal resp_1100 : std_logic_vector(32 downto 0);
    signal rval_1080 : std_logic_vector(31 downto 0);
    signal rwbar_1033 : std_logic_vector(0 downto 0);
    signal type_cast_1013_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_1015_wire : std_logic_vector(35 downto 0);
    signal type_cast_1092_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1097_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_955_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_957_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_961_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_966_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_971_wire_constant : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_982 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_990 : std_logic_vector(0 downto 0);
    signal update_server_num_998 : std_logic_vector(0 downto 0);
    signal wdata_1045 : std_logic_vector(31 downto 0);
    signal wval_1087 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1002_word_address_0 <= "000000";
    array_obj_ref_1007_word_address_0 <= "010010";
    array_obj_ref_1020_word_address_0 <= "000001";
    array_obj_ref_1079_offset_scale_factor_0 <= "000001";
    array_obj_ref_1079_resized_base_address <= "000000";
    array_obj_ref_1079_word_offset_0 <= "000000";
    konst_1052_wire_constant <= "000000";
    konst_1055_wire_constant <= "0";
    konst_1061_wire_constant <= "010010";
    konst_1064_wire_constant <= "0";
    konst_1070_wire_constant <= "000001";
    konst_1073_wire_constant <= "0";
    konst_1105_wire_constant <= "1";
    type_cast_1013_wire_constant <= "000";
    type_cast_1092_wire_constant <= "00000000000000000000000000000000";
    type_cast_1097_wire_constant <= "0";
    type_cast_955_wire_constant <= "0";
    type_cast_957_wire_constant <= "1";
    type_cast_961_wire_constant <= "0";
    type_cast_966_wire_constant <= "0";
    type_cast_971_wire_constant <= "0";
    -- logger for phi phi_stmt_952
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_952_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_952:input-0 type_cast_955_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_955_wire_constant));
          --
        end if;
        if phi_stmt_952_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_952:input-1 type_cast_957_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_957_wire_constant));
          --
        end if;
        if phi_stmt_952_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_952:sample-completed");
          --
        end if;
        if phi_stmt_952_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_952:output INIT_952= " & Convert_SLV_To_Hex_String(INIT_952));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_952: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_955_wire_constant & type_cast_957_wire_constant;
      req <= phi_stmt_952_req_0 & phi_stmt_952_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_952",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_952_ack_0,
          idata => idata,
          odata => INIT_952,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_952
    -- logger for phi phi_stmt_958
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_958_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_958:input-0 type_cast_961_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_961_wire_constant));
          --
        end if;
        if phi_stmt_958_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_958:input-1 check_control_regsiter_1058_962_buffered= " & Convert_SLV_To_Hex_String(check_control_regsiter_1058_962_buffered));
          --
        end if;
        if phi_stmt_958_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_958:sample-completed");
          --
        end if;
        if phi_stmt_958_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_958:output control_register_958= " & Convert_SLV_To_Hex_String(control_register_958));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_958: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_961_wire_constant & check_control_regsiter_1058_962_buffered;
      req <= phi_stmt_958_req_0 & phi_stmt_958_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_958",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_958_ack_0,
          idata => idata,
          odata => control_register_958,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_958
    -- logger for phi phi_stmt_963
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_963_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_963:input-0 type_cast_966_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_966_wire_constant));
          --
        end if;
        if phi_stmt_963_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_963:input-1 check_free_q_1067_967_buffered= " & Convert_SLV_To_Hex_String(check_free_q_1067_967_buffered));
          --
        end if;
        if phi_stmt_963_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_963:sample-completed");
          --
        end if;
        if phi_stmt_963_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_963:output free_q_963= " & Convert_SLV_To_Hex_String(free_q_963));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_963: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_966_wire_constant & check_free_q_1067_967_buffered;
      req <= phi_stmt_963_req_0 & phi_stmt_963_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_963",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_963_ack_0,
          idata => idata,
          odata => free_q_963,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_963
    -- logger for phi phi_stmt_968
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_968_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_968:input-0 type_cast_971_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_971_wire_constant));
          --
        end if;
        if phi_stmt_968_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_968:input-1 check_num_server_1076_972_buffered= " & Convert_SLV_To_Hex_String(check_num_server_1076_972_buffered));
          --
        end if;
        if phi_stmt_968_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_968:sample-completed");
          --
        end if;
        if phi_stmt_968_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:SoftwareRegisterAccessDaemon:DP:phi_stmt_968:output num_server_968= " & Convert_SLV_To_Hex_String(num_server_968));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_968: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_971_wire_constant & check_num_server_1076_972_buffered;
      req <= phi_stmt_968_req_0 & phi_stmt_968_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_968",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_968_ack_0,
          idata => idata,
          odata => num_server_968,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_968
    -- logger for split-operator MUX_1093_inst flow-through 
    process(rdata_1094) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:MUX_1093_inst:flowthrough inputs: " & " rwbar_1033 = "& Convert_SLV_To_Hex_String(rwbar_1033) & " rval_1080 = "& Convert_SLV_To_Hex_String(rval_1080) & " type_cast_1092_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1092_wire_constant) & " outputs:" & " rdata_1094= "  & Convert_SLV_To_Hex_String(rdata_1094));
      --
    end process; 
    -- flow-through select operator MUX_1093_inst
    rdata_1094 <= rval_1080 when (rwbar_1033(0) /=  '0') else type_cast_1092_wire_constant;
    -- logger for split-operator slice_1028_inst flow-through 
    process(lock_1029) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:slice_1028_inst:flowthrough inputs: " & " req_1024 = "& Convert_SLV_To_Hex_String(req_1024) & " outputs:" & " lock_1029= "  & Convert_SLV_To_Hex_String(lock_1029));
      --
    end process; 
    -- flow-through slice operator slice_1028_inst
    lock_1029 <= req_1024(73 downto 73);
    -- logger for split-operator slice_1032_inst flow-through 
    process(rwbar_1033) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:slice_1032_inst:flowthrough inputs: " & " req_1024 = "& Convert_SLV_To_Hex_String(req_1024) & " outputs:" & " rwbar_1033= "  & Convert_SLV_To_Hex_String(rwbar_1033));
      --
    end process; 
    -- flow-through slice operator slice_1032_inst
    rwbar_1033 <= req_1024(72 downto 72);
    -- logger for split-operator slice_1036_inst flow-through 
    process(bmask_1037) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:slice_1036_inst:flowthrough inputs: " & " req_1024 = "& Convert_SLV_To_Hex_String(req_1024) & " outputs:" & " bmask_1037= "  & Convert_SLV_To_Hex_String(bmask_1037));
      --
    end process; 
    -- flow-through slice operator slice_1036_inst
    bmask_1037 <= req_1024(71 downto 68);
    -- logger for split-operator slice_1040_inst flow-through 
    process(addr_1041) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:slice_1040_inst:flowthrough inputs: " & " req_1024 = "& Convert_SLV_To_Hex_String(req_1024) & " outputs:" & " addr_1041= "  & Convert_SLV_To_Hex_String(addr_1041));
      --
    end process; 
    -- flow-through slice operator slice_1040_inst
    addr_1041 <= req_1024(67 downto 32);
    -- logger for split-operator slice_1044_inst flow-through 
    process(wdata_1045) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:slice_1044_inst:flowthrough inputs: " & " req_1024 = "& Convert_SLV_To_Hex_String(req_1024) & " outputs:" & " wdata_1045= "  & Convert_SLV_To_Hex_String(wdata_1045));
      --
    end process; 
    -- flow-through slice operator slice_1044_inst
    wdata_1045 <= req_1024(31 downto 0);
    -- logger for split-operator slice_1048_inst flow-through 
    process(index_1049) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:slice_1048_inst:flowthrough inputs: " & " addr_1041 = "& Convert_SLV_To_Hex_String(addr_1041) & " outputs:" & " index_1049= "  & Convert_SLV_To_Hex_String(index_1049));
      --
    end process; 
    -- flow-through slice operator slice_1048_inst
    index_1049 <= addr_1041(5 downto 0);
    -- logger for split-operator check_control_regsiter_1058_962_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if check_control_regsiter_1058_962_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:check_control_regsiter_1058_962_buf:started:   inputs: " & " check_control_regsiter_1058 = "& Convert_SLV_To_Hex_String(check_control_regsiter_1058));
          --
        end if; 
        if check_control_regsiter_1058_962_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:check_control_regsiter_1058_962_buf:finished:  outputs: " & " check_control_regsiter_1058_962_buffered= "  & Convert_SLV_To_Hex_String(check_control_regsiter_1058_962_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    check_control_regsiter_1058_962_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_control_regsiter_1058_962_buf_req_0;
      check_control_regsiter_1058_962_buf_ack_0<= wack(0);
      rreq(0) <= check_control_regsiter_1058_962_buf_req_1;
      check_control_regsiter_1058_962_buf_ack_1<= rack(0);
      check_control_regsiter_1058_962_buf : InterlockBuffer generic map ( -- 
        name => "check_control_regsiter_1058_962_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_control_regsiter_1058,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_control_regsiter_1058_962_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator check_free_q_1067_967_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if check_free_q_1067_967_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:check_free_q_1067_967_buf:started:   inputs: " & " check_free_q_1067 = "& Convert_SLV_To_Hex_String(check_free_q_1067));
          --
        end if; 
        if check_free_q_1067_967_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:check_free_q_1067_967_buf:finished:  outputs: " & " check_free_q_1067_967_buffered= "  & Convert_SLV_To_Hex_String(check_free_q_1067_967_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    check_free_q_1067_967_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_free_q_1067_967_buf_req_0;
      check_free_q_1067_967_buf_ack_0<= wack(0);
      rreq(0) <= check_free_q_1067_967_buf_req_1;
      check_free_q_1067_967_buf_ack_1<= rack(0);
      check_free_q_1067_967_buf : InterlockBuffer generic map ( -- 
        name => "check_free_q_1067_967_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_free_q_1067,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_free_q_1067_967_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator check_num_server_1076_972_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if check_num_server_1076_972_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:check_num_server_1076_972_buf:started:   inputs: " & " check_num_server_1076 = "& Convert_SLV_To_Hex_String(check_num_server_1076));
          --
        end if; 
        if check_num_server_1076_972_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:check_num_server_1076_972_buf:finished:  outputs: " & " check_num_server_1076_972_buffered= "  & Convert_SLV_To_Hex_String(check_num_server_1076_972_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    check_num_server_1076_972_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_num_server_1076_972_buf_req_0;
      check_num_server_1076_972_buf_ack_0<= wack(0);
      rreq(0) <= check_num_server_1076_972_buf_req_1;
      check_num_server_1076_972_buf_ack_1<= rack(0);
      check_num_server_1076_972_buf : InterlockBuffer generic map ( -- 
        name => "check_num_server_1076_972_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_num_server_1076,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_num_server_1076_972_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1015_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1015_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:type_cast_1015_inst:started:   inputs: " & " update_free_q_pipe_990 (guard)= " & Convert_SLV_To_String(update_free_q_pipe_990) & " CONCAT_u32_u35_1014_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u35_1014_wire));
          --
        end if; 
        if type_cast_1015_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:type_cast_1015_inst:finished:  outputs: " & " type_cast_1015_wire= "  & Convert_SLV_To_Hex_String(type_cast_1015_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1015_inst_req_0;
      type_cast_1015_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1015_inst_req_1;
      type_cast_1015_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  update_free_q_pipe_990(0);
      type_cast_1015_inst_gI: SplitGuardInterface generic map(name => "type_cast_1015_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 35,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => CONCAT_u32_u35_1014_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1015_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for operator array_obj_ref_1002_gather_scatter flow-through 
    process(array_obj_ref_1002_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1002_gather_scatter:flowthrough  inputs: " & " update_control_register_pipe_982 (guard)= " & Convert_SLV_To_String(update_control_register_pipe_982) & " array_obj_ref_1002_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1002_data_0) & "outputs: " & " array_obj_ref_1002_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1002_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1002_gather_scatter
    process(array_obj_ref_1002_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1002_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1002_wire <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1007_gather_scatter flow-through 
    process(FREE_Q_32_1008) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1007_gather_scatter:flowthrough  inputs: " & " update_free_q_pipe_990 (guard)= " & Convert_SLV_To_String(update_free_q_pipe_990) & " array_obj_ref_1007_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1007_data_0) & "outputs: " & " FREE_Q_32_1008= "  & Convert_SLV_To_Hex_String(FREE_Q_32_1008));
      --
    end process; 
    -- equivalence array_obj_ref_1007_gather_scatter
    process(array_obj_ref_1007_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1007_data_0;
      ov(31 downto 0) := iv;
      FREE_Q_32_1008 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1020_gather_scatter flow-through 
    process(array_obj_ref_1020_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1020_gather_scatter:flowthrough  inputs: " & " update_server_num_998 (guard)= " & Convert_SLV_To_String(update_server_num_998) & " array_obj_ref_1020_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1020_data_0) & "outputs: " & " array_obj_ref_1020_wire= "  & Convert_SLV_To_Hex_String(array_obj_ref_1020_wire));
      --
    end process; 
    -- equivalence array_obj_ref_1020_gather_scatter
    process(array_obj_ref_1020_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1020_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1020_wire <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1079_addr_0 flow-through 
    process(array_obj_ref_1079_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_addr_0:flowthrough  inputs: " & " array_obj_ref_1079_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_1079_root_address) & "outputs: " & " array_obj_ref_1079_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1079_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_1079_addr_0
    process(array_obj_ref_1079_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1079_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_1079_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1079_gather_scatter flow-through 
    process(rval_1080) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_gather_scatter:flowthrough  inputs: " & " array_obj_ref_1079_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1079_data_0) & "outputs: " & " rval_1080= "  & Convert_SLV_To_Hex_String(rval_1080));
      --
    end process; 
    -- equivalence array_obj_ref_1079_gather_scatter
    process(array_obj_ref_1079_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1079_data_0;
      ov(31 downto 0) := iv;
      rval_1080 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1079_index_0_rename flow-through 
    process(R_index_1078_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_index_0_rename:flowthrough  inputs: " & " R_index_1078_resized = "& Convert_SLV_To_Hex_String(R_index_1078_resized) & "outputs: " & " R_index_1078_scaled= "  & Convert_SLV_To_Hex_String(R_index_1078_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_1079_index_0_rename
    process(R_index_1078_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1078_resized;
      ov(5 downto 0) := iv;
      R_index_1078_scaled <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1079_index_0_resize flow-through 
    process(R_index_1078_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_index_0_resize:flowthrough  inputs: " & " index_1049 = "& Convert_SLV_To_Hex_String(index_1049) & "outputs: " & " R_index_1078_resized= "  & Convert_SLV_To_Hex_String(R_index_1078_resized));
      --
    end process; 
    -- equivalence array_obj_ref_1079_index_0_resize
    process(index_1049) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_1049;
      ov(5 downto 0) := iv;
      R_index_1078_resized <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1079_index_offset flow-through 
    process(array_obj_ref_1079_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_index_offset:flowthrough  inputs: " & " R_index_1078_scaled = "& Convert_SLV_To_Hex_String(R_index_1078_scaled) & "outputs: " & " array_obj_ref_1079_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_1079_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_1079_index_offset
    process(R_index_1078_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_1078_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_1079_final_offset <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_1079_root_address_inst flow-through 
    process(array_obj_ref_1079_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_root_address_inst:flowthrough  inputs: " & " array_obj_ref_1079_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_1079_final_offset) & "outputs: " & " array_obj_ref_1079_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_1079_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_1079_root_address_inst
    process(array_obj_ref_1079_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1079_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_1079_root_address <= ov(5 downto 0);
      --
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_950_branch_req_0," req0 do_while_stmt_950_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_950_branch_ack_0," ack0 do_while_stmt_950_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_950_branch_ack_1," ack1 do_while_stmt_950_branch");
    do_while_stmt_950_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1105_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_950_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_950_branch_req_0,
          ack0 => do_while_stmt_950_branch_ack_0,
          ack1 => do_while_stmt_950_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator AND_u1_u1_1057_inst flow-through 
    process(check_control_regsiter_1058) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:AND_u1_u1_1057_inst:flowthrough inputs: " & " EQ_u6_u1_1053_wire = "& Convert_SLV_To_Hex_String(EQ_u6_u1_1053_wire) & " EQ_u1_u1_1056_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_1056_wire) & " outputs:" & " check_control_regsiter_1058= "  & Convert_SLV_To_Hex_String(check_control_regsiter_1058));
      --
    end process; 
    -- binary operator AND_u1_u1_1057_inst
    process(EQ_u6_u1_1053_wire, EQ_u1_u1_1056_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1053_wire, EQ_u1_u1_1056_wire, tmp_var);
      check_control_regsiter_1058 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_1066_inst flow-through 
    process(check_free_q_1067) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:AND_u1_u1_1066_inst:flowthrough inputs: " & " EQ_u6_u1_1062_wire = "& Convert_SLV_To_Hex_String(EQ_u6_u1_1062_wire) & " EQ_u1_u1_1065_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_1065_wire) & " outputs:" & " check_free_q_1067= "  & Convert_SLV_To_Hex_String(check_free_q_1067));
      --
    end process; 
    -- binary operator AND_u1_u1_1066_inst
    process(EQ_u6_u1_1062_wire, EQ_u1_u1_1065_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1062_wire, EQ_u1_u1_1065_wire, tmp_var);
      check_free_q_1067 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_1075_inst flow-through 
    process(check_num_server_1076) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:AND_u1_u1_1075_inst:flowthrough inputs: " & " EQ_u6_u1_1071_wire = "& Convert_SLV_To_Hex_String(EQ_u6_u1_1071_wire) & " EQ_u1_u1_1074_wire = "& Convert_SLV_To_Hex_String(EQ_u1_u1_1074_wire) & " outputs:" & " check_num_server_1076= "  & Convert_SLV_To_Hex_String(check_num_server_1076));
      --
    end process; 
    -- binary operator AND_u1_u1_1075_inst
    process(EQ_u6_u1_1071_wire, EQ_u1_u1_1074_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1071_wire, EQ_u1_u1_1074_wire, tmp_var);
      check_num_server_1076 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_980_inst flow-through 
    process(AND_u1_u1_980_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:AND_u1_u1_980_inst:flowthrough inputs: " & " INIT_952 = "& Convert_SLV_To_Hex_String(INIT_952) & " control_register_958 = "& Convert_SLV_To_Hex_String(control_register_958) & " outputs:" & " AND_u1_u1_980_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_980_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_980_inst
    process(INIT_952, control_register_958) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_952, control_register_958, tmp_var);
      AND_u1_u1_980_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_988_inst flow-through 
    process(AND_u1_u1_988_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:AND_u1_u1_988_inst:flowthrough inputs: " & " INIT_952 = "& Convert_SLV_To_Hex_String(INIT_952) & " free_q_963 = "& Convert_SLV_To_Hex_String(free_q_963) & " outputs:" & " AND_u1_u1_988_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_988_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_988_inst
    process(INIT_952, free_q_963) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_952, free_q_963, tmp_var);
      AND_u1_u1_988_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_996_inst flow-through 
    process(AND_u1_u1_996_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:AND_u1_u1_996_inst:flowthrough inputs: " & " INIT_952 = "& Convert_SLV_To_Hex_String(INIT_952) & " num_server_968 = "& Convert_SLV_To_Hex_String(num_server_968) & " outputs:" & " AND_u1_u1_996_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_996_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_996_inst
    process(INIT_952, num_server_968) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_952, num_server_968, tmp_var);
      AND_u1_u1_996_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u33_1099_inst flow-through 
    process(resp_1100) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:CONCAT_u1_u33_1099_inst:flowthrough inputs: " & " type_cast_1097_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1097_wire_constant) & " rdata_1094 = "& Convert_SLV_To_Hex_String(rdata_1094) & " outputs:" & " resp_1100= "  & Convert_SLV_To_Hex_String(resp_1100));
      --
    end process; 
    -- binary operator CONCAT_u1_u33_1099_inst
    process(type_cast_1097_wire_constant, rdata_1094) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1097_wire_constant, rdata_1094, tmp_var);
      resp_1100 <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u35_1014_inst flow-through 
    process(CONCAT_u32_u35_1014_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:CONCAT_u32_u35_1014_inst:flowthrough inputs: " & " update_free_q_pipe_990 (guard)= " & Convert_SLV_To_String(update_free_q_pipe_990) & " FREE_Q_32_1008 = "& Convert_SLV_To_Hex_String(FREE_Q_32_1008) & " type_cast_1013_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1013_wire_constant) & " outputs:" & " CONCAT_u32_u35_1014_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u35_1014_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u35_1014_inst
    process(FREE_Q_32_1008) -- 
      variable tmp_var : std_logic_vector(34 downto 0); -- 
    begin -- 
      ApConcat_proc(FREE_Q_32_1008, type_cast_1013_wire_constant, tmp_var);
      CONCAT_u32_u35_1014_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_1056_inst flow-through 
    process(EQ_u1_u1_1056_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:EQ_u1_u1_1056_inst:flowthrough inputs: " & " rwbar_1033 = "& Convert_SLV_To_Hex_String(rwbar_1033) & " konst_1055_wire_constant = "& Convert_SLV_To_Hex_String(konst_1055_wire_constant) & " outputs:" & " EQ_u1_u1_1056_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_1056_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_1056_inst
    process(rwbar_1033) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1033, konst_1055_wire_constant, tmp_var);
      EQ_u1_u1_1056_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_1065_inst flow-through 
    process(EQ_u1_u1_1065_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:EQ_u1_u1_1065_inst:flowthrough inputs: " & " rwbar_1033 = "& Convert_SLV_To_Hex_String(rwbar_1033) & " konst_1064_wire_constant = "& Convert_SLV_To_Hex_String(konst_1064_wire_constant) & " outputs:" & " EQ_u1_u1_1065_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_1065_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_1065_inst
    process(rwbar_1033) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1033, konst_1064_wire_constant, tmp_var);
      EQ_u1_u1_1065_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_1074_inst flow-through 
    process(EQ_u1_u1_1074_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:EQ_u1_u1_1074_inst:flowthrough inputs: " & " rwbar_1033 = "& Convert_SLV_To_Hex_String(rwbar_1033) & " konst_1073_wire_constant = "& Convert_SLV_To_Hex_String(konst_1073_wire_constant) & " outputs:" & " EQ_u1_u1_1074_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_1074_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_1074_inst
    process(rwbar_1033) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1033, konst_1073_wire_constant, tmp_var);
      EQ_u1_u1_1074_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u6_u1_1053_inst flow-through 
    process(EQ_u6_u1_1053_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:EQ_u6_u1_1053_inst:flowthrough inputs: " & " index_1049 = "& Convert_SLV_To_Hex_String(index_1049) & " konst_1052_wire_constant = "& Convert_SLV_To_Hex_String(konst_1052_wire_constant) & " outputs:" & " EQ_u6_u1_1053_wire= "  & Convert_SLV_To_Hex_String(EQ_u6_u1_1053_wire));
      --
    end process; 
    -- binary operator EQ_u6_u1_1053_inst
    process(index_1049) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1049, konst_1052_wire_constant, tmp_var);
      EQ_u6_u1_1053_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u6_u1_1062_inst flow-through 
    process(EQ_u6_u1_1062_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:EQ_u6_u1_1062_inst:flowthrough inputs: " & " index_1049 = "& Convert_SLV_To_Hex_String(index_1049) & " konst_1061_wire_constant = "& Convert_SLV_To_Hex_String(konst_1061_wire_constant) & " outputs:" & " EQ_u6_u1_1062_wire= "  & Convert_SLV_To_Hex_String(EQ_u6_u1_1062_wire));
      --
    end process; 
    -- binary operator EQ_u6_u1_1062_inst
    process(index_1049) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1049, konst_1061_wire_constant, tmp_var);
      EQ_u6_u1_1062_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u6_u1_1071_inst flow-through 
    process(EQ_u6_u1_1071_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:EQ_u6_u1_1071_inst:flowthrough inputs: " & " index_1049 = "& Convert_SLV_To_Hex_String(index_1049) & " konst_1070_wire_constant = "& Convert_SLV_To_Hex_String(konst_1070_wire_constant) & " outputs:" & " EQ_u6_u1_1071_wire= "  & Convert_SLV_To_Hex_String(EQ_u6_u1_1071_wire));
      --
    end process; 
    -- binary operator EQ_u6_u1_1071_inst
    process(index_1049) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1049, konst_1070_wire_constant, tmp_var);
      EQ_u6_u1_1071_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_977_inst flow-through 
    process(NOT_u1_u1_977_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:NOT_u1_u1_977_inst:flowthrough inputs: " & " INIT_952 = "& Convert_SLV_To_Hex_String(INIT_952) & " outputs:" & " NOT_u1_u1_977_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_977_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_977_inst
    process(INIT_952) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_952, tmp_var);
      NOT_u1_u1_977_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator NOT_u1_u1_985_inst flow-through 
    process(NOT_u1_u1_985_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:NOT_u1_u1_985_inst:flowthrough inputs: " & " INIT_952 = "& Convert_SLV_To_Hex_String(INIT_952) & " outputs:" & " NOT_u1_u1_985_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_985_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_985_inst
    process(INIT_952) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_952, tmp_var);
      NOT_u1_u1_985_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator NOT_u1_u1_993_inst flow-through 
    process(NOT_u1_u1_993_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:NOT_u1_u1_993_inst:flowthrough inputs: " & " INIT_952 = "& Convert_SLV_To_Hex_String(INIT_952) & " outputs:" & " NOT_u1_u1_993_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_993_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_993_inst
    process(INIT_952) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_952, tmp_var);
      NOT_u1_u1_993_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator OR_u1_u1_981_inst flow-through 
    process(update_control_register_pipe_982) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:OR_u1_u1_981_inst:flowthrough inputs: " & " NOT_u1_u1_977_wire = "& Convert_SLV_To_Hex_String(NOT_u1_u1_977_wire) & " AND_u1_u1_980_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_980_wire) & " outputs:" & " update_control_register_pipe_982= "  & Convert_SLV_To_Hex_String(update_control_register_pipe_982));
      --
    end process; 
    -- binary operator OR_u1_u1_981_inst
    process(NOT_u1_u1_977_wire, AND_u1_u1_980_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_977_wire, AND_u1_u1_980_wire, tmp_var);
      update_control_register_pipe_982 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_989_inst flow-through 
    process(update_free_q_pipe_990) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:OR_u1_u1_989_inst:flowthrough inputs: " & " NOT_u1_u1_985_wire = "& Convert_SLV_To_Hex_String(NOT_u1_u1_985_wire) & " AND_u1_u1_988_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_988_wire) & " outputs:" & " update_free_q_pipe_990= "  & Convert_SLV_To_Hex_String(update_free_q_pipe_990));
      --
    end process; 
    -- binary operator OR_u1_u1_989_inst
    process(NOT_u1_u1_985_wire, AND_u1_u1_988_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_985_wire, AND_u1_u1_988_wire, tmp_var);
      update_free_q_pipe_990 <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_997_inst flow-through 
    process(update_server_num_998) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:OR_u1_u1_997_inst:flowthrough inputs: " & " NOT_u1_u1_993_wire = "& Convert_SLV_To_Hex_String(NOT_u1_u1_993_wire) & " AND_u1_u1_996_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_996_wire) & " outputs:" & " update_server_num_998= "  & Convert_SLV_To_Hex_String(update_server_num_998));
      --
    end process; 
    -- binary operator OR_u1_u1_997_inst
    process(NOT_u1_u1_993_wire, AND_u1_u1_996_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_993_wire, AND_u1_u1_996_wire, tmp_var);
      update_server_num_998 <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_1002_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1002_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1002_load_0:started:   inputs: " & " update_control_register_pipe_982 (guard)= " & Convert_SLV_To_String(update_control_register_pipe_982) & " array_obj_ref_1002_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1002_word_address_0));
          --
        end if; 
        if array_obj_ref_1002_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1002_load_0:finished:  outputs: " & " array_obj_ref_1002_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1002_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1007_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1007_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1007_load_0:started:   inputs: " & " update_free_q_pipe_990 (guard)= " & Convert_SLV_To_String(update_free_q_pipe_990) & " array_obj_ref_1007_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1007_word_address_0));
          --
        end if; 
        if array_obj_ref_1007_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1007_load_0:finished:  outputs: " & " array_obj_ref_1007_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1007_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1020_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1020_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1020_load_0:started:   inputs: " & " update_server_num_998 (guard)= " & Convert_SLV_To_String(update_server_num_998) & " array_obj_ref_1020_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1020_word_address_0));
          --
        end if; 
        if array_obj_ref_1020_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1020_load_0:finished:  outputs: " & " array_obj_ref_1020_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1020_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator array_obj_ref_1079_load_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_1079_load_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_load_0:started:   inputs: " & " array_obj_ref_1079_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_1079_word_address_0));
          --
        end if; 
        if array_obj_ref_1079_load_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:array_obj_ref_1079_load_0:finished:  outputs: " & " array_obj_ref_1079_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_1079_data_0));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared load operator group (0) : array_obj_ref_1002_load_0 array_obj_ref_1007_load_0 array_obj_ref_1020_load_0 array_obj_ref_1079_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1002_load_0_req_0,
        array_obj_ref_1002_load_0_ack_0,
        array_obj_ref_1002_load_0_req_1,
        array_obj_ref_1002_load_0_ack_1,
        "array_obj_ref_1002_load_0",
        "memory_space_0" ,
        array_obj_ref_1002_data_0,
        array_obj_ref_1002_word_address_0,
        "array_obj_ref_1002_data_0",
        "array_obj_ref_1002_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1007_load_0_req_0,
        array_obj_ref_1007_load_0_ack_0,
        array_obj_ref_1007_load_0_req_1,
        array_obj_ref_1007_load_0_ack_1,
        "array_obj_ref_1007_load_0",
        "memory_space_0" ,
        array_obj_ref_1007_data_0,
        array_obj_ref_1007_word_address_0,
        "array_obj_ref_1007_data_0",
        "array_obj_ref_1007_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1020_load_0_req_0,
        array_obj_ref_1020_load_0_ack_0,
        array_obj_ref_1020_load_0_req_1,
        array_obj_ref_1020_load_0_ack_1,
        "array_obj_ref_1020_load_0",
        "memory_space_0" ,
        array_obj_ref_1020_data_0,
        array_obj_ref_1020_word_address_0,
        "array_obj_ref_1020_data_0",
        "array_obj_ref_1020_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        array_obj_ref_1079_load_0_req_0,
        array_obj_ref_1079_load_0_ack_0,
        array_obj_ref_1079_load_0_req_1,
        array_obj_ref_1079_load_0_ack_1,
        "array_obj_ref_1079_load_0",
        "memory_space_0" ,
        array_obj_ref_1079_data_0,
        array_obj_ref_1079_word_address_0,
        "array_obj_ref_1079_data_0",
        "array_obj_ref_1079_word_address_0" -- 
      );
      reqL_unguarded(3) <= array_obj_ref_1002_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1007_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1020_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1079_load_0_req_0;
      array_obj_ref_1002_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1007_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1020_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1079_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= array_obj_ref_1002_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1007_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1020_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1079_load_0_req_1;
      array_obj_ref_1002_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1007_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1020_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1079_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= update_server_num_998(0);
      guard_vector(2)  <= update_free_q_pipe_990(0);
      guard_vector(3)  <= update_control_register_pipe_982(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1002_word_address_0 & array_obj_ref_1007_word_address_0 & array_obj_ref_1020_word_address_0 & array_obj_ref_1079_word_address_0;
      array_obj_ref_1002_data_0 <= data_out(127 downto 96);
      array_obj_ref_1007_data_0 <= data_out(95 downto 64);
      array_obj_ref_1020_data_0 <= data_out(63 downto 32);
      array_obj_ref_1079_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(5 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logger for split-operator RPIPE_AFB_NIC_REQUEST_1023_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_AFB_NIC_REQUEST_1023_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:RPIPE_AFB_NIC_REQUEST_1023_inst:started:   PipeRead from AFB_NIC_REQUEST inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_AFB_NIC_REQUEST_1023_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:RPIPE_AFB_NIC_REQUEST_1023_inst:finished:  outputs: " & " req_1024= "  & Convert_SLV_To_Hex_String(req_1024));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_AFB_NIC_REQUEST_1023_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(73 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1023_inst_req_0;
      RPIPE_AFB_NIC_REQUEST_1023_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1023_inst_req_1;
      RPIPE_AFB_NIC_REQUEST_1023_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_1024 <= data_out(73 downto 0);
      AFB_NIC_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST_read_0", data_width => 74,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_REQUEST_pipe_read_req(0),
          oack => AFB_NIC_REQUEST_pipe_read_ack(0),
          odata => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_AFB_NIC_RESPONSE_1101_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_AFB_NIC_RESPONSE_1101_inst:started:   PipeWrite to AFB_NIC_RESPONSE inputs: " & " resp_1100 = "& Convert_SLV_To_Hex_String(resp_1100));
          --
        end if; 
        if WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_AFB_NIC_RESPONSE_1101_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_AFB_NIC_RESPONSE_1101_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1101_inst_req_0;
      WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_1101_inst_req_1;
      WPIPE_AFB_NIC_RESPONSE_1101_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_1100;
      AFB_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_RESPONSE_pipe_write_req(0),
          oack => AFB_NIC_RESPONSE_pipe_write_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_CONTROL_REGISTER_1000_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_CONTROL_REGISTER_1000_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_CONTROL_REGISTER_1000_inst:started:   PipeWrite to CONTROL_REGISTER inputs: " & " update_control_register_pipe_982 (guard)= " & Convert_SLV_To_String(update_control_register_pipe_982) & " array_obj_ref_1002_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1002_wire));
          --
        end if; 
        if WPIPE_CONTROL_REGISTER_1000_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_CONTROL_REGISTER_1000_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_CONTROL_REGISTER_1000_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1000_inst_req_0;
      WPIPE_CONTROL_REGISTER_1000_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1000_inst_req_1;
      WPIPE_CONTROL_REGISTER_1000_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_982(0);
      data_in <= array_obj_ref_1002_wire;
      CONTROL_REGISTER_write_1_gI: SplitGuardInterface generic map(name => "CONTROL_REGISTER_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      CONTROL_REGISTER_write_1: OutputPortRevised -- 
        generic map ( name => "CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => CONTROL_REGISTER_pipe_write_req(0),
          oack => CONTROL_REGISTER_pipe_write_ack(0),
          odata => CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator WPIPE_FREE_Q_1010_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_FREE_Q_1010_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_FREE_Q_1010_inst:started:   PipeWrite to FREE_Q inputs: " & " update_free_q_pipe_990 (guard)= " & Convert_SLV_To_String(update_free_q_pipe_990) & " type_cast_1015_wire = "& Convert_SLV_To_Hex_String(type_cast_1015_wire));
          --
        end if; 
        if WPIPE_FREE_Q_1010_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_FREE_Q_1010_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (2) : WPIPE_FREE_Q_1010_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_FREE_Q_1010_inst_req_0;
      WPIPE_FREE_Q_1010_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_FREE_Q_1010_inst_req_1;
      WPIPE_FREE_Q_1010_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_free_q_pipe_990(0);
      data_in <= type_cast_1015_wire;
      FREE_Q_write_2_gI: SplitGuardInterface generic map(name => "FREE_Q_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      FREE_Q_write_2: OutputPortRevised -- 
        generic map ( name => "FREE_Q", data_width => 36, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => FREE_Q_pipe_write_req(0),
          oack => FREE_Q_pipe_write_ack(0),
          odata => FREE_Q_pipe_write_data(35 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logger for split-operator WPIPE_NUMBER_OF_SERVERS_1018_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_NUMBER_OF_SERVERS_1018_inst:started:   PipeWrite to NUMBER_OF_SERVERS inputs: " & " update_server_num_998 (guard)= " & Convert_SLV_To_String(update_server_num_998) & " array_obj_ref_1020_wire = "& Convert_SLV_To_Hex_String(array_obj_ref_1020_wire));
          --
        end if; 
        if WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:WPIPE_NUMBER_OF_SERVERS_1018_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (3) : WPIPE_NUMBER_OF_SERVERS_1018_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1018_inst_req_0;
      WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1018_inst_req_1;
      WPIPE_NUMBER_OF_SERVERS_1018_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_server_num_998(0);
      data_in <= array_obj_ref_1020_wire;
      NUMBER_OF_SERVERS_write_3_gI: SplitGuardInterface generic map(name => "NUMBER_OF_SERVERS_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NUMBER_OF_SERVERS_write_3: OutputPortRevised -- 
        generic map ( name => "NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- logger for split-operator call_stmt_1087_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1087_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:call_stmt_1087_call:started:  Call to module UpdateRegister inputs: " & " rwbar_1033 (guard complement )= " & Convert_SLV_To_String(rwbar_1033) & " bmask_1037 = "& Convert_SLV_To_Hex_String(bmask_1037) & " rval_1080 = "& Convert_SLV_To_Hex_String(rval_1080) & " wdata_1045 = "& Convert_SLV_To_Hex_String(wdata_1045) & " index_1049 = "& Convert_SLV_To_Hex_String(index_1049));
          --
        end if; 
        if call_stmt_1087_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:SoftwareRegisterAccessDaemon:DP:call_stmt_1087_call:finished:  outputs: " & " wval_1087= "  & Convert_SLV_To_Hex_String(wval_1087));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1087_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1087_call_req_0;
      call_stmt_1087_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1087_call_req_1;
      call_stmt_1087_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_1033(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_1037 & rval_1080 & wdata_1045 & index_1049;
      wval_1087 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end SoftwareRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity UpdateRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    bmask : in  std_logic_vector(3 downto 0);
    rval : in  std_logic_vector(31 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    index : in  std_logic_vector(5 downto 0);
    wval : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity UpdateRegister;
architecture UpdateRegister_arch of UpdateRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 74)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal rval_buffer :  std_logic_vector(31 downto 0);
  signal rval_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(5 downto 0);
  signal index_update_enable: Boolean;
  -- output port buffer signals
  signal wval_buffer :  std_logic_vector(31 downto 0);
  signal wval_update_enable: Boolean;
  signal UpdateRegister_CP_34_start: Boolean;
  signal UpdateRegister_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u16_u32_181_inst_req_0 : boolean;
  signal CONCAT_u16_u32_181_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_181_inst_req_1 : boolean;
  signal CONCAT_u16_u32_181_inst_ack_1 : boolean;
  signal array_obj_ref_184_store_0_req_0 : boolean;
  signal array_obj_ref_184_store_0_ack_0 : boolean;
  signal array_obj_ref_184_store_0_req_1 : boolean;
  signal array_obj_ref_184_store_0_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "UpdateRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 74) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(3 downto 0) <= bmask;
  bmask_buffer <= in_buffer_data_out(3 downto 0);
  in_buffer_data_in(35 downto 4) <= rval;
  rval_buffer <= in_buffer_data_out(35 downto 4);
  in_buffer_data_in(67 downto 36) <= wdata;
  wdata_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(73 downto 68) <= index;
  index_buffer <= in_buffer_data_out(73 downto 68);
  in_buffer_data_in(tag_length + 73 downto 74) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 73 downto 74);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  UpdateRegister_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "UpdateRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wval_buffer;
  wval <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,UpdateRegister_CP_34_start,"UpdateRegister cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,UpdateRegister_CP_34_symbol, "UpdateRegister cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  UpdateRegister_CP_34: Block -- control-path 
    signal UpdateRegister_CP_34_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    UpdateRegister_CP_34_elements(0) <= UpdateRegister_CP_34_start;
    UpdateRegister_CP_34_symbol <= UpdateRegister_CP_34_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (39) 
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_word_addrgen/root_register_ack
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_sample_start_
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_update_start_
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Sample/rr
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Update/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Update/cr
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_update_start_
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_offset_calculated
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_resized_0
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_computed_0
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/word_access_complete/word_0/cr
      -- 
    -- logger for CP element group UpdateRegister_CP_34_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and UpdateRegister_CP_34_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:UpdateRegister_CP_34_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:CONCAT_u16_u32_181_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:CONCAT_u16_u32_181_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:array_obj_ref_184_store_0_req_1 fired."); 
        -- 
      end if; --
    end process; 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_181_inst_req_0); -- 
    cr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => CONCAT_u16_u32_181_inst_req_1); -- 
    cr_114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(0), ack => array_obj_ref_184_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_sample_completed_
      -- CP-element group 1: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Sample/ra
      -- 
    -- logger for CP element group UpdateRegister_CP_34_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and UpdateRegister_CP_34_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:UpdateRegister_CP_34_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:CONCAT_u16_u32_181_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_181_inst_ack_0, ack => UpdateRegister_CP_34_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_update_completed_
      -- CP-element group 2: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Update/$exit
      -- CP-element group 2: 	 assign_stmt_117_to_assign_stmt_186/CONCAT_u16_u32_181_Update/ca
      -- 
    -- logger for CP element group UpdateRegister_CP_34_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and UpdateRegister_CP_34_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:UpdateRegister_CP_34_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:CONCAT_u16_u32_181_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_181_inst_ack_1, ack => UpdateRegister_CP_34_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/array_obj_ref_184_Split/$entry
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/array_obj_ref_184_Split/$exit
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_sample_start_
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/array_obj_ref_184_Split/split_req
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/array_obj_ref_184_Split/split_ack
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/word_access_start/word_0/rr
      -- 
    -- logger for CP element group UpdateRegister_CP_34_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and UpdateRegister_CP_34_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:UpdateRegister_CP_34_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:array_obj_ref_184_store_0_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_34_elements(3), ack => array_obj_ref_184_store_0_req_0); -- 
    UpdateRegister_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "UpdateRegister_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= UpdateRegister_CP_34_elements(0) & UpdateRegister_CP_34_elements(2);
      gj_UpdateRegister_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => UpdateRegister_CP_34_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_sample_completed_
      -- CP-element group 4: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Sample/word_access_start/word_0/ra
      -- 
    -- logger for CP element group UpdateRegister_CP_34_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and UpdateRegister_CP_34_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:UpdateRegister_CP_34_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:array_obj_ref_184_store_0_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_184_store_0_ack_0, ack => UpdateRegister_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_117_to_assign_stmt_186/$exit
      -- CP-element group 5: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_update_completed_
      -- CP-element group 5: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/$exit
      -- CP-element group 5: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_117_to_assign_stmt_186/array_obj_ref_184_Update/word_access_complete/word_0/ca
      -- 
    -- logger for CP element group UpdateRegister_CP_34_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and UpdateRegister_CP_34_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:UpdateRegister_CP_34_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:UpdateRegister:CP:array_obj_ref_184_store_0_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_184_store_0_ack_1, ack => UpdateRegister_CP_34_elements(5)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_171_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_180_wire : std_logic_vector(15 downto 0);
    signal MUX_166_wire : std_logic_vector(7 downto 0);
    signal MUX_170_wire : std_logic_vector(7 downto 0);
    signal MUX_175_wire : std_logic_vector(7 downto 0);
    signal MUX_179_wire : std_logic_vector(7 downto 0);
    signal R_index_183_resized : std_logic_vector(5 downto 0);
    signal R_index_183_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_184_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_184_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_184_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_184_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_184_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_184_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_184_word_offset_0 : std_logic_vector(5 downto 0);
    signal b0_117 : std_logic_vector(0 downto 0);
    signal b1_121 : std_logic_vector(0 downto 0);
    signal b2_125 : std_logic_vector(0 downto 0);
    signal b3_129 : std_logic_vector(0 downto 0);
    signal r0_133 : std_logic_vector(7 downto 0);
    signal r1_137 : std_logic_vector(7 downto 0);
    signal r2_141 : std_logic_vector(7 downto 0);
    signal r3_145 : std_logic_vector(7 downto 0);
    signal w0_149 : std_logic_vector(7 downto 0);
    signal w1_153 : std_logic_vector(7 downto 0);
    signal w2_157 : std_logic_vector(7 downto 0);
    signal w3_161 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_184_offset_scale_factor_0 <= "000001";
    array_obj_ref_184_resized_base_address <= "000000";
    array_obj_ref_184_word_offset_0 <= "000000";
    -- logger for split-operator MUX_166_inst flow-through 
    process(MUX_166_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:MUX_166_inst:flowthrough inputs: " & " b0_117 = "& Convert_SLV_To_Hex_String(b0_117) & " w0_149 = "& Convert_SLV_To_Hex_String(w0_149) & " r0_133 = "& Convert_SLV_To_Hex_String(r0_133) & " outputs:" & " MUX_166_wire= "  & Convert_SLV_To_Hex_String(MUX_166_wire));
      --
    end process; 
    -- flow-through select operator MUX_166_inst
    MUX_166_wire <= w0_149 when (b0_117(0) /=  '0') else r0_133;
    -- logger for split-operator MUX_170_inst flow-through 
    process(MUX_170_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:MUX_170_inst:flowthrough inputs: " & " b1_121 = "& Convert_SLV_To_Hex_String(b1_121) & " w1_153 = "& Convert_SLV_To_Hex_String(w1_153) & " r1_137 = "& Convert_SLV_To_Hex_String(r1_137) & " outputs:" & " MUX_170_wire= "  & Convert_SLV_To_Hex_String(MUX_170_wire));
      --
    end process; 
    -- flow-through select operator MUX_170_inst
    MUX_170_wire <= w1_153 when (b1_121(0) /=  '0') else r1_137;
    -- logger for split-operator MUX_175_inst flow-through 
    process(MUX_175_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:MUX_175_inst:flowthrough inputs: " & " b2_125 = "& Convert_SLV_To_Hex_String(b2_125) & " w2_157 = "& Convert_SLV_To_Hex_String(w2_157) & " r2_141 = "& Convert_SLV_To_Hex_String(r2_141) & " outputs:" & " MUX_175_wire= "  & Convert_SLV_To_Hex_String(MUX_175_wire));
      --
    end process; 
    -- flow-through select operator MUX_175_inst
    MUX_175_wire <= w2_157 when (b2_125(0) /=  '0') else r2_141;
    -- logger for split-operator MUX_179_inst flow-through 
    process(MUX_179_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:MUX_179_inst:flowthrough inputs: " & " b3_129 = "& Convert_SLV_To_Hex_String(b3_129) & " w3_161 = "& Convert_SLV_To_Hex_String(w3_161) & " r3_145 = "& Convert_SLV_To_Hex_String(r3_145) & " outputs:" & " MUX_179_wire= "  & Convert_SLV_To_Hex_String(MUX_179_wire));
      --
    end process; 
    -- flow-through select operator MUX_179_inst
    MUX_179_wire <= w3_161 when (b3_129(0) /=  '0') else r3_145;
    -- logger for split-operator slice_116_inst flow-through 
    process(b0_117) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_116_inst:flowthrough inputs: " & " bmask_buffer = "& Convert_SLV_To_Hex_String(bmask_buffer) & " outputs:" & " b0_117= "  & Convert_SLV_To_Hex_String(b0_117));
      --
    end process; 
    -- flow-through slice operator slice_116_inst
    b0_117 <= bmask_buffer(3 downto 3);
    -- logger for split-operator slice_120_inst flow-through 
    process(b1_121) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_120_inst:flowthrough inputs: " & " bmask_buffer = "& Convert_SLV_To_Hex_String(bmask_buffer) & " outputs:" & " b1_121= "  & Convert_SLV_To_Hex_String(b1_121));
      --
    end process; 
    -- flow-through slice operator slice_120_inst
    b1_121 <= bmask_buffer(2 downto 2);
    -- logger for split-operator slice_124_inst flow-through 
    process(b2_125) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_124_inst:flowthrough inputs: " & " bmask_buffer = "& Convert_SLV_To_Hex_String(bmask_buffer) & " outputs:" & " b2_125= "  & Convert_SLV_To_Hex_String(b2_125));
      --
    end process; 
    -- flow-through slice operator slice_124_inst
    b2_125 <= bmask_buffer(1 downto 1);
    -- logger for split-operator slice_128_inst flow-through 
    process(b3_129) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_128_inst:flowthrough inputs: " & " bmask_buffer = "& Convert_SLV_To_Hex_String(bmask_buffer) & " outputs:" & " b3_129= "  & Convert_SLV_To_Hex_String(b3_129));
      --
    end process; 
    -- flow-through slice operator slice_128_inst
    b3_129 <= bmask_buffer(0 downto 0);
    -- logger for split-operator slice_132_inst flow-through 
    process(r0_133) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_132_inst:flowthrough inputs: " & " rval_buffer = "& Convert_SLV_To_Hex_String(rval_buffer) & " outputs:" & " r0_133= "  & Convert_SLV_To_Hex_String(r0_133));
      --
    end process; 
    -- flow-through slice operator slice_132_inst
    r0_133 <= rval_buffer(31 downto 24);
    -- logger for split-operator slice_136_inst flow-through 
    process(r1_137) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_136_inst:flowthrough inputs: " & " rval_buffer = "& Convert_SLV_To_Hex_String(rval_buffer) & " outputs:" & " r1_137= "  & Convert_SLV_To_Hex_String(r1_137));
      --
    end process; 
    -- flow-through slice operator slice_136_inst
    r1_137 <= rval_buffer(23 downto 16);
    -- logger for split-operator slice_140_inst flow-through 
    process(r2_141) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_140_inst:flowthrough inputs: " & " rval_buffer = "& Convert_SLV_To_Hex_String(rval_buffer) & " outputs:" & " r2_141= "  & Convert_SLV_To_Hex_String(r2_141));
      --
    end process; 
    -- flow-through slice operator slice_140_inst
    r2_141 <= rval_buffer(15 downto 8);
    -- logger for split-operator slice_144_inst flow-through 
    process(r3_145) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_144_inst:flowthrough inputs: " & " rval_buffer = "& Convert_SLV_To_Hex_String(rval_buffer) & " outputs:" & " r3_145= "  & Convert_SLV_To_Hex_String(r3_145));
      --
    end process; 
    -- flow-through slice operator slice_144_inst
    r3_145 <= rval_buffer(7 downto 0);
    -- logger for split-operator slice_148_inst flow-through 
    process(w0_149) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_148_inst:flowthrough inputs: " & " wdata_buffer = "& Convert_SLV_To_Hex_String(wdata_buffer) & " outputs:" & " w0_149= "  & Convert_SLV_To_Hex_String(w0_149));
      --
    end process; 
    -- flow-through slice operator slice_148_inst
    w0_149 <= wdata_buffer(31 downto 24);
    -- logger for split-operator slice_152_inst flow-through 
    process(w1_153) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_152_inst:flowthrough inputs: " & " wdata_buffer = "& Convert_SLV_To_Hex_String(wdata_buffer) & " outputs:" & " w1_153= "  & Convert_SLV_To_Hex_String(w1_153));
      --
    end process; 
    -- flow-through slice operator slice_152_inst
    w1_153 <= wdata_buffer(23 downto 16);
    -- logger for split-operator slice_156_inst flow-through 
    process(w2_157) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_156_inst:flowthrough inputs: " & " wdata_buffer = "& Convert_SLV_To_Hex_String(wdata_buffer) & " outputs:" & " w2_157= "  & Convert_SLV_To_Hex_String(w2_157));
      --
    end process; 
    -- flow-through slice operator slice_156_inst
    w2_157 <= wdata_buffer(15 downto 8);
    -- logger for split-operator slice_160_inst flow-through 
    process(w3_161) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:slice_160_inst:flowthrough inputs: " & " wdata_buffer = "& Convert_SLV_To_Hex_String(wdata_buffer) & " outputs:" & " w3_161= "  & Convert_SLV_To_Hex_String(w3_161));
      --
    end process; 
    -- flow-through slice operator slice_160_inst
    w3_161 <= wdata_buffer(7 downto 0);
    -- logger for operator array_obj_ref_184_addr_0 flow-through 
    process(array_obj_ref_184_word_address_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_addr_0:flowthrough  inputs: " & " array_obj_ref_184_root_address = "& Convert_SLV_To_Hex_String(array_obj_ref_184_root_address) & "outputs: " & " array_obj_ref_184_word_address_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_184_word_address_0));
      --
    end process; 
    -- equivalence array_obj_ref_184_addr_0
    process(array_obj_ref_184_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_184_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_184_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_184_gather_scatter flow-through 
    process(array_obj_ref_184_data_0) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_gather_scatter:flowthrough  inputs: " & " wval_buffer = "& Convert_SLV_To_Hex_String(wval_buffer) & "outputs: " & " array_obj_ref_184_data_0= "  & Convert_SLV_To_Hex_String(array_obj_ref_184_data_0));
      --
    end process; 
    -- equivalence array_obj_ref_184_gather_scatter
    process(wval_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := wval_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_184_data_0 <= ov(31 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_184_index_0_rename flow-through 
    process(R_index_183_scaled) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_index_0_rename:flowthrough  inputs: " & " R_index_183_resized = "& Convert_SLV_To_Hex_String(R_index_183_resized) & "outputs: " & " R_index_183_scaled= "  & Convert_SLV_To_Hex_String(R_index_183_scaled));
      --
    end process; 
    -- equivalence array_obj_ref_184_index_0_rename
    process(R_index_183_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_183_resized;
      ov(5 downto 0) := iv;
      R_index_183_scaled <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_184_index_0_resize flow-through 
    process(R_index_183_resized) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_index_0_resize:flowthrough  inputs: " & " index_buffer = "& Convert_SLV_To_Hex_String(index_buffer) & "outputs: " & " R_index_183_resized= "  & Convert_SLV_To_Hex_String(R_index_183_resized));
      --
    end process; 
    -- equivalence array_obj_ref_184_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(5 downto 0) := iv;
      R_index_183_resized <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_184_index_offset flow-through 
    process(array_obj_ref_184_final_offset) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_index_offset:flowthrough  inputs: " & " R_index_183_scaled = "& Convert_SLV_To_Hex_String(R_index_183_scaled) & "outputs: " & " array_obj_ref_184_final_offset= "  & Convert_SLV_To_Hex_String(array_obj_ref_184_final_offset));
      --
    end process; 
    -- equivalence array_obj_ref_184_index_offset
    process(R_index_183_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_183_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_184_final_offset <= ov(5 downto 0);
      --
    end process;
    -- logger for operator array_obj_ref_184_root_address_inst flow-through 
    process(array_obj_ref_184_root_address) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_root_address_inst:flowthrough  inputs: " & " array_obj_ref_184_final_offset = "& Convert_SLV_To_Hex_String(array_obj_ref_184_final_offset) & "outputs: " & " array_obj_ref_184_root_address= "  & Convert_SLV_To_Hex_String(array_obj_ref_184_root_address));
      --
    end process; 
    -- equivalence array_obj_ref_184_root_address_inst
    process(array_obj_ref_184_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_184_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_184_root_address <= ov(5 downto 0);
      --
    end process;
    -- logger for split-operator CONCAT_u16_u32_181_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u16_u32_181_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:CONCAT_u16_u32_181_inst:started:   inputs: " & " CONCAT_u8_u16_171_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_171_wire) & " CONCAT_u8_u16_180_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_180_wire));
          --
        end if; 
        if CONCAT_u16_u32_181_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:CONCAT_u16_u32_181_inst:finished:  outputs: " & " wval_buffer= "  & Convert_SLV_To_Hex_String(wval_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : CONCAT_u16_u32_181_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_171_wire & CONCAT_u8_u16_180_wire;
      wval_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_181_inst_req_0;
      CONCAT_u16_u32_181_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_181_inst_req_1;
      CONCAT_u16_u32_181_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator CONCAT_u8_u16_171_inst flow-through 
    process(CONCAT_u8_u16_171_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:CONCAT_u8_u16_171_inst:flowthrough inputs: " & " MUX_166_wire = "& Convert_SLV_To_Hex_String(MUX_166_wire) & " MUX_170_wire = "& Convert_SLV_To_Hex_String(MUX_170_wire) & " outputs:" & " CONCAT_u8_u16_171_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_171_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_171_inst
    process(MUX_166_wire, MUX_170_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_166_wire, MUX_170_wire, tmp_var);
      CONCAT_u8_u16_171_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u8_u16_180_inst flow-through 
    process(CONCAT_u8_u16_180_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:CONCAT_u8_u16_180_inst:flowthrough inputs: " & " MUX_175_wire = "& Convert_SLV_To_Hex_String(MUX_175_wire) & " MUX_179_wire = "& Convert_SLV_To_Hex_String(MUX_179_wire) & " outputs:" & " CONCAT_u8_u16_180_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_180_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_180_inst
    process(MUX_175_wire, MUX_179_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_175_wire, MUX_179_wire, tmp_var);
      CONCAT_u8_u16_180_wire <= tmp_var; --
    end process;
    -- logger for split-operator array_obj_ref_184_store_0
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if array_obj_ref_184_store_0_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_store_0:started:   inputs: " & " array_obj_ref_184_word_address_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_184_word_address_0) & " array_obj_ref_184_data_0 = "& Convert_SLV_To_Hex_String(array_obj_ref_184_data_0));
          --
        end if; 
        if array_obj_ref_184_store_0_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:UpdateRegister:DP:array_obj_ref_184_store_0:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      array_obj_ref_184_store_0_req_0,
      array_obj_ref_184_store_0_ack_0,
      array_obj_ref_184_store_0_req_1,
      array_obj_ref_184_store_0_ack_1,
      "array_obj_ref_184_store_0",
      "memory_space_0" ,
      array_obj_ref_184_data_0,
      array_obj_ref_184_word_address_0,
      "array_obj_ref_184_data_0",
      "array_obj_ref_184_word_address_0" -- 
    );
    -- shared store operator group (0) : array_obj_ref_184_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_184_store_0_req_0;
      array_obj_ref_184_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_184_store_0_req_1;
      array_obj_ref_184_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_184_word_address_0;
      data_in <= array_obj_ref_184_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(5 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end UpdateRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity accessMemory is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(7 downto 0);
    addr : in  std_logic_vector(35 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemory;
architecture accessMemory_arch of accessMemory is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 110)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(7 downto 0);
  signal bmask_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemory_CP_259_start: Boolean;
  signal accessMemory_CP_259_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemory_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 110) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(9 downto 2) <= bmask;
  bmask_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(45 downto 10) <= addr;
  addr_buffer <= in_buffer_data_out(45 downto 10);
  in_buffer_data_in(109 downto 46) <= wdata;
  wdata_buffer <= in_buffer_data_out(109 downto 46);
  in_buffer_data_in(tag_length + 109 downto 110) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 109 downto 110);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= lock_update_enable & rwbar_update_enable & bmask_update_enable & addr_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemory_CP_259_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemory_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_259_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemory_CP_259_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_259_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMemory_CP_259_start,"accessMemory cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,accessMemory_CP_259_symbol, "accessMemory cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemory_CP_259: Block -- control-path 
    signal accessMemory_CP_259_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    accessMemory_CP_259_elements(0) <= accessMemory_CP_259_start;
    accessMemory_CP_259_symbol <= accessMemory_CP_259_elements(22);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	8 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_259_to_assign_stmt_273/$entry
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(1) <= accessMemory_CP_259_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_259_to_assign_stmt_273/lock_update_enable
      -- CP-element group 2: 	 assign_stmt_259_to_assign_stmt_273/lock_update_enable_out
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_259_elements(9);
      gj_accessMemory_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	9 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	17 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_259_to_assign_stmt_273/rwbar_update_enable
      -- CP-element group 3: 	 assign_stmt_259_to_assign_stmt_273/rwbar_update_enable_out
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_259_elements(9);
      gj_accessMemory_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	9 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	18 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_259_to_assign_stmt_273/bmask_update_enable
      -- CP-element group 4: 	 assign_stmt_259_to_assign_stmt_273/bmask_update_enable_out
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_259_elements(9);
      gj_accessMemory_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	9 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_259_to_assign_stmt_273/addr_update_enable
      -- CP-element group 5: 	 assign_stmt_259_to_assign_stmt_273/addr_update_enable_out
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_259_elements(9);
      gj_accessMemory_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	20 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_259_to_assign_stmt_273/wdata_update_enable
      -- CP-element group 6: 	 assign_stmt_259_to_assign_stmt_273/wdata_update_enable_out
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessMemory_CP_259_elements(9);
      gj_accessMemory_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	21 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_259_to_assign_stmt_273/rdata_update_enable
      -- CP-element group 7: 	 assign_stmt_259_to_assign_stmt_273/rdata_update_enable_in
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(7) <= accessMemory_CP_259_elements(21);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_sample_start_
      -- CP-element group 8: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Sample/$entry
      -- CP-element group 8: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Sample/req
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_259_elements(8), ack => WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_0); -- 
    accessMemory_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessMemory_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_259_elements(1) & accessMemory_CP_259_elements(10);
      gj_accessMemory_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: 	3 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	5 
    -- CP-element group 9: 	6 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_sample_completed_
      -- CP-element group 9: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_update_start_
      -- CP-element group 9: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Sample/$exit
      -- CP-element group 9: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Sample/ack
      -- CP-element group 9: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Update/$entry
      -- CP-element group 9: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Update/req
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_0, ack => accessMemory_CP_259_elements(9)); -- 
    req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_259_elements(9), ack => WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_update_completed_
      -- CP-element group 10: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Update/$exit
      -- CP-element group 10: 	 assign_stmt_259_to_assign_stmt_273/WPIPE_NIC_TO_MEMORY_REQUEST_260_Update/ack
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_1, ack => accessMemory_CP_259_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_sample_start_
      -- CP-element group 11: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Sample/rr
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_259_elements(11), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_0); -- 
    accessMemory_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_259_elements(1) & accessMemory_CP_259_elements(14);
      gj_accessMemory_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	7 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_update_start_
      -- CP-element group 12: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Update/$entry
      -- CP-element group 12: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Update/cr
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_259_elements(12), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_1); -- 
    accessMemory_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_259_elements(13) & accessMemory_CP_259_elements(7);
      gj_accessMemory_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	12 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_sample_completed_
      -- CP-element group 13: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Sample/$exit
      -- CP-element group 13: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Sample/ra
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_0, ack => accessMemory_CP_259_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_update_completed_
      -- CP-element group 14: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Update/$exit
      -- CP-element group 14: 	 assign_stmt_259_to_assign_stmt_273/RPIPE_MEMORY_TO_NIC_RESPONSE_264_Update/ca
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_1, ack => accessMemory_CP_259_elements(14)); -- 
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 assign_stmt_259_to_assign_stmt_273/$exit
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_259_elements(14) & accessMemory_CP_259_elements(10);
      gj_accessMemory_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_259_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 lock_update_enable
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(16) <= accessMemory_CP_259_elements(2);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	3 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 rwbar_update_enable
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(17) <= accessMemory_CP_259_elements(3);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	4 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 bmask_update_enable
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(18) <= accessMemory_CP_259_elements(4);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 addr_update_enable
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(19) <= accessMemory_CP_259_elements(5);
    -- CP-element group 20:  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	6 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 wdata_update_enable
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(20) <= accessMemory_CP_259_elements(6);
    -- CP-element group 21:  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	7 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 rdata_update_enable
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 22:  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 $exit
      -- 
    -- logger for CP element group accessMemory_CP_259_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and accessMemory_CP_259_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:accessMemory:CP:accessMemory_CP_259_elements(22) fired."); 
        -- 
      end if; --
    end process; 
    accessMemory_CP_259_elements(22) <= accessMemory_CP_259_elements(15);
    --  hookup: inputs to control-path 
    accessMemory_CP_259_elements(21) <= rdata_update_enable;
    -- hookup: output from control-path 
    lock_update_enable <= accessMemory_CP_259_elements(16);
    rwbar_update_enable <= accessMemory_CP_259_elements(17);
    bmask_update_enable <= accessMemory_CP_259_elements(18);
    addr_update_enable <= accessMemory_CP_259_elements(19);
    wdata_update_enable <= accessMemory_CP_259_elements(20);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_252_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_254_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_257_wire : std_logic_vector(99 downto 0);
    signal err_269 : std_logic_vector(0 downto 0);
    signal request_259 : std_logic_vector(109 downto 0);
    signal response_265 : std_logic_vector(64 downto 0);
    -- 
  begin -- 
    -- logger for split-operator slice_268_inst flow-through 
    process(err_269) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:slice_268_inst:flowthrough inputs: " & " response_265 = "& Convert_SLV_To_Hex_String(response_265) & " outputs:" & " err_269= "  & Convert_SLV_To_Hex_String(err_269));
      --
    end process; 
    -- flow-through slice operator slice_268_inst
    err_269 <= response_265(64 downto 64);
    -- logger for split-operator slice_272_inst flow-through 
    process(rdata_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:slice_272_inst:flowthrough inputs: " & " response_265 = "& Convert_SLV_To_Hex_String(response_265) & " outputs:" & " rdata_buffer= "  & Convert_SLV_To_Hex_String(rdata_buffer));
      --
    end process; 
    -- flow-through slice operator slice_272_inst
    rdata_buffer <= response_265(63 downto 0);
    -- logger for split-operator CONCAT_u10_u110_258_inst flow-through 
    process(request_259) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:CONCAT_u10_u110_258_inst:flowthrough inputs: " & " CONCAT_u2_u10_254_wire = "& Convert_SLV_To_Hex_String(CONCAT_u2_u10_254_wire) & " CONCAT_u36_u100_257_wire = "& Convert_SLV_To_Hex_String(CONCAT_u36_u100_257_wire) & " outputs:" & " request_259= "  & Convert_SLV_To_Hex_String(request_259));
      --
    end process; 
    -- binary operator CONCAT_u10_u110_258_inst
    process(CONCAT_u2_u10_254_wire, CONCAT_u36_u100_257_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_254_wire, CONCAT_u36_u100_257_wire, tmp_var);
      request_259 <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u2_252_inst flow-through 
    process(CONCAT_u1_u2_252_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:CONCAT_u1_u2_252_inst:flowthrough inputs: " & " lock_buffer = "& Convert_SLV_To_Hex_String(lock_buffer) & " rwbar_buffer = "& Convert_SLV_To_Hex_String(rwbar_buffer) & " outputs:" & " CONCAT_u1_u2_252_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u2_252_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u2_252_inst
    process(lock_buffer, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(lock_buffer, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_252_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u2_u10_254_inst flow-through 
    process(CONCAT_u2_u10_254_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:CONCAT_u2_u10_254_inst:flowthrough inputs: " & " CONCAT_u1_u2_252_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u2_252_wire) & " bmask_buffer = "& Convert_SLV_To_Hex_String(bmask_buffer) & " outputs:" & " CONCAT_u2_u10_254_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u2_u10_254_wire));
      --
    end process; 
    -- binary operator CONCAT_u2_u10_254_inst
    process(CONCAT_u1_u2_252_wire, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_252_wire, bmask_buffer, tmp_var);
      CONCAT_u2_u10_254_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u36_u100_257_inst flow-through 
    process(CONCAT_u36_u100_257_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:CONCAT_u36_u100_257_inst:flowthrough inputs: " & " addr_buffer = "& Convert_SLV_To_Hex_String(addr_buffer) & " wdata_buffer = "& Convert_SLV_To_Hex_String(wdata_buffer) & " outputs:" & " CONCAT_u36_u100_257_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u36_u100_257_wire));
      --
    end process; 
    -- binary operator CONCAT_u36_u100_257_inst
    process(addr_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_buffer, wdata_buffer, tmp_var);
      CONCAT_u36_u100_257_wire <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst:started:   PipeRead from MEMORY_TO_NIC_RESPONSE inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst:finished:  outputs: " & " response_265= "  & Convert_SLV_To_Hex_String(response_265));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_0;
      RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_req_1;
      RPIPE_MEMORY_TO_NIC_RESPONSE_264_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_265 <= data_out(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE_read_0", data_width => 65,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_NIC_TO_MEMORY_REQUEST_260_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:WPIPE_NIC_TO_MEMORY_REQUEST_260_inst:started:   PipeWrite to NIC_TO_MEMORY_REQUEST inputs: " & " request_259 = "& Convert_SLV_To_Hex_String(request_259));
          --
        end if; 
        if WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:accessMemory:DP:WPIPE_NIC_TO_MEMORY_REQUEST_260_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_NIC_TO_MEMORY_REQUEST_260_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_0;
      WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_req_1;
      WPIPE_NIC_TO_MEMORY_REQUEST_260_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_259;
      NIC_TO_MEMORY_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_write_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemory_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity acquireMutex is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    m_ok : out  std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity acquireMutex;
architecture acquireMutex_arch of acquireMutex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal m_ok_buffer :  std_logic_vector(0 downto 0);
  signal acquireMutex_CP_311_start: Boolean;
  signal acquireMutex_CP_311_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_296_call_req_0 : boolean;
  signal call_stmt_296_call_ack_0 : boolean;
  signal call_stmt_296_call_req_1 : boolean;
  signal call_stmt_296_call_ack_1 : boolean;
  signal call_stmt_320_call_req_0 : boolean;
  signal call_stmt_320_call_ack_0 : boolean;
  signal call_stmt_320_call_req_1 : boolean;
  signal call_stmt_320_call_ack_1 : boolean;
  signal if_stmt_323_branch_req_0 : boolean;
  signal if_stmt_323_branch_ack_1 : boolean;
  signal if_stmt_323_branch_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "acquireMutex_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  acquireMutex_CP_311_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "acquireMutex_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  m_ok_buffer <= "1";
  out_buffer_data_in(0 downto 0) <= m_ok_buffer;
  m_ok <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireMutex_CP_311_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= acquireMutex_CP_311_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireMutex_CP_311_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,acquireMutex_CP_311_start,"acquireMutex cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,acquireMutex_CP_311_symbol, "acquireMutex cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  acquireMutex_CP_311: Block -- control-path 
    signal acquireMutex_CP_311_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    acquireMutex_CP_311_elements(0) <= acquireMutex_CP_311_start;
    acquireMutex_CP_311_symbol <= acquireMutex_CP_311_elements(6);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_278/$entry
      -- CP-element group 0: 	 branch_block_stmt_278/branch_block_stmt_278__entry__
      -- CP-element group 0: 	 branch_block_stmt_278/assign_stmt_281__entry__
      -- CP-element group 0: 	 branch_block_stmt_278/assign_stmt_281__exit__
      -- CP-element group 0: 	 branch_block_stmt_278/merge_stmt_283__entry__
      -- CP-element group 0: 	 branch_block_stmt_278/assign_stmt_281/$entry
      -- CP-element group 0: 	 branch_block_stmt_278/assign_stmt_281/$exit
      -- CP-element group 0: 	 branch_block_stmt_278/merge_stmt_283_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_278/merge_stmt_283__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_278/merge_stmt_283__entry___PhiReq/$exit
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	7 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Sample/cra
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_296_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_296_call_ack_0, ack => acquireMutex_CP_311_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Sample/crr
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_296_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_320_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_296_call_ack_1, ack => acquireMutex_CP_311_elements(2)); -- 
    crr_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_311_elements(2), ack => call_stmt_320_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Sample/cra
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_320_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_320_call_ack_0, ack => acquireMutex_CP_311_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	7 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320__exit__
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323__entry__
      -- CP-element group 4: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/NEQ_u32_u1_326_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/NEQ_u32_u1_326_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/NEQ_u32_u1_326/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_278/NEQ_u32_u1_326_place
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_278/if_stmt_323_else_link/$entry
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_320_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:if_stmt_323_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_320_call_ack_1, ack => acquireMutex_CP_311_elements(4)); -- 
    branch_req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_311_elements(4), ack => if_stmt_323_branch_req_0); -- 
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_278/if_stmt_323_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_278/if_stmt_323_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_278/loopback
      -- CP-element group 5: 	 branch_block_stmt_278/loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_278/loopback_PhiReq/$exit
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:if_stmt_323_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_323_branch_ack_1, ack => acquireMutex_CP_311_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (8) 
      -- CP-element group 6: 	 $exit
      -- CP-element group 6: 	 branch_block_stmt_278/$exit
      -- CP-element group 6: 	 branch_block_stmt_278/branch_block_stmt_278__exit__
      -- CP-element group 6: 	 branch_block_stmt_278/if_stmt_323__exit__
      -- CP-element group 6: 	 branch_block_stmt_278/if_stmt_323_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_278/if_stmt_323_else_link/else_choice_transition
      -- CP-element group 6: 	 assign_stmt_333/$entry
      -- CP-element group 6: 	 assign_stmt_333/$exit
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:if_stmt_323_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_323_branch_ack_0, ack => acquireMutex_CP_311_elements(6)); -- 
    -- CP-element group 7:  merge  fork  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	4 
    -- CP-element group 7:  members (16) 
      -- CP-element group 7: 	 branch_block_stmt_278/merge_stmt_283__exit__
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320__entry__
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/$entry
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_update_start_
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Sample/crr
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_296_Update/ccr
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_update_start_
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_278/call_stmt_296_to_call_stmt_320/call_stmt_320_Update/ccr
      -- CP-element group 7: 	 branch_block_stmt_278/merge_stmt_283_PhiReqMerge
      -- CP-element group 7: 	 branch_block_stmt_278/merge_stmt_283_PhiAck/$entry
      -- CP-element group 7: 	 branch_block_stmt_278/merge_stmt_283_PhiAck/$exit
      -- CP-element group 7: 	 branch_block_stmt_278/merge_stmt_283_PhiAck/dummy
      -- 
    -- logger for CP element group acquireMutex_CP_311_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and acquireMutex_CP_311_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:acquireMutex_CP_311_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_296_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_296_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:acquireMutex:CP:call_stmt_320_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_311_elements(7), ack => call_stmt_296_call_req_0); -- 
    ccr_345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_311_elements(7), ack => call_stmt_296_call_req_1); -- 
    ccr_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireMutex_CP_311_elements(7), ack => call_stmt_320_call_req_1); -- 
    acquireMutex_CP_311_elements(7) <= OrReduce(acquireMutex_CP_311_elements(5) & acquireMutex_CP_311_elements(0));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NEQ_u32_u1_326_wire : std_logic_vector(0 downto 0);
    signal NOT_u8_u8_291_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_316_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_320 : std_logic_vector(63 downto 0);
    signal konst_325_wire_constant : std_logic_vector(31 downto 0);
    signal mutex_address_281 : std_logic_vector(35 downto 0);
    signal mutex_plus_nentries_296 : std_logic_vector(63 downto 0);
    signal mutex_val_301 : std_logic_vector(31 downto 0);
    signal slice_306_wire : std_logic_vector(31 downto 0);
    signal type_cast_286_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_288_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_294_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_304_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_311_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_313_wire_constant : std_logic_vector(0 downto 0);
    signal wval_308 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_291_wire_constant <= "11111111";
    NOT_u8_u8_316_wire_constant <= "11111111";
    konst_325_wire_constant <= "00000000000000000000000000000000";
    type_cast_286_wire_constant <= "1";
    type_cast_288_wire_constant <= "1";
    type_cast_294_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_304_wire_constant <= "00000000000000000000000000000001";
    type_cast_311_wire_constant <= "0";
    type_cast_313_wire_constant <= "0";
    -- logger for split-operator slice_300_inst flow-through 
    process(mutex_val_301) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:slice_300_inst:flowthrough inputs: " & " mutex_plus_nentries_296 = "& Convert_SLV_To_Hex_String(mutex_plus_nentries_296) & " outputs:" & " mutex_val_301= "  & Convert_SLV_To_Hex_String(mutex_val_301));
      --
    end process; 
    -- flow-through slice operator slice_300_inst
    mutex_val_301 <= mutex_plus_nentries_296(63 downto 32);
    -- logger for split-operator slice_306_inst flow-through 
    process(slice_306_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:slice_306_inst:flowthrough inputs: " & " mutex_plus_nentries_296 = "& Convert_SLV_To_Hex_String(mutex_plus_nentries_296) & " outputs:" & " slice_306_wire= "  & Convert_SLV_To_Hex_String(slice_306_wire));
      --
    end process; 
    -- flow-through slice operator slice_306_inst
    slice_306_wire <= mutex_plus_nentries_296(31 downto 0);
    -- logger for split-operator W_mutex_address_279_inst flow-through 
    process(mutex_address_281) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:W_mutex_address_279_inst:flowthrough inputs: " & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " outputs:" & " mutex_address_281= "  & Convert_SLV_To_Hex_String(mutex_address_281));
      --
    end process; 
    -- interlock W_mutex_address_279_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 35 downto 0) := q_base_address_buffer(35 downto 0);
      mutex_address_281 <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_323_branch_req_0," req0 if_stmt_323_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_323_branch_ack_0," ack0 if_stmt_323_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_323_branch_ack_1," ack1 if_stmt_323_branch");
    if_stmt_323_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u32_u1_326_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_323_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_323_branch_req_0,
          ack0 => if_stmt_323_branch_ack_0,
          ack1 => if_stmt_323_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator CONCAT_u32_u64_307_inst flow-through 
    process(wval_308) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:CONCAT_u32_u64_307_inst:flowthrough inputs: " & " type_cast_304_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_304_wire_constant) & " slice_306_wire = "& Convert_SLV_To_Hex_String(slice_306_wire) & " outputs:" & " wval_308= "  & Convert_SLV_To_Hex_String(wval_308));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_307_inst
    process(type_cast_304_wire_constant, slice_306_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_304_wire_constant, slice_306_wire, tmp_var);
      wval_308 <= tmp_var; --
    end process;
    -- logger for split-operator NEQ_u32_u1_326_inst flow-through 
    process(NEQ_u32_u1_326_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:NEQ_u32_u1_326_inst:flowthrough inputs: " & " mutex_val_301 = "& Convert_SLV_To_Hex_String(mutex_val_301) & " konst_325_wire_constant = "& Convert_SLV_To_Hex_String(konst_325_wire_constant) & " outputs:" & " NEQ_u32_u1_326_wire= "  & Convert_SLV_To_Hex_String(NEQ_u32_u1_326_wire));
      --
    end process; 
    -- binary operator NEQ_u32_u1_326_inst
    process(mutex_val_301) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(mutex_val_301, konst_325_wire_constant, tmp_var);
      NEQ_u32_u1_326_wire <= tmp_var; --
    end process;
    -- logger for split-operator call_stmt_320_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_320_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:call_stmt_320_call:started:  Call to module accessMemory inputs: " & " type_cast_311_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_311_wire_constant) & " type_cast_313_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_313_wire_constant) & " NOT_u8_u8_316_wire_constant = "& Convert_SLV_To_Hex_String(NOT_u8_u8_316_wire_constant) & " mutex_address_281 = "& Convert_SLV_To_Hex_String(mutex_address_281) & " wval_308 = "& Convert_SLV_To_Hex_String(wval_308));
          --
        end if; 
        if call_stmt_320_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:call_stmt_320_call:finished:  outputs: " & " ignore_320= "  & Convert_SLV_To_Hex_String(ignore_320));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_296_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_296_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:call_stmt_296_call:started:  Call to module accessMemory inputs: " & " type_cast_286_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_286_wire_constant) & " type_cast_288_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_288_wire_constant) & " NOT_u8_u8_291_wire_constant = "& Convert_SLV_To_Hex_String(NOT_u8_u8_291_wire_constant) & " mutex_address_281 = "& Convert_SLV_To_Hex_String(mutex_address_281) & " type_cast_294_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_294_wire_constant));
          --
        end if; 
        if call_stmt_296_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:acquireMutex:DP:call_stmt_296_call:finished:  outputs: " & " mutex_plus_nentries_296= "  & Convert_SLV_To_Hex_String(mutex_plus_nentries_296));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_320_call call_stmt_296_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_320_call_req_0;
      reqL_unguarded(0) <= call_stmt_296_call_req_0;
      call_stmt_320_call_ack_0 <= ackL_unguarded(1);
      call_stmt_296_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_320_call_req_1;
      reqR_unguarded(0) <= call_stmt_296_call_req_1;
      call_stmt_320_call_ack_1 <= ackR_unguarded(1);
      call_stmt_296_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_311_wire_constant & type_cast_313_wire_constant & NOT_u8_u8_316_wire_constant & mutex_address_281 & wval_308 & type_cast_286_wire_constant & type_cast_288_wire_constant & NOT_u8_u8_291_wire_constant & mutex_address_281 & type_cast_294_wire_constant;
      ignore_320 <= data_out(127 downto 64);
      mutex_plus_nentries_296 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end acquireMutex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity delay_time_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    T : in  std_logic_vector(31 downto 0);
    delay_done : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity delay_time_Operator;
architecture delay_time_Operator_arch of delay_time_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal T_buffer :  std_logic_vector(31 downto 0);
  signal T_update_enable: Boolean;
  signal T_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal delay_done_buffer :  std_logic_vector(0 downto 0);
  signal delay_time_CP_1095_start: Boolean;
  signal delay_time_CP_1095_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_785_branch_req_0 : boolean;
  signal phi_stmt_787_req_1 : boolean;
  signal phi_stmt_787_req_0 : boolean;
  signal phi_stmt_787_ack_0 : boolean;
  signal T_789_buf_req_0 : boolean;
  signal T_789_buf_ack_0 : boolean;
  signal T_789_buf_req_1 : boolean;
  signal T_789_buf_ack_1 : boolean;
  signal nR_796_790_buf_req_0 : boolean;
  signal nR_796_790_buf_ack_0 : boolean;
  signal nR_796_790_buf_req_1 : boolean;
  signal nR_796_790_buf_ack_1 : boolean;
  signal do_while_stmt_785_branch_ack_0 : boolean;
  signal do_while_stmt_785_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  sample_ack <= delay_time_CP_1095_symbol;
  -- input handling ------------------------------------------------
  T_buffer <= T;
  delay_time_CP_1095_start <= sample_req;
  -- output handling  -------------------------------------------------------
  delay_done_buffer <= "1";
  delay_done <= delay_done_buffer;
  update_ack_symbol <= delay_time_CP_1095_symbol;
  update_ack <= update_ack_symbol;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,delay_time_CP_1095_start,"delay_time cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,delay_time_CP_1095_symbol, "delay_time cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  delay_time_CP_1095: Block -- control-path 
    signal delay_time_CP_1095_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    delay_time_CP_1095_elements(0) <= delay_time_CP_1095_start;
    delay_time_CP_1095_symbol <= delay_time_CP_1095_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_784/$entry
      -- CP-element group 0: 	 branch_block_stmt_784/branch_block_stmt_784__entry__
      -- CP-element group 0: 	 branch_block_stmt_784/do_while_stmt_785__entry__
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	32 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (8) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_784/$exit
      -- CP-element group 1: 	 branch_block_stmt_784/branch_block_stmt_784__exit__
      -- CP-element group 1: 	 branch_block_stmt_784/do_while_stmt_785__exit__
      -- CP-element group 1: 	 branch_block_stmt_784/assign_stmt_803__entry__
      -- CP-element group 1: 	 branch_block_stmt_784/assign_stmt_803__exit__
      -- CP-element group 1: 	 branch_block_stmt_784/assign_stmt_803/$entry
      -- CP-element group 1: 	 branch_block_stmt_784/assign_stmt_803/$exit
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(1) <= delay_time_CP_1095_elements(32);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_784/do_while_stmt_785/$entry
      -- CP-element group 2: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785__entry__
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(2) <= delay_time_CP_1095_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	32 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785__exit__
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group delay_time_CP_1095_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_784/do_while_stmt_785/loop_back
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group delay_time_CP_1095_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	31 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_784/do_while_stmt_785/condition_done
      -- CP-element group 5: 	 branch_block_stmt_784/do_while_stmt_785/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_784/do_while_stmt_785/loop_taken/$entry
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(5) <= delay_time_CP_1095_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	14 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_784/do_while_stmt_785/loop_body_done
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(6) <= delay_time_CP_1095_elements(14);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(7) <= delay_time_CP_1095_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(8) <= delay_time_CP_1095_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	29 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/loop_body_start
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group delay_time_CP_1095_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	29 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/condition_evaluated
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:do_while_stmt_785_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_1121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1095_elements(10), ack => do_while_stmt_785_branch_req_0); -- 
    delay_time_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1095_elements(29) & delay_time_CP_1095_elements(15);
      gj_delay_time_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1095_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_sample_start__ps
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1095_elements(12) & delay_time_CP_1095_elements(15);
      gj_delay_time_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1095_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_sample_start_
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1095_elements(9) & delay_time_CP_1095_elements(14);
      gj_delay_time_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1095_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_update_start_
      -- CP-element group 13: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_update_start__ps
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_1095_elements(9) & delay_time_CP_1095_elements(15);
      gj_delay_time_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_1095_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/$exit
      -- CP-element group 14: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_sample_completed__ps
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group delay_time_CP_1095_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_update_completed__ps
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group delay_time_CP_1095_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_loopback_trigger
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(16) <= delay_time_CP_1095_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_loopback_sample_req_ps
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:phi_stmt_787_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_787_loopback_sample_req_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_787_loopback_sample_req_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1095_elements(17), ack => phi_stmt_787_req_1); -- 
    -- Element group delay_time_CP_1095_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_entry_trigger
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(18) <= delay_time_CP_1095_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_entry_sample_req_ps
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:phi_stmt_787_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_787_entry_sample_req_1139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_787_entry_sample_req_1139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1095_elements(19), ack => phi_stmt_787_req_0); -- 
    -- Element group delay_time_CP_1095_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/phi_stmt_787_phi_mux_ack_ps
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:phi_stmt_787_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_787_phi_mux_ack_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_787_ack_0, ack => delay_time_CP_1095_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Sample/req
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:T_789_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1095_elements(21), ack => T_789_buf_req_0); -- 
    -- Element group delay_time_CP_1095_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_update_start_
      -- CP-element group 22: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Update/req
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:T_789_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1095_elements(22), ack => T_789_buf_req_1); -- 
    -- Element group delay_time_CP_1095_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_sample_completed__ps
      -- CP-element group 23: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Sample/ack
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:T_789_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_789_buf_ack_0, ack => delay_time_CP_1095_elements(23)); -- 
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_T_789_Update/ack
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:T_789_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_789_buf_ack_1, ack => delay_time_CP_1095_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Sample/req
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:nR_796_790_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_1173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1095_elements(25), ack => nR_796_790_buf_req_0); -- 
    -- Element group delay_time_CP_1095_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_update_start_
      -- CP-element group 26: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Update/req
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:nR_796_790_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_1095_elements(26), ack => nR_796_790_buf_req_1); -- 
    -- Element group delay_time_CP_1095_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Sample/ack
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:nR_796_790_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_796_790_buf_ack_0, ack => delay_time_CP_1095_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/R_nR_790_Update/ack
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:nR_796_790_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_796_790_buf_ack_1, ack => delay_time_CP_1095_elements(28)); -- 
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	9 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	10 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_784/do_while_stmt_785/do_while_stmt_785_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group delay_time_CP_1095_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => delay_time_CP_1095_elements(9), ack => delay_time_CP_1095_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_784/do_while_stmt_785/loop_exit/$exit
      -- CP-element group 30: 	 branch_block_stmt_784/do_while_stmt_785/loop_exit/ack
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:do_while_stmt_785_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_785_branch_ack_0, ack => delay_time_CP_1095_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_784/do_while_stmt_785/loop_taken/$exit
      -- CP-element group 31: 	 branch_block_stmt_784/do_while_stmt_785/loop_taken/ack
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:do_while_stmt_785_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_785_branch_ack_1, ack => delay_time_CP_1095_elements(31)); -- 
    -- CP-element group 32:  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	3 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	1 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_784/do_while_stmt_785/$exit
      -- 
    -- logger for CP element group delay_time_CP_1095_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and delay_time_CP_1095_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:delay_time:CP:delay_time_CP_1095_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    delay_time_CP_1095_elements(32) <= delay_time_CP_1095_elements(3);
    delay_time_do_while_stmt_785_terminator_1190: loop_terminator -- 
      generic map (name => " delay_time_do_while_stmt_785_terminator_1190", max_iterations_in_flight =>7) 
      port map(loop_body_exit => delay_time_CP_1095_elements(6),loop_continue => delay_time_CP_1095_elements(31),loop_terminate => delay_time_CP_1095_elements(30),loop_back => delay_time_CP_1095_elements(4),loop_exit => delay_time_CP_1095_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_787_phi_seq_1180_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= delay_time_CP_1095_elements(18);
      delay_time_CP_1095_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= delay_time_CP_1095_elements(23);
      delay_time_CP_1095_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= delay_time_CP_1095_elements(24);
      delay_time_CP_1095_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= delay_time_CP_1095_elements(16);
      delay_time_CP_1095_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= delay_time_CP_1095_elements(27);
      delay_time_CP_1095_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= delay_time_CP_1095_elements(28);
      delay_time_CP_1095_elements(17) <= phi_mux_reqs(1);
      phi_stmt_787_phi_seq_1180 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_787_phi_seq_1180") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => delay_time_CP_1095_elements(11), 
          phi_sample_ack => delay_time_CP_1095_elements(14), 
          phi_update_req => delay_time_CP_1095_elements(13), 
          phi_update_ack => delay_time_CP_1095_elements(15), 
          phi_mux_ack => delay_time_CP_1095_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1122_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= delay_time_CP_1095_elements(7);
        preds(1)  <= delay_time_CP_1095_elements(8);
        entry_tmerge_1122 : transition_merge -- 
          generic map(name => " entry_tmerge_1122")
          port map (preds => preds, symbol_out => delay_time_CP_1095_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_787 : std_logic_vector(31 downto 0);
    signal T_789_buffered : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_800_wire : std_logic_vector(0 downto 0);
    signal konst_794_wire_constant : std_logic_vector(31 downto 0);
    signal konst_799_wire_constant : std_logic_vector(31 downto 0);
    signal nR_796 : std_logic_vector(31 downto 0);
    signal nR_796_790_buffered : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_794_wire_constant <= "00000000000000000000000000000001";
    konst_799_wire_constant <= "00000000000000000000000000000000";
    -- logger for phi phi_stmt_787
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_787_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:delay_time:DP:phi_stmt_787:input-0 T_789_buffered= " & Convert_SLV_To_Hex_String(T_789_buffered));
          --
        end if;
        if phi_stmt_787_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:delay_time:DP:phi_stmt_787:input-1 nR_796_790_buffered= " & Convert_SLV_To_Hex_String(nR_796_790_buffered));
          --
        end if;
        if phi_stmt_787_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:delay_time:DP:phi_stmt_787:sample-completed");
          --
        end if;
        if phi_stmt_787_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:delay_time:DP:phi_stmt_787:output R_787= " & Convert_SLV_To_Hex_String(R_787));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_787: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= T_789_buffered & nR_796_790_buffered;
      req <= phi_stmt_787_req_0 & phi_stmt_787_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_787",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_787_ack_0,
          idata => idata,
          odata => R_787,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_787
    -- logger for split-operator T_789_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if T_789_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:delay_time:DP:T_789_buf:started:   inputs: " & " T_buffer = "& Convert_SLV_To_Hex_String(T_buffer));
          --
        end if; 
        if T_789_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:delay_time:DP:T_789_buf:finished:  outputs: " & " T_789_buffered= "  & Convert_SLV_To_Hex_String(T_789_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    T_789_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= T_789_buf_req_0;
      T_789_buf_ack_0<= wack(0);
      rreq(0) <= T_789_buf_req_1;
      T_789_buf_ack_1<= rack(0);
      T_789_buf : InterlockBuffer generic map ( -- 
        name => "T_789_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_789_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nR_796_790_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nR_796_790_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:delay_time:DP:nR_796_790_buf:started:   inputs: " & " nR_796 = "& Convert_SLV_To_Hex_String(nR_796));
          --
        end if; 
        if nR_796_790_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:delay_time:DP:nR_796_790_buf:finished:  outputs: " & " nR_796_790_buffered= "  & Convert_SLV_To_Hex_String(nR_796_790_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nR_796_790_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_796_790_buf_req_0;
      nR_796_790_buf_ack_0<= wack(0);
      rreq(0) <= nR_796_790_buf_req_1;
      nR_796_790_buf_ack_1<= rack(0);
      nR_796_790_buf : InterlockBuffer generic map ( -- 
        name => "nR_796_790_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_796_790_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_785_branch_req_0," req0 do_while_stmt_785_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_785_branch_ack_0," ack0 do_while_stmt_785_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_785_branch_ack_1," ack1 do_while_stmt_785_branch");
    do_while_stmt_785_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u32_u1_800_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_785_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_785_branch_req_0,
          ack0 => do_while_stmt_785_branch_ack_0,
          ack1 => do_while_stmt_785_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator SUB_u32_u32_795_inst flow-through 
    process(nR_796) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:delay_time:DP:SUB_u32_u32_795_inst:flowthrough inputs: " & " R_787 = "& Convert_SLV_To_Hex_String(R_787) & " konst_794_wire_constant = "& Convert_SLV_To_Hex_String(konst_794_wire_constant) & " outputs:" & " nR_796= "  & Convert_SLV_To_Hex_String(nR_796));
      --
    end process; 
    -- binary operator SUB_u32_u32_795_inst
    process(R_787) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_787, konst_794_wire_constant, tmp_var);
      nR_796 <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u32_u1_800_inst flow-through 
    process(UGT_u32_u1_800_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:delay_time:DP:UGT_u32_u1_800_inst:flowthrough inputs: " & " R_787 = "& Convert_SLV_To_Hex_String(R_787) & " konst_799_wire_constant = "& Convert_SLV_To_Hex_String(konst_799_wire_constant) & " outputs:" & " UGT_u32_u1_800_wire= "  & Convert_SLV_To_Hex_String(UGT_u32_u1_800_wire));
      --
    end process; 
    -- binary operator UGT_u32_u1_800_inst
    process(R_787) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(R_787, konst_799_wire_constant, tmp_var);
      UGT_u32_u1_800_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end delay_time_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity getQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    read_pointer : in  std_logic_vector(31 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueElement;
architecture getQueueElement_arch of getQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal read_pointer_buffer :  std_logic_vector(31 downto 0);
  signal read_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal getQueueElement_CP_436_start: Boolean;
  signal getQueueElement_CP_436_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal MUX_411_inst_ack_1 : boolean;
  signal call_stmt_396_call_req_1 : boolean;
  signal MUX_411_inst_req_1 : boolean;
  signal call_stmt_396_call_ack_1 : boolean;
  signal MUX_411_inst_ack_0 : boolean;
  signal MUX_411_inst_req_0 : boolean;
  signal call_stmt_396_call_ack_0 : boolean;
  signal call_stmt_396_call_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= read_pointer;
  read_pointer_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueElement_CP_436_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_436_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueElement_CP_436_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_436_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,getQueueElement_CP_436_start,"getQueueElement cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,getQueueElement_CP_436_symbol, "getQueueElement cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueElement_CP_436: Block -- control-path 
    signal getQueueElement_CP_436_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueElement_CP_436_elements(0) <= getQueueElement_CP_436_start;
    getQueueElement_CP_436_symbol <= getQueueElement_CP_436_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_update_start_
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_update_start_
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_sample_start_
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Update/ccr
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_complete/req
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_complete/$entry
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Update/$entry
      -- CP-element group 0: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Sample/crr
      -- 
    -- logger for CP element group getQueueElement_CP_436_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueueElement_CP_436_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:getQueueElement_CP_436_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:call_stmt_396_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:call_stmt_396_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:MUX_411_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_436_elements(0), ack => call_stmt_396_call_req_0); -- 
    ccr_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_436_elements(0), ack => call_stmt_396_call_req_1); -- 
    req_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_436_elements(0), ack => MUX_411_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_sample_completed_
      -- CP-element group 1: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Sample/cra
      -- 
    -- logger for CP element group getQueueElement_CP_436_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueueElement_CP_436_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:getQueueElement_CP_436_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:call_stmt_396_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_396_call_ack_0, ack => getQueueElement_CP_436_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_update_completed_
      -- CP-element group 2: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_start/$entry
      -- CP-element group 2: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_sample_start_
      -- CP-element group 2: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Update/cca
      -- CP-element group 2: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_start/req
      -- CP-element group 2: 	 assign_stmt_371_to_assign_stmt_412/call_stmt_396_Update/$exit
      -- 
    -- logger for CP element group getQueueElement_CP_436_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueueElement_CP_436_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:getQueueElement_CP_436_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:call_stmt_396_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:MUX_411_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_396_call_ack_1, ack => getQueueElement_CP_436_elements(2)); -- 
    req_463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_436_elements(2), ack => MUX_411_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_sample_completed_
      -- CP-element group 3: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_start/ack
      -- CP-element group 3: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_start/$exit
      -- 
    -- logger for CP element group getQueueElement_CP_436_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueueElement_CP_436_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:getQueueElement_CP_436_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:MUX_411_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_411_inst_ack_0, ack => getQueueElement_CP_436_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_complete/ack
      -- CP-element group 4: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_update_completed_
      -- CP-element group 4: 	 assign_stmt_371_to_assign_stmt_412/MUX_411_complete/$exit
      -- CP-element group 4: 	 assign_stmt_371_to_assign_stmt_412/$exit
      -- CP-element group 4: 	 $exit
      -- 
    -- logger for CP element group getQueueElement_CP_436_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueueElement_CP_436_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:getQueueElement_CP_436_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueueElement:CP:MUX_411_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_411_inst_ack_1, ack => getQueueElement_CP_436_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_408_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_380_wire : std_logic_vector(33 downto 0);
    signal NOT_u8_u8_391_wire_constant : std_logic_vector(7 downto 0);
    signal buffer_address_371 : std_logic_vector(35 downto 0);
    signal e0_400 : std_logic_vector(31 downto 0);
    signal e1_404 : std_logic_vector(31 downto 0);
    signal element_pair_396 : std_logic_vector(63 downto 0);
    signal element_pair_address_384 : std_logic_vector(35 downto 0);
    signal konst_407_wire_constant : std_logic_vector(31 downto 0);
    signal slice_376_wire : std_logic_vector(30 downto 0);
    signal type_cast_369_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_379_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_382_wire : std_logic_vector(35 downto 0);
    signal type_cast_386_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_388_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_394_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_391_wire_constant <= "11111111";
    konst_407_wire_constant <= "00000000000000000000000000000000";
    type_cast_369_wire_constant <= "000000000000000000000000000000010000";
    type_cast_379_wire_constant <= "000";
    type_cast_386_wire_constant <= "0";
    type_cast_388_wire_constant <= "1";
    type_cast_394_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- logger for split-operator MUX_411_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_411_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:MUX_411_inst:started:   inputs: " & " BITSEL_u32_u1_408_wire = "& Convert_SLV_To_Hex_String(BITSEL_u32_u1_408_wire) & " e1_404 = "& Convert_SLV_To_Hex_String(e1_404) & " e0_400 = "& Convert_SLV_To_Hex_String(e0_400));
          --
        end if; 
        if MUX_411_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:MUX_411_inst:finished:  outputs: " & " q_r_data_buffer= "  & Convert_SLV_To_Hex_String(q_r_data_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_411_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_411_inst_req_0;
      MUX_411_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_411_inst_req_1;
      MUX_411_inst_ack_1<= update_ack(0);
      MUX_411_inst: SelectSplitProtocol generic map(name => "MUX_411_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => e1_404, y => e0_400, sel => BITSEL_u32_u1_408_wire, z => q_r_data_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_376_inst flow-through 
    process(slice_376_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:slice_376_inst:flowthrough inputs: " & " read_pointer_buffer = "& Convert_SLV_To_Hex_String(read_pointer_buffer) & " outputs:" & " slice_376_wire= "  & Convert_SLV_To_Hex_String(slice_376_wire));
      --
    end process; 
    -- flow-through slice operator slice_376_inst
    slice_376_wire <= read_pointer_buffer(31 downto 1);
    -- logger for split-operator slice_399_inst flow-through 
    process(e0_400) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:slice_399_inst:flowthrough inputs: " & " element_pair_396 = "& Convert_SLV_To_Hex_String(element_pair_396) & " outputs:" & " e0_400= "  & Convert_SLV_To_Hex_String(e0_400));
      --
    end process; 
    -- flow-through slice operator slice_399_inst
    e0_400 <= element_pair_396(63 downto 32);
    -- logger for split-operator slice_403_inst flow-through 
    process(e1_404) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:slice_403_inst:flowthrough inputs: " & " element_pair_396 = "& Convert_SLV_To_Hex_String(element_pair_396) & " outputs:" & " e1_404= "  & Convert_SLV_To_Hex_String(e1_404));
      --
    end process; 
    -- flow-through slice operator slice_403_inst
    e1_404 <= element_pair_396(31 downto 0);
    -- logger for split-operator type_cast_382_inst flow-through 
    process(type_cast_382_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:type_cast_382_inst:flowthrough inputs: " & " CONCAT_u31_u34_380_wire = "& Convert_SLV_To_Hex_String(CONCAT_u31_u34_380_wire) & " outputs:" & " type_cast_382_wire= "  & Convert_SLV_To_Hex_String(type_cast_382_wire));
      --
    end process; 
    -- interlock type_cast_382_inst
    process(CONCAT_u31_u34_380_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_380_wire(33 downto 0);
      type_cast_382_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ADD_u36_u36_370_inst flow-through 
    process(buffer_address_371) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:ADD_u36_u36_370_inst:flowthrough inputs: " & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " type_cast_369_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_369_wire_constant) & " outputs:" & " buffer_address_371= "  & Convert_SLV_To_Hex_String(buffer_address_371));
      --
    end process; 
    -- binary operator ADD_u36_u36_370_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_369_wire_constant, tmp_var);
      buffer_address_371 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u36_u36_383_inst flow-through 
    process(element_pair_address_384) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:ADD_u36_u36_383_inst:flowthrough inputs: " & " buffer_address_371 = "& Convert_SLV_To_Hex_String(buffer_address_371) & " type_cast_382_wire = "& Convert_SLV_To_Hex_String(type_cast_382_wire) & " outputs:" & " element_pair_address_384= "  & Convert_SLV_To_Hex_String(element_pair_address_384));
      --
    end process; 
    -- binary operator ADD_u36_u36_383_inst
    process(buffer_address_371, type_cast_382_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_371, type_cast_382_wire, tmp_var);
      element_pair_address_384 <= tmp_var; --
    end process;
    -- logger for split-operator BITSEL_u32_u1_408_inst flow-through 
    process(BITSEL_u32_u1_408_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:BITSEL_u32_u1_408_inst:flowthrough inputs: " & " read_pointer_buffer = "& Convert_SLV_To_Hex_String(read_pointer_buffer) & " konst_407_wire_constant = "& Convert_SLV_To_Hex_String(konst_407_wire_constant) & " outputs:" & " BITSEL_u32_u1_408_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u32_u1_408_wire));
      --
    end process; 
    -- binary operator BITSEL_u32_u1_408_inst
    process(read_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(read_pointer_buffer, konst_407_wire_constant, tmp_var);
      BITSEL_u32_u1_408_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u31_u34_380_inst flow-through 
    process(CONCAT_u31_u34_380_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:CONCAT_u31_u34_380_inst:flowthrough inputs: " & " slice_376_wire = "& Convert_SLV_To_Hex_String(slice_376_wire) & " type_cast_379_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_379_wire_constant) & " outputs:" & " CONCAT_u31_u34_380_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u31_u34_380_wire));
      --
    end process; 
    -- binary operator CONCAT_u31_u34_380_inst
    process(slice_376_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_376_wire, type_cast_379_wire_constant, tmp_var);
      CONCAT_u31_u34_380_wire <= tmp_var; --
    end process;
    -- logger for split-operator call_stmt_396_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_396_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:call_stmt_396_call:started:  Call to module accessMemory inputs: " & " type_cast_386_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_386_wire_constant) & " type_cast_388_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_388_wire_constant) & " NOT_u8_u8_391_wire_constant = "& Convert_SLV_To_Hex_String(NOT_u8_u8_391_wire_constant) & " element_pair_address_384 = "& Convert_SLV_To_Hex_String(element_pair_address_384) & " type_cast_394_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_394_wire_constant));
          --
        end if; 
        if call_stmt_396_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getQueueElement:DP:call_stmt_396_call:finished:  outputs: " & " element_pair_396= "  & Convert_SLV_To_Hex_String(element_pair_396));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_396_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_396_call_req_0;
      call_stmt_396_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_396_call_req_1;
      call_stmt_396_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_386_wire_constant & type_cast_388_wire_constant & NOT_u8_u8_391_wire_constant & element_pair_address_384 & type_cast_394_wire_constant;
      element_pair_396 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity getQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : out  std_logic_vector(31 downto 0);
    rp : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointers;
architecture getQueuePointers_arch of getQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  signal getQueuePointers_CP_416_start: Boolean;
  signal getQueuePointers_CP_416_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_352_call_ack_1 : boolean;
  signal call_stmt_352_call_req_1 : boolean;
  signal call_stmt_352_call_req_0 : boolean;
  signal call_stmt_352_call_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointers_CP_416_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wp_buffer;
  wp <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= rp_buffer;
  rp <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_416_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointers_CP_416_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_416_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,getQueuePointers_CP_416_start,"getQueuePointers cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,getQueuePointers_CP_416_symbol, "getQueuePointers cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointers_CP_416: Block -- control-path 
    signal getQueuePointers_CP_416_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    getQueuePointers_CP_416_elements(0) <= getQueuePointers_CP_416_start;
    getQueuePointers_CP_416_symbol <= getQueuePointers_CP_416_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Update/ccr
      -- CP-element group 0: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Update/$entry
      -- CP-element group 0: 	 call_stmt_352_to_assign_stmt_360/$entry
      -- CP-element group 0: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Sample/crr
      -- CP-element group 0: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_update_start_
      -- CP-element group 0: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_sample_start_
      -- 
    -- logger for CP element group getQueuePointers_CP_416_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueuePointers_CP_416_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueuePointers:CP:getQueuePointers_CP_416_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueuePointers:CP:call_stmt_352_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueuePointers:CP:call_stmt_352_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_416_elements(0), ack => call_stmt_352_call_req_0); -- 
    ccr_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_416_elements(0), ack => call_stmt_352_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Sample/$exit
      -- CP-element group 1: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Sample/cra
      -- CP-element group 1: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_sample_completed_
      -- 
    -- logger for CP element group getQueuePointers_CP_416_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueuePointers_CP_416_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueuePointers:CP:getQueuePointers_CP_416_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueuePointers:CP:call_stmt_352_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_352_call_ack_0, ack => getQueuePointers_CP_416_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Update/cca
      -- CP-element group 2: 	 call_stmt_352_to_assign_stmt_360/$exit
      -- CP-element group 2: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_Update/$exit
      -- CP-element group 2: 	 call_stmt_352_to_assign_stmt_360/call_stmt_352_update_completed_
      -- CP-element group 2: 	 $exit
      -- 
    -- logger for CP element group getQueuePointers_CP_416_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getQueuePointers_CP_416_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueuePointers:CP:getQueuePointers_CP_416_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getQueuePointers:CP:call_stmt_352_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_352_call_ack_1, ack => getQueuePointers_CP_416_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_348_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_345_wire_constant : std_logic_vector(7 downto 0);
    signal konst_347_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_340_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_342_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(63 downto 0);
    signal wp_rp_352 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_345_wire_constant <= "11111111";
    konst_347_wire_constant <= "000000000000000000000000000000001000";
    type_cast_340_wire_constant <= "0";
    type_cast_342_wire_constant <= "1";
    type_cast_350_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- logger for split-operator slice_355_inst flow-through 
    process(wp_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueuePointers:DP:slice_355_inst:flowthrough inputs: " & " wp_rp_352 = "& Convert_SLV_To_Hex_String(wp_rp_352) & " outputs:" & " wp_buffer= "  & Convert_SLV_To_Hex_String(wp_buffer));
      --
    end process; 
    -- flow-through slice operator slice_355_inst
    wp_buffer <= wp_rp_352(63 downto 32);
    -- logger for split-operator slice_359_inst flow-through 
    process(rp_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueuePointers:DP:slice_359_inst:flowthrough inputs: " & " wp_rp_352 = "& Convert_SLV_To_Hex_String(wp_rp_352) & " outputs:" & " rp_buffer= "  & Convert_SLV_To_Hex_String(rp_buffer));
      --
    end process; 
    -- flow-through slice operator slice_359_inst
    rp_buffer <= wp_rp_352(31 downto 0);
    -- logger for split-operator ADD_u36_u36_348_inst flow-through 
    process(ADD_u36_u36_348_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getQueuePointers:DP:ADD_u36_u36_348_inst:flowthrough inputs: " & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " konst_347_wire_constant = "& Convert_SLV_To_Hex_String(konst_347_wire_constant) & " outputs:" & " ADD_u36_u36_348_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_348_wire));
      --
    end process; 
    -- binary operator ADD_u36_u36_348_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_347_wire_constant, tmp_var);
      ADD_u36_u36_348_wire <= tmp_var; --
    end process;
    -- logger for split-operator call_stmt_352_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_352_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getQueuePointers:DP:call_stmt_352_call:started:  Call to module accessMemory inputs: " & " type_cast_340_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_340_wire_constant) & " type_cast_342_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_342_wire_constant) & " NOT_u8_u8_345_wire_constant = "& Convert_SLV_To_Hex_String(NOT_u8_u8_345_wire_constant) & " ADD_u36_u36_348_wire = "& Convert_SLV_To_Hex_String(ADD_u36_u36_348_wire) & " type_cast_350_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_350_wire_constant));
          --
        end if; 
        if call_stmt_352_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getQueuePointers:DP:call_stmt_352_call:finished:  outputs: " & " wp_rp_352= "  & Convert_SLV_To_Hex_String(wp_rp_352));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_352_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_352_call_req_0;
      call_stmt_352_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_352_call_req_1;
      call_stmt_352_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_340_wire_constant & type_cast_342_wire_constant & NOT_u8_u8_345_wire_constant & ADD_u36_u36_348_wire & type_cast_350_wire_constant;
      wp_rp_352 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity getTxPacketPointerFromServer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_index : in  std_logic_vector(5 downto 0);
    pkt_pointer : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTxPacketPointerFromServer;
architecture getTxPacketPointerFromServer_arch of getTxPacketPointerFromServer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 6)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_index_buffer :  std_logic_vector(5 downto 0);
  signal queue_index_update_enable: Boolean;
  -- output port buffer signals
  signal pkt_pointer_buffer :  std_logic_vector(31 downto 0);
  signal pkt_pointer_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal getTxPacketPointerFromServer_CP_2107_start: Boolean;
  signal getTxPacketPointerFromServer_CP_2107_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1126_call_req_0 : boolean;
  signal call_stmt_1126_call_ack_0 : boolean;
  signal call_stmt_1126_call_req_1 : boolean;
  signal call_stmt_1126_call_ack_1 : boolean;
  signal call_stmt_1138_call_req_0 : boolean;
  signal call_stmt_1138_call_ack_0 : boolean;
  signal call_stmt_1138_call_req_1 : boolean;
  signal call_stmt_1138_call_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 6) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= queue_index;
  queue_index_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(tag_length + 5 downto 6) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 5 downto 6);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 7);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= queue_index_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTxPacketPointerFromServer_CP_2107_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= pkt_pointer_buffer;
  pkt_pointer <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2107_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  pkt_pointer_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "pkt_pointer_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_pkt_pointer_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => pkt_pointer_update_enable, clk => clk, reset => reset); --
  end block;
  status_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "status_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_status_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => status_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2107_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_2107_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,getTxPacketPointerFromServer_CP_2107_start,"getTxPacketPointerFromServer cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,getTxPacketPointerFromServer_CP_2107_symbol, "getTxPacketPointerFromServer cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTxPacketPointerFromServer_CP_2107: Block -- control-path 
    signal getTxPacketPointerFromServer_CP_2107_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    getTxPacketPointerFromServer_CP_2107_elements(0) <= getTxPacketPointerFromServer_CP_2107_start;
    getTxPacketPointerFromServer_CP_2107_symbol <= getTxPacketPointerFromServer_CP_2107_elements(16);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_1117_to_call_stmt_1138/$entry
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    getTxPacketPointerFromServer_CP_2107_elements(1) <= getTxPacketPointerFromServer_CP_2107_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_1117_to_call_stmt_1138/queue_index_update_enable
      -- CP-element group 2: 	 assign_stmt_1117_to_call_stmt_1138/queue_index_update_enable_out
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    getTxPacketPointerFromServer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_2107_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2107_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	14 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_1117_to_call_stmt_1138/pkt_pointer_update_enable
      -- CP-element group 3: 	 assign_stmt_1117_to_call_stmt_1138/pkt_pointer_update_enable_in
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    getTxPacketPointerFromServer_CP_2107_elements(3) <= getTxPacketPointerFromServer_CP_2107_elements(14);
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_1117_to_call_stmt_1138/status_update_enable
      -- CP-element group 4: 	 assign_stmt_1117_to_call_stmt_1138/status_update_enable_in
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    getTxPacketPointerFromServer_CP_2107_elements(4) <= getTxPacketPointerFromServer_CP_2107_elements(15);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_sample_start_
      -- CP-element group 5: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Sample/crr
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1126_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2107_elements(5), ack => call_stmt_1126_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2107_elements(1) & getTxPacketPointerFromServer_CP_2107_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2107_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	11 
    -- CP-element group 6: 	8 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_update_start_
      -- CP-element group 6: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Update/$entry
      -- CP-element group 6: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Update/ccr
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1126_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_2131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2107_elements(6), ack => call_stmt_1126_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2107_elements(11) & getTxPacketPointerFromServer_CP_2107_elements(8);
      gj_getTxPacketPointerFromServer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2107_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_sample_completed_
      -- CP-element group 7: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Sample/cra
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1126_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1126_call_ack_0, ack => getTxPacketPointerFromServer_CP_2107_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_update_completed_
      -- CP-element group 8: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Update/$exit
      -- CP-element group 8: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1126_Update/cca
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1126_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1126_call_ack_1, ack => getTxPacketPointerFromServer_CP_2107_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_sample_start_
      -- CP-element group 9: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Sample/crr
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1138_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2107_elements(9), ack => call_stmt_1138_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2107_elements(8) & getTxPacketPointerFromServer_CP_2107_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2107_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_update_start_
      -- CP-element group 10: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Update/$entry
      -- CP-element group 10: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Update/ccr
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1138_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_2145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_2107_elements(10), ack => call_stmt_1138_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "getTxPacketPointerFromServer_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_2107_elements(3) & getTxPacketPointerFromServer_CP_2107_elements(4) & getTxPacketPointerFromServer_CP_2107_elements(12);
      gj_getTxPacketPointerFromServer_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_2107_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_sample_completed_
      -- CP-element group 11: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Sample/cra
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1138_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1138_call_ack_0, ack => getTxPacketPointerFromServer_CP_2107_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 assign_stmt_1117_to_call_stmt_1138/$exit
      -- CP-element group 12: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_update_completed_
      -- CP-element group 12: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Update/$exit
      -- CP-element group 12: 	 assign_stmt_1117_to_call_stmt_1138/call_stmt_1138_Update/cca
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:call_stmt_1138_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1138_call_ack_1, ack => getTxPacketPointerFromServer_CP_2107_elements(12)); -- 
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 queue_index_update_enable
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    getTxPacketPointerFromServer_CP_2107_elements(13) <= getTxPacketPointerFromServer_CP_2107_elements(2);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 pkt_pointer_update_enable
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 status_update_enable
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 16:  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 $exit
      -- 
    -- logger for CP element group getTxPacketPointerFromServer_CP_2107_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and getTxPacketPointerFromServer_CP_2107_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:getTxPacketPointerFromServer:CP:getTxPacketPointerFromServer_CP_2107_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    getTxPacketPointerFromServer_CP_2107_elements(16) <= getTxPacketPointerFromServer_CP_2107_elements(12);
    --  hookup: inputs to control-path 
    getTxPacketPointerFromServer_CP_2107_elements(14) <= pkt_pointer_update_enable;
    getTxPacketPointerFromServer_CP_2107_elements(15) <= status_update_enable;
    -- hookup: output from control-path 
    queue_index_update_enable <= getTxPacketPointerFromServer_CP_2107_elements(13);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1115_wire : std_logic_vector(5 downto 0);
    signal R_TX_QUEUES_REG_START_OFFSET_1114_wire_constant : std_logic_vector(5 downto 0);
    signal register_index_1117 : std_logic_vector(5 downto 0);
    signal tx_queue_pointer_32_1126 : std_logic_vector(31 downto 0);
    signal tx_queue_pointer_36_1132 : std_logic_vector(35 downto 0);
    signal type_cast_1119_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1121_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1124_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1130_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1134_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_TX_QUEUES_REG_START_OFFSET_1114_wire_constant <= "001010";
    type_cast_1119_wire_constant <= "1";
    type_cast_1121_wire_constant <= "0001";
    type_cast_1124_wire_constant <= "00000000000000000000000000000000";
    type_cast_1130_wire_constant <= "0000";
    type_cast_1134_wire_constant <= "0";
    -- logger for split-operator type_cast_1116_inst flow-through 
    process(register_index_1117) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getTxPacketPointerFromServer:DP:type_cast_1116_inst:flowthrough inputs: " & " ADD_u6_u6_1115_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_1115_wire) & " outputs:" & " register_index_1117= "  & Convert_SLV_To_Hex_String(register_index_1117));
      --
    end process; 
    -- interlock type_cast_1116_inst
    process(ADD_u6_u6_1115_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1115_wire(5 downto 0);
      register_index_1117 <= tmp_var; -- 
    end process;
    -- logger for split-operator ADD_u6_u6_1115_inst flow-through 
    process(ADD_u6_u6_1115_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getTxPacketPointerFromServer:DP:ADD_u6_u6_1115_inst:flowthrough inputs: " & " queue_index_buffer = "& Convert_SLV_To_Hex_String(queue_index_buffer) & " R_TX_QUEUES_REG_START_OFFSET_1114_wire_constant = "& Convert_SLV_To_Hex_String(R_TX_QUEUES_REG_START_OFFSET_1114_wire_constant) & " outputs:" & " ADD_u6_u6_1115_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_1115_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_1115_inst
    process(queue_index_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(queue_index_buffer, R_TX_QUEUES_REG_START_OFFSET_1114_wire_constant, tmp_var);
      ADD_u6_u6_1115_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u36_1131_inst flow-through 
    process(tx_queue_pointer_36_1132) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:getTxPacketPointerFromServer:DP:CONCAT_u32_u36_1131_inst:flowthrough inputs: " & " tx_queue_pointer_32_1126 = "& Convert_SLV_To_Hex_String(tx_queue_pointer_32_1126) & " type_cast_1130_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1130_wire_constant) & " outputs:" & " tx_queue_pointer_36_1132= "  & Convert_SLV_To_Hex_String(tx_queue_pointer_36_1132));
      --
    end process; 
    -- binary operator CONCAT_u32_u36_1131_inst
    process(tx_queue_pointer_32_1126) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(tx_queue_pointer_32_1126, type_cast_1130_wire_constant, tmp_var);
      tx_queue_pointer_36_1132 <= tmp_var; --
    end process;
    -- logger for split-operator call_stmt_1126_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1126_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getTxPacketPointerFromServer:DP:call_stmt_1126_call:started:  Call to module AccessRegister inputs: " & " type_cast_1119_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1119_wire_constant) & " type_cast_1121_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1121_wire_constant) & " register_index_1117 = "& Convert_SLV_To_Hex_String(register_index_1117) & " type_cast_1124_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1124_wire_constant));
          --
        end if; 
        if call_stmt_1126_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getTxPacketPointerFromServer:DP:call_stmt_1126_call:finished:  outputs: " & " tx_queue_pointer_32_1126= "  & Convert_SLV_To_Hex_String(tx_queue_pointer_32_1126));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1126_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1126_call_req_0;
      call_stmt_1126_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1126_call_req_1;
      call_stmt_1126_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1119_wire_constant & type_cast_1121_wire_constant & register_index_1117 & type_cast_1124_wire_constant;
      tx_queue_pointer_32_1126 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_1138_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1138_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getTxPacketPointerFromServer:DP:call_stmt_1138_call:started:  Call to module popFromQueue inputs: " & " type_cast_1134_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1134_wire_constant) & " tx_queue_pointer_36_1132 = "& Convert_SLV_To_Hex_String(tx_queue_pointer_36_1132));
          --
        end if; 
        if call_stmt_1138_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:getTxPacketPointerFromServer:DP:call_stmt_1138_call:finished:  outputs: " & " pkt_pointer_buffer= "  & Convert_SLV_To_Hex_String(pkt_pointer_buffer) & " status_buffer= "  & Convert_SLV_To_Hex_String(status_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_1138_call 
    popFromQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1138_call_req_0;
      call_stmt_1138_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1138_call_req_1;
      call_stmt_1138_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_1_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1134_wire_constant & tx_queue_pointer_36_1132;
      pkt_pointer_buffer <= data_out(32 downto 1);
      status_buffer <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getTxPacketPointerFromServer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadBuffer is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
    writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
    writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
    writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadBuffer;
architecture loadBuffer_arch of loadBuffer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal loadBuffer_CP_925_start: Boolean;
  signal loadBuffer_CP_925_symbol: Boolean;
  -- volatile/operator module components. 
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_672_call_req_1 : boolean;
  signal call_stmt_667_call_req_0 : boolean;
  signal call_stmt_667_call_ack_0 : boolean;
  signal call_stmt_661_call_req_0 : boolean;
  signal call_stmt_667_call_req_1 : boolean;
  signal call_stmt_661_call_ack_0 : boolean;
  signal call_stmt_672_call_ack_0 : boolean;
  signal call_stmt_667_call_ack_1 : boolean;
  signal call_stmt_672_call_ack_1 : boolean;
  signal call_stmt_672_call_req_0 : boolean;
  signal call_stmt_661_call_ack_1 : boolean;
  signal call_stmt_661_call_req_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadBuffer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 31);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_buffer_pointer_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadBuffer_CP_925_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadBuffer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_925_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  bad_packet_identifier_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 40) := "bad_packet_identifier_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_bad_packet_identifier_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => bad_packet_identifier_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 31,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadBuffer_CP_925_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_925_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,loadBuffer_CP_925_start,"loadBuffer cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,loadBuffer_CP_925_symbol, "loadBuffer cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadBuffer_CP_925: Block -- control-path 
    signal loadBuffer_CP_925_elements: BooleanArray(18 downto 0);
    -- 
  begin -- 
    loadBuffer_CP_925_elements(0) <= loadBuffer_CP_925_start;
    loadBuffer_CP_925_symbol <= loadBuffer_CP_925_elements(18);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	8 
    -- CP-element group 1: 	12 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_661_to_call_stmt_672/$entry
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    loadBuffer_CP_925_elements(1) <= loadBuffer_CP_925_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	14 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_661_to_call_stmt_672/rx_buffer_pointer_update_enable
      -- CP-element group 2: 	 call_stmt_661_to_call_stmt_672/rx_buffer_pointer_update_enable_out
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    loadBuffer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_925_elements(6) & loadBuffer_CP_925_elements(10) & loadBuffer_CP_925_elements(14);
      gj_loadBuffer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_925_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	17 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	9 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_661_to_call_stmt_672/bad_packet_identifier_update_enable_in
      -- CP-element group 3: 	 call_stmt_661_to_call_stmt_672/bad_packet_identifier_update_enable
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    loadBuffer_CP_925_elements(3) <= loadBuffer_CP_925_elements(17);
    -- CP-element group 4:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Sample/crr
      -- CP-element group 4: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_sample_start_
      -- CP-element group 4: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Sample/$entry
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_661_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_925_elements(4), ack => call_stmt_661_call_req_0); -- 
    loadBuffer_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_925_elements(1) & loadBuffer_CP_925_elements(6) & loadBuffer_CP_925_elements(15);
      gj_loadBuffer_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_925_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: 	10 
    -- CP-element group 5: 	15 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_update_start_
      -- CP-element group 5: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Update/ccr
      -- CP-element group 5: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Update/$entry
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_661_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_925_elements(5), ack => call_stmt_661_call_req_1); -- 
    loadBuffer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_925_elements(7) & loadBuffer_CP_925_elements(10) & loadBuffer_CP_925_elements(15);
      gj_loadBuffer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_925_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: marked-successors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: 	4 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Sample/$exit
      -- CP-element group 6: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Sample/cra
      -- CP-element group 6: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_sample_completed_
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_661_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_661_call_ack_0, ack => loadBuffer_CP_925_elements(6)); -- 
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_update_completed_
      -- CP-element group 7: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Update/cca
      -- CP-element group 7: 	 call_stmt_661_to_call_stmt_672/call_stmt_661_Update/$exit
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_661_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_661_call_ack_1, ack => loadBuffer_CP_925_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: 	7 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Sample/$entry
      -- CP-element group 8: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Sample/crr
      -- CP-element group 8: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_sample_start_
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_667_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_925_elements(8), ack => call_stmt_667_call_req_0); -- 
    loadBuffer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_925_elements(1) & loadBuffer_CP_925_elements(7) & loadBuffer_CP_925_elements(10);
      gj_loadBuffer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_925_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	3 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_update_start_
      -- CP-element group 9: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Update/$entry
      -- CP-element group 9: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Update/ccr
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_667_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_925_elements(9), ack => call_stmt_667_call_req_1); -- 
    loadBuffer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_925_elements(3) & loadBuffer_CP_925_elements(11) & loadBuffer_CP_925_elements(14);
      gj_loadBuffer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_925_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: 	5 
    -- CP-element group 10: 	8 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_sample_completed_
      -- CP-element group 10: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Sample/$exit
      -- CP-element group 10: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Sample/cra
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_667_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_667_call_ack_0, ack => loadBuffer_CP_925_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Update/$exit
      -- CP-element group 11: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_update_completed_
      -- CP-element group 11: 	 call_stmt_661_to_call_stmt_672/call_stmt_667_Update/cca
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_667_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_667_call_ack_1, ack => loadBuffer_CP_925_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	1 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_sample_start_
      -- CP-element group 12: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Sample/crr
      -- CP-element group 12: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Sample/$entry
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_672_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_925_elements(12), ack => call_stmt_672_call_req_0); -- 
    loadBuffer_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_925_elements(1) & loadBuffer_CP_925_elements(11) & loadBuffer_CP_925_elements(14);
      gj_loadBuffer_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_925_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Update/ccr
      -- CP-element group 13: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Update/$entry
      -- CP-element group 13: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_update_start_
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_672_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_925_elements(13), ack => call_stmt_672_call_req_1); -- 
    loadBuffer_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadBuffer_CP_925_elements(15);
      gj_loadBuffer_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_925_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_sample_completed_
      -- CP-element group 14: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Sample/cra
      -- CP-element group 14: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Sample/$exit
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_672_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_672_call_ack_0, ack => loadBuffer_CP_925_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	5 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (4) 
      -- CP-element group 15: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Update/$exit
      -- CP-element group 15: 	 call_stmt_661_to_call_stmt_672/$exit
      -- CP-element group 15: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_Update/cca
      -- CP-element group 15: 	 call_stmt_661_to_call_stmt_672/call_stmt_672_update_completed_
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:call_stmt_672_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_672_call_ack_1, ack => loadBuffer_CP_925_elements(15)); -- 
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 rx_buffer_pointer_update_enable
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    loadBuffer_CP_925_elements(16) <= loadBuffer_CP_925_elements(2);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	3 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 bad_packet_identifier_update_enable
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 18:  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 $exit
      -- 
    -- logger for CP element group loadBuffer_CP_925_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and loadBuffer_CP_925_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:loadBuffer:CP:loadBuffer_CP_925_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    loadBuffer_CP_925_elements(18) <= loadBuffer_CP_925_elements(15);
    --  hookup: inputs to control-path 
    loadBuffer_CP_925_elements(17) <= bad_packet_identifier_update_enable;
    -- hookup: output from control-path 
    rx_buffer_pointer_update_enable <= loadBuffer_CP_925_elements(16);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal last_keep_667 : std_logic_vector(7 downto 0);
    signal new_buf_pointer_661 : std_logic_vector(35 downto 0);
    signal packet_size_667 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    -- logger for split-operator call_stmt_661_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_661_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadBuffer:DP:call_stmt_661_call:started:  Call to module writeEthernetHeaderToMem inputs: " & " rx_buffer_pointer_buffer = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_buffer));
          --
        end if; 
        if call_stmt_661_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadBuffer:DP:call_stmt_661_call:finished:  outputs: " & " new_buf_pointer_661= "  & Convert_SLV_To_Hex_String(new_buf_pointer_661));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_661_call 
    writeEthernetHeaderToMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_661_call_req_0;
      call_stmt_661_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_661_call_req_1;
      call_stmt_661_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeEthernetHeaderToMem_call_group_0_gI: SplitGuardInterface generic map(name => "writeEthernetHeaderToMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer;
      new_buf_pointer_661 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeEthernetHeaderToMem_call_reqs(0),
          ackR => writeEthernetHeaderToMem_call_acks(0),
          dataR => writeEthernetHeaderToMem_call_data(35 downto 0),
          tagR => writeEthernetHeaderToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeEthernetHeaderToMem_return_acks(0), -- cross-over
          ackL => writeEthernetHeaderToMem_return_reqs(0), -- cross-over
          dataL => writeEthernetHeaderToMem_return_data(35 downto 0),
          tagL => writeEthernetHeaderToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_667_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_667_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadBuffer:DP:call_stmt_667_call:started:  Call to module writePayloadToMem inputs: " & " rx_buffer_pointer_buffer = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_buffer) & " new_buf_pointer_661 = "& Convert_SLV_To_Hex_String(new_buf_pointer_661));
          --
        end if; 
        if call_stmt_667_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadBuffer:DP:call_stmt_667_call:finished:  outputs: " & " packet_size_667= "  & Convert_SLV_To_Hex_String(packet_size_667) & " bad_packet_identifier_buffer= "  & Convert_SLV_To_Hex_String(bad_packet_identifier_buffer) & " last_keep_667= "  & Convert_SLV_To_Hex_String(last_keep_667));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_667_call 
    writePayloadToMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(16 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_667_call_req_0;
      call_stmt_667_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_667_call_req_1;
      call_stmt_667_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writePayloadToMem_call_group_1_gI: SplitGuardInterface generic map(name => "writePayloadToMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer & new_buf_pointer_661;
      packet_size_667 <= data_out(16 downto 9);
      bad_packet_identifier_buffer <= data_out(8 downto 8);
      last_keep_667 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writePayloadToMem_call_reqs(0),
          ackR => writePayloadToMem_call_acks(0),
          dataR => writePayloadToMem_call_data(71 downto 0),
          tagR => writePayloadToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 17,
          owidth => 17,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writePayloadToMem_return_acks(0), -- cross-over
          ackL => writePayloadToMem_return_reqs(0), -- cross-over
          dataL => writePayloadToMem_return_data(16 downto 0),
          tagL => writePayloadToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_672_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_672_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadBuffer:DP:call_stmt_672_call:started:  Call to module writeControlInformationToMem inputs: " & " bad_packet_identifier_buffer (guard complement )= " & Convert_SLV_To_String(bad_packet_identifier_buffer) & " rx_buffer_pointer_buffer = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_buffer) & " packet_size_667 = "& Convert_SLV_To_Hex_String(packet_size_667) & " last_keep_667 = "& Convert_SLV_To_Hex_String(last_keep_667));
          --
        end if; 
        if call_stmt_672_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:loadBuffer:DP:call_stmt_672_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_672_call 
    writeControlInformationToMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(51 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_672_call_req_0;
      call_stmt_672_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_672_call_req_1;
      call_stmt_672_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not bad_packet_identifier_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeControlInformationToMem_call_group_2_gI: SplitGuardInterface generic map(name => "writeControlInformationToMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer & packet_size_667 & last_keep_667;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 52,
        owidth => 52,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeControlInformationToMem_call_reqs(0),
          ackR => writeControlInformationToMem_call_acks(0),
          dataR => writeControlInformationToMem_call_data(51 downto 0),
          tagR => writeControlInformationToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeControlInformationToMem_return_acks(0), -- cross-over
          ackL => writeControlInformationToMem_return_reqs(0), -- cross-over
          tagL => writeControlInformationToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end loadBuffer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity macToNicInterface is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_0_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_0_pipe_read_data : in   std_logic_vector(63 downto 0);
    mac_to_nic_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_1_pipe_read_data : in   std_logic_vector(15 downto 0);
    mac_to_nic_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_data : out  std_logic_vector(72 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity macToNicInterface;
architecture macToNicInterface_arch of macToNicInterface is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal macToNicInterface_CP_2153_start: Boolean;
  signal macToNicInterface_CP_2153_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1145_branch_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_0_1149_inst_req_0 : boolean;
  signal WPIPE_mac_to_nic_data_1157_inst_ack_1 : boolean;
  signal do_while_stmt_1145_branch_ack_1 : boolean;
  signal RPIPE_mac_to_nic_data_0_1149_inst_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_0_1149_inst_req_1 : boolean;
  signal do_while_stmt_1145_branch_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_0_1149_inst_ack_1 : boolean;
  signal RPIPE_mac_to_nic_data_1_1152_inst_ack_1 : boolean;
  signal RPIPE_mac_to_nic_data_1_1152_inst_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_1_1152_inst_ack_0 : boolean;
  signal WPIPE_mac_to_nic_data_1157_inst_req_1 : boolean;
  signal WPIPE_mac_to_nic_data_1157_inst_ack_0 : boolean;
  signal CONCAT_u9_u73_1162_inst_ack_1 : boolean;
  signal CONCAT_u9_u73_1162_inst_req_1 : boolean;
  signal CONCAT_u9_u73_1162_inst_ack_0 : boolean;
  signal CONCAT_u9_u73_1162_inst_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_1_1152_inst_req_1 : boolean;
  signal WPIPE_mac_to_nic_data_1157_inst_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "macToNicInterface_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  macToNicInterface_CP_2153_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "macToNicInterface_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= macToNicInterface_CP_2153_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= macToNicInterface_CP_2153_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= macToNicInterface_CP_2153_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,macToNicInterface_CP_2153_start,"macToNicInterface cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,macToNicInterface_CP_2153_symbol, "macToNicInterface cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  macToNicInterface_CP_2153: Block -- control-path 
    signal macToNicInterface_CP_2153_elements: BooleanArray(35 downto 0);
    -- 
  begin -- 
    macToNicInterface_CP_2153_elements(0) <= macToNicInterface_CP_2153_start;
    macToNicInterface_CP_2153_symbol <= macToNicInterface_CP_2153_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1144/do_while_stmt_1145__entry__
      -- CP-element group 0: 	 branch_block_stmt_1144/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1144/branch_block_stmt_1144__entry__
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	34 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1144/branch_block_stmt_1144__exit__
      -- CP-element group 1: 	 branch_block_stmt_1144/do_while_stmt_1145__exit__
      -- CP-element group 1: 	 branch_block_stmt_1144/$exit
      -- CP-element group 1: 	 $exit
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_CP_2153_elements(1) <= macToNicInterface_CP_2153_elements(34);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145__entry__
      -- CP-element group 2: 	 branch_block_stmt_1144/do_while_stmt_1145/$entry
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_CP_2153_elements(2) <= macToNicInterface_CP_2153_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	34 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145__exit__
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group macToNicInterface_CP_2153_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_back
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group macToNicInterface_CP_2153_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	32 
    -- CP-element group 5: 	33 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1144/do_while_stmt_1145/condition_done
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_CP_2153_elements(5) <= macToNicInterface_CP_2153_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	35 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_body_done
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_CP_2153_elements(6) <= macToNicInterface_CP_2153_elements(35);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_CP_2153_elements(7) <= macToNicInterface_CP_2153_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_CP_2153_elements(8) <= macToNicInterface_CP_2153_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	19 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1147_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1150_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/$entry
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group macToNicInterface_CP_2153_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	31 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/condition_evaluated
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:do_while_stmt_1145_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(10), ack => do_while_stmt_1145_branch_req_0); -- 
    macToNicInterface_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(31) & macToNicInterface_CP_2153_elements(13);
      gj_macToNicInterface_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	20 
    -- CP-element group 11: 	15 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(9) & macToNicInterface_CP_2153_elements(13);
      gj_macToNicInterface_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	21 
    -- CP-element group 12: 	16 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(19) & macToNicInterface_CP_2153_elements(14);
      gj_macToNicInterface_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	23 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(18) & macToNicInterface_CP_2153_elements(23);
      gj_macToNicInterface_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	26 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1147_update_start_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(9) & macToNicInterface_CP_2153_elements(26);
      gj_macToNicInterface_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_sample_start_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_0_1149_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(15), ack => RPIPE_mac_to_nic_data_0_1149_inst_req_0); -- 
    macToNicInterface_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(11) & macToNicInterface_CP_2153_elements(18);
      gj_macToNicInterface_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: 	17 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_update_start_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_0_1149_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(16), ack => RPIPE_mac_to_nic_data_0_1149_inst_req_1); -- 
    macToNicInterface_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(12) & macToNicInterface_CP_2153_elements(17);
      gj_macToNicInterface_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: 	35 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_sample_completed_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_0_1149_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_0_1149_inst_ack_0, ack => macToNicInterface_CP_2153_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	13 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_0_1149_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1147_update_completed_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_0_1149_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_0_1149_inst_ack_1, ack => macToNicInterface_CP_2153_elements(18)); -- 
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	9 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	26 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1150_update_start_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(9) & macToNicInterface_CP_2153_elements(26);
      gj_macToNicInterface_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	11 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_sample_start_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_1_1152_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(20), ack => RPIPE_mac_to_nic_data_1_1152_inst_req_0); -- 
    macToNicInterface_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(11) & macToNicInterface_CP_2153_elements(23);
      gj_macToNicInterface_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	12 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Update/$entry
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_1_1152_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(21), ack => RPIPE_mac_to_nic_data_1_1152_inst_req_1); -- 
    macToNicInterface_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(22) & macToNicInterface_CP_2153_elements(12);
      gj_macToNicInterface_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	35 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Sample/ra
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_1_1152_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1_1152_inst_ack_0, ack => macToNicInterface_CP_2153_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	13 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1150_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/RPIPE_mac_to_nic_data_1_1152_Update/$exit
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:RPIPE_mac_to_nic_data_1_1152_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1_1152_inst_ack_1, ack => macToNicInterface_CP_2153_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_sample_start_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:CONCAT_u9_u73_1162_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(24), ack => CONCAT_u9_u73_1162_inst_req_0); -- 
    macToNicInterface_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(18) & macToNicInterface_CP_2153_elements(23) & macToNicInterface_CP_2153_elements(26);
      gj_macToNicInterface_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_update_start_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:CONCAT_u9_u73_1162_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(25), ack => CONCAT_u9_u73_1162_inst_req_1); -- 
    macToNicInterface_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= macToNicInterface_CP_2153_elements(29);
      gj_macToNicInterface_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	19 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	14 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_sample_completed_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:CONCAT_u9_u73_1162_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u9_u73_1162_inst_ack_0, ack => macToNicInterface_CP_2153_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/CONCAT_u9_u73_1162_update_completed_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:CONCAT_u9_u73_1162_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u9_u73_1162_inst_ack_1, ack => macToNicInterface_CP_2153_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Sample/$entry
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:WPIPE_mac_to_nic_data_1157_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(28), ack => WPIPE_mac_to_nic_data_1157_inst_req_0); -- 
    macToNicInterface_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(27) & macToNicInterface_CP_2153_elements(30);
      gj_macToNicInterface_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Sample/$exit
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:WPIPE_mac_to_nic_data_1157_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:WPIPE_mac_to_nic_data_1157_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mac_to_nic_data_1157_inst_ack_0, ack => macToNicInterface_CP_2153_elements(29)); -- 
    req_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => macToNicInterface_CP_2153_elements(29), ack => WPIPE_mac_to_nic_data_1157_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Update/ack
      -- CP-element group 30: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/WPIPE_mac_to_nic_data_1157_update_completed_
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:WPIPE_mac_to_nic_data_1157_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mac_to_nic_data_1157_inst_ack_1, ack => macToNicInterface_CP_2153_elements(30)); -- 
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	10 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group macToNicInterface_CP_2153_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => macToNicInterface_CP_2153_elements(9), ack => macToNicInterface_CP_2153_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	5 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_exit/$exit
      -- CP-element group 32: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_exit/ack
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:do_while_stmt_1145_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1145_branch_ack_0, ack => macToNicInterface_CP_2153_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	5 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_taken/$exit
      -- CP-element group 33: 	 branch_block_stmt_1144/do_while_stmt_1145/loop_taken/ack
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:do_while_stmt_1145_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1145_branch_ack_1, ack => macToNicInterface_CP_2153_elements(33)); -- 
    -- CP-element group 34:  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	3 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	1 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1144/do_while_stmt_1145/$exit
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_CP_2153_elements(34) <= macToNicInterface_CP_2153_elements(3);
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	22 
    -- CP-element group 35: 	30 
    -- CP-element group 35: 	17 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	6 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/aggregated_phi_sample_ack
      -- CP-element group 35: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1150_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/phi_stmt_1147_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1144/do_while_stmt_1145/do_while_stmt_1145_loop_body/$exit
      -- 
    -- logger for CP element group macToNicInterface_CP_2153_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and macToNicInterface_CP_2153_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:macToNicInterface:CP:macToNicInterface_CP_2153_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    macToNicInterface_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "macToNicInterface_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= macToNicInterface_CP_2153_elements(22) & macToNicInterface_CP_2153_elements(30) & macToNicInterface_CP_2153_elements(17);
      gj_macToNicInterface_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => macToNicInterface_CP_2153_elements(35), clk => clk, reset => reset); --
    end block;
    macToNicInterface_do_while_stmt_1145_terminator_2256: loop_terminator -- 
      generic map (name => " macToNicInterface_do_while_stmt_1145_terminator_2256", max_iterations_in_flight =>7) 
      port map(loop_body_exit => macToNicInterface_CP_2153_elements(6),loop_continue => macToNicInterface_CP_2153_elements(33),loop_terminate => macToNicInterface_CP_2153_elements(32),loop_back => macToNicInterface_CP_2153_elements(4),loop_exit => macToNicInterface_CP_2153_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_2178_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= macToNicInterface_CP_2153_elements(7);
        preds(1)  <= macToNicInterface_CP_2153_elements(8);
        entry_tmerge_2178 : transition_merge -- 
          generic map(name => " entry_tmerge_2178")
          port map (preds => preds, symbol_out => macToNicInterface_CP_2153_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u9_u73_1162_wire : std_logic_vector(72 downto 0);
    signal RPIPE_mac_to_nic_data_0_1149_wire : std_logic_vector(63 downto 0);
    signal RPIPE_mac_to_nic_data_1_1152_wire : std_logic_vector(15 downto 0);
    signal konst_1165_wire_constant : std_logic_vector(0 downto 0);
    signal rdata0_1147 : std_logic_vector(63 downto 0);
    signal rdata1_1150 : std_logic_vector(15 downto 0);
    signal slice_1160_wire : std_logic_vector(8 downto 0);
    -- 
  begin -- 
    konst_1165_wire_constant <= "1";
    -- logger for split-operator slice_1160_inst flow-through 
    process(slice_1160_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:slice_1160_inst:flowthrough inputs: " & " rdata1_1150 = "& Convert_SLV_To_Hex_String(rdata1_1150) & " outputs:" & " slice_1160_wire= "  & Convert_SLV_To_Hex_String(slice_1160_wire));
      --
    end process; 
    -- flow-through slice operator slice_1160_inst
    slice_1160_wire <= rdata1_1150(8 downto 0);
    -- logger for split-operator ssrc_phi_stmt_1147 flow-through 
    process(rdata0_1147) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:ssrc_phi_stmt_1147:flowthrough inputs: " & " RPIPE_mac_to_nic_data_0_1149_wire = "& Convert_SLV_To_Hex_String(RPIPE_mac_to_nic_data_0_1149_wire) & " outputs:" & " rdata0_1147= "  & Convert_SLV_To_Hex_String(rdata0_1147));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1147
    process(RPIPE_mac_to_nic_data_0_1149_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := RPIPE_mac_to_nic_data_0_1149_wire(63 downto 0);
      rdata0_1147 <= tmp_var; -- 
    end process;
    -- logger for split-operator ssrc_phi_stmt_1150 flow-through 
    process(rdata1_1150) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:ssrc_phi_stmt_1150:flowthrough inputs: " & " RPIPE_mac_to_nic_data_1_1152_wire = "& Convert_SLV_To_Hex_String(RPIPE_mac_to_nic_data_1_1152_wire) & " outputs:" & " rdata1_1150= "  & Convert_SLV_To_Hex_String(rdata1_1150));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1150
    process(RPIPE_mac_to_nic_data_1_1152_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := RPIPE_mac_to_nic_data_1_1152_wire(15 downto 0);
      rdata1_1150 <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1145_branch_req_0," req0 do_while_stmt_1145_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1145_branch_ack_0," ack0 do_while_stmt_1145_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1145_branch_ack_1," ack1 do_while_stmt_1145_branch");
    do_while_stmt_1145_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1165_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1145_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1145_branch_req_0,
          ack0 => do_while_stmt_1145_branch_ack_0,
          ack1 => do_while_stmt_1145_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator CONCAT_u9_u73_1162_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u9_u73_1162_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:CONCAT_u9_u73_1162_inst:started:   inputs: " & " slice_1160_wire = "& Convert_SLV_To_Hex_String(slice_1160_wire) & " rdata0_1147 = "& Convert_SLV_To_Hex_String(rdata0_1147));
          --
        end if; 
        if CONCAT_u9_u73_1162_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:CONCAT_u9_u73_1162_inst:finished:  outputs: " & " CONCAT_u9_u73_1162_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u9_u73_1162_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : CONCAT_u9_u73_1162_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_1160_wire & rdata0_1147;
      CONCAT_u9_u73_1162_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u9_u73_1162_inst_req_0;
      CONCAT_u9_u73_1162_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u9_u73_1162_inst_req_1;
      CONCAT_u9_u73_1162_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator RPIPE_mac_to_nic_data_0_1149_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_mac_to_nic_data_0_1149_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:RPIPE_mac_to_nic_data_0_1149_inst:started:   PipeRead from mac_to_nic_data_0 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_mac_to_nic_data_0_1149_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:RPIPE_mac_to_nic_data_0_1149_inst:finished:  outputs: " & " RPIPE_mac_to_nic_data_0_1149_wire= "  & Convert_SLV_To_Hex_String(RPIPE_mac_to_nic_data_0_1149_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_mac_to_nic_data_0_1149_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_0_1149_inst_req_0;
      RPIPE_mac_to_nic_data_0_1149_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_0_1149_inst_req_1;
      RPIPE_mac_to_nic_data_0_1149_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_0_1149_wire <= data_out(63 downto 0);
      mac_to_nic_data_0_read_0_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_0_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_0_read_0: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_0_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_0_pipe_read_req(0),
          oack => mac_to_nic_data_0_pipe_read_ack(0),
          odata => mac_to_nic_data_0_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator RPIPE_mac_to_nic_data_1_1152_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_mac_to_nic_data_1_1152_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:RPIPE_mac_to_nic_data_1_1152_inst:started:   PipeRead from mac_to_nic_data_1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_mac_to_nic_data_1_1152_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:RPIPE_mac_to_nic_data_1_1152_inst:finished:  outputs: " & " RPIPE_mac_to_nic_data_1_1152_wire= "  & Convert_SLV_To_Hex_String(RPIPE_mac_to_nic_data_1_1152_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (1) : RPIPE_mac_to_nic_data_1_1152_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_1_1152_inst_req_0;
      RPIPE_mac_to_nic_data_1_1152_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_1_1152_inst_req_1;
      RPIPE_mac_to_nic_data_1_1152_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_1_1152_wire <= data_out(15 downto 0);
      mac_to_nic_data_1_read_1_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_1_read_1: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_1_pipe_read_req(0),
          oack => mac_to_nic_data_1_pipe_read_ack(0),
          odata => mac_to_nic_data_1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- logger for split-operator WPIPE_mac_to_nic_data_1157_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_mac_to_nic_data_1157_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:WPIPE_mac_to_nic_data_1157_inst:started:   PipeWrite to mac_to_nic_data inputs: " & " CONCAT_u9_u73_1162_wire = "& Convert_SLV_To_Hex_String(CONCAT_u9_u73_1162_wire));
          --
        end if; 
        if WPIPE_mac_to_nic_data_1157_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:macToNicInterface:DP:WPIPE_mac_to_nic_data_1157_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_mac_to_nic_data_1157_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_mac_to_nic_data_1157_inst_req_0;
      WPIPE_mac_to_nic_data_1157_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_mac_to_nic_data_1157_inst_req_1;
      WPIPE_mac_to_nic_data_1157_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u9_u73_1162_wire;
      mac_to_nic_data_write_0_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_write_0: OutputPortRevised -- 
        generic map ( name => "mac_to_nic_data", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => mac_to_nic_data_pipe_write_req(0),
          oack => mac_to_nic_data_pipe_write_ack(0),
          odata => mac_to_nic_data_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end macToNicInterface_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity memoryToNicInterface is -- 
  generic (tag_length : integer); 
  port ( -- 
    mem_resp0_pipe0_pipe_read_req : out  std_logic_vector(0 downto 0);
    mem_resp0_pipe0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mem_resp0_pipe0_pipe_read_data : in   std_logic_vector(63 downto 0);
    mem_resp0_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    mem_resp0_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mem_resp0_pipe1_pipe_read_data : in   std_logic_vector(7 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(64 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity memoryToNicInterface;
architecture memoryToNicInterface_arch of memoryToNicInterface is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal memoryToNicInterface_CP_2257_start: Boolean;
  signal memoryToNicInterface_CP_2257_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_mem_resp0_pipe0_1174_inst_ack_0 : boolean;
  signal RPIPE_mem_resp0_pipe0_1174_inst_ack_1 : boolean;
  signal RPIPE_mem_resp0_pipe0_1174_inst_req_1 : boolean;
  signal CONCAT_u1_u65_1184_inst_req_1 : boolean;
  signal CONCAT_u1_u65_1184_inst_ack_0 : boolean;
  signal WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_0 : boolean;
  signal RPIPE_mem_resp0_pipe1_1177_inst_req_0 : boolean;
  signal RPIPE_mem_resp0_pipe1_1177_inst_ack_0 : boolean;
  signal RPIPE_mem_resp0_pipe0_1174_inst_req_0 : boolean;
  signal RPIPE_mem_resp0_pipe1_1177_inst_req_1 : boolean;
  signal do_while_stmt_1170_branch_ack_0 : boolean;
  signal RPIPE_mem_resp0_pipe1_1177_inst_ack_1 : boolean;
  signal CONCAT_u1_u65_1184_inst_ack_1 : boolean;
  signal CONCAT_u1_u65_1184_inst_req_0 : boolean;
  signal WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_0 : boolean;
  signal do_while_stmt_1170_branch_ack_1 : boolean;
  signal do_while_stmt_1170_branch_req_0 : boolean;
  signal WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_1 : boolean;
  signal WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "memoryToNicInterface_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  memoryToNicInterface_CP_2257_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "memoryToNicInterface_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memoryToNicInterface_CP_2257_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= memoryToNicInterface_CP_2257_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= memoryToNicInterface_CP_2257_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,memoryToNicInterface_CP_2257_start,"memoryToNicInterface cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,memoryToNicInterface_CP_2257_symbol, "memoryToNicInterface cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  memoryToNicInterface_CP_2257: Block -- control-path 
    signal memoryToNicInterface_CP_2257_elements: BooleanArray(35 downto 0);
    -- 
  begin -- 
    memoryToNicInterface_CP_2257_elements(0) <= memoryToNicInterface_CP_2257_start;
    memoryToNicInterface_CP_2257_symbol <= memoryToNicInterface_CP_2257_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1169/do_while_stmt_1170__entry__
      -- CP-element group 0: 	 branch_block_stmt_1169/$entry
      -- CP-element group 0: 	 branch_block_stmt_1169/branch_block_stmt_1169__entry__
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	34 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1169/$exit
      -- CP-element group 1: 	 branch_block_stmt_1169/do_while_stmt_1170__exit__
      -- CP-element group 1: 	 branch_block_stmt_1169/branch_block_stmt_1169__exit__
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_CP_2257_elements(1) <= memoryToNicInterface_CP_2257_elements(34);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1169/do_while_stmt_1170/$entry
      -- CP-element group 2: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170__entry__
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_CP_2257_elements(2) <= memoryToNicInterface_CP_2257_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	34 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170__exit__
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memoryToNicInterface_CP_2257_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_back
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memoryToNicInterface_CP_2257_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	32 
    -- CP-element group 5: 	33 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1169/do_while_stmt_1170/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_exit/$entry
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_CP_2257_elements(5) <= memoryToNicInterface_CP_2257_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	35 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_body_done
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_CP_2257_elements(6) <= memoryToNicInterface_CP_2257_elements(35);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_CP_2257_elements(7) <= memoryToNicInterface_CP_2257_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_CP_2257_elements(8) <= memoryToNicInterface_CP_2257_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	19 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1172_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1175_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/loop_body_start
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memoryToNicInterface_CP_2257_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	31 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/condition_evaluated
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:do_while_stmt_1170_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(10), ack => do_while_stmt_1170_branch_req_0); -- 
    memoryToNicInterface_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(13) & memoryToNicInterface_CP_2257_elements(31);
      gj_memoryToNicInterface_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	20 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(9) & memoryToNicInterface_CP_2257_elements(13);
      gj_memoryToNicInterface_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	19 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	21 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(14) & memoryToNicInterface_CP_2257_elements(19);
      gj_memoryToNicInterface_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	23 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(18) & memoryToNicInterface_CP_2257_elements(23);
      gj_memoryToNicInterface_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	26 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1172_update_start_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(9) & memoryToNicInterface_CP_2257_elements(26);
      gj_memoryToNicInterface_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_sample_start_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe0_1174_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(15), ack => RPIPE_mem_resp0_pipe0_1174_inst_req_0); -- 
    memoryToNicInterface_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(11) & memoryToNicInterface_CP_2257_elements(18);
      gj_memoryToNicInterface_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: 	17 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Update/$entry
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe0_1174_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(16), ack => RPIPE_mem_resp0_pipe0_1174_inst_req_1); -- 
    memoryToNicInterface_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(12) & memoryToNicInterface_CP_2257_elements(17);
      gj_memoryToNicInterface_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: 	35 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Sample/$exit
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe0_1174_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mem_resp0_pipe0_1174_inst_ack_0, ack => memoryToNicInterface_CP_2257_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	24 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1172_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe0_1174_Update/$exit
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe0_1174_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mem_resp0_pipe0_1174_inst_ack_1, ack => memoryToNicInterface_CP_2257_elements(18)); -- 
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	9 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	26 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1175_update_start_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(9) & memoryToNicInterface_CP_2257_elements(26);
      gj_memoryToNicInterface_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	11 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_sample_start_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe1_1177_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(20), ack => RPIPE_mem_resp0_pipe1_1177_inst_req_0); -- 
    memoryToNicInterface_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(11) & memoryToNicInterface_CP_2257_elements(23);
      gj_memoryToNicInterface_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	12 
    -- CP-element group 21: 	22 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Update/cr
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe1_1177_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(21), ack => RPIPE_mem_resp0_pipe1_1177_inst_req_1); -- 
    memoryToNicInterface_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(12) & memoryToNicInterface_CP_2257_elements(22);
      gj_memoryToNicInterface_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	35 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_sample_completed_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe1_1177_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mem_resp0_pipe1_1177_inst_ack_0, ack => memoryToNicInterface_CP_2257_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	13 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/RPIPE_mem_resp0_pipe1_1177_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1175_update_completed_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:RPIPE_mem_resp0_pipe1_1177_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mem_resp0_pipe1_1177_inst_ack_1, ack => memoryToNicInterface_CP_2257_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: 	23 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Sample/rr
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:CONCAT_u1_u65_1184_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(24), ack => CONCAT_u1_u65_1184_inst_req_0); -- 
    memoryToNicInterface_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(18) & memoryToNicInterface_CP_2257_elements(23) & memoryToNicInterface_CP_2257_elements(26);
      gj_memoryToNicInterface_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_update_start_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:CONCAT_u1_u65_1184_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(25), ack => CONCAT_u1_u65_1184_inst_req_1); -- 
    memoryToNicInterface_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= memoryToNicInterface_CP_2257_elements(29);
      gj_memoryToNicInterface_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: 	19 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_sample_completed_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:CONCAT_u1_u65_1184_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u65_1184_inst_ack_0, ack => memoryToNicInterface_CP_2257_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/CONCAT_u1_u65_1184_update_completed_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:CONCAT_u1_u65_1184_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u1_u65_1184_inst_ack_1, ack => memoryToNicInterface_CP_2257_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Sample/$entry
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(28), ack => WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_0); -- 
    memoryToNicInterface_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(27) & memoryToNicInterface_CP_2257_elements(30);
      gj_memoryToNicInterface_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Update/req
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_0, ack => memoryToNicInterface_CP_2257_elements(29)); -- 
    req_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => memoryToNicInterface_CP_2257_elements(29), ack => WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_Update/ack
      -- CP-element group 30: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/WPIPE_MEMORY_TO_NIC_RESPONSE_1179_update_completed_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_1, ack => memoryToNicInterface_CP_2257_elements(30)); -- 
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	10 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group memoryToNicInterface_CP_2257_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => memoryToNicInterface_CP_2257_elements(9), ack => memoryToNicInterface_CP_2257_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	5 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_exit/ack
      -- CP-element group 32: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_exit/$exit
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:do_while_stmt_1170_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1170_branch_ack_0, ack => memoryToNicInterface_CP_2257_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	5 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_taken/$exit
      -- CP-element group 33: 	 branch_block_stmt_1169/do_while_stmt_1170/loop_taken/ack
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:do_while_stmt_1170_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1170_branch_ack_1, ack => memoryToNicInterface_CP_2257_elements(33)); -- 
    -- CP-element group 34:  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	3 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	1 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1169/do_while_stmt_1170/$exit
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_CP_2257_elements(34) <= memoryToNicInterface_CP_2257_elements(3);
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	17 
    -- CP-element group 35: 	22 
    -- CP-element group 35: 	30 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	6 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/aggregated_phi_sample_ack
      -- CP-element group 35: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/$exit
      -- CP-element group 35: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1175_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1169/do_while_stmt_1170/do_while_stmt_1170_loop_body/phi_stmt_1172_sample_completed_
      -- 
    -- logger for CP element group memoryToNicInterface_CP_2257_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and memoryToNicInterface_CP_2257_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:memoryToNicInterface:CP:memoryToNicInterface_CP_2257_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    memoryToNicInterface_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "memoryToNicInterface_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= memoryToNicInterface_CP_2257_elements(17) & memoryToNicInterface_CP_2257_elements(22) & memoryToNicInterface_CP_2257_elements(30);
      gj_memoryToNicInterface_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(35), clk => clk, reset => reset); --
    end block;
    memoryToNicInterface_do_while_stmt_1170_terminator_2360: loop_terminator -- 
      generic map (name => " memoryToNicInterface_do_while_stmt_1170_terminator_2360", max_iterations_in_flight =>7) 
      port map(loop_body_exit => memoryToNicInterface_CP_2257_elements(6),loop_continue => memoryToNicInterface_CP_2257_elements(33),loop_terminate => memoryToNicInterface_CP_2257_elements(32),loop_back => memoryToNicInterface_CP_2257_elements(4),loop_exit => memoryToNicInterface_CP_2257_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_2282_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= memoryToNicInterface_CP_2257_elements(7);
        preds(1)  <= memoryToNicInterface_CP_2257_elements(8);
        entry_tmerge_2282 : transition_merge -- 
          generic map(name => " entry_tmerge_2282")
          port map (preds => preds, symbol_out => memoryToNicInterface_CP_2257_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u8_u1_1182_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u1_u65_1184_wire : std_logic_vector(64 downto 0);
    signal RPIPE_mem_resp0_pipe0_1174_wire : std_logic_vector(63 downto 0);
    signal RPIPE_mem_resp0_pipe1_1177_wire : std_logic_vector(7 downto 0);
    signal konst_1181_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1187_wire_constant : std_logic_vector(0 downto 0);
    signal rdata0_1172 : std_logic_vector(63 downto 0);
    signal rdata1_1175 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1181_wire_constant <= "00000000";
    konst_1187_wire_constant <= "1";
    -- logger for split-operator ssrc_phi_stmt_1172 flow-through 
    process(rdata0_1172) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:ssrc_phi_stmt_1172:flowthrough inputs: " & " RPIPE_mem_resp0_pipe0_1174_wire = "& Convert_SLV_To_Hex_String(RPIPE_mem_resp0_pipe0_1174_wire) & " outputs:" & " rdata0_1172= "  & Convert_SLV_To_Hex_String(rdata0_1172));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1172
    process(RPIPE_mem_resp0_pipe0_1174_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := RPIPE_mem_resp0_pipe0_1174_wire(63 downto 0);
      rdata0_1172 <= tmp_var; -- 
    end process;
    -- logger for split-operator ssrc_phi_stmt_1175 flow-through 
    process(rdata1_1175) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:ssrc_phi_stmt_1175:flowthrough inputs: " & " RPIPE_mem_resp0_pipe1_1177_wire = "& Convert_SLV_To_Hex_String(RPIPE_mem_resp0_pipe1_1177_wire) & " outputs:" & " rdata1_1175= "  & Convert_SLV_To_Hex_String(rdata1_1175));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1175
    process(RPIPE_mem_resp0_pipe1_1177_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := RPIPE_mem_resp0_pipe1_1177_wire(7 downto 0);
      rdata1_1175 <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1170_branch_req_0," req0 do_while_stmt_1170_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1170_branch_ack_0," ack0 do_while_stmt_1170_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1170_branch_ack_1," ack1 do_while_stmt_1170_branch");
    do_while_stmt_1170_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1187_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1170_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1170_branch_req_0,
          ack0 => do_while_stmt_1170_branch_ack_0,
          ack1 => do_while_stmt_1170_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator BITSEL_u8_u1_1182_inst flow-through 
    process(BITSEL_u8_u1_1182_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:BITSEL_u8_u1_1182_inst:flowthrough inputs: " & " rdata1_1175 = "& Convert_SLV_To_Hex_String(rdata1_1175) & " konst_1181_wire_constant = "& Convert_SLV_To_Hex_String(konst_1181_wire_constant) & " outputs:" & " BITSEL_u8_u1_1182_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u8_u1_1182_wire));
      --
    end process; 
    -- binary operator BITSEL_u8_u1_1182_inst
    process(rdata1_1175) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(rdata1_1175, konst_1181_wire_constant, tmp_var);
      BITSEL_u8_u1_1182_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u65_1184_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u1_u65_1184_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:CONCAT_u1_u65_1184_inst:started:   inputs: " & " BITSEL_u8_u1_1182_wire = "& Convert_SLV_To_Hex_String(BITSEL_u8_u1_1182_wire) & " rdata0_1172 = "& Convert_SLV_To_Hex_String(rdata0_1172));
          --
        end if; 
        if CONCAT_u1_u65_1184_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:CONCAT_u1_u65_1184_inst:finished:  outputs: " & " CONCAT_u1_u65_1184_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u65_1184_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : CONCAT_u1_u65_1184_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(64 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= BITSEL_u8_u1_1182_wire & rdata0_1172;
      CONCAT_u1_u65_1184_wire <= data_out(64 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u1_u65_1184_inst_req_0;
      CONCAT_u1_u65_1184_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u1_u65_1184_inst_req_1;
      CONCAT_u1_u65_1184_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 65,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator RPIPE_mem_resp0_pipe0_1174_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_mem_resp0_pipe0_1174_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:RPIPE_mem_resp0_pipe0_1174_inst:started:   PipeRead from mem_resp0_pipe0 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_mem_resp0_pipe0_1174_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:RPIPE_mem_resp0_pipe0_1174_inst:finished:  outputs: " & " RPIPE_mem_resp0_pipe0_1174_wire= "  & Convert_SLV_To_Hex_String(RPIPE_mem_resp0_pipe0_1174_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_mem_resp0_pipe0_1174_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mem_resp0_pipe0_1174_inst_req_0;
      RPIPE_mem_resp0_pipe0_1174_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mem_resp0_pipe0_1174_inst_req_1;
      RPIPE_mem_resp0_pipe0_1174_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mem_resp0_pipe0_1174_wire <= data_out(63 downto 0);
      mem_resp0_pipe0_read_0_gI: SplitGuardInterface generic map(name => "mem_resp0_pipe0_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mem_resp0_pipe0_read_0: InputPortRevised -- 
        generic map ( name => "mem_resp0_pipe0_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mem_resp0_pipe0_pipe_read_req(0),
          oack => mem_resp0_pipe0_pipe_read_ack(0),
          odata => mem_resp0_pipe0_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator RPIPE_mem_resp0_pipe1_1177_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_mem_resp0_pipe1_1177_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:RPIPE_mem_resp0_pipe1_1177_inst:started:   PipeRead from mem_resp0_pipe1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_mem_resp0_pipe1_1177_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:RPIPE_mem_resp0_pipe1_1177_inst:finished:  outputs: " & " RPIPE_mem_resp0_pipe1_1177_wire= "  & Convert_SLV_To_Hex_String(RPIPE_mem_resp0_pipe1_1177_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (1) : RPIPE_mem_resp0_pipe1_1177_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mem_resp0_pipe1_1177_inst_req_0;
      RPIPE_mem_resp0_pipe1_1177_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mem_resp0_pipe1_1177_inst_req_1;
      RPIPE_mem_resp0_pipe1_1177_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mem_resp0_pipe1_1177_wire <= data_out(7 downto 0);
      mem_resp0_pipe1_read_1_gI: SplitGuardInterface generic map(name => "mem_resp0_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mem_resp0_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "mem_resp0_pipe1_read_1", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mem_resp0_pipe1_pipe_read_req(0),
          oack => mem_resp0_pipe1_pipe_read_ack(0),
          odata => mem_resp0_pipe1_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- logger for split-operator WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst:started:   PipeWrite to MEMORY_TO_NIC_RESPONSE inputs: " & " CONCAT_u1_u65_1184_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u65_1184_wire));
          --
        end if; 
        if WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:memoryToNicInterface:DP:WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_0;
      WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_req_1;
      WPIPE_MEMORY_TO_NIC_RESPONSE_1179_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u1_u65_1184_wire;
      MEMORY_TO_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE", data_width => 65, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_write_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_write_data(64 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end memoryToNicInterface_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity nextLSTATE_Volatile is -- 
  port ( -- 
    clk, reset: in std_logic; 
    RX : in  std_logic_vector(72 downto 0);
    LSTATE : in  std_logic_vector(1 downto 0);
    nLSTATE : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity nextLSTATE_Volatile;
architecture nextLSTATE_Volatile_arch of nextLSTATE_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal RX_buffer :  std_logic_vector(72 downto 0);
  signal LSTATE_buffer :  std_logic_vector(1 downto 0);
  -- output port buffer signals
  signal nLSTATE_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  RX_buffer <= RX;
  LSTATE_buffer <= LSTATE;
  -- output handling  -------------------------------------------------------
  nLSTATE <= nLSTATE_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1230_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1238_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1214_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1220_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1227_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1236_wire : std_logic_vector(0 downto 0);
    signal MUX_1217_wire : std_logic_vector(1 downto 0);
    signal MUX_1223_wire : std_logic_vector(1 downto 0);
    signal MUX_1233_wire : std_logic_vector(1 downto 0);
    signal MUX_1241_wire : std_logic_vector(1 downto 0);
    signal NOT_u1_u1_1229_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_1224_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_1242_wire : std_logic_vector(1 downto 0);
    signal R_S0_1213_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1239_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1215_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1219_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1221_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1226_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1231_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_1235_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1208_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1216_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1222_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1232_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1240_wire_constant : std_logic_vector(1 downto 0);
    signal last_word_1210 : std_logic_vector(0 downto 0);
    signal tdata_1201 : std_logic_vector(63 downto 0);
    signal tkeep_1205 : std_logic_vector(7 downto 0);
    signal tlast_1197 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_S0_1213_wire_constant <= "00";
    R_S0_1239_wire_constant <= "00";
    R_S1_1215_wire_constant <= "01";
    R_S1_1219_wire_constant <= "01";
    R_S2_1221_wire_constant <= "10";
    R_S2_1226_wire_constant <= "10";
    R_S2_1231_wire_constant <= "10";
    R_S2_1235_wire_constant <= "10";
    konst_1208_wire_constant <= "1";
    konst_1216_wire_constant <= "00";
    konst_1222_wire_constant <= "00";
    konst_1232_wire_constant <= "00";
    konst_1240_wire_constant <= "00";
    -- logger for split-operator MUX_1217_inst flow-through 
    process(MUX_1217_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:MUX_1217_inst:flowthrough inputs: " & " EQ_u2_u1_1214_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_1214_wire) & " R_S1_1215_wire_constant = "& Convert_SLV_To_Hex_String(R_S1_1215_wire_constant) & " konst_1216_wire_constant = "& Convert_SLV_To_Hex_String(konst_1216_wire_constant) & " outputs:" & " MUX_1217_wire= "  & Convert_SLV_To_Hex_String(MUX_1217_wire));
      --
    end process; 
    -- flow-through select operator MUX_1217_inst
    MUX_1217_wire <= R_S1_1215_wire_constant when (EQ_u2_u1_1214_wire(0) /=  '0') else konst_1216_wire_constant;
    -- logger for split-operator MUX_1223_inst flow-through 
    process(MUX_1223_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:MUX_1223_inst:flowthrough inputs: " & " EQ_u2_u1_1220_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_1220_wire) & " R_S2_1221_wire_constant = "& Convert_SLV_To_Hex_String(R_S2_1221_wire_constant) & " konst_1222_wire_constant = "& Convert_SLV_To_Hex_String(konst_1222_wire_constant) & " outputs:" & " MUX_1223_wire= "  & Convert_SLV_To_Hex_String(MUX_1223_wire));
      --
    end process; 
    -- flow-through select operator MUX_1223_inst
    MUX_1223_wire <= R_S2_1221_wire_constant when (EQ_u2_u1_1220_wire(0) /=  '0') else konst_1222_wire_constant;
    -- logger for split-operator MUX_1233_inst flow-through 
    process(MUX_1233_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:MUX_1233_inst:flowthrough inputs: " & " AND_u1_u1_1230_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_1230_wire) & " R_S2_1231_wire_constant = "& Convert_SLV_To_Hex_String(R_S2_1231_wire_constant) & " konst_1232_wire_constant = "& Convert_SLV_To_Hex_String(konst_1232_wire_constant) & " outputs:" & " MUX_1233_wire= "  & Convert_SLV_To_Hex_String(MUX_1233_wire));
      --
    end process; 
    -- flow-through select operator MUX_1233_inst
    MUX_1233_wire <= R_S2_1231_wire_constant when (AND_u1_u1_1230_wire(0) /=  '0') else konst_1232_wire_constant;
    -- logger for split-operator MUX_1241_inst flow-through 
    process(MUX_1241_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:MUX_1241_inst:flowthrough inputs: " & " AND_u1_u1_1238_wire = "& Convert_SLV_To_Hex_String(AND_u1_u1_1238_wire) & " R_S0_1239_wire_constant = "& Convert_SLV_To_Hex_String(R_S0_1239_wire_constant) & " konst_1240_wire_constant = "& Convert_SLV_To_Hex_String(konst_1240_wire_constant) & " outputs:" & " MUX_1241_wire= "  & Convert_SLV_To_Hex_String(MUX_1241_wire));
      --
    end process; 
    -- flow-through select operator MUX_1241_inst
    MUX_1241_wire <= R_S0_1239_wire_constant when (AND_u1_u1_1238_wire(0) /=  '0') else konst_1240_wire_constant;
    -- logger for split-operator slice_1196_inst flow-through 
    process(tlast_1197) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:slice_1196_inst:flowthrough inputs: " & " RX_buffer = "& Convert_SLV_To_Hex_String(RX_buffer) & " outputs:" & " tlast_1197= "  & Convert_SLV_To_Hex_String(tlast_1197));
      --
    end process; 
    -- flow-through slice operator slice_1196_inst
    tlast_1197 <= RX_buffer(72 downto 72);
    -- logger for split-operator slice_1200_inst flow-through 
    process(tdata_1201) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:slice_1200_inst:flowthrough inputs: " & " RX_buffer = "& Convert_SLV_To_Hex_String(RX_buffer) & " outputs:" & " tdata_1201= "  & Convert_SLV_To_Hex_String(tdata_1201));
      --
    end process; 
    -- flow-through slice operator slice_1200_inst
    tdata_1201 <= RX_buffer(71 downto 8);
    -- logger for split-operator slice_1204_inst flow-through 
    process(tkeep_1205) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:slice_1204_inst:flowthrough inputs: " & " RX_buffer = "& Convert_SLV_To_Hex_String(RX_buffer) & " outputs:" & " tkeep_1205= "  & Convert_SLV_To_Hex_String(tkeep_1205));
      --
    end process; 
    -- flow-through slice operator slice_1204_inst
    tkeep_1205 <= RX_buffer(7 downto 0);
    -- logger for split-operator AND_u1_u1_1230_inst flow-through 
    process(AND_u1_u1_1230_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:AND_u1_u1_1230_inst:flowthrough inputs: " & " EQ_u2_u1_1227_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_1227_wire) & " NOT_u1_u1_1229_wire = "& Convert_SLV_To_Hex_String(NOT_u1_u1_1229_wire) & " outputs:" & " AND_u1_u1_1230_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_1230_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_1230_inst
    process(EQ_u2_u1_1227_wire, NOT_u1_u1_1229_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1227_wire, NOT_u1_u1_1229_wire, tmp_var);
      AND_u1_u1_1230_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_1238_inst flow-through 
    process(AND_u1_u1_1238_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:AND_u1_u1_1238_inst:flowthrough inputs: " & " EQ_u2_u1_1236_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_1236_wire) & " last_word_1210 = "& Convert_SLV_To_Hex_String(last_word_1210) & " outputs:" & " AND_u1_u1_1238_wire= "  & Convert_SLV_To_Hex_String(AND_u1_u1_1238_wire));
      --
    end process; 
    -- binary operator AND_u1_u1_1238_inst
    process(EQ_u2_u1_1236_wire, last_word_1210) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_1236_wire, last_word_1210, tmp_var);
      AND_u1_u1_1238_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_1209_inst flow-through 
    process(last_word_1210) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:EQ_u1_u1_1209_inst:flowthrough inputs: " & " tlast_1197 = "& Convert_SLV_To_Hex_String(tlast_1197) & " konst_1208_wire_constant = "& Convert_SLV_To_Hex_String(konst_1208_wire_constant) & " outputs:" & " last_word_1210= "  & Convert_SLV_To_Hex_String(last_word_1210));
      --
    end process; 
    -- binary operator EQ_u1_u1_1209_inst
    process(tlast_1197) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tlast_1197, konst_1208_wire_constant, tmp_var);
      last_word_1210 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1214_inst flow-through 
    process(EQ_u2_u1_1214_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:EQ_u2_u1_1214_inst:flowthrough inputs: " & " LSTATE_buffer = "& Convert_SLV_To_Hex_String(LSTATE_buffer) & " R_S0_1213_wire_constant = "& Convert_SLV_To_Hex_String(R_S0_1213_wire_constant) & " outputs:" & " EQ_u2_u1_1214_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1214_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1214_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S0_1213_wire_constant, tmp_var);
      EQ_u2_u1_1214_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1220_inst flow-through 
    process(EQ_u2_u1_1220_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:EQ_u2_u1_1220_inst:flowthrough inputs: " & " LSTATE_buffer = "& Convert_SLV_To_Hex_String(LSTATE_buffer) & " R_S1_1219_wire_constant = "& Convert_SLV_To_Hex_String(R_S1_1219_wire_constant) & " outputs:" & " EQ_u2_u1_1220_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1220_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1220_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S1_1219_wire_constant, tmp_var);
      EQ_u2_u1_1220_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1227_inst flow-through 
    process(EQ_u2_u1_1227_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:EQ_u2_u1_1227_inst:flowthrough inputs: " & " LSTATE_buffer = "& Convert_SLV_To_Hex_String(LSTATE_buffer) & " R_S2_1226_wire_constant = "& Convert_SLV_To_Hex_String(R_S2_1226_wire_constant) & " outputs:" & " EQ_u2_u1_1227_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1227_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1227_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1226_wire_constant, tmp_var);
      EQ_u2_u1_1227_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1236_inst flow-through 
    process(EQ_u2_u1_1236_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:EQ_u2_u1_1236_inst:flowthrough inputs: " & " LSTATE_buffer = "& Convert_SLV_To_Hex_String(LSTATE_buffer) & " R_S2_1235_wire_constant = "& Convert_SLV_To_Hex_String(R_S2_1235_wire_constant) & " outputs:" & " EQ_u2_u1_1236_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1236_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1236_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_1235_wire_constant, tmp_var);
      EQ_u2_u1_1236_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_1229_inst flow-through 
    process(NOT_u1_u1_1229_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:NOT_u1_u1_1229_inst:flowthrough inputs: " & " last_word_1210 = "& Convert_SLV_To_Hex_String(last_word_1210) & " outputs:" & " NOT_u1_u1_1229_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_1229_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_1229_inst
    process(last_word_1210) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_word_1210, tmp_var);
      NOT_u1_u1_1229_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator OR_u2_u2_1224_inst flow-through 
    process(OR_u2_u2_1224_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:OR_u2_u2_1224_inst:flowthrough inputs: " & " MUX_1217_wire = "& Convert_SLV_To_Hex_String(MUX_1217_wire) & " MUX_1223_wire = "& Convert_SLV_To_Hex_String(MUX_1223_wire) & " outputs:" & " OR_u2_u2_1224_wire= "  & Convert_SLV_To_Hex_String(OR_u2_u2_1224_wire));
      --
    end process; 
    -- binary operator OR_u2_u2_1224_inst
    process(MUX_1217_wire, MUX_1223_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1217_wire, MUX_1223_wire, tmp_var);
      OR_u2_u2_1224_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u2_u2_1242_inst flow-through 
    process(OR_u2_u2_1242_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:OR_u2_u2_1242_inst:flowthrough inputs: " & " MUX_1233_wire = "& Convert_SLV_To_Hex_String(MUX_1233_wire) & " MUX_1241_wire = "& Convert_SLV_To_Hex_String(MUX_1241_wire) & " outputs:" & " OR_u2_u2_1242_wire= "  & Convert_SLV_To_Hex_String(OR_u2_u2_1242_wire));
      --
    end process; 
    -- binary operator OR_u2_u2_1242_inst
    process(MUX_1233_wire, MUX_1241_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1233_wire, MUX_1241_wire, tmp_var);
      OR_u2_u2_1242_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u2_u2_1243_inst flow-through 
    process(nLSTATE_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nextLSTATE:DP:OR_u2_u2_1243_inst:flowthrough inputs: " & " OR_u2_u2_1224_wire = "& Convert_SLV_To_Hex_String(OR_u2_u2_1224_wire) & " OR_u2_u2_1242_wire = "& Convert_SLV_To_Hex_String(OR_u2_u2_1242_wire) & " outputs:" & " nLSTATE_buffer= "  & Convert_SLV_To_Hex_String(nLSTATE_buffer));
      --
    end process; 
    -- binary operator OR_u2_u2_1243_inst
    process(OR_u2_u2_1224_wire, OR_u2_u2_1242_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_1224_wire, OR_u2_u2_1242_wire, tmp_var);
      nLSTATE_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end nextLSTATE_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity nicRxFromMacDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
    nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
    nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicRxFromMacDaemon;
architecture nicRxFromMacDaemon_arch of nicRxFromMacDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicRxFromMacDaemon_CP_2364_start: Boolean;
  signal nicRxFromMacDaemon_CP_2364_symbol: Boolean;
  -- volatile/operator module components. 
  component nextLSTATE_Volatile is -- 
    port ( -- 
      clk, reset: in std_logic; 
      RX : in  std_logic_vector(72 downto 0);
      LSTATE : in  std_logic_vector(1 downto 0);
      nLSTATE : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal do_while_stmt_1248_branch_req_0 : boolean;
  signal phi_stmt_1250_req_0 : boolean;
  signal phi_stmt_1250_req_1 : boolean;
  signal phi_stmt_1250_ack_0 : boolean;
  signal nLSTATE_1264_1252_buf_req_0 : boolean;
  signal nLSTATE_1264_1252_buf_ack_0 : boolean;
  signal nLSTATE_1264_1252_buf_req_1 : boolean;
  signal nLSTATE_1264_1252_buf_ack_1 : boolean;
  signal RPIPE_mac_to_nic_data_1256_inst_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_1256_inst_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_1256_inst_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_1256_inst_ack_1 : boolean;
  signal MUX_1284_inst_req_0 : boolean;
  signal MUX_1284_inst_ack_0 : boolean;
  signal MUX_1284_inst_req_1 : boolean;
  signal MUX_1284_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_1275_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_header_1275_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_header_1275_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_header_1275_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_packet_1286_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1286_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_1286_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_packet_1286_inst_ack_1 : boolean;
  signal do_while_stmt_1248_branch_ack_0 : boolean;
  signal do_while_stmt_1248_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicRxFromMacDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicRxFromMacDaemon_CP_2364_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicRxFromMacDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2364_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2364_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_2364_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,nicRxFromMacDaemon_CP_2364_start,"nicRxFromMacDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,nicRxFromMacDaemon_CP_2364_symbol, "nicRxFromMacDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicRxFromMacDaemon_CP_2364: Block -- control-path 
    signal nicRxFromMacDaemon_CP_2364_elements: BooleanArray(51 downto 0);
    -- 
  begin -- 
    nicRxFromMacDaemon_CP_2364_elements(0) <= nicRxFromMacDaemon_CP_2364_start;
    nicRxFromMacDaemon_CP_2364_symbol <= nicRxFromMacDaemon_CP_2364_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1247/$entry
      -- CP-element group 0: 	 branch_block_stmt_1247/branch_block_stmt_1247__entry__
      -- CP-element group 0: 	 branch_block_stmt_1247/do_while_stmt_1248__entry__
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	51 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1247/$exit
      -- CP-element group 1: 	 branch_block_stmt_1247/branch_block_stmt_1247__exit__
      -- CP-element group 1: 	 branch_block_stmt_1247/do_while_stmt_1248__exit__
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(1) <= nicRxFromMacDaemon_CP_2364_elements(51);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1247/do_while_stmt_1248/$entry
      -- CP-element group 2: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248__entry__
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(2) <= nicRxFromMacDaemon_CP_2364_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	51 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248__exit__
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_back
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	49 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1247/do_while_stmt_1248/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_taken/$entry
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(5) <= nicRxFromMacDaemon_CP_2364_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	48 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_body_done
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(6) <= nicRxFromMacDaemon_CP_2364_elements(48);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(7) <= nicRxFromMacDaemon_CP_2364_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(8) <= nicRxFromMacDaemon_CP_2364_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	47 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1254_sample_start_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	47 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/condition_evaluated
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:do_while_stmt_1248_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(10), ack => do_while_stmt_1248_branch_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(14) & nicRxFromMacDaemon_CP_2364_elements(47);
      gj_nicRxFromMacDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_sample_start__ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(9) & nicRxFromMacDaemon_CP_2364_elements(15) & nicRxFromMacDaemon_CP_2364_elements(14);
      gj_nicRxFromMacDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	48 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1254_sample_completed_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(35) & nicRxFromMacDaemon_CP_2364_elements(17);
      gj_nicRxFromMacDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_update_start__ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(32) & nicRxFromMacDaemon_CP_2364_elements(16);
      gj_nicRxFromMacDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(36) & nicRxFromMacDaemon_CP_2364_elements(18);
      gj_nicRxFromMacDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_sample_start_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(9) & nicRxFromMacDaemon_CP_2364_elements(12);
      gj_nicRxFromMacDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	42 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_update_start_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(9) & nicRxFromMacDaemon_CP_2364_elements(39) & nicRxFromMacDaemon_CP_2364_elements(42);
      gj_nicRxFromMacDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_sample_completed__ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18: 	41 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_update_completed__ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_loopback_trigger
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(19) <= nicRxFromMacDaemon_CP_2364_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_loopback_sample_req_ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:phi_stmt_1250_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1250_loopback_sample_req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1250_loopback_sample_req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(20), ack => phi_stmt_1250_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_entry_trigger
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(21) <= nicRxFromMacDaemon_CP_2364_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_entry_sample_req_ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:phi_stmt_1250_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1250_entry_sample_req_2406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1250_entry_sample_req_2406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(22), ack => phi_stmt_1250_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1250_phi_mux_ack_ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:phi_stmt_1250_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1250_phi_mux_ack_2409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1250_ack_0, ack => nicRxFromMacDaemon_CP_2364_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Sample/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nLSTATE_1264_1252_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(24), ack => nLSTATE_1264_1252_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Update/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nLSTATE_1264_1252_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(25), ack => nLSTATE_1264_1252_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Sample/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nLSTATE_1264_1252_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1264_1252_buf_ack_0, ack => nicRxFromMacDaemon_CP_2364_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_nLSTATE_1252_Update/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nLSTATE_1264_1252_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_1264_1252_buf_ack_1, ack => nicRxFromMacDaemon_CP_2364_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_sample_completed_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_update_start_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_update_completed__ps
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(30) <= nicRxFromMacDaemon_CP_2364_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/R_S0_1253_update_completed_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2364_elements(29), ack => nicRxFromMacDaemon_CP_2364_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	39 
    -- CP-element group 32: 	45 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1254_update_start_
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(9) & nicRxFromMacDaemon_CP_2364_elements(39) & nicRxFromMacDaemon_CP_2364_elements(45);
      gj_nicRxFromMacDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Sample/rr
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:RPIPE_mac_to_nic_data_1256_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(33), ack => RPIPE_mac_to_nic_data_1256_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(11) & nicRxFromMacDaemon_CP_2364_elements(36);
      gj_nicRxFromMacDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Update/cr
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:RPIPE_mac_to_nic_data_1256_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(34), ack => RPIPE_mac_to_nic_data_1256_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(13) & nicRxFromMacDaemon_CP_2364_elements(35);
      gj_nicRxFromMacDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Sample/ra
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:RPIPE_mac_to_nic_data_1256_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1256_inst_ack_0, ack => nicRxFromMacDaemon_CP_2364_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	44 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/phi_stmt_1254_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/RPIPE_mac_to_nic_data_1256_Update/ca
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:RPIPE_mac_to_nic_data_1256_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_1256_inst_ack_1, ack => nicRxFromMacDaemon_CP_2364_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_start/$entry
      -- CP-element group 37: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_start/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:MUX_1284_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(37), ack => MUX_1284_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(36) & nicRxFromMacDaemon_CP_2364_elements(18) & nicRxFromMacDaemon_CP_2364_elements(39);
      gj_nicRxFromMacDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	42 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_complete/$entry
      -- CP-element group 38: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_complete/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:MUX_1284_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(38), ack => MUX_1284_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicRxFromMacDaemon_CP_2364_elements(42);
      gj_nicRxFromMacDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: 	32 
    -- CP-element group 39: 	16 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_start/$exit
      -- CP-element group 39: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_start/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:MUX_1284_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1284_inst_ack_0, ack => nicRxFromMacDaemon_CP_2364_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_complete/$exit
      -- CP-element group 40: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/MUX_1284_complete/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:MUX_1284_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1284_inst_ack_1, ack => nicRxFromMacDaemon_CP_2364_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Sample/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_header_1275_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(41), ack => WPIPE_nic_rx_to_header_1275_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(40) & nicRxFromMacDaemon_CP_2364_elements(18) & nicRxFromMacDaemon_CP_2364_elements(43);
      gj_nicRxFromMacDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	38 
    -- CP-element group 42: 	16 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_update_start_
      -- CP-element group 42: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Update/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_header_1275_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_header_1275_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1275_inst_ack_0, ack => nicRxFromMacDaemon_CP_2364_elements(42)); -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(42), ack => WPIPE_nic_rx_to_header_1275_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	48 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_header_1275_Update/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_header_1275_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_1275_inst_ack_1, ack => nicRxFromMacDaemon_CP_2364_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	36 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Sample/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_packet_1286_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(44), ack => WPIPE_nic_rx_to_packet_1286_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(36) & nicRxFromMacDaemon_CP_2364_elements(46);
      gj_nicRxFromMacDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	32 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Update/req
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_packet_1286_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_packet_1286_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1286_inst_ack_0, ack => nicRxFromMacDaemon_CP_2364_elements(45)); -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_2364_elements(45), ack => WPIPE_nic_rx_to_packet_1286_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/WPIPE_nic_rx_to_packet_1286_Update/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:WPIPE_nic_rx_to_packet_1286_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_1286_inst_ack_1, ack => nicRxFromMacDaemon_CP_2364_elements(46)); -- 
    -- CP-element group 47:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	9 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	10 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(47) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicRxFromMacDaemon_CP_2364_elements(47) is a control-delay.
    cp_element_47_delay: control_delay_element  generic map(name => " 47_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_2364_elements(9), ack => nicRxFromMacDaemon_CP_2364_elements(47), clk => clk, reset =>reset);
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	12 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	6 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1247/do_while_stmt_1248/do_while_stmt_1248_loop_body/$exit
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_2364_elements(12) & nicRxFromMacDaemon_CP_2364_elements(43) & nicRxFromMacDaemon_CP_2364_elements(46);
      gj_nicRxFromMacDaemon_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	5 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_exit/$exit
      -- CP-element group 49: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_exit/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:do_while_stmt_1248_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1248_branch_ack_0, ack => nicRxFromMacDaemon_CP_2364_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_taken/$exit
      -- CP-element group 50: 	 branch_block_stmt_1247/do_while_stmt_1248/loop_taken/ack
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:do_while_stmt_1248_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1248_branch_ack_1, ack => nicRxFromMacDaemon_CP_2364_elements(50)); -- 
    -- CP-element group 51:  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	3 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	1 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1247/do_while_stmt_1248/$exit
      -- 
    -- logger for CP element group nicRxFromMacDaemon_CP_2364_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicRxFromMacDaemon_CP_2364_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicRxFromMacDaemon:CP:nicRxFromMacDaemon_CP_2364_elements(51) fired."); 
        -- 
      end if; --
    end process; 
    nicRxFromMacDaemon_CP_2364_elements(51) <= nicRxFromMacDaemon_CP_2364_elements(3);
    nicRxFromMacDaemon_do_while_stmt_1248_terminator_2507: loop_terminator -- 
      generic map (name => " nicRxFromMacDaemon_do_while_stmt_1248_terminator_2507", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicRxFromMacDaemon_CP_2364_elements(6),loop_continue => nicRxFromMacDaemon_CP_2364_elements(50),loop_terminate => nicRxFromMacDaemon_CP_2364_elements(49),loop_back => nicRxFromMacDaemon_CP_2364_elements(4),loop_exit => nicRxFromMacDaemon_CP_2364_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1250_phi_seq_2437_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_2364_elements(19);
      nicRxFromMacDaemon_CP_2364_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_2364_elements(26);
      nicRxFromMacDaemon_CP_2364_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_2364_elements(27);
      nicRxFromMacDaemon_CP_2364_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_2364_elements(21);
      nicRxFromMacDaemon_CP_2364_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_2364_elements(28);
      nicRxFromMacDaemon_CP_2364_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_2364_elements(30);
      nicRxFromMacDaemon_CP_2364_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1250_phi_seq_2437 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1250_phi_seq_2437") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_2364_elements(11), 
          phi_sample_ack => nicRxFromMacDaemon_CP_2364_elements(17), 
          phi_update_req => nicRxFromMacDaemon_CP_2364_elements(13), 
          phi_update_ack => nicRxFromMacDaemon_CP_2364_elements(18), 
          phi_mux_ack => nicRxFromMacDaemon_CP_2364_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2389_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicRxFromMacDaemon_CP_2364_elements(7);
        preds(1)  <= nicRxFromMacDaemon_CP_2364_elements(8);
        entry_tmerge_2389 : transition_merge -- 
          generic map(name => " entry_tmerge_2389")
          port map (preds => preds, symbol_out => nicRxFromMacDaemon_CP_2364_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u65_u73_1282_wire : std_logic_vector(72 downto 0);
    signal EQ_u2_u1_1268_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1271_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1278_wire : std_logic_vector(0 downto 0);
    signal LSTATE_1250 : std_logic_vector(1 downto 0);
    signal MUX_1284_wire : std_logic_vector(72 downto 0);
    signal RPIPE_mac_to_nic_data_1256_wire : std_logic_vector(72 downto 0);
    signal RX_1254 : std_logic_vector(72 downto 0);
    signal R_HEADER_TKEEP_1281_wire_constant : std_logic_vector(7 downto 0);
    signal R_S0_1253_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_1267_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1270_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_1277_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1292_wire_constant : std_logic_vector(0 downto 0);
    signal nLSTATE_1264 : std_logic_vector(1 downto 0);
    signal nLSTATE_1264_1252_buffered : std_logic_vector(1 downto 0);
    signal slice_1280_wire : std_logic_vector(64 downto 0);
    signal write_to_header_1273 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_HEADER_TKEEP_1281_wire_constant <= "00111111";
    R_S0_1253_wire_constant <= "00";
    R_S0_1267_wire_constant <= "00";
    R_S1_1270_wire_constant <= "01";
    R_S1_1277_wire_constant <= "01";
    konst_1292_wire_constant <= "1";
    -- logger for phi phi_stmt_1250
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1250_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:nicRxFromMacDaemon:DP:phi_stmt_1250:input-0 nLSTATE_1264_1252_buffered= " & Convert_SLV_To_Hex_String(nLSTATE_1264_1252_buffered));
          --
        end if;
        if phi_stmt_1250_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:nicRxFromMacDaemon:DP:phi_stmt_1250:input-1 R_S0_1253_wire_constant= " & Convert_SLV_To_Hex_String(R_S0_1253_wire_constant));
          --
        end if;
        if phi_stmt_1250_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:nicRxFromMacDaemon:DP:phi_stmt_1250:sample-completed");
          --
        end if;
        if phi_stmt_1250_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:nicRxFromMacDaemon:DP:phi_stmt_1250:output LSTATE_1250= " & Convert_SLV_To_Hex_String(LSTATE_1250));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1250: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nLSTATE_1264_1252_buffered & R_S0_1253_wire_constant;
      req <= phi_stmt_1250_req_0 & phi_stmt_1250_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1250",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1250_ack_0,
          idata => idata,
          odata => LSTATE_1250,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1250
    -- logger for split-operator MUX_1284_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if MUX_1284_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:MUX_1284_inst:started:   inputs: " & " write_to_header_1273 (guard)= " & Convert_SLV_To_String(write_to_header_1273) & " EQ_u2_u1_1278_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_1278_wire) & " CONCAT_u65_u73_1282_wire = "& Convert_SLV_To_Hex_String(CONCAT_u65_u73_1282_wire) & " RX_1254 = "& Convert_SLV_To_Hex_String(RX_1254));
          --
        end if; 
        if MUX_1284_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:MUX_1284_inst:finished:  outputs: " & " MUX_1284_wire= "  & Convert_SLV_To_Hex_String(MUX_1284_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    MUX_1284_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= MUX_1284_inst_req_0;
      MUX_1284_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= MUX_1284_inst_req_1;
      MUX_1284_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  write_to_header_1273(0);
      MUX_1284_inst_gI: SplitGuardInterface generic map(name => "MUX_1284_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      MUX_1284_inst: SelectSplitProtocol generic map(name => "MUX_1284_inst", data_width => 73, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u65_u73_1282_wire, y => RX_1254, sel => EQ_u2_u1_1278_wire, z => MUX_1284_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_1280_inst flow-through 
    process(slice_1280_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:slice_1280_inst:flowthrough inputs: " & " write_to_header_1273 (guard)= " & Convert_SLV_To_String(write_to_header_1273) & " RX_1254 = "& Convert_SLV_To_Hex_String(RX_1254) & " outputs:" & " slice_1280_wire= "  & Convert_SLV_To_Hex_String(slice_1280_wire));
      --
    end process; 
    -- flow-through slice operator slice_1280_inst
    slice_1280_wire <= RX_1254(72 downto 8);
    -- logger for split-operator nLSTATE_1264_1252_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nLSTATE_1264_1252_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:nLSTATE_1264_1252_buf:started:   inputs: " & " nLSTATE_1264 = "& Convert_SLV_To_Hex_String(nLSTATE_1264));
          --
        end if; 
        if nLSTATE_1264_1252_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:nLSTATE_1264_1252_buf:finished:  outputs: " & " nLSTATE_1264_1252_buffered= "  & Convert_SLV_To_Hex_String(nLSTATE_1264_1252_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nLSTATE_1264_1252_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nLSTATE_1264_1252_buf_req_0;
      nLSTATE_1264_1252_buf_ack_0<= wack(0);
      rreq(0) <= nLSTATE_1264_1252_buf_req_1;
      nLSTATE_1264_1252_buf_ack_1<= rack(0);
      nLSTATE_1264_1252_buf : InterlockBuffer generic map ( -- 
        name => "nLSTATE_1264_1252_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nLSTATE_1264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nLSTATE_1264_1252_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator ssrc_phi_stmt_1254 flow-through 
    process(RX_1254) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:ssrc_phi_stmt_1254:flowthrough inputs: " & " RPIPE_mac_to_nic_data_1256_wire = "& Convert_SLV_To_Hex_String(RPIPE_mac_to_nic_data_1256_wire) & " outputs:" & " RX_1254= "  & Convert_SLV_To_Hex_String(RX_1254));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1254
    process(RPIPE_mac_to_nic_data_1256_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_mac_to_nic_data_1256_wire(72 downto 0);
      RX_1254 <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1248_branch_req_0," req0 do_while_stmt_1248_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1248_branch_ack_0," ack0 do_while_stmt_1248_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1248_branch_ack_1," ack1 do_while_stmt_1248_branch");
    do_while_stmt_1248_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1292_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1248_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1248_branch_req_0,
          ack0 => do_while_stmt_1248_branch_ack_0,
          ack1 => do_while_stmt_1248_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator CONCAT_u65_u73_1282_inst flow-through 
    process(CONCAT_u65_u73_1282_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:CONCAT_u65_u73_1282_inst:flowthrough inputs: " & " write_to_header_1273 (guard)= " & Convert_SLV_To_String(write_to_header_1273) & " slice_1280_wire = "& Convert_SLV_To_Hex_String(slice_1280_wire) & " R_HEADER_TKEEP_1281_wire_constant = "& Convert_SLV_To_Hex_String(R_HEADER_TKEEP_1281_wire_constant) & " outputs:" & " CONCAT_u65_u73_1282_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u65_u73_1282_wire));
      --
    end process; 
    -- binary operator CONCAT_u65_u73_1282_inst
    process(slice_1280_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1280_wire, R_HEADER_TKEEP_1281_wire_constant, tmp_var);
      CONCAT_u65_u73_1282_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1268_inst flow-through 
    process(EQ_u2_u1_1268_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:EQ_u2_u1_1268_inst:flowthrough inputs: " & " LSTATE_1250 = "& Convert_SLV_To_Hex_String(LSTATE_1250) & " R_S0_1267_wire_constant = "& Convert_SLV_To_Hex_String(R_S0_1267_wire_constant) & " outputs:" & " EQ_u2_u1_1268_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1268_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1268_inst
    process(LSTATE_1250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1250, R_S0_1267_wire_constant, tmp_var);
      EQ_u2_u1_1268_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1271_inst flow-through 
    process(EQ_u2_u1_1271_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:EQ_u2_u1_1271_inst:flowthrough inputs: " & " LSTATE_1250 = "& Convert_SLV_To_Hex_String(LSTATE_1250) & " R_S1_1270_wire_constant = "& Convert_SLV_To_Hex_String(R_S1_1270_wire_constant) & " outputs:" & " EQ_u2_u1_1271_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1271_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1271_inst
    process(LSTATE_1250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1250, R_S1_1270_wire_constant, tmp_var);
      EQ_u2_u1_1271_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u2_u1_1278_inst flow-through 
    process(EQ_u2_u1_1278_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:EQ_u2_u1_1278_inst:flowthrough inputs: " & " write_to_header_1273 (guard)= " & Convert_SLV_To_String(write_to_header_1273) & " LSTATE_1250 = "& Convert_SLV_To_Hex_String(LSTATE_1250) & " R_S1_1277_wire_constant = "& Convert_SLV_To_Hex_String(R_S1_1277_wire_constant) & " outputs:" & " EQ_u2_u1_1278_wire= "  & Convert_SLV_To_Hex_String(EQ_u2_u1_1278_wire));
      --
    end process; 
    -- binary operator EQ_u2_u1_1278_inst
    process(LSTATE_1250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_1250, R_S1_1277_wire_constant, tmp_var);
      EQ_u2_u1_1278_wire <= tmp_var; --
    end process;
    -- logger for split-operator OR_u1_u1_1272_inst flow-through 
    process(write_to_header_1273) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:OR_u1_u1_1272_inst:flowthrough inputs: " & " EQ_u2_u1_1268_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_1268_wire) & " EQ_u2_u1_1271_wire = "& Convert_SLV_To_Hex_String(EQ_u2_u1_1271_wire) & " outputs:" & " write_to_header_1273= "  & Convert_SLV_To_Hex_String(write_to_header_1273));
      --
    end process; 
    -- binary operator OR_u1_u1_1272_inst
    process(EQ_u2_u1_1268_wire, EQ_u2_u1_1271_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_1268_wire, EQ_u2_u1_1271_wire, tmp_var);
      write_to_header_1273 <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_mac_to_nic_data_1256_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_mac_to_nic_data_1256_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:RPIPE_mac_to_nic_data_1256_inst:started:   PipeRead from mac_to_nic_data inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_mac_to_nic_data_1256_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:RPIPE_mac_to_nic_data_1256_inst:finished:  outputs: " & " RPIPE_mac_to_nic_data_1256_wire= "  & Convert_SLV_To_Hex_String(RPIPE_mac_to_nic_data_1256_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_mac_to_nic_data_1256_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_1256_inst_req_0;
      RPIPE_mac_to_nic_data_1256_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_1256_inst_req_1;
      RPIPE_mac_to_nic_data_1256_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_1256_wire <= data_out(72 downto 0);
      mac_to_nic_data_read_0_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_read_0: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_pipe_read_req(0),
          oack => mac_to_nic_data_pipe_read_ack(0),
          odata => mac_to_nic_data_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_nic_rx_to_header_1275_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_nic_rx_to_header_1275_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:WPIPE_nic_rx_to_header_1275_inst:started:   PipeWrite to nic_rx_to_header inputs: " & " write_to_header_1273 (guard)= " & Convert_SLV_To_String(write_to_header_1273) & " MUX_1284_wire = "& Convert_SLV_To_Hex_String(MUX_1284_wire));
          --
        end if; 
        if WPIPE_nic_rx_to_header_1275_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:WPIPE_nic_rx_to_header_1275_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_nic_rx_to_header_1275_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_header_1275_inst_req_0;
      WPIPE_nic_rx_to_header_1275_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_header_1275_inst_req_1;
      WPIPE_nic_rx_to_header_1275_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_to_header_1273(0);
      data_in <= MUX_1284_wire;
      nic_rx_to_header_write_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_write_0: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_header", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_header_pipe_write_req(0),
          oack => nic_rx_to_header_pipe_write_ack(0),
          odata => nic_rx_to_header_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_nic_rx_to_packet_1286_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_nic_rx_to_packet_1286_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:WPIPE_nic_rx_to_packet_1286_inst:started:   PipeWrite to nic_rx_to_packet inputs: " & " RX_1254 = "& Convert_SLV_To_Hex_String(RX_1254));
          --
        end if; 
        if WPIPE_nic_rx_to_packet_1286_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:WPIPE_nic_rx_to_packet_1286_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_nic_rx_to_packet_1286_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1286_inst_req_0;
      WPIPE_nic_rx_to_packet_1286_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_packet_1286_inst_req_1;
      WPIPE_nic_rx_to_packet_1286_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= RX_1254;
      nic_rx_to_packet_write_1_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_write_1: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_packet", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_packet_pipe_write_req(0),
          oack => nic_rx_to_packet_pipe_write_ack(0),
          odata => nic_rx_to_packet_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator call_stmt_1264_call flow-through 
    process(nLSTATE_1264) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicRxFromMacDaemon:DP:call_stmt_1264_call:flowthrough inputs: " & " RX_1254 = "& Convert_SLV_To_Hex_String(RX_1254) & " LSTATE_1250 = "& Convert_SLV_To_Hex_String(LSTATE_1250) & " outputs:" & " nLSTATE_1264= "  & Convert_SLV_To_Hex_String(nLSTATE_1264));
      --
    end process; 
    volatile_operator_nextLSTATE_3543: nextLSTATE_Volatile port map(RX => RX_1254, LSTATE => LSTATE_1250, nLSTATE => nLSTATE_1264, clk => clk, reset => reset); 
    -- 
  end Block; -- data_path
  -- 
end nicRxFromMacDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity nicToMacInterface is -- 
  generic (tag_length : integer); 
  port ( -- 
    nic_to_mac_transmit_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_data : in   std_logic_vector(72 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicToMacInterface;
architecture nicToMacInterface_arch of nicToMacInterface is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicToMacInterface_CP_2508_start: Boolean;
  signal nicToMacInterface_CP_2508_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_1 : boolean;
  signal type_cast_1310_inst_ack_0 : boolean;
  signal RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_1 : boolean;
  signal do_while_stmt_1297_branch_ack_0 : boolean;
  signal type_cast_1310_inst_req_0 : boolean;
  signal do_while_stmt_1297_branch_ack_1 : boolean;
  signal type_cast_1310_inst_req_1 : boolean;
  signal slice_1305_inst_ack_1 : boolean;
  signal slice_1305_inst_req_1 : boolean;
  signal slice_1305_inst_ack_0 : boolean;
  signal type_cast_1310_inst_ack_1 : boolean;
  signal RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_0 : boolean;
  signal slice_1305_inst_req_0 : boolean;
  signal do_while_stmt_1297_branch_req_0 : boolean;
  signal RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicToMacInterface_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicToMacInterface_CP_2508_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicToMacInterface_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicToMacInterface_CP_2508_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicToMacInterface_CP_2508_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicToMacInterface_CP_2508_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,nicToMacInterface_CP_2508_start,"nicToMacInterface cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,nicToMacInterface_CP_2508_symbol, "nicToMacInterface cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicToMacInterface_CP_2508: Block -- control-path 
    signal nicToMacInterface_CP_2508_elements: BooleanArray(29 downto 0);
    -- 
  begin -- 
    nicToMacInterface_CP_2508_elements(0) <= nicToMacInterface_CP_2508_start;
    nicToMacInterface_CP_2508_symbol <= nicToMacInterface_CP_2508_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1296/do_while_stmt_1297__entry__
      -- CP-element group 0: 	 branch_block_stmt_1296/branch_block_stmt_1296__entry__
      -- CP-element group 0: 	 branch_block_stmt_1296/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	29 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1296/do_while_stmt_1297__exit__
      -- CP-element group 1: 	 branch_block_stmt_1296/$exit
      -- CP-element group 1: 	 branch_block_stmt_1296/branch_block_stmt_1296__exit__
      -- CP-element group 1: 	 $exit
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_CP_2508_elements(1) <= nicToMacInterface_CP_2508_elements(29);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1296/do_while_stmt_1297/$entry
      -- CP-element group 2: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297__entry__
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_CP_2508_elements(2) <= nicToMacInterface_CP_2508_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	29 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297__exit__
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMacInterface_CP_2508_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_back
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMacInterface_CP_2508_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	27 
    -- CP-element group 5: 	28 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1296/do_while_stmt_1297/condition_done
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_CP_2508_elements(5) <= nicToMacInterface_CP_2508_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	26 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_body_done
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_CP_2508_elements(6) <= nicToMacInterface_CP_2508_elements(26);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_CP_2508_elements(7) <= nicToMacInterface_CP_2508_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_CP_2508_elements(8) <= nicToMacInterface_CP_2508_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	25 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/phi_stmt_1299_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/loop_body_start
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMacInterface_CP_2508_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	25 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/condition_evaluated
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:do_while_stmt_1297_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMacInterface_CP_2508_elements(10), ack => do_while_stmt_1297_branch_req_0); -- 
    nicToMacInterface_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(16) & nicToMacInterface_CP_2508_elements(25);
      gj_nicToMacInterface_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(9) & nicToMacInterface_CP_2508_elements(16);
      gj_nicToMacInterface_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	23 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/phi_stmt_1299_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(9) & nicToMacInterface_CP_2508_elements(19) & nicToMacInterface_CP_2508_elements(23);
      gj_nicToMacInterface_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Sample/rr
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMacInterface_CP_2508_elements(13), ack => RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_0); -- 
    nicToMacInterface_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(11) & nicToMacInterface_CP_2508_elements(16);
      gj_nicToMacInterface_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_update_start_
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMacInterface_CP_2508_elements(14), ack => RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_1); -- 
    nicToMacInterface_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(15) & nicToMacInterface_CP_2508_elements(12);
      gj_nicToMacInterface_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	14 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/phi_stmt_1299_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/aggregated_phi_sample_ack
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_0, ack => nicToMacInterface_CP_2508_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16: 	21 
    -- CP-element group 16: 	10 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/RPIPE_nic_to_mac_transmit_pipe_1301_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/phi_stmt_1299_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_1, ack => nicToMacInterface_CP_2508_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_sample_start_
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:slice_1305_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMacInterface_CP_2508_elements(17), ack => slice_1305_inst_req_0); -- 
    nicToMacInterface_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(16) & nicToMacInterface_CP_2508_elements(19);
      gj_nicToMacInterface_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_update_start_
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:slice_1305_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMacInterface_CP_2508_elements(18), ack => slice_1305_inst_req_1); -- 
    nicToMacInterface_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicToMacInterface_CP_2508_elements(20);
      gj_nicToMacInterface_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_sample_completed_
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:slice_1305_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1305_inst_ack_0, ack => nicToMacInterface_CP_2508_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	26 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/slice_1305_update_completed_
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:slice_1305_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1305_inst_ack_1, ack => nicToMacInterface_CP_2508_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_sample_start_
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:type_cast_1310_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMacInterface_CP_2508_elements(21), ack => type_cast_1310_inst_req_0); -- 
    nicToMacInterface_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(16) & nicToMacInterface_CP_2508_elements(23);
      gj_nicToMacInterface_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Update/cr
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:type_cast_1310_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMacInterface_CP_2508_elements(22), ack => type_cast_1310_inst_req_1); -- 
    nicToMacInterface_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicToMacInterface_CP_2508_elements(24);
      gj_nicToMacInterface_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	12 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_sample_completed_
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:type_cast_1310_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_0, ack => nicToMacInterface_CP_2508_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/type_cast_1310_Update/ca
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:type_cast_1310_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1310_inst_ack_1, ack => nicToMacInterface_CP_2508_elements(24)); -- 
    -- CP-element group 25:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	9 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	10 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMacInterface_CP_2508_elements(25) is a control-delay.
    cp_element_25_delay: control_delay_element  generic map(name => " 25_delay", delay_value => 1)  port map(req => nicToMacInterface_CP_2508_elements(9), ack => nicToMacInterface_CP_2508_elements(25), clk => clk, reset =>reset);
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: 	15 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	6 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1296/do_while_stmt_1297/do_while_stmt_1297_loop_body/$exit
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(26) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "nicToMacInterface_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicToMacInterface_CP_2508_elements(20) & nicToMacInterface_CP_2508_elements(15) & nicToMacInterface_CP_2508_elements(24);
      gj_nicToMacInterface_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	5 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_exit/ack
      -- CP-element group 27: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_exit/$exit
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:do_while_stmt_1297_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1297_branch_ack_0, ack => nicToMacInterface_CP_2508_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	5 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_taken/$exit
      -- CP-element group 28: 	 branch_block_stmt_1296/do_while_stmt_1297/loop_taken/ack
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:do_while_stmt_1297_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1297_branch_ack_1, ack => nicToMacInterface_CP_2508_elements(28)); -- 
    -- CP-element group 29:  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	3 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	1 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1296/do_while_stmt_1297/$exit
      -- 
    -- logger for CP element group nicToMacInterface_CP_2508_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMacInterface_CP_2508_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMacInterface:CP:nicToMacInterface_CP_2508_elements(29) fired."); 
        -- 
      end if; --
    end process; 
    nicToMacInterface_CP_2508_elements(29) <= nicToMacInterface_CP_2508_elements(3);
    nicToMacInterface_do_while_stmt_1297_terminator_2593: loop_terminator -- 
      generic map (name => " nicToMacInterface_do_while_stmt_1297_terminator_2593", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicToMacInterface_CP_2508_elements(6),loop_continue => nicToMacInterface_CP_2508_elements(28),loop_terminate => nicToMacInterface_CP_2508_elements(27),loop_back => nicToMacInterface_CP_2508_elements(4),loop_exit => nicToMacInterface_CP_2508_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_2533_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicToMacInterface_CP_2508_elements(7);
        preds(1)  <= nicToMacInterface_CP_2508_elements(8);
        entry_tmerge_2533 : transition_merge -- 
          generic map(name => " entry_tmerge_2533")
          port map (preds => preds, symbol_out => nicToMacInterface_CP_2508_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_nic_to_mac_transmit_pipe_1301_wire : std_logic_vector(72 downto 0);
    signal konst_1313_wire_constant : std_logic_vector(0 downto 0);
    signal nic_to_mac_data0_1306 : std_logic_vector(63 downto 0);
    signal nic_to_mac_data1_1311 : std_logic_vector(15 downto 0);
    signal rdata_1299 : std_logic_vector(72 downto 0);
    signal slice_1309_wire : std_logic_vector(8 downto 0);
    -- 
  begin -- 
    konst_1313_wire_constant <= "1";
    -- logger for split-operator slice_1305_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_1305_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:slice_1305_inst:started:   inputs: " & " rdata_1299 = "& Convert_SLV_To_Hex_String(rdata_1299));
          --
        end if; 
        if slice_1305_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:slice_1305_inst:finished:  outputs: " & " nic_to_mac_data0_1306= "  & Convert_SLV_To_Hex_String(nic_to_mac_data0_1306));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_1305_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1305_inst_req_0;
      slice_1305_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1305_inst_req_1;
      slice_1305_inst_ack_1<= update_ack(0);
      slice_1305_inst: SliceSplitProtocol generic map(name => "slice_1305_inst", in_data_width => 73, high_index => 63, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdata_1299, dout => nic_to_mac_data0_1306, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_1309_inst flow-through 
    process(slice_1309_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:slice_1309_inst:flowthrough inputs: " & " rdata_1299 = "& Convert_SLV_To_Hex_String(rdata_1299) & " outputs:" & " slice_1309_wire= "  & Convert_SLV_To_Hex_String(slice_1309_wire));
      --
    end process; 
    -- flow-through slice operator slice_1309_inst
    slice_1309_wire <= rdata_1299(8 downto 0);
    -- logger for split-operator ssrc_phi_stmt_1299 flow-through 
    process(rdata_1299) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:ssrc_phi_stmt_1299:flowthrough inputs: " & " RPIPE_nic_to_mac_transmit_pipe_1301_wire = "& Convert_SLV_To_Hex_String(RPIPE_nic_to_mac_transmit_pipe_1301_wire) & " outputs:" & " rdata_1299= "  & Convert_SLV_To_Hex_String(rdata_1299));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1299
    process(RPIPE_nic_to_mac_transmit_pipe_1301_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_to_mac_transmit_pipe_1301_wire(72 downto 0);
      rdata_1299 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1310_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1310_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:type_cast_1310_inst:started:   inputs: " & " slice_1309_wire = "& Convert_SLV_To_Hex_String(slice_1309_wire));
          --
        end if; 
        if type_cast_1310_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:type_cast_1310_inst:finished:  outputs: " & " nic_to_mac_data1_1311= "  & Convert_SLV_To_Hex_String(nic_to_mac_data1_1311));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1310_inst_req_0;
      type_cast_1310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1310_inst_req_1;
      type_cast_1310_inst_ack_1<= rack(0);
      type_cast_1310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 9,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => slice_1309_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nic_to_mac_data1_1311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1297_branch_req_0," req0 do_while_stmt_1297_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1297_branch_ack_0," ack0 do_while_stmt_1297_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1297_branch_ack_1," ack1 do_while_stmt_1297_branch");
    do_while_stmt_1297_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1313_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1297_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1297_branch_req_0,
          ack0 => do_while_stmt_1297_branch_ack_0,
          ack1 => do_while_stmt_1297_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_nic_to_mac_transmit_pipe_1301_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:RPIPE_nic_to_mac_transmit_pipe_1301_inst:started:   PipeRead from nic_to_mac_transmit_pipe inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMacInterface:DP:RPIPE_nic_to_mac_transmit_pipe_1301_inst:finished:  outputs: " & " RPIPE_nic_to_mac_transmit_pipe_1301_wire= "  & Convert_SLV_To_Hex_String(RPIPE_nic_to_mac_transmit_pipe_1301_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_nic_to_mac_transmit_pipe_1301_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_0;
      RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_to_mac_transmit_pipe_1301_inst_req_1;
      RPIPE_nic_to_mac_transmit_pipe_1301_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_to_mac_transmit_pipe_1301_wire <= data_out(72 downto 0);
      nic_to_mac_transmit_pipe_read_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_read_0: InputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_to_mac_transmit_pipe_pipe_read_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_read_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end nicToMacInterface_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity nicToMemoryInterface is -- 
  generic (tag_length : integer); 
  port ( -- 
    NIC_TO_MEMORY_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_data : in   std_logic_vector(109 downto 0);
    mem_req0_pipe0_pipe_write_req : out  std_logic_vector(0 downto 0);
    mem_req0_pipe0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    mem_req0_pipe0_pipe_write_data : out  std_logic_vector(63 downto 0);
    mem_req0_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    mem_req0_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    mem_req0_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicToMemoryInterface;
architecture nicToMemoryInterface_arch of nicToMemoryInterface is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicToMemoryInterface_CP_2594_start: Boolean;
  signal nicToMemoryInterface_CP_2594_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_mem_req0_pipe0_1324_inst_req_0 : boolean;
  signal WPIPE_mem_req0_pipe0_1324_inst_ack_0 : boolean;
  signal RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_0 : boolean;
  signal type_cast_1332_inst_req_0 : boolean;
  signal type_cast_1332_inst_ack_0 : boolean;
  signal WPIPE_mem_req0_pipe0_1324_inst_ack_1 : boolean;
  signal WPIPE_mem_req0_pipe0_1324_inst_req_1 : boolean;
  signal do_while_stmt_1318_branch_ack_1 : boolean;
  signal do_while_stmt_1318_branch_ack_0 : boolean;
  signal WPIPE_mem_req0_pipe1_1328_inst_ack_1 : boolean;
  signal WPIPE_mem_req0_pipe1_1328_inst_req_1 : boolean;
  signal do_while_stmt_1318_branch_req_0 : boolean;
  signal WPIPE_mem_req0_pipe1_1328_inst_ack_0 : boolean;
  signal WPIPE_mem_req0_pipe1_1328_inst_req_0 : boolean;
  signal slice_1326_inst_ack_1 : boolean;
  signal slice_1326_inst_req_1 : boolean;
  signal type_cast_1332_inst_ack_1 : boolean;
  signal type_cast_1332_inst_req_1 : boolean;
  signal slice_1326_inst_ack_0 : boolean;
  signal slice_1326_inst_req_0 : boolean;
  signal RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_1 : boolean;
  signal RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_1 : boolean;
  signal RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicToMemoryInterface_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicToMemoryInterface_CP_2594_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicToMemoryInterface_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicToMemoryInterface_CP_2594_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicToMemoryInterface_CP_2594_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicToMemoryInterface_CP_2594_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,nicToMemoryInterface_CP_2594_start,"nicToMemoryInterface cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,nicToMemoryInterface_CP_2594_symbol, "nicToMemoryInterface cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicToMemoryInterface_CP_2594: Block -- control-path 
    signal nicToMemoryInterface_CP_2594_elements: BooleanArray(35 downto 0);
    -- 
  begin -- 
    nicToMemoryInterface_CP_2594_elements(0) <= nicToMemoryInterface_CP_2594_start;
    nicToMemoryInterface_CP_2594_symbol <= nicToMemoryInterface_CP_2594_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1317/do_while_stmt_1318__entry__
      -- CP-element group 0: 	 branch_block_stmt_1317/branch_block_stmt_1317__entry__
      -- CP-element group 0: 	 branch_block_stmt_1317/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	35 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1317/do_while_stmt_1318__exit__
      -- CP-element group 1: 	 branch_block_stmt_1317/branch_block_stmt_1317__exit__
      -- CP-element group 1: 	 branch_block_stmt_1317/$exit
      -- CP-element group 1: 	 $exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_CP_2594_elements(1) <= nicToMemoryInterface_CP_2594_elements(35);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1317/do_while_stmt_1318/$entry
      -- CP-element group 2: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318__entry__
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_CP_2594_elements(2) <= nicToMemoryInterface_CP_2594_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	35 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318__exit__
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMemoryInterface_CP_2594_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_back
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMemoryInterface_CP_2594_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	34 
    -- CP-element group 5: 	33 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1317/do_while_stmt_1318/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_exit/$entry
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_CP_2594_elements(5) <= nicToMemoryInterface_CP_2594_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	32 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_body_done
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_CP_2594_elements(6) <= nicToMemoryInterface_CP_2594_elements(32);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_CP_2594_elements(7) <= nicToMemoryInterface_CP_2594_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_CP_2594_elements(8) <= nicToMemoryInterface_CP_2594_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/phi_stmt_1320_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/$entry
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMemoryInterface_CP_2594_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	31 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/condition_evaluated
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:do_while_stmt_1318_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(10), ack => do_while_stmt_1318_branch_req_0); -- 
    nicToMemoryInterface_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(16) & nicToMemoryInterface_CP_2594_elements(31);
      gj_nicToMemoryInterface_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(9) & nicToMemoryInterface_CP_2594_elements(16);
      gj_nicToMemoryInterface_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	26 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/phi_stmt_1320_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(9) & nicToMemoryInterface_CP_2594_elements(19) & nicToMemoryInterface_CP_2594_elements(26);
      gj_nicToMemoryInterface_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_sample_start_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(13), ack => RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_0); -- 
    nicToMemoryInterface_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(11) & nicToMemoryInterface_CP_2594_elements(16);
      gj_nicToMemoryInterface_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Update/$entry
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(14), ack => RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_1); -- 
    nicToMemoryInterface_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(15) & nicToMemoryInterface_CP_2594_elements(12);
      gj_nicToMemoryInterface_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	32 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/phi_stmt_1320_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/aggregated_phi_sample_ack
      -- CP-element group 15: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Sample/ra
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_0, ack => nicToMemoryInterface_CP_2594_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16: 	24 
    -- CP-element group 16: 	10 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/phi_stmt_1320_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/aggregated_phi_update_ack
      -- CP-element group 16: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/RPIPE_NIC_TO_MEMORY_REQUEST_1322_Update/$exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_1, ack => nicToMemoryInterface_CP_2594_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_sample_start_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:slice_1326_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(17), ack => slice_1326_inst_req_0); -- 
    nicToMemoryInterface_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(16) & nicToMemoryInterface_CP_2594_elements(19);
      gj_nicToMemoryInterface_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_update_start_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:slice_1326_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(18), ack => slice_1326_inst_req_1); -- 
    nicToMemoryInterface_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicToMemoryInterface_CP_2594_elements(22);
      gj_nicToMemoryInterface_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_sample_completed_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:slice_1326_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1326_inst_ack_0, ack => nicToMemoryInterface_CP_2594_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/slice_1326_update_completed_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:slice_1326_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1326_inst_ack_1, ack => nicToMemoryInterface_CP_2594_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Sample/req
      -- CP-element group 21: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_sample_start_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe0_1324_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(21), ack => WPIPE_mem_req0_pipe0_1324_inst_req_0); -- 
    nicToMemoryInterface_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(20) & nicToMemoryInterface_CP_2594_elements(23);
      gj_nicToMemoryInterface_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Sample/ack
      -- CP-element group 22: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Update/req
      -- CP-element group 22: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Update/$entry
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe0_1324_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe0_1324_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mem_req0_pipe0_1324_inst_ack_0, ack => nicToMemoryInterface_CP_2594_elements(22)); -- 
    req_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(22), ack => WPIPE_mem_req0_pipe0_1324_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	32 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Update/ack
      -- CP-element group 23: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe0_1324_Update/$exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe0_1324_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mem_req0_pipe0_1324_inst_ack_1, ack => nicToMemoryInterface_CP_2594_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	16 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_sample_start_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:type_cast_1332_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(24), ack => type_cast_1332_inst_req_0); -- 
    nicToMemoryInterface_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(16) & nicToMemoryInterface_CP_2594_elements(26);
      gj_nicToMemoryInterface_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Update/$entry
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:type_cast_1332_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(25), ack => type_cast_1332_inst_req_1); -- 
    nicToMemoryInterface_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicToMemoryInterface_CP_2594_elements(29);
      gj_nicToMemoryInterface_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	12 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Sample/ra
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:type_cast_1332_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_0, ack => nicToMemoryInterface_CP_2594_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/type_cast_1332_Update/$exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:type_cast_1332_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1332_inst_ack_1, ack => nicToMemoryInterface_CP_2594_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Sample/$entry
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe1_1328_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(28), ack => WPIPE_mem_req0_pipe1_1328_inst_req_0); -- 
    nicToMemoryInterface_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(27) & nicToMemoryInterface_CP_2594_elements(30);
      gj_nicToMemoryInterface_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Update/req
      -- CP-element group 29: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_update_start_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe1_1328_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe1_1328_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mem_req0_pipe1_1328_inst_ack_0, ack => nicToMemoryInterface_CP_2594_elements(29)); -- 
    req_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToMemoryInterface_CP_2594_elements(29), ack => WPIPE_mem_req0_pipe1_1328_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Update/ack
      -- CP-element group 30: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/WPIPE_mem_req0_pipe1_1328_update_completed_
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:WPIPE_mem_req0_pipe1_1328_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_mem_req0_pipe1_1328_inst_ack_1, ack => nicToMemoryInterface_CP_2594_elements(30)); -- 
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	10 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToMemoryInterface_CP_2594_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => nicToMemoryInterface_CP_2594_elements(9), ack => nicToMemoryInterface_CP_2594_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	15 
    -- CP-element group 32: 	30 
    -- CP-element group 32: 	23 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	6 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1317/do_while_stmt_1318/do_while_stmt_1318_loop_body/$exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(32) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "nicToMemoryInterface_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicToMemoryInterface_CP_2594_elements(15) & nicToMemoryInterface_CP_2594_elements(30) & nicToMemoryInterface_CP_2594_elements(23);
      gj_nicToMemoryInterface_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	5 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_exit/ack
      -- CP-element group 33: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_exit/$exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:do_while_stmt_1318_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1318_branch_ack_0, ack => nicToMemoryInterface_CP_2594_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	5 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_taken/ack
      -- CP-element group 34: 	 branch_block_stmt_1317/do_while_stmt_1318/loop_taken/$exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:do_while_stmt_1318_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1318_branch_ack_1, ack => nicToMemoryInterface_CP_2594_elements(34)); -- 
    -- CP-element group 35:  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	3 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	1 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1317/do_while_stmt_1318/$exit
      -- 
    -- logger for CP element group nicToMemoryInterface_CP_2594_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToMemoryInterface_CP_2594_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToMemoryInterface:CP:nicToMemoryInterface_CP_2594_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    nicToMemoryInterface_CP_2594_elements(35) <= nicToMemoryInterface_CP_2594_elements(3);
    nicToMemoryInterface_do_while_stmt_1318_terminator_2707: loop_terminator -- 
      generic map (name => " nicToMemoryInterface_do_while_stmt_1318_terminator_2707", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicToMemoryInterface_CP_2594_elements(6),loop_continue => nicToMemoryInterface_CP_2594_elements(34),loop_terminate => nicToMemoryInterface_CP_2594_elements(33),loop_back => nicToMemoryInterface_CP_2594_elements(4),loop_exit => nicToMemoryInterface_CP_2594_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_2619_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicToMemoryInterface_CP_2594_elements(7);
        preds(1)  <= nicToMemoryInterface_CP_2594_elements(8);
        entry_tmerge_2619 : transition_merge -- 
          generic map(name => " entry_tmerge_2619")
          port map (preds => preds, symbol_out => nicToMemoryInterface_CP_2594_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire : std_logic_vector(109 downto 0);
    signal konst_1335_wire_constant : std_logic_vector(0 downto 0);
    signal rdata_1320 : std_logic_vector(109 downto 0);
    signal slice_1326_wire : std_logic_vector(63 downto 0);
    signal slice_1331_wire : std_logic_vector(45 downto 0);
    signal type_cast_1332_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1335_wire_constant <= "1";
    -- logger for split-operator slice_1326_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if slice_1326_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:slice_1326_inst:started:   inputs: " & " rdata_1320 = "& Convert_SLV_To_Hex_String(rdata_1320));
          --
        end if; 
        if slice_1326_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:slice_1326_inst:finished:  outputs: " & " slice_1326_wire= "  & Convert_SLV_To_Hex_String(slice_1326_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    slice_1326_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1326_inst_req_0;
      slice_1326_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1326_inst_req_1;
      slice_1326_inst_ack_1<= update_ack(0);
      slice_1326_inst: SliceSplitProtocol generic map(name => "slice_1326_inst", in_data_width => 110, high_index => 63, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => rdata_1320, dout => slice_1326_wire, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- logger for split-operator slice_1331_inst flow-through 
    process(slice_1331_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:slice_1331_inst:flowthrough inputs: " & " rdata_1320 = "& Convert_SLV_To_Hex_String(rdata_1320) & " outputs:" & " slice_1331_wire= "  & Convert_SLV_To_Hex_String(slice_1331_wire));
      --
    end process; 
    -- flow-through slice operator slice_1331_inst
    slice_1331_wire <= rdata_1320(45 downto 0);
    -- logger for split-operator ssrc_phi_stmt_1320 flow-through 
    process(rdata_1320) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:ssrc_phi_stmt_1320:flowthrough inputs: " & " RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire = "& Convert_SLV_To_Hex_String(RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire) & " outputs:" & " rdata_1320= "  & Convert_SLV_To_Hex_String(rdata_1320));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1320
    process(RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 109 downto 0) := RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire(109 downto 0);
      rdata_1320 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1332_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1332_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:type_cast_1332_inst:started:   inputs: " & " slice_1331_wire = "& Convert_SLV_To_Hex_String(slice_1331_wire));
          --
        end if; 
        if type_cast_1332_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:type_cast_1332_inst:finished:  outputs: " & " type_cast_1332_wire= "  & Convert_SLV_To_Hex_String(type_cast_1332_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1332_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1332_inst_req_0;
      type_cast_1332_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1332_inst_req_1;
      type_cast_1332_inst_ack_1<= rack(0);
      type_cast_1332_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1332_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 46,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => slice_1331_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1332_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1318_branch_req_0," req0 do_while_stmt_1318_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1318_branch_ack_0," ack0 do_while_stmt_1318_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1318_branch_ack_1," ack1 do_while_stmt_1318_branch");
    do_while_stmt_1318_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1335_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1318_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1318_branch_req_0,
          ack0 => do_while_stmt_1318_branch_ack_0,
          ack1 => do_while_stmt_1318_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst:started:   PipeRead from NIC_TO_MEMORY_REQUEST inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst:finished:  outputs: " & " RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire= "  & Convert_SLV_To_Hex_String(RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(109 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_0;
      RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_req_1;
      RPIPE_NIC_TO_MEMORY_REQUEST_1322_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_NIC_TO_MEMORY_REQUEST_1322_wire <= data_out(109 downto 0);
      NIC_TO_MEMORY_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST_read_0", data_width => 110,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_read_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_read_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_read_data(109 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_mem_req0_pipe0_1324_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_mem_req0_pipe0_1324_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:WPIPE_mem_req0_pipe0_1324_inst:started:   PipeWrite to mem_req0_pipe0 inputs: " & " slice_1326_wire = "& Convert_SLV_To_Hex_String(slice_1326_wire));
          --
        end if; 
        if WPIPE_mem_req0_pipe0_1324_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:WPIPE_mem_req0_pipe0_1324_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_mem_req0_pipe0_1324_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_mem_req0_pipe0_1324_inst_req_0;
      WPIPE_mem_req0_pipe0_1324_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_mem_req0_pipe0_1324_inst_req_1;
      WPIPE_mem_req0_pipe0_1324_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= slice_1326_wire;
      mem_req0_pipe0_write_0_gI: SplitGuardInterface generic map(name => "mem_req0_pipe0_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      mem_req0_pipe0_write_0: OutputPortRevised -- 
        generic map ( name => "mem_req0_pipe0", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => mem_req0_pipe0_pipe_write_req(0),
          oack => mem_req0_pipe0_pipe_write_ack(0),
          odata => mem_req0_pipe0_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_mem_req0_pipe1_1328_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_mem_req0_pipe1_1328_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:WPIPE_mem_req0_pipe1_1328_inst:started:   PipeWrite to mem_req0_pipe1 inputs: " & " type_cast_1332_wire = "& Convert_SLV_To_Hex_String(type_cast_1332_wire));
          --
        end if; 
        if WPIPE_mem_req0_pipe1_1328_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToMemoryInterface:DP:WPIPE_mem_req0_pipe1_1328_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_mem_req0_pipe1_1328_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_mem_req0_pipe1_1328_inst_req_0;
      WPIPE_mem_req0_pipe1_1328_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_mem_req0_pipe1_1328_inst_req_1;
      WPIPE_mem_req0_pipe1_1328_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1332_wire;
      mem_req0_pipe1_write_1_gI: SplitGuardInterface generic map(name => "mem_req0_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      mem_req0_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "mem_req0_pipe1", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => mem_req0_pipe1_pipe_write_req(0),
          oack => mem_req0_pipe1_pipe_write_ack(0),
          odata => mem_req0_pipe1_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end nicToMemoryInterface_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity nicToProcessorInterface is -- 
  generic (tag_length : integer); 
  port ( -- 
    AFB_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(32 downto 0);
    control_word_response_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    control_word_response_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    control_word_response_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicToProcessorInterface;
architecture nicToProcessorInterface_arch of nicToProcessorInterface is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicToProcessorInterface_CP_2708_start: Boolean;
  signal nicToProcessorInterface_CP_2708_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_AFB_NIC_RESPONSE_1344_inst_req_1 : boolean;
  signal do_while_stmt_1340_branch_ack_1 : boolean;
  signal WPIPE_control_word_response_pipe_1346_inst_req_1 : boolean;
  signal WPIPE_control_word_response_pipe_1346_inst_ack_1 : boolean;
  signal RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_RESPONSE_1344_inst_req_0 : boolean;
  signal type_cast_1348_inst_req_0 : boolean;
  signal WPIPE_control_word_response_pipe_1346_inst_ack_0 : boolean;
  signal do_while_stmt_1340_branch_req_0 : boolean;
  signal type_cast_1348_inst_ack_0 : boolean;
  signal type_cast_1348_inst_ack_1 : boolean;
  signal do_while_stmt_1340_branch_ack_0 : boolean;
  signal type_cast_1348_inst_req_1 : boolean;
  signal WPIPE_control_word_response_pipe_1346_inst_req_0 : boolean;
  signal RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicToProcessorInterface_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicToProcessorInterface_CP_2708_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicToProcessorInterface_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicToProcessorInterface_CP_2708_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicToProcessorInterface_CP_2708_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicToProcessorInterface_CP_2708_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,nicToProcessorInterface_CP_2708_start,"nicToProcessorInterface cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,nicToProcessorInterface_CP_2708_symbol, "nicToProcessorInterface cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicToProcessorInterface_CP_2708: Block -- control-path 
    signal nicToProcessorInterface_CP_2708_elements: BooleanArray(28 downto 0);
    -- 
  begin -- 
    nicToProcessorInterface_CP_2708_elements(0) <= nicToProcessorInterface_CP_2708_start;
    nicToProcessorInterface_CP_2708_symbol <= nicToProcessorInterface_CP_2708_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1339/$entry
      -- CP-element group 0: 	 branch_block_stmt_1339/branch_block_stmt_1339__entry__
      -- CP-element group 0: 	 branch_block_stmt_1339/do_while_stmt_1340__entry__
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	28 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1339/$exit
      -- CP-element group 1: 	 branch_block_stmt_1339/do_while_stmt_1340__exit__
      -- CP-element group 1: 	 branch_block_stmt_1339/branch_block_stmt_1339__exit__
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_CP_2708_elements(1) <= nicToProcessorInterface_CP_2708_elements(28);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1339/do_while_stmt_1340/$entry
      -- CP-element group 2: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340__entry__
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_CP_2708_elements(2) <= nicToProcessorInterface_CP_2708_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	28 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340__exit__
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToProcessorInterface_CP_2708_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_back
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToProcessorInterface_CP_2708_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	26 
    -- CP-element group 5: 	27 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1339/do_while_stmt_1340/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_taken/$entry
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_CP_2708_elements(5) <= nicToProcessorInterface_CP_2708_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	25 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_body_done
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_CP_2708_elements(6) <= nicToProcessorInterface_CP_2708_elements(25);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_CP_2708_elements(7) <= nicToProcessorInterface_CP_2708_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_CP_2708_elements(8) <= nicToProcessorInterface_CP_2708_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	24 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/phi_stmt_1342_sample_start_
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToProcessorInterface_CP_2708_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	24 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/condition_evaluated
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:do_while_stmt_1340_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToProcessorInterface_CP_2708_elements(10), ack => do_while_stmt_1340_branch_req_0); -- 
    nicToProcessorInterface_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(16) & nicToProcessorInterface_CP_2708_elements(24);
      gj_nicToProcessorInterface_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(9) & nicToProcessorInterface_CP_2708_elements(16);
      gj_nicToProcessorInterface_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	19 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/aggregated_phi_update_req
      -- CP-element group 12: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/phi_stmt_1342_update_start_
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(9) & nicToProcessorInterface_CP_2708_elements(19);
      gj_nicToProcessorInterface_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_sample_start_
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:RPIPE_AFB_NIC_RESPONSE_1344_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToProcessorInterface_CP_2708_elements(13), ack => RPIPE_AFB_NIC_RESPONSE_1344_inst_req_0); -- 
    nicToProcessorInterface_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(11) & nicToProcessorInterface_CP_2708_elements(16);
      gj_nicToProcessorInterface_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: 	15 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_update_start_
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:RPIPE_AFB_NIC_RESPONSE_1344_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToProcessorInterface_CP_2708_elements(14), ack => RPIPE_AFB_NIC_RESPONSE_1344_inst_req_1); -- 
    nicToProcessorInterface_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(12) & nicToProcessorInterface_CP_2708_elements(15);
      gj_nicToProcessorInterface_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	14 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/aggregated_phi_sample_ack
      -- CP-element group 15: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/phi_stmt_1342_sample_completed_
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_0, ack => nicToProcessorInterface_CP_2708_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: 	17 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/aggregated_phi_update_ack
      -- CP-element group 16: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/phi_stmt_1342_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/RPIPE_AFB_NIC_RESPONSE_1344_Update/ca
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_1, ack => nicToProcessorInterface_CP_2708_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_sample_start_
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:type_cast_1348_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToProcessorInterface_CP_2708_elements(17), ack => type_cast_1348_inst_req_0); -- 
    nicToProcessorInterface_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(16) & nicToProcessorInterface_CP_2708_elements(19);
      gj_nicToProcessorInterface_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Update/cr
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:type_cast_1348_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToProcessorInterface_CP_2708_elements(18), ack => type_cast_1348_inst_req_1); -- 
    nicToProcessorInterface_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicToProcessorInterface_CP_2708_elements(22);
      gj_nicToProcessorInterface_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_sample_completed_
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:type_cast_1348_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1348_inst_ack_0, ack => nicToProcessorInterface_CP_2708_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/type_cast_1348_Update/ca
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:type_cast_1348_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1348_inst_ack_1, ack => nicToProcessorInterface_CP_2708_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Sample/req
      -- CP-element group 21: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Sample/$entry
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:WPIPE_control_word_response_pipe_1346_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToProcessorInterface_CP_2708_elements(21), ack => WPIPE_control_word_response_pipe_1346_inst_req_0); -- 
    nicToProcessorInterface_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(20) & nicToProcessorInterface_CP_2708_elements(23);
      gj_nicToProcessorInterface_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Update/req
      -- CP-element group 22: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Sample/ack
      -- CP-element group 22: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Sample/$exit
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:WPIPE_control_word_response_pipe_1346_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:WPIPE_control_word_response_pipe_1346_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_control_word_response_pipe_1346_inst_ack_0, ack => nicToProcessorInterface_CP_2708_elements(22)); -- 
    req_2782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicToProcessorInterface_CP_2708_elements(22), ack => WPIPE_control_word_response_pipe_1346_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/WPIPE_control_word_response_pipe_1346_Update/ack
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:WPIPE_control_word_response_pipe_1346_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_control_word_response_pipe_1346_inst_ack_1, ack => nicToProcessorInterface_CP_2708_elements(23)); -- 
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	9 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	10 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group nicToProcessorInterface_CP_2708_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => nicToProcessorInterface_CP_2708_elements(9), ack => nicToProcessorInterface_CP_2708_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	6 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1339/do_while_stmt_1340/do_while_stmt_1340_loop_body/$exit
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "nicToProcessorInterface_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicToProcessorInterface_CP_2708_elements(15) & nicToProcessorInterface_CP_2708_elements(23);
      gj_nicToProcessorInterface_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	5 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_exit/$exit
      -- CP-element group 26: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_exit/ack
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:do_while_stmt_1340_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1340_branch_ack_0, ack => nicToProcessorInterface_CP_2708_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	5 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_taken/ack
      -- CP-element group 27: 	 branch_block_stmt_1339/do_while_stmt_1340/loop_taken/$exit
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:do_while_stmt_1340_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1340_branch_ack_1, ack => nicToProcessorInterface_CP_2708_elements(27)); -- 
    -- CP-element group 28:  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	3 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	1 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1339/do_while_stmt_1340/$exit
      -- 
    -- logger for CP element group nicToProcessorInterface_CP_2708_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and nicToProcessorInterface_CP_2708_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:nicToProcessorInterface:CP:nicToProcessorInterface_CP_2708_elements(28) fired."); 
        -- 
      end if; --
    end process; 
    nicToProcessorInterface_CP_2708_elements(28) <= nicToProcessorInterface_CP_2708_elements(3);
    nicToProcessorInterface_do_while_stmt_1340_terminator_2793: loop_terminator -- 
      generic map (name => " nicToProcessorInterface_do_while_stmt_1340_terminator_2793", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicToProcessorInterface_CP_2708_elements(6),loop_continue => nicToProcessorInterface_CP_2708_elements(27),loop_terminate => nicToProcessorInterface_CP_2708_elements(26),loop_back => nicToProcessorInterface_CP_2708_elements(4),loop_exit => nicToProcessorInterface_CP_2708_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_2733_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicToProcessorInterface_CP_2708_elements(7);
        preds(1)  <= nicToProcessorInterface_CP_2708_elements(8);
        entry_tmerge_2733 : transition_merge -- 
          generic map(name => " entry_tmerge_2733")
          port map (preds => preds, symbol_out => nicToProcessorInterface_CP_2708_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_AFB_NIC_RESPONSE_1344_wire : std_logic_vector(32 downto 0);
    signal konst_1351_wire_constant : std_logic_vector(0 downto 0);
    signal rdata_1342 : std_logic_vector(32 downto 0);
    signal type_cast_1348_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1351_wire_constant <= "1";
    -- logger for split-operator ssrc_phi_stmt_1342 flow-through 
    process(rdata_1342) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:nicToProcessorInterface:DP:ssrc_phi_stmt_1342:flowthrough inputs: " & " RPIPE_AFB_NIC_RESPONSE_1344_wire = "& Convert_SLV_To_Hex_String(RPIPE_AFB_NIC_RESPONSE_1344_wire) & " outputs:" & " rdata_1342= "  & Convert_SLV_To_Hex_String(rdata_1342));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1342
    process(RPIPE_AFB_NIC_RESPONSE_1344_wire) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 32 downto 0) := RPIPE_AFB_NIC_RESPONSE_1344_wire(32 downto 0);
      rdata_1342 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1348_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if type_cast_1348_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToProcessorInterface:DP:type_cast_1348_inst:started:   inputs: " & " rdata_1342 = "& Convert_SLV_To_Hex_String(rdata_1342));
          --
        end if; 
        if type_cast_1348_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToProcessorInterface:DP:type_cast_1348_inst:finished:  outputs: " & " type_cast_1348_wire= "  & Convert_SLV_To_Hex_String(type_cast_1348_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    type_cast_1348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1348_inst_req_0;
      type_cast_1348_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1348_inst_req_1;
      type_cast_1348_inst_ack_1<= rack(0);
      type_cast_1348_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 33,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rdata_1342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1348_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1340_branch_req_0," req0 do_while_stmt_1340_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1340_branch_ack_0," ack0 do_while_stmt_1340_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1340_branch_ack_1," ack1 do_while_stmt_1340_branch");
    do_while_stmt_1340_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1351_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1340_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1340_branch_req_0,
          ack0 => do_while_stmt_1340_branch_ack_0,
          ack1 => do_while_stmt_1340_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator RPIPE_AFB_NIC_RESPONSE_1344_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToProcessorInterface:DP:RPIPE_AFB_NIC_RESPONSE_1344_inst:started:   PipeRead from AFB_NIC_RESPONSE inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToProcessorInterface:DP:RPIPE_AFB_NIC_RESPONSE_1344_inst:finished:  outputs: " & " RPIPE_AFB_NIC_RESPONSE_1344_wire= "  & Convert_SLV_To_Hex_String(RPIPE_AFB_NIC_RESPONSE_1344_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_AFB_NIC_RESPONSE_1344_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_RESPONSE_1344_inst_req_0;
      RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_RESPONSE_1344_inst_req_1;
      RPIPE_AFB_NIC_RESPONSE_1344_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_AFB_NIC_RESPONSE_1344_wire <= data_out(32 downto 0);
      AFB_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_RESPONSE_pipe_read_req(0),
          oack => AFB_NIC_RESPONSE_pipe_read_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator WPIPE_control_word_response_pipe_1346_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_control_word_response_pipe_1346_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToProcessorInterface:DP:WPIPE_control_word_response_pipe_1346_inst:started:   PipeWrite to control_word_response_pipe inputs: " & " type_cast_1348_wire = "& Convert_SLV_To_Hex_String(type_cast_1348_wire));
          --
        end if; 
        if WPIPE_control_word_response_pipe_1346_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:nicToProcessorInterface:DP:WPIPE_control_word_response_pipe_1346_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_control_word_response_pipe_1346_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_control_word_response_pipe_1346_inst_req_0;
      WPIPE_control_word_response_pipe_1346_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_control_word_response_pipe_1346_inst_req_1;
      WPIPE_control_word_response_pipe_1346_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1348_wire;
      control_word_response_pipe_write_0_gI: SplitGuardInterface generic map(name => "control_word_response_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      control_word_response_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "control_word_response_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => control_word_response_pipe_pipe_write_req(0),
          oack => control_word_response_pipe_pipe_write_ack(0),
          odata => control_word_response_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end nicToProcessorInterface_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity popFromQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_call_data : out  std_logic_vector(67 downto 0);
    getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_return_data : in   std_logic_vector(31 downto 0);
    getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_call_data : out  std_logic_vector(35 downto 0);
    releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
    acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_call_data : out  std_logic_vector(35 downto 0);
    acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_return_data : in   std_logic_vector(0 downto 0);
    acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity popFromQueue;
architecture popFromQueue_arch of popFromQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 37)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal popFromQueue_CP_510_start: Boolean;
  signal popFromQueue_CP_510_symbol: Boolean;
  -- volatile/operator module components. 
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_pointer : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_462_call_ack_1 : boolean;
  signal call_stmt_492_call_req_0 : boolean;
  signal call_stmt_462_call_req_0 : boolean;
  signal call_stmt_498_call_ack_0 : boolean;
  signal call_stmt_498_call_ack_1 : boolean;
  signal call_stmt_487_call_req_0 : boolean;
  signal call_stmt_498_call_req_1 : boolean;
  signal NOT_u1_u1_501_inst_req_1 : boolean;
  signal call_stmt_462_call_req_1 : boolean;
  signal call_stmt_467_call_ack_1 : boolean;
  signal call_stmt_467_call_req_1 : boolean;
  signal call_stmt_467_call_ack_0 : boolean;
  signal call_stmt_467_call_req_0 : boolean;
  signal call_stmt_487_call_ack_1 : boolean;
  signal call_stmt_498_call_req_0 : boolean;
  signal call_stmt_492_call_ack_0 : boolean;
  signal call_stmt_487_call_ack_0 : boolean;
  signal call_stmt_462_call_ack_0 : boolean;
  signal call_stmt_487_call_req_1 : boolean;
  signal call_stmt_492_call_ack_1 : boolean;
  signal call_stmt_492_call_req_1 : boolean;
  signal NOT_u1_u1_501_inst_ack_0 : boolean;
  signal NOT_u1_u1_501_inst_req_0 : boolean;
  signal NOT_u1_u1_501_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "popFromQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 37) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(tag_length + 36 downto 37) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 36 downto 37);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  popFromQueue_CP_510_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "popFromQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_510_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= popFromQueue_CP_510_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_510_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,popFromQueue_CP_510_start,"popFromQueue cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,popFromQueue_CP_510_symbol, "popFromQueue cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  popFromQueue_CP_510: Block -- control-path 
    signal popFromQueue_CP_510_elements: BooleanArray(14 downto 0);
    -- 
  begin -- 
    popFromQueue_CP_510_elements(0) <= popFromQueue_CP_510_start;
    popFromQueue_CP_510_symbol <= popFromQueue_CP_510_elements(14);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_462/call_stmt_462_Sample/crr
      -- CP-element group 0: 	 call_stmt_462/call_stmt_462_sample_start_
      -- CP-element group 0: 	 call_stmt_462/call_stmt_462_Update/ccr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_462/$entry
      -- CP-element group 0: 	 call_stmt_462/call_stmt_462_Sample/$entry
      -- CP-element group 0: 	 call_stmt_462/call_stmt_462_Update/$entry
      -- CP-element group 0: 	 call_stmt_462/call_stmt_462_update_start_
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_462_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_462_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ccr_528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(0), ack => call_stmt_462_call_req_1); -- 
    crr_523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(0), ack => call_stmt_462_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_462/call_stmt_462_Sample/$exit
      -- CP-element group 1: 	 call_stmt_462/call_stmt_462_Sample/cra
      -- CP-element group 1: 	 call_stmt_462/call_stmt_462_sample_completed_
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_462_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_462_call_ack_0, ack => popFromQueue_CP_510_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (17) 
      -- CP-element group 2: 	 call_stmt_462/call_stmt_462_Update/cca
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/$entry
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Update/ccr
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Update/$entry
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Sample/crr
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Sample/$entry
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_update_start_
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_update_start_
      -- CP-element group 2: 	 call_stmt_462/call_stmt_462_update_completed_
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_update_start_
      -- CP-element group 2: 	 call_stmt_462/$exit
      -- CP-element group 2: 	 call_stmt_462/call_stmt_462_Update/$exit
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_sample_start_
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Update/$entry
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Update/ccr
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Update/ccr
      -- CP-element group 2: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Update/$entry
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_462_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_487_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_492_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_467_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_467_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_462_call_ack_1, ack => popFromQueue_CP_510_elements(2)); -- 
    ccr_559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(2), ack => call_stmt_487_call_req_1); -- 
    ccr_573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(2), ack => call_stmt_492_call_req_1); -- 
    crr_540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(2), ack => call_stmt_467_call_req_0); -- 
    ccr_545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(2), ack => call_stmt_467_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Sample/cra
      -- CP-element group 3: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Sample/$exit
      -- CP-element group 3: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_sample_completed_
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_467_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_467_call_ack_0, ack => popFromQueue_CP_510_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_sample_start_
      -- CP-element group 4: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Sample/crr
      -- CP-element group 4: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Update/cca
      -- CP-element group 4: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_Update/$exit
      -- CP-element group 4: 	 call_stmt_467_to_call_stmt_492/call_stmt_467_update_completed_
      -- CP-element group 4: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Sample/$entry
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_467_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_487_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_467_call_ack_1, ack => popFromQueue_CP_510_elements(4)); -- 
    crr_554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(4), ack => call_stmt_487_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Sample/$exit
      -- CP-element group 5: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Sample/cra
      -- CP-element group 5: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_sample_completed_
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_487_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_487_call_ack_0, ack => popFromQueue_CP_510_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_update_completed_
      -- CP-element group 6: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Update/$exit
      -- CP-element group 6: 	 call_stmt_467_to_call_stmt_492/call_stmt_487_Update/cca
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_487_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_487_call_ack_1, ack => popFromQueue_CP_510_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Sample/crr
      -- CP-element group 7: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Sample/$entry
      -- CP-element group 7: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_sample_start_
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_492_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(7), ack => call_stmt_492_call_req_0); -- 
    popFromQueue_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "popFromQueue_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_510_elements(4) & popFromQueue_CP_510_elements(6);
      gj_popFromQueue_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_510_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Sample/$exit
      -- CP-element group 8: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_sample_completed_
      -- CP-element group 8: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Sample/cra
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_492_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_492_call_ack_0, ack => popFromQueue_CP_510_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (17) 
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Update/ccr
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Update/cr
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Update/$entry
      -- CP-element group 9: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_update_completed_
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_update_start_
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/$entry
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Sample/crr
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_sample_start_
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_sample_start_
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Sample/$entry
      -- CP-element group 9: 	 call_stmt_467_to_call_stmt_492/$exit
      -- CP-element group 9: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Update/cca
      -- CP-element group 9: 	 call_stmt_467_to_call_stmt_492/call_stmt_492_Update/$exit
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Sample/rr
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Sample/$entry
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_update_start_
      -- CP-element group 9: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Update/$entry
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_492_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:NOT_u1_u1_501_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_498_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_498_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:NOT_u1_u1_501_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_492_call_ack_1, ack => popFromQueue_CP_510_elements(9)); -- 
    rr_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(9), ack => NOT_u1_u1_501_inst_req_0); -- 
    crr_585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(9), ack => call_stmt_498_call_req_0); -- 
    ccr_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(9), ack => call_stmt_498_call_req_1); -- 
    cr_604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_510_elements(9), ack => NOT_u1_u1_501_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Sample/cra
      -- CP-element group 10: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_sample_completed_
      -- CP-element group 10: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Sample/$exit
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_498_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_498_call_ack_0, ack => popFromQueue_CP_510_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_update_completed_
      -- CP-element group 11: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Update/cca
      -- CP-element group 11: 	 call_stmt_498_to_assign_stmt_502/call_stmt_498_Update/$exit
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:call_stmt_498_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_498_call_ack_1, ack => popFromQueue_CP_510_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Sample/ra
      -- CP-element group 12: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_sample_completed_
      -- CP-element group 12: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Sample/$exit
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:NOT_u1_u1_501_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_501_inst_ack_0, ack => popFromQueue_CP_510_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Update/$exit
      -- CP-element group 13: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_update_completed_
      -- CP-element group 13: 	 call_stmt_498_to_assign_stmt_502/NOT_u1_u1_501_Update/ca
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:NOT_u1_u1_501_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_501_inst_ack_1, ack => popFromQueue_CP_510_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 $exit
      -- CP-element group 14: 	 call_stmt_498_to_assign_stmt_502/$exit
      -- 
    -- logger for CP element group popFromQueue_CP_510_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and popFromQueue_CP_510_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:popFromQueue:CP:popFromQueue_CP_510_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    popFromQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_510_elements(11) & popFromQueue_CP_510_elements(13);
      gj_popFromQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_510_elements(14), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_479_wire : std_logic_vector(31 downto 0);
    signal R_QUEUE_SIZE_MASK_480_wire_constant : std_logic_vector(31 downto 0);
    signal konst_478_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_462 : std_logic_vector(0 downto 0);
    signal next_rp_482 : std_logic_vector(31 downto 0);
    signal q_empty_475 : std_logic_vector(0 downto 0);
    signal read_pointer_467 : std_logic_vector(31 downto 0);
    signal write_pointer_467 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_QUEUE_SIZE_MASK_480_wire_constant <= "00000000000000000000000100000000";
    konst_478_wire_constant <= "00000000000000000000000000000001";
    -- logger for split-operator ADD_u32_u32_479_inst flow-through 
    process(ADD_u32_u32_479_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:ADD_u32_u32_479_inst:flowthrough inputs: " & " read_pointer_467 = "& Convert_SLV_To_Hex_String(read_pointer_467) & " konst_478_wire_constant = "& Convert_SLV_To_Hex_String(konst_478_wire_constant) & " outputs:" & " ADD_u32_u32_479_wire= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_479_wire));
      --
    end process; 
    -- binary operator ADD_u32_u32_479_inst
    process(read_pointer_467) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(read_pointer_467, konst_478_wire_constant, tmp_var);
      ADD_u32_u32_479_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_481_inst flow-through 
    process(next_rp_482) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:AND_u32_u32_481_inst:flowthrough inputs: " & " ADD_u32_u32_479_wire = "& Convert_SLV_To_Hex_String(ADD_u32_u32_479_wire) & " R_QUEUE_SIZE_MASK_480_wire_constant = "& Convert_SLV_To_Hex_String(R_QUEUE_SIZE_MASK_480_wire_constant) & " outputs:" & " next_rp_482= "  & Convert_SLV_To_Hex_String(next_rp_482));
      --
    end process; 
    -- binary operator AND_u32_u32_481_inst
    process(ADD_u32_u32_479_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ADD_u32_u32_479_wire, R_QUEUE_SIZE_MASK_480_wire_constant, tmp_var);
      next_rp_482 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_474_inst flow-through 
    process(q_empty_475) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:EQ_u32_u1_474_inst:flowthrough inputs: " & " write_pointer_467 = "& Convert_SLV_To_Hex_String(write_pointer_467) & " read_pointer_467 = "& Convert_SLV_To_Hex_String(read_pointer_467) & " outputs:" & " q_empty_475= "  & Convert_SLV_To_Hex_String(q_empty_475));
      --
    end process; 
    -- binary operator EQ_u32_u1_474_inst
    process(write_pointer_467, read_pointer_467) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_pointer_467, read_pointer_467, tmp_var);
      q_empty_475 <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_501_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NOT_u1_u1_501_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:NOT_u1_u1_501_inst:started:   inputs: " & " q_empty_475 = "& Convert_SLV_To_Hex_String(q_empty_475));
          --
        end if; 
        if NOT_u1_u1_501_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:NOT_u1_u1_501_inst:finished:  outputs: " & " status_buffer= "  & Convert_SLV_To_Hex_String(status_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (3) : NOT_u1_u1_501_inst 
    ApIntNot_group_3: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= q_empty_475;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_501_inst_req_0;
      NOT_u1_u1_501_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_501_inst_req_1;
      NOT_u1_u1_501_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_3_gI: SplitGuardInterface generic map(name => "ApIntNot_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- logger for split-operator call_stmt_462_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_462_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_462_call:started:  Call to module acquireMutex inputs: " & " lock_buffer (guard)= " & Convert_SLV_To_String(lock_buffer) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer));
          --
        end if; 
        if call_stmt_462_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_462_call:finished:  outputs: " & " m_ok_462= "  & Convert_SLV_To_Hex_String(m_ok_462));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_462_call 
    acquireMutex_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_462_call_req_0;
      call_stmt_462_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_462_call_req_1;
      call_stmt_462_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireMutex_call_group_0_gI: SplitGuardInterface generic map(name => "acquireMutex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_462 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireMutex_call_reqs(0),
          ackR => acquireMutex_call_acks(0),
          dataR => acquireMutex_call_data(35 downto 0),
          tagR => acquireMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireMutex_return_acks(0), -- cross-over
          ackL => acquireMutex_return_reqs(0), -- cross-over
          dataL => acquireMutex_return_data(0 downto 0),
          tagL => acquireMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_467_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_467_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_467_call:started:  Call to module getQueuePointers inputs: " & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer));
          --
        end if; 
        if call_stmt_467_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_467_call:finished:  outputs: " & " write_pointer_467= "  & Convert_SLV_To_Hex_String(write_pointer_467) & " read_pointer_467= "  & Convert_SLV_To_Hex_String(read_pointer_467));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_467_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_467_call_req_0;
      call_stmt_467_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_467_call_req_1;
      call_stmt_467_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_pointer_467 <= data_out(63 downto 32);
      read_pointer_467 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_487_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_487_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_487_call:started:  Call to module getQueueElement inputs: " & " q_empty_475 (guard complement )= " & Convert_SLV_To_String(q_empty_475) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " read_pointer_467 = "& Convert_SLV_To_Hex_String(read_pointer_467));
          --
        end if; 
        if call_stmt_487_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_487_call:finished:  outputs: " & " q_r_data_buffer= "  & Convert_SLV_To_Hex_String(q_r_data_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_487_call 
    getQueueElement_call_group_2: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_487_call_req_0;
      call_stmt_487_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_487_call_req_1;
      call_stmt_487_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_475(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueElement_call_group_2_gI: SplitGuardInterface generic map(name => "getQueueElement_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & read_pointer_467;
      q_r_data_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueElement_call_reqs(0),
          ackR => getQueueElement_call_acks(0),
          dataR => getQueueElement_call_data(67 downto 0),
          tagR => getQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueElement_return_acks(0), -- cross-over
          ackL => getQueueElement_return_reqs(0), -- cross-over
          dataL => getQueueElement_return_data(31 downto 0),
          tagL => getQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- logger for split-operator call_stmt_492_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_492_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_492_call:started:  Call to module setQueuePointers inputs: " & " q_empty_475 (guard complement )= " & Convert_SLV_To_String(q_empty_475) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " write_pointer_467 = "& Convert_SLV_To_Hex_String(write_pointer_467) & " next_rp_482 = "& Convert_SLV_To_Hex_String(next_rp_482));
          --
        end if; 
        if call_stmt_492_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_492_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (3) : call_stmt_492_call 
    setQueuePointers_call_group_3: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_492_call_req_0;
      call_stmt_492_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_492_call_req_1;
      call_stmt_492_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_475(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_3_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_pointer_467 & next_rp_482;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- logger for split-operator call_stmt_498_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_498_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_498_call:started:  Call to module releaseMutex inputs: " & " lock_buffer (guard)= " & Convert_SLV_To_String(lock_buffer) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer));
          --
        end if; 
        if call_stmt_498_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:popFromQueue:DP:call_stmt_498_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (4) : call_stmt_498_call 
    releaseMutex_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_498_call_req_0;
      call_stmt_498_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_498_call_req_1;
      call_stmt_498_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseMutex_call_group_4_gI: SplitGuardInterface generic map(name => "releaseMutex_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseMutex_call_reqs(0),
          ackR => releaseMutex_call_acks(0),
          dataR => releaseMutex_call_data(35 downto 0),
          tagR => releaseMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseMutex_return_acks(0), -- cross-over
          ackL => releaseMutex_return_reqs(0), -- cross-over
          tagL => releaseMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end popFromQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity populateRxQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity populateRxQueue;
architecture populateRxQueue_arch of populateRxQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal populateRxQueue_CP_1194_start: Boolean;
  signal populateRxQueue_CP_1194_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component delay_time_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      T : in  std_logic_vector(31 downto 0);
      delay_done : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u6_u6_814_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_0 : boolean;
  signal n_q_index_854_815_buf_req_0 : boolean;
  signal ADD_u6_u6_814_inst_ack_0 : boolean;
  signal ADD_u6_u6_814_inst_req_0 : boolean;
  signal W_selected_q_index_871_inst_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_1 : boolean;
  signal call_stmt_860_call_req_0 : boolean;
  signal n_q_index_854_815_buf_ack_0 : boolean;
  signal call_stmt_860_call_ack_0 : boolean;
  signal ADD_u6_u6_814_inst_ack_1 : boolean;
  signal phi_stmt_810_req_0 : boolean;
  signal n_q_index_854_815_buf_req_1 : boolean;
  signal if_stmt_861_branch_ack_0 : boolean;
  signal n_q_index_854_815_buf_ack_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_1 : boolean;
  signal call_stmt_860_call_req_1 : boolean;
  signal phi_stmt_810_req_1 : boolean;
  signal W_selected_q_index_871_inst_req_0 : boolean;
  signal call_stmt_860_call_ack_1 : boolean;
  signal phi_stmt_810_ack_0 : boolean;
  signal W_selected_q_index_871_inst_req_1 : boolean;
  signal if_stmt_861_branch_ack_1 : boolean;
  signal W_selected_q_index_871_inst_ack_0 : boolean;
  signal if_stmt_861_branch_req_0 : boolean;
  signal call_stmt_831_call_req_0 : boolean;
  signal call_stmt_831_call_ack_0 : boolean;
  signal call_stmt_831_call_req_1 : boolean;
  signal call_stmt_831_call_ack_1 : boolean;
  signal call_stmt_844_call_req_0 : boolean;
  signal call_stmt_844_call_ack_0 : boolean;
  signal call_stmt_844_call_req_1 : boolean;
  signal call_stmt_844_call_ack_1 : boolean;
  signal AND_u6_u6_853_inst_req_0 : boolean;
  signal AND_u6_u6_853_inst_ack_0 : boolean;
  signal AND_u6_u6_853_inst_req_1 : boolean;
  signal AND_u6_u6_853_inst_ack_1 : boolean;
  signal if_stmt_855_branch_req_0 : boolean;
  signal if_stmt_855_branch_ack_1 : boolean;
  signal if_stmt_855_branch_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "populateRxQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  populateRxQueue_CP_1194_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "populateRxQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1194_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= populateRxQueue_CP_1194_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_1194_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,populateRxQueue_CP_1194_start,"populateRxQueue cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,populateRxQueue_CP_1194_symbol, "populateRxQueue cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  populateRxQueue_CP_1194: Block -- control-path 
    signal populateRxQueue_CP_1194_elements: BooleanArray(28 downto 0);
    -- 
  begin -- 
    populateRxQueue_CP_1194_elements(0) <= populateRxQueue_CP_1194_start;
    populateRxQueue_CP_1194_symbol <= populateRxQueue_CP_1194_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	20 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 branch_block_stmt_808/merge_stmt_809_dead_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_808/$entry
      -- CP-element group 0: 	 branch_block_stmt_808/branch_block_stmt_808__entry__
      -- CP-element group 0: 	 branch_block_stmt_808/merge_stmt_809__entry__
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  merge  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	19 
    -- CP-element group 1: 	14 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_808/$exit
      -- CP-element group 1: 	 branch_block_stmt_808/branch_block_stmt_808__exit__
      -- CP-element group 1: 	 branch_block_stmt_808/if_stmt_855__exit__
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    populateRxQueue_CP_1194_elements(1) <= OrReduce(populateRxQueue_CP_1194_elements(19) & populateRxQueue_CP_1194_elements(14));
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	28 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Sample/cra
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_831_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_831_call_ack_0, ack => populateRxQueue_CP_1194_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	28 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Sample/crr
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_831_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_844_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_1224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_831_call_ack_1, ack => populateRxQueue_CP_1194_elements(3)); -- 
    crr_1232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(3), ack => call_stmt_844_call_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Sample/cra
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_844_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_844_call_ack_0, ack => populateRxQueue_CP_1194_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	28 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Update/cca
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_844_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_844_call_ack_1, ack => populateRxQueue_CP_1194_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	28 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Sample/ra
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:AND_u6_u6_853_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_853_inst_ack_0, ack => populateRxQueue_CP_1194_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	28 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Update/ca
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:AND_u6_u6_853_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_853_inst_ack_1, ack => populateRxQueue_CP_1194_elements(7)); -- 
    -- CP-element group 8:  branch  join  transition  place  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: 	5 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (22) 
      -- CP-element group 8: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854__exit__
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855__entry__
      -- CP-element group 8: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/$exit
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_dead_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/$entry
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/$exit
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/$entry
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/$exit
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/$entry
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/$exit
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Update/cr
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/NOT_u1_u1_857/SplitProtocol/Update/ca
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_eval_test/branch_req
      -- CP-element group 8: 	 branch_block_stmt_808/NOT_u1_u1_857_place
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_if_link/$entry
      -- CP-element group 8: 	 branch_block_stmt_808/if_stmt_855_else_link/$entry
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:if_stmt_855_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(8), ack => if_stmt_855_branch_req_0); -- 
    populateRxQueue_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "populateRxQueue_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1194_elements(7) & populateRxQueue_CP_1194_elements(5);
      gj_populateRxQueue_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1194_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  fork  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (10) 
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Sample/crr
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_update_start_
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Update/ccr
      -- CP-element group 9: 	 branch_block_stmt_808/if_stmt_855_if_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_808/if_stmt_855_if_link/if_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860__entry__
      -- CP-element group 9: 	 branch_block_stmt_808/call_stmt_860/$entry
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:if_stmt_855_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_860_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_860_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_855_branch_ack_1, ack => populateRxQueue_CP_1194_elements(9)); -- 
    crr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(9), ack => call_stmt_860_call_req_0); -- 
    ccr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(9), ack => call_stmt_860_call_req_1); -- 
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	18 
    -- CP-element group 10:  members (13) 
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Sample/req
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873__entry__
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/$entry
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_update_start_
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Sample/req
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Update/req
      -- CP-element group 10: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_808/if_stmt_855_else_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_808/if_stmt_855_else_link/else_choice_transition
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:if_stmt_855_branch_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:W_selected_q_index_871_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:W_selected_q_index_871_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_855_branch_ack_0, ack => populateRxQueue_CP_1194_elements(10)); -- 
    req_1356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(10), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_0); -- 
    req_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(10), ack => W_selected_q_index_871_inst_req_0); -- 
    req_1375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(10), ack => W_selected_q_index_871_inst_req_1); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Sample/cra
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_860_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_860_call_ack_0, ack => populateRxQueue_CP_1194_elements(11)); -- 
    -- CP-element group 12:  branch  transition  place  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (27) 
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/$exit
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/$exit
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Sample/rr
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/EQ_u1_u1_864_inputs/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/EQ_u1_u1_864_inputs/$exit
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_808/call_stmt_860/call_stmt_860_Update/cca
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_else_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/EQ_u1_u1_864_place
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Update/ca
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861_eval_test/EQ_u1_u1_864/SplitProtocol/Update/cr
      -- CP-element group 12: 	 branch_block_stmt_808/call_stmt_860__exit__
      -- CP-element group 12: 	 branch_block_stmt_808/if_stmt_861__entry__
      -- CP-element group 12: 	 branch_block_stmt_808/call_stmt_860/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_860_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:if_stmt_861_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_1306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_860_call_ack_1, ack => populateRxQueue_CP_1194_elements(12)); -- 
    branch_req_1333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(12), ack => if_stmt_861_branch_req_0); -- 
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	24 
    -- CP-element group 13: 	25 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Sample/req
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/$entry
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/$entry
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Update/req
      -- CP-element group 13: 	 branch_block_stmt_808/loopback
      -- CP-element group 13: 	 branch_block_stmt_808/if_stmt_861_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_808/if_stmt_861_if_link/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:if_stmt_861_branch_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:n_q_index_854_815_buf_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:n_q_index_854_815_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_861_branch_ack_1, ack => populateRxQueue_CP_1194_elements(13)); -- 
    req_1438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(13), ack => n_q_index_854_815_buf_req_0); -- 
    req_1443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(13), ack => n_q_index_854_815_buf_req_1); -- 
    -- CP-element group 14:  merge  transition  place  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	1 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_808/if_stmt_861_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_808/if_stmt_861_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_808/if_stmt_861__exit__
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(14) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:if_stmt_861_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_1342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_861_branch_ack_0, ack => populateRxQueue_CP_1194_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Sample/ack
      -- CP-element group 15: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Update/req
      -- CP-element group 15: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_update_start_
      -- CP-element group 15: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Sample/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_0, ack => populateRxQueue_CP_1194_elements(15)); -- 
    req_1361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(15), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	19 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_Update/ack
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_1, ack => populateRxQueue_CP_1194_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Sample/ack
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:W_selected_q_index_871_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_selected_q_index_871_inst_ack_0, ack => populateRxQueue_CP_1194_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	10 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Update/ack
      -- CP-element group 18: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/assign_stmt_873_Update/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:W_selected_q_index_871_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_selected_q_index_871_inst_ack_1, ack => populateRxQueue_CP_1194_elements(18)); -- 
    -- CP-element group 19:  join  transition  place  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	16 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	1 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873__exit__
      -- CP-element group 19: 	 branch_block_stmt_808/assign_stmt_870_to_assign_stmt_873/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    populateRxQueue_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1194_elements(16) & populateRxQueue_CP_1194_elements(18);
      gj_populateRxQueue_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1194_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (21) 
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Update/cr
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/$exit
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Update/ack
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Update/req
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Sample/ack
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Sample/req
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/$exit
      -- CP-element group 20: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/ADD_u6_u6_814_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812/$entry
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:ADD_u6_u6_814_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:ADD_u6_u6_814_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cr_1420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(20), ack => ADD_u6_u6_814_inst_req_1); -- 
    rr_1415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(20), ack => ADD_u6_u6_814_inst_req_0); -- 
    populateRxQueue_CP_1194_elements(20) <= populateRxQueue_CP_1194_elements(0);
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Sample/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:ADD_u6_u6_814_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u6_u6_814_inst_ack_0, ack => populateRxQueue_CP_1194_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Update/ca
      -- CP-element group 22: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/Update/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:ADD_u6_u6_814_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u6_u6_814_inst_ack_1, ack => populateRxQueue_CP_1194_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	27 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/$exit
      -- CP-element group 23: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/$exit
      -- CP-element group 23: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/$exit
      -- CP-element group 23: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/$exit
      -- CP-element group 23: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_req
      -- CP-element group 23: 	 branch_block_stmt_808/merge_stmt_809__entry___PhiReq/phi_stmt_810/phi_stmt_810_sources/ADD_u6_u6_814/SplitProtocol/$exit
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:phi_stmt_810_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_810_req_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_810_req_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(23), ack => phi_stmt_810_req_0); -- 
    populateRxQueue_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1194_elements(22) & populateRxQueue_CP_1194_elements(21);
      gj_populateRxQueue_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1194_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	13 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Sample/ack
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:n_q_index_854_815_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_1439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_854_815_buf_ack_0, ack => populateRxQueue_CP_1194_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	13 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/Update/ack
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:n_q_index_854_815_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_1444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_854_815_buf_ack_1, ack => populateRxQueue_CP_1194_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/$exit
      -- CP-element group 26: 	 branch_block_stmt_808/loopback_PhiReq/$exit
      -- CP-element group 26: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/$exit
      -- CP-element group 26: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_sources/Interlock/$exit
      -- CP-element group 26: 	 branch_block_stmt_808/loopback_PhiReq/phi_stmt_810/phi_stmt_810_req
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:phi_stmt_810_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_810_req_1445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_810_req_1445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(26), ack => phi_stmt_810_req_1); -- 
    populateRxQueue_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_1194_elements(24) & populateRxQueue_CP_1194_elements(25);
      gj_populateRxQueue_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_1194_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  merge  transition  place  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_808/merge_stmt_809_PhiReqMerge
      -- CP-element group 27: 	 branch_block_stmt_808/merge_stmt_809_PhiAck/$entry
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(27) fired."); 
        -- 
      end if; --
    end process; 
    populateRxQueue_CP_1194_elements(27) <= OrReduce(populateRxQueue_CP_1194_elements(23) & populateRxQueue_CP_1194_elements(26));
    -- CP-element group 28:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: 	6 
    -- CP-element group 28: 	7 
    -- CP-element group 28: 	3 
    -- CP-element group 28: 	5 
    -- CP-element group 28:  members (20) 
      -- CP-element group 28: 	 branch_block_stmt_808/merge_stmt_809_PhiAck/$exit
      -- CP-element group 28: 	 branch_block_stmt_808/merge_stmt_809_PhiAck/phi_stmt_810_ack
      -- CP-element group 28: 	 branch_block_stmt_808/merge_stmt_809__exit__
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854__entry__
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/$entry
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_update_start_
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Sample/crr
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_831_Update/ccr
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_update_start_
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/call_stmt_844_Update/ccr
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_update_start_
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_808/assign_stmt_822_to_assign_stmt_854/AND_u6_u6_853_Update/cr
      -- 
    -- logger for CP element group populateRxQueue_CP_1194_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and populateRxQueue_CP_1194_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:populateRxQueue_CP_1194_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:phi_stmt_810_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_831_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_831_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:call_stmt_844_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:AND_u6_u6_853_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:populateRxQueue:CP:AND_u6_u6_853_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_810_ack_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_810_ack_0, ack => populateRxQueue_CP_1194_elements(28)); -- 
    crr_1218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(28), ack => call_stmt_831_call_req_0); -- 
    ccr_1223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(28), ack => call_stmt_831_call_req_1); -- 
    ccr_1237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(28), ack => call_stmt_844_call_req_1); -- 
    rr_1246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(28), ack => AND_u6_u6_853_inst_req_0); -- 
    cr_1251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_1194_elements(28), ack => AND_u6_u6_853_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_814_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_820_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_848_wire : std_logic_vector(5 downto 0);
    signal EQ_u1_u1_864_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_857_wire : std_logic_vector(0 downto 0);
    signal RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_849_wire : std_logic_vector(31 downto 0);
    signal R_RX_QUEUES_REG_START_OFFSET_819_wire_constant : std_logic_vector(5 downto 0);
    signal SUB_u32_u32_851_wire : std_logic_vector(31 downto 0);
    signal konst_813_wire_constant : std_logic_vector(5 downto 0);
    signal konst_847_wire_constant : std_logic_vector(5 downto 0);
    signal konst_850_wire_constant : std_logic_vector(31 downto 0);
    signal konst_858_wire_constant : std_logic_vector(31 downto 0);
    signal konst_863_wire_constant : std_logic_vector(0 downto 0);
    signal n_q_index_854 : std_logic_vector(5 downto 0);
    signal n_q_index_854_815_buffered : std_logic_vector(5 downto 0);
    signal push_status_844 : std_logic_vector(0 downto 0);
    signal q_index_810 : std_logic_vector(5 downto 0);
    signal register_index_822 : std_logic_vector(5 downto 0);
    signal rx_queue_pointer_32_831 : std_logic_vector(31 downto 0);
    signal rx_queue_pointer_36_837 : std_logic_vector(35 downto 0);
    signal selected_q_index_873 : std_logic_vector(5 downto 0);
    signal slice_842_wire : std_logic_vector(31 downto 0);
    signal status_860 : std_logic_vector(0 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_826_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_829_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_835_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_839_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_852_wire : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    R_RX_QUEUES_REG_START_OFFSET_819_wire_constant <= "000010";
    konst_813_wire_constant <= "000001";
    konst_847_wire_constant <= "000001";
    konst_850_wire_constant <= "00000000000000000000000000000001";
    konst_858_wire_constant <= "00000000000000000000000000100000";
    konst_863_wire_constant <= "0";
    type_cast_824_wire_constant <= "1";
    type_cast_826_wire_constant <= "0001";
    type_cast_829_wire_constant <= "00000000000000000000000000000000";
    type_cast_835_wire_constant <= "0000";
    type_cast_839_wire_constant <= "0";
    -- logger for phi phi_stmt_810
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_810_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:populateRxQueue:DP:phi_stmt_810:input-0 ADD_u6_u6_814_wire= " & Convert_SLV_To_Hex_String(ADD_u6_u6_814_wire));
          --
        end if;
        if phi_stmt_810_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:populateRxQueue:DP:phi_stmt_810:input-1 n_q_index_854_815_buffered= " & Convert_SLV_To_Hex_String(n_q_index_854_815_buffered));
          --
        end if;
        if phi_stmt_810_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:populateRxQueue:DP:phi_stmt_810:sample-completed");
          --
        end if;
        if phi_stmt_810_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:populateRxQueue:DP:phi_stmt_810:output q_index_810= " & Convert_SLV_To_Hex_String(q_index_810));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_810: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u6_u6_814_wire & n_q_index_854_815_buffered;
      req <= phi_stmt_810_req_0 & phi_stmt_810_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_810",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_810_ack_0,
          idata => idata,
          odata => q_index_810,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_810
    -- logger for split-operator slice_842_inst flow-through 
    process(slice_842_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:slice_842_inst:flowthrough inputs: " & " rx_buffer_pointer_buffer = "& Convert_SLV_To_Hex_String(rx_buffer_pointer_buffer) & " outputs:" & " slice_842_wire= "  & Convert_SLV_To_Hex_String(slice_842_wire));
      --
    end process; 
    -- flow-through slice operator slice_842_inst
    slice_842_wire <= rx_buffer_pointer_buffer(35 downto 4);
    -- logger for split-operator W_selected_q_index_871_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if W_selected_q_index_871_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:W_selected_q_index_871_inst:started:   inputs: " & " q_index_810 = "& Convert_SLV_To_Hex_String(q_index_810));
          --
        end if; 
        if W_selected_q_index_871_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:W_selected_q_index_871_inst:finished:  outputs: " & " selected_q_index_873= "  & Convert_SLV_To_Hex_String(selected_q_index_873));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    W_selected_q_index_871_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_selected_q_index_871_inst_req_0;
      W_selected_q_index_871_inst_ack_0<= wack(0);
      rreq(0) <= W_selected_q_index_871_inst_req_1;
      W_selected_q_index_871_inst_ack_1<= rack(0);
      W_selected_q_index_871_inst : InterlockBuffer generic map ( -- 
        name => "W_selected_q_index_871_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_index_810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => selected_q_index_873,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator n_q_index_854_815_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if n_q_index_854_815_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:n_q_index_854_815_buf:started:   inputs: " & " n_q_index_854 = "& Convert_SLV_To_Hex_String(n_q_index_854));
          --
        end if; 
        if n_q_index_854_815_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:n_q_index_854_815_buf:finished:  outputs: " & " n_q_index_854_815_buffered= "  & Convert_SLV_To_Hex_String(n_q_index_854_815_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    n_q_index_854_815_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_q_index_854_815_buf_req_0;
      n_q_index_854_815_buf_ack_0<= wack(0);
      rreq(0) <= n_q_index_854_815_buf_req_1;
      n_q_index_854_815_buf_ack_1<= rack(0);
      n_q_index_854_815_buf : InterlockBuffer generic map ( -- 
        name => "n_q_index_854_815_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_q_index_854,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_q_index_854_815_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_821_inst flow-through 
    process(register_index_822) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:type_cast_821_inst:flowthrough inputs: " & " ADD_u6_u6_820_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_820_wire) & " outputs:" & " register_index_822= "  & Convert_SLV_To_Hex_String(register_index_822));
      --
    end process; 
    -- interlock type_cast_821_inst
    process(ADD_u6_u6_820_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_820_wire(5 downto 0);
      register_index_822 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_852_inst flow-through 
    process(type_cast_852_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:type_cast_852_inst:flowthrough inputs: " & " SUB_u32_u32_851_wire = "& Convert_SLV_To_Hex_String(SUB_u32_u32_851_wire) & " outputs:" & " type_cast_852_wire= "  & Convert_SLV_To_Hex_String(type_cast_852_wire));
      --
    end process; 
    -- interlock type_cast_852_inst
    process(SUB_u32_u32_851_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_851_wire(5 downto 0);
      type_cast_852_wire <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_855_branch_req_0," req0 if_stmt_855_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_855_branch_ack_0," ack0 if_stmt_855_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_855_branch_ack_1," ack1 if_stmt_855_branch");
    if_stmt_855_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_857_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_855_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_855_branch_req_0,
          ack0 => if_stmt_855_branch_ack_0,
          ack1 => if_stmt_855_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_861_branch_req_0," req0 if_stmt_861_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_861_branch_ack_0," ack0 if_stmt_861_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_861_branch_ack_1," ack1 if_stmt_861_branch");
    if_stmt_861_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_864_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_861_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_861_branch_req_0,
          ack0 => if_stmt_861_branch_ack_0,
          ack1 => if_stmt_861_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u6_u6_814_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u6_u6_814_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:ADD_u6_u6_814_inst:started:   inputs: " & " RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire = "& Convert_SLV_To_Hex_String(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire) & " konst_813_wire_constant = "& Convert_SLV_To_Hex_String(konst_813_wire_constant));
          --
        end if; 
        if ADD_u6_u6_814_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:ADD_u6_u6_814_inst:finished:  outputs: " & " ADD_u6_u6_814_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_814_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u6_u6_814_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire;
      ADD_u6_u6_814_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u6_u6_814_inst_req_0;
      ADD_u6_u6_814_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u6_u6_814_inst_req_1;
      ADD_u6_u6_814_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "000001",
          constant_width => 6,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator ADD_u6_u6_820_inst flow-through 
    process(ADD_u6_u6_820_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:ADD_u6_u6_820_inst:flowthrough inputs: " & " q_index_810 = "& Convert_SLV_To_Hex_String(q_index_810) & " R_RX_QUEUES_REG_START_OFFSET_819_wire_constant = "& Convert_SLV_To_Hex_String(R_RX_QUEUES_REG_START_OFFSET_819_wire_constant) & " outputs:" & " ADD_u6_u6_820_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_820_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_820_inst
    process(q_index_810) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_810, R_RX_QUEUES_REG_START_OFFSET_819_wire_constant, tmp_var);
      ADD_u6_u6_820_wire <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u6_u6_848_inst flow-through 
    process(ADD_u6_u6_848_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:ADD_u6_u6_848_inst:flowthrough inputs: " & " q_index_810 = "& Convert_SLV_To_Hex_String(q_index_810) & " konst_847_wire_constant = "& Convert_SLV_To_Hex_String(konst_847_wire_constant) & " outputs:" & " ADD_u6_u6_848_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_848_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_848_inst
    process(q_index_810) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_810, konst_847_wire_constant, tmp_var);
      ADD_u6_u6_848_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u6_u6_853_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if AND_u6_u6_853_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:AND_u6_u6_853_inst:started:   inputs: " & " ADD_u6_u6_848_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_848_wire) & " type_cast_852_wire = "& Convert_SLV_To_Hex_String(type_cast_852_wire));
          --
        end if; 
        if AND_u6_u6_853_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:AND_u6_u6_853_inst:finished:  outputs: " & " n_q_index_854= "  & Convert_SLV_To_Hex_String(n_q_index_854));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (3) : AND_u6_u6_853_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_848_wire & type_cast_852_wire;
      n_q_index_854 <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_853_inst_req_0;
      AND_u6_u6_853_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_853_inst_req_1;
      AND_u6_u6_853_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- logger for split-operator CONCAT_u32_u36_836_inst flow-through 
    process(rx_queue_pointer_36_837) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:CONCAT_u32_u36_836_inst:flowthrough inputs: " & " rx_queue_pointer_32_831 = "& Convert_SLV_To_Hex_String(rx_queue_pointer_32_831) & " type_cast_835_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_835_wire_constant) & " outputs:" & " rx_queue_pointer_36_837= "  & Convert_SLV_To_Hex_String(rx_queue_pointer_36_837));
      --
    end process; 
    -- binary operator CONCAT_u32_u36_836_inst
    process(rx_queue_pointer_32_831) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(rx_queue_pointer_32_831, type_cast_835_wire_constant, tmp_var);
      rx_queue_pointer_36_837 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u1_u1_864_inst flow-through 
    process(EQ_u1_u1_864_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:EQ_u1_u1_864_inst:flowthrough inputs: " & " status_860 = "& Convert_SLV_To_Hex_String(status_860) & " konst_863_wire_constant = "& Convert_SLV_To_Hex_String(konst_863_wire_constant) & " outputs:" & " EQ_u1_u1_864_wire= "  & Convert_SLV_To_Hex_String(EQ_u1_u1_864_wire));
      --
    end process; 
    -- binary operator EQ_u1_u1_864_inst
    process(status_860) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(status_860, konst_863_wire_constant, tmp_var);
      EQ_u1_u1_864_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_857_inst flow-through 
    process(NOT_u1_u1_857_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:NOT_u1_u1_857_inst:flowthrough inputs: " & " push_status_844 = "& Convert_SLV_To_Hex_String(push_status_844) & " outputs:" & " NOT_u1_u1_857_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_857_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_857_inst
    process(push_status_844) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", push_status_844, tmp_var);
      NOT_u1_u1_857_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator SUB_u32_u32_851_inst flow-through 
    process(SUB_u32_u32_851_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:SUB_u32_u32_851_inst:flowthrough inputs: " & " RPIPE_NUMBER_OF_SERVERS_849_wire = "& Convert_SLV_To_Hex_String(RPIPE_NUMBER_OF_SERVERS_849_wire) & " konst_850_wire_constant = "& Convert_SLV_To_Hex_String(konst_850_wire_constant) & " outputs:" & " SUB_u32_u32_851_wire= "  & Convert_SLV_To_Hex_String(SUB_u32_u32_851_wire));
      --
    end process; 
    -- binary operator SUB_u32_u32_851_inst
    process(RPIPE_NUMBER_OF_SERVERS_849_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_849_wire, konst_850_wire_constant, tmp_var);
      SUB_u32_u32_851_wire <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_inst flow-through 
    process(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire= "  & Convert_SLV_To_Hex_String(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire));
      --
    end process; 
    -- read from input-signal LAST_WRITTEN_RX_QUEUE_INDEX
    RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_812_wire <= LAST_WRITTEN_RX_QUEUE_INDEX;
    -- logger for split-operator RPIPE_NUMBER_OF_SERVERS_849_inst flow-through 
    process(RPIPE_NUMBER_OF_SERVERS_849_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:RPIPE_NUMBER_OF_SERVERS_849_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_NUMBER_OF_SERVERS_849_wire= "  & Convert_SLV_To_Hex_String(RPIPE_NUMBER_OF_SERVERS_849_wire));
      --
    end process; 
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_849_wire <= NUMBER_OF_SERVERS;
    -- logger for split-operator WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst:started:   PipeWrite to LAST_WRITTEN_RX_QUEUE_INDEX inputs: " & " q_index_810 = "& Convert_SLV_To_Hex_String(q_index_810));
          --
        end if; 
        if WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_868_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= q_index_810;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_831_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_831_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:call_stmt_831_call:started:  Call to module AccessRegister inputs: " & " type_cast_824_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_824_wire_constant) & " type_cast_826_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_826_wire_constant) & " register_index_822 = "& Convert_SLV_To_Hex_String(register_index_822) & " type_cast_829_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_829_wire_constant));
          --
        end if; 
        if call_stmt_831_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:call_stmt_831_call:finished:  outputs: " & " rx_queue_pointer_32_831= "  & Convert_SLV_To_Hex_String(rx_queue_pointer_32_831));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_831_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_831_call_req_0;
      call_stmt_831_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_831_call_req_1;
      call_stmt_831_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_824_wire_constant & type_cast_826_wire_constant & register_index_822 & type_cast_829_wire_constant;
      rx_queue_pointer_32_831 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_844_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_844_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:call_stmt_844_call:started:  Call to module pushIntoQueue inputs: " & " type_cast_839_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_839_wire_constant) & " rx_queue_pointer_36_837 = "& Convert_SLV_To_Hex_String(rx_queue_pointer_36_837) & " slice_842_wire = "& Convert_SLV_To_Hex_String(slice_842_wire));
          --
        end if; 
        if call_stmt_844_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:call_stmt_844_call:finished:  outputs: " & " push_status_844= "  & Convert_SLV_To_Hex_String(push_status_844));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_844_call 
    pushIntoQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_844_call_req_0;
      call_stmt_844_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_844_call_req_1;
      call_stmt_844_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_1_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_839_wire_constant & rx_queue_pointer_36_837 & slice_842_wire;
      push_status_844 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_860_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_860_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:call_stmt_860_call:started:  Call to module delay_time inputs: " & " konst_858_wire_constant = "& Convert_SLV_To_Hex_String(konst_858_wire_constant));
          --
        end if; 
        if call_stmt_860_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:populateRxQueue:DP:call_stmt_860_call:finished:  outputs: " & " status_860= "  & Convert_SLV_To_Hex_String(status_860));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    operator_delay_time_2117_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_860_call_req_0;
      call_stmt_860_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_860_call_req_1;
      call_stmt_860_call_ack_1<= update_ack(0);
      call_stmt_860_call: delay_time_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        T => konst_858_wire_constant,
        delay_done => status_860,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end populateRxQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity processorToNicInterface is -- 
  generic (tag_length : integer); 
  port ( -- 
    control_word_request_pipe_1_pipe_read_req : out  std_logic_vector(0 downto 0);
    control_word_request_pipe_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    control_word_request_pipe_1_pipe_read_data : in   std_logic_vector(63 downto 0);
    control_word_request_pipe_0_pipe_read_req : out  std_logic_vector(0 downto 0);
    control_word_request_pipe_0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    control_word_request_pipe_0_pipe_read_data : in   std_logic_vector(31 downto 0);
    AFB_NIC_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_data : out  std_logic_vector(73 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity processorToNicInterface;
architecture processorToNicInterface_arch of processorToNicInterface is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal processorToNicInterface_CP_2794_start: Boolean;
  signal processorToNicInterface_CP_2794_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1356_branch_req_0 : boolean;
  signal RPIPE_control_word_request_pipe_0_1360_inst_req_0 : boolean;
  signal RPIPE_control_word_request_pipe_0_1360_inst_ack_0 : boolean;
  signal RPIPE_control_word_request_pipe_0_1360_inst_req_1 : boolean;
  signal RPIPE_control_word_request_pipe_0_1360_inst_ack_1 : boolean;
  signal RPIPE_control_word_request_pipe_1_1363_inst_req_0 : boolean;
  signal RPIPE_control_word_request_pipe_1_1363_inst_ack_0 : boolean;
  signal RPIPE_control_word_request_pipe_1_1363_inst_req_1 : boolean;
  signal RPIPE_control_word_request_pipe_1_1363_inst_ack_1 : boolean;
  signal CONCAT_u42_u74_1373_inst_req_0 : boolean;
  signal CONCAT_u42_u74_1373_inst_ack_0 : boolean;
  signal CONCAT_u42_u74_1373_inst_req_1 : boolean;
  signal CONCAT_u42_u74_1373_inst_ack_1 : boolean;
  signal WPIPE_AFB_NIC_REQUEST_1368_inst_req_0 : boolean;
  signal WPIPE_AFB_NIC_REQUEST_1368_inst_ack_0 : boolean;
  signal WPIPE_AFB_NIC_REQUEST_1368_inst_req_1 : boolean;
  signal WPIPE_AFB_NIC_REQUEST_1368_inst_ack_1 : boolean;
  signal do_while_stmt_1356_branch_ack_0 : boolean;
  signal do_while_stmt_1356_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "processorToNicInterface_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  processorToNicInterface_CP_2794_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "processorToNicInterface_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= processorToNicInterface_CP_2794_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= processorToNicInterface_CP_2794_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= processorToNicInterface_CP_2794_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,processorToNicInterface_CP_2794_start,"processorToNicInterface cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,processorToNicInterface_CP_2794_symbol, "processorToNicInterface cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  processorToNicInterface_CP_2794: Block -- control-path 
    signal processorToNicInterface_CP_2794_elements: BooleanArray(35 downto 0);
    -- 
  begin -- 
    processorToNicInterface_CP_2794_elements(0) <= processorToNicInterface_CP_2794_start;
    processorToNicInterface_CP_2794_symbol <= processorToNicInterface_CP_2794_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1355/$entry
      -- CP-element group 0: 	 branch_block_stmt_1355/branch_block_stmt_1355__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1355/do_while_stmt_1356__entry__
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	34 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1355/$exit
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1355/branch_block_stmt_1355__exit__
      -- CP-element group 1: 	 branch_block_stmt_1355/do_while_stmt_1356__exit__
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_CP_2794_elements(1) <= processorToNicInterface_CP_2794_elements(34);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1355/do_while_stmt_1356/$entry
      -- CP-element group 2: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356__entry__
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_CP_2794_elements(2) <= processorToNicInterface_CP_2794_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	34 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356__exit__
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processorToNicInterface_CP_2794_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_back
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processorToNicInterface_CP_2794_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	32 
    -- CP-element group 5: 	33 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1355/do_while_stmt_1356/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_taken/$entry
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_CP_2794_elements(5) <= processorToNicInterface_CP_2794_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	35 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_body_done
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_CP_2794_elements(6) <= processorToNicInterface_CP_2794_elements(35);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_CP_2794_elements(7) <= processorToNicInterface_CP_2794_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_CP_2794_elements(8) <= processorToNicInterface_CP_2794_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	19 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1358_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1361_sample_start_
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processorToNicInterface_CP_2794_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	31 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/condition_evaluated
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:do_while_stmt_1356_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(10), ack => do_while_stmt_1356_branch_req_0); -- 
    processorToNicInterface_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(31) & processorToNicInterface_CP_2794_elements(13);
      gj_processorToNicInterface_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	20 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(9) & processorToNicInterface_CP_2794_elements(13);
      gj_processorToNicInterface_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	19 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	21 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(14) & processorToNicInterface_CP_2794_elements(19);
      gj_processorToNicInterface_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	23 
    -- CP-element group 13: 	18 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(23) & processorToNicInterface_CP_2794_elements(18);
      gj_processorToNicInterface_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	26 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1358_update_start_
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(9) & processorToNicInterface_CP_2794_elements(26);
      gj_processorToNicInterface_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Sample/rr
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_0_1360_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(15), ack => RPIPE_control_word_request_pipe_0_1360_inst_req_0); -- 
    processorToNicInterface_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(11) & processorToNicInterface_CP_2794_elements(18);
      gj_processorToNicInterface_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: 	17 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Update/cr
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(16) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_0_1360_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(16), ack => RPIPE_control_word_request_pipe_0_1360_inst_req_1); -- 
    processorToNicInterface_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(12) & processorToNicInterface_CP_2794_elements(17);
      gj_processorToNicInterface_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	35 
    -- CP-element group 17: 	16 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Sample/ra
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(17) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_0_1360_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_control_word_request_pipe_0_1360_inst_ack_0, ack => processorToNicInterface_CP_2794_elements(17)); -- 
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: 	24 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1358_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_0_1360_Update/ca
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_0_1360_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_control_word_request_pipe_0_1360_inst_ack_1, ack => processorToNicInterface_CP_2794_elements(18)); -- 
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	9 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	26 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	12 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1361_update_start_
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(9) & processorToNicInterface_CP_2794_elements(26);
      gj_processorToNicInterface_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	11 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Sample/rr
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_1_1363_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(20), ack => RPIPE_control_word_request_pipe_1_1363_inst_req_0); -- 
    processorToNicInterface_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(11) & processorToNicInterface_CP_2794_elements(23);
      gj_processorToNicInterface_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	12 
    -- CP-element group 21: 	22 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Update/cr
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_1_1363_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(21), ack => RPIPE_control_word_request_pipe_1_1363_inst_req_1); -- 
    processorToNicInterface_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(12) & processorToNicInterface_CP_2794_elements(22);
      gj_processorToNicInterface_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	35 
    -- CP-element group 22: 	21 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Sample/ra
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_1_1363_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_control_word_request_pipe_1_1363_inst_ack_0, ack => processorToNicInterface_CP_2794_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	13 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1361_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/RPIPE_control_word_request_pipe_1_1363_Update/ca
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:RPIPE_control_word_request_pipe_1_1363_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_control_word_request_pipe_1_1363_inst_ack_1, ack => processorToNicInterface_CP_2794_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Sample/rr
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:CONCAT_u42_u74_1373_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_2867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(24), ack => CONCAT_u42_u74_1373_inst_req_0); -- 
    processorToNicInterface_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(23) & processorToNicInterface_CP_2794_elements(18) & processorToNicInterface_CP_2794_elements(26);
      gj_processorToNicInterface_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Update/cr
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:CONCAT_u42_u74_1373_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(25), ack => CONCAT_u42_u74_1373_inst_req_1); -- 
    processorToNicInterface_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= processorToNicInterface_CP_2794_elements(29);
      gj_processorToNicInterface_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	19 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Sample/ra
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:CONCAT_u42_u74_1373_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_2868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u42_u74_1373_inst_ack_0, ack => processorToNicInterface_CP_2794_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/CONCAT_u42_u74_1373_Update/ca
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:CONCAT_u42_u74_1373_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u42_u74_1373_inst_ack_1, ack => processorToNicInterface_CP_2794_elements(27)); -- 
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Sample/req
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:WPIPE_AFB_NIC_REQUEST_1368_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(28), ack => WPIPE_AFB_NIC_REQUEST_1368_inst_req_0); -- 
    processorToNicInterface_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(27) & processorToNicInterface_CP_2794_elements(30);
      gj_processorToNicInterface_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Update/req
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:WPIPE_AFB_NIC_REQUEST_1368_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:WPIPE_AFB_NIC_REQUEST_1368_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_REQUEST_1368_inst_ack_0, ack => processorToNicInterface_CP_2794_elements(29)); -- 
    req_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => processorToNicInterface_CP_2794_elements(29), ack => WPIPE_AFB_NIC_REQUEST_1368_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/WPIPE_AFB_NIC_REQUEST_1368_Update/ack
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:WPIPE_AFB_NIC_REQUEST_1368_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_REQUEST_1368_inst_ack_1, ack => processorToNicInterface_CP_2794_elements(30)); -- 
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	10 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group processorToNicInterface_CP_2794_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => processorToNicInterface_CP_2794_elements(9), ack => processorToNicInterface_CP_2794_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	5 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_exit/$exit
      -- CP-element group 32: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_exit/ack
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:do_while_stmt_1356_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1356_branch_ack_0, ack => processorToNicInterface_CP_2794_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	5 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_taken/$exit
      -- CP-element group 33: 	 branch_block_stmt_1355/do_while_stmt_1356/loop_taken/ack
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:do_while_stmt_1356_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1356_branch_ack_1, ack => processorToNicInterface_CP_2794_elements(33)); -- 
    -- CP-element group 34:  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	3 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	1 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1355/do_while_stmt_1356/$exit
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_CP_2794_elements(34) <= processorToNicInterface_CP_2794_elements(3);
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: 	17 
    -- CP-element group 35: 	22 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	6 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/$exit
      -- CP-element group 35: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/aggregated_phi_sample_ack
      -- CP-element group 35: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1358_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1355/do_while_stmt_1356/do_while_stmt_1356_loop_body/phi_stmt_1361_sample_completed_
      -- 
    -- logger for CP element group processorToNicInterface_CP_2794_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and processorToNicInterface_CP_2794_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:processorToNicInterface:CP:processorToNicInterface_CP_2794_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    processorToNicInterface_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "processorToNicInterface_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= processorToNicInterface_CP_2794_elements(30) & processorToNicInterface_CP_2794_elements(17) & processorToNicInterface_CP_2794_elements(22);
      gj_processorToNicInterface_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(35), clk => clk, reset => reset); --
    end block;
    processorToNicInterface_do_while_stmt_1356_terminator_2897: loop_terminator -- 
      generic map (name => " processorToNicInterface_do_while_stmt_1356_terminator_2897", max_iterations_in_flight =>7) 
      port map(loop_body_exit => processorToNicInterface_CP_2794_elements(6),loop_continue => processorToNicInterface_CP_2794_elements(33),loop_terminate => processorToNicInterface_CP_2794_elements(32),loop_back => processorToNicInterface_CP_2794_elements(4),loop_exit => processorToNicInterface_CP_2794_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_2819_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= processorToNicInterface_CP_2794_elements(7);
        preds(1)  <= processorToNicInterface_CP_2794_elements(8);
        entry_tmerge_2819 : transition_merge -- 
          generic map(name => " entry_tmerge_2819")
          port map (preds => preds, symbol_out => processorToNicInterface_CP_2794_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u42_u74_1373_wire : std_logic_vector(73 downto 0);
    signal RPIPE_control_word_request_pipe_0_1360_wire : std_logic_vector(31 downto 0);
    signal RPIPE_control_word_request_pipe_1_1363_wire : std_logic_vector(63 downto 0);
    signal konst_1376_wire_constant : std_logic_vector(0 downto 0);
    signal rdata0_1358 : std_logic_vector(31 downto 0);
    signal rdata1_1361 : std_logic_vector(63 downto 0);
    signal slice_1371_wire : std_logic_vector(41 downto 0);
    -- 
  begin -- 
    konst_1376_wire_constant <= "1";
    -- logger for split-operator slice_1371_inst flow-through 
    process(slice_1371_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:slice_1371_inst:flowthrough inputs: " & " rdata1_1361 = "& Convert_SLV_To_Hex_String(rdata1_1361) & " outputs:" & " slice_1371_wire= "  & Convert_SLV_To_Hex_String(slice_1371_wire));
      --
    end process; 
    -- flow-through slice operator slice_1371_inst
    slice_1371_wire <= rdata1_1361(41 downto 0);
    -- logger for split-operator ssrc_phi_stmt_1358 flow-through 
    process(rdata0_1358) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:ssrc_phi_stmt_1358:flowthrough inputs: " & " RPIPE_control_word_request_pipe_0_1360_wire = "& Convert_SLV_To_Hex_String(RPIPE_control_word_request_pipe_0_1360_wire) & " outputs:" & " rdata0_1358= "  & Convert_SLV_To_Hex_String(rdata0_1358));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1358
    process(RPIPE_control_word_request_pipe_0_1360_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := RPIPE_control_word_request_pipe_0_1360_wire(31 downto 0);
      rdata0_1358 <= tmp_var; -- 
    end process;
    -- logger for split-operator ssrc_phi_stmt_1361 flow-through 
    process(rdata1_1361) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:ssrc_phi_stmt_1361:flowthrough inputs: " & " RPIPE_control_word_request_pipe_1_1363_wire = "& Convert_SLV_To_Hex_String(RPIPE_control_word_request_pipe_1_1363_wire) & " outputs:" & " rdata1_1361= "  & Convert_SLV_To_Hex_String(rdata1_1361));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1361
    process(RPIPE_control_word_request_pipe_1_1363_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := RPIPE_control_word_request_pipe_1_1363_wire(63 downto 0);
      rdata1_1361 <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1356_branch_req_0," req0 do_while_stmt_1356_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1356_branch_ack_0," ack0 do_while_stmt_1356_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1356_branch_ack_1," ack1 do_while_stmt_1356_branch");
    do_while_stmt_1356_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1376_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1356_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1356_branch_req_0,
          ack0 => do_while_stmt_1356_branch_ack_0,
          ack1 => do_while_stmt_1356_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator CONCAT_u42_u74_1373_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u42_u74_1373_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:CONCAT_u42_u74_1373_inst:started:   inputs: " & " slice_1371_wire = "& Convert_SLV_To_Hex_String(slice_1371_wire) & " rdata0_1358 = "& Convert_SLV_To_Hex_String(rdata0_1358));
          --
        end if; 
        if CONCAT_u42_u74_1373_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:CONCAT_u42_u74_1373_inst:finished:  outputs: " & " CONCAT_u42_u74_1373_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u42_u74_1373_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : CONCAT_u42_u74_1373_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(73 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_1371_wire & rdata0_1358;
      CONCAT_u42_u74_1373_wire <= data_out(73 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u42_u74_1373_inst_req_0;
      CONCAT_u42_u74_1373_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u42_u74_1373_inst_req_1;
      CONCAT_u42_u74_1373_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 42,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 74,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator RPIPE_control_word_request_pipe_0_1360_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_control_word_request_pipe_0_1360_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:RPIPE_control_word_request_pipe_0_1360_inst:started:   PipeRead from control_word_request_pipe_0 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_control_word_request_pipe_0_1360_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:RPIPE_control_word_request_pipe_0_1360_inst:finished:  outputs: " & " RPIPE_control_word_request_pipe_0_1360_wire= "  & Convert_SLV_To_Hex_String(RPIPE_control_word_request_pipe_0_1360_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_control_word_request_pipe_0_1360_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_control_word_request_pipe_0_1360_inst_req_0;
      RPIPE_control_word_request_pipe_0_1360_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_control_word_request_pipe_0_1360_inst_req_1;
      RPIPE_control_word_request_pipe_0_1360_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_control_word_request_pipe_0_1360_wire <= data_out(31 downto 0);
      control_word_request_pipe_0_read_0_gI: SplitGuardInterface generic map(name => "control_word_request_pipe_0_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      control_word_request_pipe_0_read_0: InputPortRevised -- 
        generic map ( name => "control_word_request_pipe_0_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => control_word_request_pipe_0_pipe_read_req(0),
          oack => control_word_request_pipe_0_pipe_read_ack(0),
          odata => control_word_request_pipe_0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator RPIPE_control_word_request_pipe_1_1363_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_control_word_request_pipe_1_1363_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:RPIPE_control_word_request_pipe_1_1363_inst:started:   PipeRead from control_word_request_pipe_1 inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_control_word_request_pipe_1_1363_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:RPIPE_control_word_request_pipe_1_1363_inst:finished:  outputs: " & " RPIPE_control_word_request_pipe_1_1363_wire= "  & Convert_SLV_To_Hex_String(RPIPE_control_word_request_pipe_1_1363_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (1) : RPIPE_control_word_request_pipe_1_1363_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_control_word_request_pipe_1_1363_inst_req_0;
      RPIPE_control_word_request_pipe_1_1363_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_control_word_request_pipe_1_1363_inst_req_1;
      RPIPE_control_word_request_pipe_1_1363_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_control_word_request_pipe_1_1363_wire <= data_out(63 downto 0);
      control_word_request_pipe_1_read_1_gI: SplitGuardInterface generic map(name => "control_word_request_pipe_1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      control_word_request_pipe_1_read_1: InputPortRevised -- 
        generic map ( name => "control_word_request_pipe_1_read_1", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => control_word_request_pipe_1_pipe_read_req(0),
          oack => control_word_request_pipe_1_pipe_read_ack(0),
          odata => control_word_request_pipe_1_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- logger for split-operator WPIPE_AFB_NIC_REQUEST_1368_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_AFB_NIC_REQUEST_1368_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:WPIPE_AFB_NIC_REQUEST_1368_inst:started:   PipeWrite to AFB_NIC_REQUEST inputs: " & " CONCAT_u42_u74_1373_wire = "& Convert_SLV_To_Hex_String(CONCAT_u42_u74_1373_wire));
          --
        end if; 
        if WPIPE_AFB_NIC_REQUEST_1368_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:processorToNicInterface:DP:WPIPE_AFB_NIC_REQUEST_1368_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_AFB_NIC_REQUEST_1368_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_REQUEST_1368_inst_req_0;
      WPIPE_AFB_NIC_REQUEST_1368_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_REQUEST_1368_inst_req_1;
      WPIPE_AFB_NIC_REQUEST_1368_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u42_u74_1373_wire;
      AFB_NIC_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST", data_width => 74, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_REQUEST_pipe_write_req(0),
          oack => AFB_NIC_REQUEST_pipe_write_ack(0),
          odata => AFB_NIC_REQUEST_pipe_write_data(73 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end processorToNicInterface_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity pushIntoQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_call_data : out  std_logic_vector(99 downto 0);
    setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_call_data : out  std_logic_vector(35 downto 0);
    releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
    releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
    releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
    acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_call_data : out  std_logic_vector(35 downto 0);
    acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
    acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
    acquireMutex_return_data : in   std_logic_vector(0 downto 0);
    acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity pushIntoQueue;
architecture pushIntoQueue_arch of pushIntoQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 69)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal pushIntoQueue_CP_999_start: Boolean;
  signal pushIntoQueue_CP_999_symbol: Boolean;
  -- volatile/operator module components. 
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_pointer : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_749_call_ack_0 : boolean;
  signal call_stmt_744_call_ack_1 : boolean;
  signal call_stmt_749_call_req_0 : boolean;
  signal call_stmt_766_call_req_0 : boolean;
  signal call_stmt_766_call_req_1 : boolean;
  signal call_stmt_744_call_ack_0 : boolean;
  signal call_stmt_744_call_req_0 : boolean;
  signal call_stmt_749_call_req_1 : boolean;
  signal call_stmt_771_call_ack_1 : boolean;
  signal call_stmt_744_call_req_1 : boolean;
  signal call_stmt_766_call_ack_1 : boolean;
  signal call_stmt_766_call_ack_0 : boolean;
  signal call_stmt_771_call_req_0 : boolean;
  signal call_stmt_771_call_ack_0 : boolean;
  signal call_stmt_771_call_req_1 : boolean;
  signal call_stmt_749_call_ack_1 : boolean;
  signal call_stmt_775_call_req_0 : boolean;
  signal call_stmt_775_call_ack_0 : boolean;
  signal call_stmt_775_call_req_1 : boolean;
  signal call_stmt_775_call_ack_1 : boolean;
  signal NOT_u1_u1_778_inst_req_0 : boolean;
  signal NOT_u1_u1_778_inst_ack_0 : boolean;
  signal NOT_u1_u1_778_inst_req_1 : boolean;
  signal NOT_u1_u1_778_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "pushIntoQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 69) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(68 downto 37) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(68 downto 37);
  in_buffer_data_in(tag_length + 68 downto 69) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 68 downto 69);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  pushIntoQueue_CP_999_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "pushIntoQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_999_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= pushIntoQueue_CP_999_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_999_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,pushIntoQueue_CP_999_start,"pushIntoQueue cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,pushIntoQueue_CP_999_symbol, "pushIntoQueue cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  pushIntoQueue_CP_999: Block -- control-path 
    signal pushIntoQueue_CP_999_elements: BooleanArray(14 downto 0);
    -- 
  begin -- 
    pushIntoQueue_CP_999_elements(0) <= pushIntoQueue_CP_999_start;
    pushIntoQueue_CP_999_symbol <= pushIntoQueue_CP_999_elements(14);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_744/$entry
      -- CP-element group 0: 	 call_stmt_744/call_stmt_744_update_start_
      -- CP-element group 0: 	 call_stmt_744/call_stmt_744_Update/$entry
      -- CP-element group 0: 	 call_stmt_744/call_stmt_744_Sample/crr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_744/call_stmt_744_Update/ccr
      -- CP-element group 0: 	 call_stmt_744/call_stmt_744_Sample/$entry
      -- CP-element group 0: 	 call_stmt_744/call_stmt_744_sample_start_
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_744_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_744_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(0), ack => call_stmt_744_call_req_0); -- 
    ccr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(0), ack => call_stmt_744_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_744/call_stmt_744_Sample/cra
      -- CP-element group 1: 	 call_stmt_744/call_stmt_744_sample_completed_
      -- CP-element group 1: 	 call_stmt_744/call_stmt_744_Sample/$exit
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_744_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_744_call_ack_0, ack => pushIntoQueue_CP_999_elements(1)); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2:  members (17) 
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_update_start_
      -- CP-element group 2: 	 call_stmt_744/call_stmt_744_Update/cca
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Sample/crr
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Update/$entry
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Update/$entry
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_update_start_
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/$entry
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_sample_start_
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Update/ccr
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Update/ccr
      -- CP-element group 2: 	 call_stmt_744/call_stmt_744_Update/$exit
      -- CP-element group 2: 	 call_stmt_744/$exit
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Sample/$entry
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Update/$entry
      -- CP-element group 2: 	 call_stmt_744/call_stmt_744_update_completed_
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Update/ccr
      -- CP-element group 2: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_update_start_
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_744_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_749_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_749_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_771_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_766_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_744_call_ack_1, ack => pushIntoQueue_CP_999_elements(2)); -- 
    crr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(2), ack => call_stmt_749_call_req_0); -- 
    ccr_1034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(2), ack => call_stmt_749_call_req_1); -- 
    ccr_1062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(2), ack => call_stmt_771_call_req_1); -- 
    ccr_1048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(2), ack => call_stmt_766_call_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_sample_completed_
      -- CP-element group 3: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Sample/cra
      -- CP-element group 3: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Sample/$exit
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_749_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_749_call_ack_0, ack => pushIntoQueue_CP_999_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Sample/crr
      -- CP-element group 4: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_update_completed_
      -- CP-element group 4: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Update/$exit
      -- CP-element group 4: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Sample/$entry
      -- CP-element group 4: 	 call_stmt_749_to_call_stmt_771/call_stmt_749_Update/cca
      -- CP-element group 4: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_sample_start_
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(4) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_749_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_766_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_1035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_749_call_ack_1, ack => pushIntoQueue_CP_999_elements(4)); -- 
    crr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(4), ack => call_stmt_766_call_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Sample/$exit
      -- CP-element group 5: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Sample/cra
      -- CP-element group 5: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_sample_completed_
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_766_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_766_call_ack_0, ack => pushIntoQueue_CP_999_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_update_completed_
      -- CP-element group 6: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Update/cca
      -- CP-element group 6: 	 call_stmt_749_to_call_stmt_771/call_stmt_766_Update/$exit
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_766_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_766_call_ack_1, ack => pushIntoQueue_CP_999_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Sample/$entry
      -- CP-element group 7: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_sample_start_
      -- CP-element group 7: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Sample/crr
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(7) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_771_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(7), ack => call_stmt_771_call_req_0); -- 
    pushIntoQueue_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "pushIntoQueue_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_999_elements(4) & pushIntoQueue_CP_999_elements(6);
      gj_pushIntoQueue_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_999_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Sample/$exit
      -- CP-element group 8: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_sample_completed_
      -- CP-element group 8: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Sample/cra
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(8) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_771_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_771_call_ack_0, ack => pushIntoQueue_CP_999_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (17) 
      -- CP-element group 9: 	 call_stmt_749_to_call_stmt_771/$exit
      -- CP-element group 9: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_update_completed_
      -- CP-element group 9: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Update/cca
      -- CP-element group 9: 	 call_stmt_749_to_call_stmt_771/call_stmt_771_Update/$exit
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/$entry
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_sample_start_
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_update_start_
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Sample/$entry
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Sample/crr
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Update/$entry
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Update/ccr
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_sample_start_
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_update_start_
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Sample/$entry
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Sample/rr
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Update/$entry
      -- CP-element group 9: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Update/cr
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(9) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_771_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:NOT_u1_u1_778_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:NOT_u1_u1_778_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_775_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_775_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_771_call_ack_1, ack => pushIntoQueue_CP_999_elements(9)); -- 
    rr_1088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(9), ack => NOT_u1_u1_778_inst_req_0); -- 
    cr_1093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(9), ack => NOT_u1_u1_778_inst_req_1); -- 
    crr_1074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(9), ack => call_stmt_775_call_req_0); -- 
    ccr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_999_elements(9), ack => call_stmt_775_call_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_sample_completed_
      -- CP-element group 10: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Sample/$exit
      -- CP-element group 10: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Sample/cra
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_775_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_1075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_775_call_ack_0, ack => pushIntoQueue_CP_999_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_update_completed_
      -- CP-element group 11: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Update/$exit
      -- CP-element group 11: 	 call_stmt_775_to_assign_stmt_779/call_stmt_775_Update/cca
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(11) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:call_stmt_775_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_775_call_ack_1, ack => pushIntoQueue_CP_999_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_sample_completed_
      -- CP-element group 12: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Sample/$exit
      -- CP-element group 12: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Sample/ra
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:NOT_u1_u1_778_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_1089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_778_inst_ack_0, ack => pushIntoQueue_CP_999_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_update_completed_
      -- CP-element group 13: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Update/$exit
      -- CP-element group 13: 	 call_stmt_775_to_assign_stmt_779/NOT_u1_u1_778_Update/ca
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(13) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:NOT_u1_u1_778_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_1094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_778_inst_ack_1, ack => pushIntoQueue_CP_999_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 $exit
      -- CP-element group 14: 	 call_stmt_775_to_assign_stmt_779/$exit
      -- 
    -- logger for CP element group pushIntoQueue_CP_999_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and pushIntoQueue_CP_999_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:pushIntoQueue:CP:pushIntoQueue_CP_999_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    pushIntoQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_999_elements(11) & pushIntoQueue_CP_999_elements(13);
      gj_pushIntoQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_999_elements(14), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_753_wire : std_logic_vector(31 downto 0);
    signal R_QUEUE_SIZE_MASK_754_wire_constant : std_logic_vector(31 downto 0);
    signal konst_752_wire_constant : std_logic_vector(31 downto 0);
    signal m_ok_744 : std_logic_vector(0 downto 0);
    signal next_wp_756 : std_logic_vector(31 downto 0);
    signal q_full_761 : std_logic_vector(0 downto 0);
    signal read_pointer_749 : std_logic_vector(31 downto 0);
    signal write_pointer_749 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    R_QUEUE_SIZE_MASK_754_wire_constant <= "00000000000000000000000100000000";
    konst_752_wire_constant <= "00000000000000000000000000000001";
    -- logger for split-operator ADD_u32_u32_753_inst flow-through 
    process(ADD_u32_u32_753_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:ADD_u32_u32_753_inst:flowthrough inputs: " & " write_pointer_749 = "& Convert_SLV_To_Hex_String(write_pointer_749) & " konst_752_wire_constant = "& Convert_SLV_To_Hex_String(konst_752_wire_constant) & " outputs:" & " ADD_u32_u32_753_wire= "  & Convert_SLV_To_Hex_String(ADD_u32_u32_753_wire));
      --
    end process; 
    -- binary operator ADD_u32_u32_753_inst
    process(write_pointer_749) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(write_pointer_749, konst_752_wire_constant, tmp_var);
      ADD_u32_u32_753_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u32_u32_755_inst flow-through 
    process(next_wp_756) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:AND_u32_u32_755_inst:flowthrough inputs: " & " ADD_u32_u32_753_wire = "& Convert_SLV_To_Hex_String(ADD_u32_u32_753_wire) & " R_QUEUE_SIZE_MASK_754_wire_constant = "& Convert_SLV_To_Hex_String(R_QUEUE_SIZE_MASK_754_wire_constant) & " outputs:" & " next_wp_756= "  & Convert_SLV_To_Hex_String(next_wp_756));
      --
    end process; 
    -- binary operator AND_u32_u32_755_inst
    process(ADD_u32_u32_753_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ADD_u32_u32_753_wire, R_QUEUE_SIZE_MASK_754_wire_constant, tmp_var);
      next_wp_756 <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u32_u1_760_inst flow-through 
    process(q_full_761) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:EQ_u32_u1_760_inst:flowthrough inputs: " & " next_wp_756 = "& Convert_SLV_To_Hex_String(next_wp_756) & " read_pointer_749 = "& Convert_SLV_To_Hex_String(read_pointer_749) & " outputs:" & " q_full_761= "  & Convert_SLV_To_Hex_String(q_full_761));
      --
    end process; 
    -- binary operator EQ_u32_u1_760_inst
    process(next_wp_756, read_pointer_749) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_wp_756, read_pointer_749, tmp_var);
      q_full_761 <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_778_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if NOT_u1_u1_778_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:NOT_u1_u1_778_inst:started:   inputs: " & " q_full_761 = "& Convert_SLV_To_Hex_String(q_full_761));
          --
        end if; 
        if NOT_u1_u1_778_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:NOT_u1_u1_778_inst:finished:  outputs: " & " status_buffer= "  & Convert_SLV_To_Hex_String(status_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (3) : NOT_u1_u1_778_inst 
    ApIntNot_group_3: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= q_full_761;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_778_inst_req_0;
      NOT_u1_u1_778_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_778_inst_req_1;
      NOT_u1_u1_778_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_3_gI: SplitGuardInterface generic map(name => "ApIntNot_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- logger for split-operator call_stmt_744_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_744_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_744_call:started:  Call to module acquireMutex inputs: " & " lock_buffer (guard)= " & Convert_SLV_To_String(lock_buffer) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer));
          --
        end if; 
        if call_stmt_744_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_744_call:finished:  outputs: " & " m_ok_744= "  & Convert_SLV_To_Hex_String(m_ok_744));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_744_call 
    acquireMutex_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_744_call_req_0;
      call_stmt_744_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_744_call_req_1;
      call_stmt_744_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireMutex_call_group_0_gI: SplitGuardInterface generic map(name => "acquireMutex_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_744 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireMutex_call_reqs(0),
          ackR => acquireMutex_call_acks(0),
          dataR => acquireMutex_call_data(35 downto 0),
          tagR => acquireMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireMutex_return_acks(0), -- cross-over
          ackL => acquireMutex_return_reqs(0), -- cross-over
          dataL => acquireMutex_return_data(0 downto 0),
          tagL => acquireMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_749_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_749_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_749_call:started:  Call to module getQueuePointers inputs: " & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer));
          --
        end if; 
        if call_stmt_749_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_749_call:finished:  outputs: " & " write_pointer_749= "  & Convert_SLV_To_Hex_String(write_pointer_749) & " read_pointer_749= "  & Convert_SLV_To_Hex_String(read_pointer_749));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_749_call 
    getQueuePointers_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_749_call_req_0;
      call_stmt_749_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_749_call_req_1;
      call_stmt_749_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_1_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_pointer_749 <= data_out(63 downto 32);
      read_pointer_749 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_766_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_766_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_766_call:started:  Call to module setQueueElement inputs: " & " q_full_761 (guard complement )= " & Convert_SLV_To_String(q_full_761) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " write_pointer_749 = "& Convert_SLV_To_Hex_String(write_pointer_749) & " q_w_data_buffer = "& Convert_SLV_To_Hex_String(q_w_data_buffer));
          --
        end if; 
        if call_stmt_766_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_766_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_766_call 
    setQueueElement_call_group_2: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_766_call_req_0;
      call_stmt_766_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_766_call_req_1;
      call_stmt_766_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_761(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueueElement_call_group_2_gI: SplitGuardInterface generic map(name => "setQueueElement_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_pointer_749 & q_w_data_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueueElement_call_reqs(0),
          ackR => setQueueElement_call_acks(0),
          dataR => setQueueElement_call_data(99 downto 0),
          tagR => setQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueueElement_return_acks(0), -- cross-over
          ackL => setQueueElement_return_reqs(0), -- cross-over
          tagL => setQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- logger for split-operator call_stmt_771_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_771_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_771_call:started:  Call to module setQueuePointers inputs: " & " q_full_761 (guard complement )= " & Convert_SLV_To_String(q_full_761) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " write_pointer_749 = "& Convert_SLV_To_Hex_String(write_pointer_749) & " next_wp_756 = "& Convert_SLV_To_Hex_String(next_wp_756));
          --
        end if; 
        if call_stmt_771_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_771_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (3) : call_stmt_771_call 
    setQueuePointers_call_group_3: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_771_call_req_0;
      call_stmt_771_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_771_call_req_1;
      call_stmt_771_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_761(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_3_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_pointer_749 & next_wp_756;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- logger for split-operator call_stmt_775_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_775_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_775_call:started:  Call to module releaseMutex inputs: " & " lock_buffer (guard)= " & Convert_SLV_To_String(lock_buffer) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer));
          --
        end if; 
        if call_stmt_775_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:pushIntoQueue:DP:call_stmt_775_call:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (4) : call_stmt_775_call 
    releaseMutex_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_775_call_req_0;
      call_stmt_775_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_775_call_req_1;
      call_stmt_775_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_buffer(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseMutex_call_group_4_gI: SplitGuardInterface generic map(name => "releaseMutex_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseMutex_call_reqs(0),
          ackR => releaseMutex_call_acks(0),
          dataR => releaseMutex_call_data(35 downto 0),
          tagR => releaseMutex_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseMutex_return_acks(0), -- cross-over
          ackL => releaseMutex_return_reqs(0), -- cross-over
          tagL => releaseMutex_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end pushIntoQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity releaseMutex is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity releaseMutex;
architecture releaseMutex_arch of releaseMutex is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal releaseMutex_CP_490_start: Boolean;
  signal releaseMutex_CP_490_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_450_call_ack_1 : boolean;
  signal call_stmt_450_call_req_1 : boolean;
  signal call_stmt_450_call_ack_0 : boolean;
  signal call_stmt_450_call_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "releaseMutex_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  releaseMutex_CP_490_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "releaseMutex_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseMutex_CP_490_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= releaseMutex_CP_490_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseMutex_CP_490_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,releaseMutex_CP_490_start,"releaseMutex cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,releaseMutex_CP_490_symbol, "releaseMutex cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  releaseMutex_CP_490: Block -- control-path 
    signal releaseMutex_CP_490_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    releaseMutex_CP_490_elements(0) <= releaseMutex_CP_490_start;
    releaseMutex_CP_490_symbol <= releaseMutex_CP_490_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_450/call_stmt_450_Update/ccr
      -- CP-element group 0: 	 call_stmt_450/call_stmt_450_Update/$entry
      -- CP-element group 0: 	 call_stmt_450/call_stmt_450_update_start_
      -- CP-element group 0: 	 call_stmt_450/$entry
      -- CP-element group 0: 	 call_stmt_450/call_stmt_450_Sample/crr
      -- CP-element group 0: 	 call_stmt_450/call_stmt_450_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_450/call_stmt_450_sample_start_
      -- 
    -- logger for CP element group releaseMutex_CP_490_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and releaseMutex_CP_490_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:releaseMutex:CP:releaseMutex_CP_490_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:releaseMutex:CP:call_stmt_450_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:releaseMutex:CP:call_stmt_450_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseMutex_CP_490_elements(0), ack => call_stmt_450_call_req_0); -- 
    ccr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseMutex_CP_490_elements(0), ack => call_stmt_450_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_450/call_stmt_450_Sample/cra
      -- CP-element group 1: 	 call_stmt_450/call_stmt_450_Sample/$exit
      -- CP-element group 1: 	 call_stmt_450/call_stmt_450_sample_completed_
      -- 
    -- logger for CP element group releaseMutex_CP_490_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and releaseMutex_CP_490_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:releaseMutex:CP:releaseMutex_CP_490_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:releaseMutex:CP:call_stmt_450_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_450_call_ack_0, ack => releaseMutex_CP_490_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_450/call_stmt_450_Update/cca
      -- CP-element group 2: 	 call_stmt_450/call_stmt_450_Update/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_450/$exit
      -- CP-element group 2: 	 call_stmt_450/call_stmt_450_update_completed_
      -- 
    -- logger for CP element group releaseMutex_CP_490_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and releaseMutex_CP_490_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:releaseMutex:CP:releaseMutex_CP_490_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:releaseMutex:CP:call_stmt_450_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_450_call_ack_1, ack => releaseMutex_CP_490_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u4_u8_445_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_450 : std_logic_vector(63 downto 0);
    signal type_cast_437_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_439_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_448_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_445_wire_constant <= "11110000";
    type_cast_437_wire_constant <= "0";
    type_cast_439_wire_constant <= "0";
    type_cast_448_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- logger for split-operator call_stmt_450_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_450_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:releaseMutex:DP:call_stmt_450_call:started:  Call to module accessMemory inputs: " & " type_cast_437_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_437_wire_constant) & " type_cast_439_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_439_wire_constant) & " CONCAT_u4_u8_445_wire_constant = "& Convert_SLV_To_Hex_String(CONCAT_u4_u8_445_wire_constant) & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " type_cast_448_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_448_wire_constant));
          --
        end if; 
        if call_stmt_450_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:releaseMutex:DP:call_stmt_450_call:finished:  outputs: " & " ignore_450= "  & Convert_SLV_To_Hex_String(ignore_450));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_450_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_450_call_req_0;
      call_stmt_450_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_450_call_req_1;
      call_stmt_450_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_437_wire_constant & type_cast_439_wire_constant & CONCAT_u4_u8_445_wire_constant & q_base_address_buffer & type_cast_448_wire_constant;
      ignore_450 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end releaseMutex_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity setQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    write_pointer : in  std_logic_vector(31 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueueElement;
architecture setQueueElement_arch of setQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal write_pointer_buffer :  std_logic_vector(31 downto 0);
  signal write_pointer_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal setQueueElement_CP_979_start: Boolean;
  signal setQueueElement_CP_979_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_734_call_req_0 : boolean;
  signal call_stmt_734_call_ack_0 : boolean;
  signal call_stmt_734_call_ack_1 : boolean;
  signal call_stmt_734_call_req_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= write_pointer;
  write_pointer_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueueElement_CP_979_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_979_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueueElement_CP_979_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_979_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,setQueueElement_CP_979_start,"setQueueElement cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,setQueueElement_CP_979_symbol, "setQueueElement cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueueElement_CP_979: Block -- control-path 
    signal setQueueElement_CP_979_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueueElement_CP_979_elements(0) <= setQueueElement_CP_979_start;
    setQueueElement_CP_979_symbol <= setQueueElement_CP_979_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Sample/crr
      -- CP-element group 0: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_update_start_
      -- CP-element group 0: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_sample_start_
      -- CP-element group 0: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_683_to_call_stmt_734/$entry
      -- CP-element group 0: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Update/ccr
      -- 
    -- logger for CP element group setQueueElement_CP_979_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and setQueueElement_CP_979_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueueElement:CP:setQueueElement_CP_979_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueueElement:CP:call_stmt_734_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueueElement:CP:call_stmt_734_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_979_elements(0), ack => call_stmt_734_call_req_0); -- 
    ccr_997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_979_elements(0), ack => call_stmt_734_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_sample_completed_
      -- CP-element group 1: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Sample/cra
      -- 
    -- logger for CP element group setQueueElement_CP_979_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and setQueueElement_CP_979_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueueElement:CP:setQueueElement_CP_979_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueueElement:CP:call_stmt_734_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_734_call_ack_0, ack => setQueueElement_CP_979_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_update_completed_
      -- CP-element group 2: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Update/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_683_to_call_stmt_734/call_stmt_734_Update/cca
      -- CP-element group 2: 	 assign_stmt_683_to_call_stmt_734/$exit
      -- 
    -- logger for CP element group setQueueElement_CP_979_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and setQueueElement_CP_979_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueueElement:CP:setQueueElement_CP_979_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueueElement:CP:call_stmt_734_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_734_call_ack_1, ack => setQueueElement_CP_979_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_697_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_715_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_690_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u32_u64_719_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_723_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_703_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_709_wire_constant : std_logic_vector(7 downto 0);
    signal bmask_711 : std_logic_vector(7 downto 0);
    signal buffer_address_683 : std_logic_vector(35 downto 0);
    signal element_pair_address_693 : std_logic_vector(35 downto 0);
    signal ignore_734 : std_logic_vector(63 downto 0);
    signal konst_696_wire_constant : std_logic_vector(31 downto 0);
    signal konst_714_wire_constant : std_logic_vector(31 downto 0);
    signal slice_687_wire : std_logic_vector(30 downto 0);
    signal type_cast_681_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_689_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_691_wire : std_logic_vector(35 downto 0);
    signal type_cast_717_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_722_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_727_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_729_wire_constant : std_logic_vector(0 downto 0);
    signal wval_725 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_703_wire_constant <= "00001111";
    CONCAT_u4_u8_709_wire_constant <= "11110000";
    konst_696_wire_constant <= "00000000000000000000000000000000";
    konst_714_wire_constant <= "00000000000000000000000000000000";
    type_cast_681_wire_constant <= "000000000000000000000000000000010000";
    type_cast_689_wire_constant <= "000";
    type_cast_717_wire_constant <= "00000000000000000000000000000000";
    type_cast_722_wire_constant <= "00000000000000000000000000000000";
    type_cast_727_wire_constant <= "0";
    type_cast_729_wire_constant <= "0";
    -- logger for split-operator MUX_710_inst flow-through 
    process(bmask_711) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:MUX_710_inst:flowthrough inputs: " & " BITSEL_u32_u1_697_wire = "& Convert_SLV_To_Hex_String(BITSEL_u32_u1_697_wire) & " CONCAT_u4_u8_703_wire_constant = "& Convert_SLV_To_Hex_String(CONCAT_u4_u8_703_wire_constant) & " CONCAT_u4_u8_709_wire_constant = "& Convert_SLV_To_Hex_String(CONCAT_u4_u8_709_wire_constant) & " outputs:" & " bmask_711= "  & Convert_SLV_To_Hex_String(bmask_711));
      --
    end process; 
    -- flow-through select operator MUX_710_inst
    bmask_711 <= CONCAT_u4_u8_703_wire_constant when (BITSEL_u32_u1_697_wire(0) /=  '0') else CONCAT_u4_u8_709_wire_constant;
    -- logger for split-operator MUX_724_inst flow-through 
    process(wval_725) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:MUX_724_inst:flowthrough inputs: " & " BITSEL_u32_u1_715_wire = "& Convert_SLV_To_Hex_String(BITSEL_u32_u1_715_wire) & " CONCAT_u32_u64_719_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_719_wire) & " CONCAT_u32_u64_723_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_723_wire) & " outputs:" & " wval_725= "  & Convert_SLV_To_Hex_String(wval_725));
      --
    end process; 
    -- flow-through select operator MUX_724_inst
    wval_725 <= CONCAT_u32_u64_719_wire when (BITSEL_u32_u1_715_wire(0) /=  '0') else CONCAT_u32_u64_723_wire;
    -- logger for split-operator slice_687_inst flow-through 
    process(slice_687_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:slice_687_inst:flowthrough inputs: " & " write_pointer_buffer = "& Convert_SLV_To_Hex_String(write_pointer_buffer) & " outputs:" & " slice_687_wire= "  & Convert_SLV_To_Hex_String(slice_687_wire));
      --
    end process; 
    -- flow-through slice operator slice_687_inst
    slice_687_wire <= write_pointer_buffer(31 downto 1);
    -- logger for split-operator type_cast_691_inst flow-through 
    process(type_cast_691_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:type_cast_691_inst:flowthrough inputs: " & " CONCAT_u31_u34_690_wire = "& Convert_SLV_To_Hex_String(CONCAT_u31_u34_690_wire) & " outputs:" & " type_cast_691_wire= "  & Convert_SLV_To_Hex_String(type_cast_691_wire));
      --
    end process; 
    -- interlock type_cast_691_inst
    process(CONCAT_u31_u34_690_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_690_wire(33 downto 0);
      type_cast_691_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator ADD_u36_u36_682_inst flow-through 
    process(buffer_address_683) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:ADD_u36_u36_682_inst:flowthrough inputs: " & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " type_cast_681_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_681_wire_constant) & " outputs:" & " buffer_address_683= "  & Convert_SLV_To_Hex_String(buffer_address_683));
      --
    end process; 
    -- binary operator ADD_u36_u36_682_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_681_wire_constant, tmp_var);
      buffer_address_683 <= tmp_var; --
    end process;
    -- logger for split-operator ADD_u36_u36_692_inst flow-through 
    process(element_pair_address_693) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:ADD_u36_u36_692_inst:flowthrough inputs: " & " buffer_address_683 = "& Convert_SLV_To_Hex_String(buffer_address_683) & " type_cast_691_wire = "& Convert_SLV_To_Hex_String(type_cast_691_wire) & " outputs:" & " element_pair_address_693= "  & Convert_SLV_To_Hex_String(element_pair_address_693));
      --
    end process; 
    -- binary operator ADD_u36_u36_692_inst
    process(buffer_address_683, type_cast_691_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_683, type_cast_691_wire, tmp_var);
      element_pair_address_693 <= tmp_var; --
    end process;
    -- logger for split-operator BITSEL_u32_u1_697_inst flow-through 
    process(BITSEL_u32_u1_697_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:BITSEL_u32_u1_697_inst:flowthrough inputs: " & " write_pointer_buffer = "& Convert_SLV_To_Hex_String(write_pointer_buffer) & " konst_696_wire_constant = "& Convert_SLV_To_Hex_String(konst_696_wire_constant) & " outputs:" & " BITSEL_u32_u1_697_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u32_u1_697_wire));
      --
    end process; 
    -- binary operator BITSEL_u32_u1_697_inst
    process(write_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_pointer_buffer, konst_696_wire_constant, tmp_var);
      BITSEL_u32_u1_697_wire <= tmp_var; --
    end process;
    -- logger for split-operator BITSEL_u32_u1_715_inst flow-through 
    process(BITSEL_u32_u1_715_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:BITSEL_u32_u1_715_inst:flowthrough inputs: " & " write_pointer_buffer = "& Convert_SLV_To_Hex_String(write_pointer_buffer) & " konst_714_wire_constant = "& Convert_SLV_To_Hex_String(konst_714_wire_constant) & " outputs:" & " BITSEL_u32_u1_715_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u32_u1_715_wire));
      --
    end process; 
    -- binary operator BITSEL_u32_u1_715_inst
    process(write_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_pointer_buffer, konst_714_wire_constant, tmp_var);
      BITSEL_u32_u1_715_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u31_u34_690_inst flow-through 
    process(CONCAT_u31_u34_690_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:CONCAT_u31_u34_690_inst:flowthrough inputs: " & " slice_687_wire = "& Convert_SLV_To_Hex_String(slice_687_wire) & " type_cast_689_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_689_wire_constant) & " outputs:" & " CONCAT_u31_u34_690_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u31_u34_690_wire));
      --
    end process; 
    -- binary operator CONCAT_u31_u34_690_inst
    process(slice_687_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_687_wire, type_cast_689_wire_constant, tmp_var);
      CONCAT_u31_u34_690_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_719_inst flow-through 
    process(CONCAT_u32_u64_719_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:CONCAT_u32_u64_719_inst:flowthrough inputs: " & " type_cast_717_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_717_wire_constant) & " q_w_data_buffer = "& Convert_SLV_To_Hex_String(q_w_data_buffer) & " outputs:" & " CONCAT_u32_u64_719_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_719_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_719_inst
    process(type_cast_717_wire_constant, q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_717_wire_constant, q_w_data_buffer, tmp_var);
      CONCAT_u32_u64_719_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_723_inst flow-through 
    process(CONCAT_u32_u64_723_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:CONCAT_u32_u64_723_inst:flowthrough inputs: " & " q_w_data_buffer = "& Convert_SLV_To_Hex_String(q_w_data_buffer) & " type_cast_722_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_722_wire_constant) & " outputs:" & " CONCAT_u32_u64_723_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_723_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_723_inst
    process(q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(q_w_data_buffer, type_cast_722_wire_constant, tmp_var);
      CONCAT_u32_u64_723_wire <= tmp_var; --
    end process;
    -- logger for split-operator call_stmt_734_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_734_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:call_stmt_734_call:started:  Call to module accessMemory inputs: " & " type_cast_727_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_727_wire_constant) & " type_cast_729_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_729_wire_constant) & " bmask_711 = "& Convert_SLV_To_Hex_String(bmask_711) & " element_pair_address_693 = "& Convert_SLV_To_Hex_String(element_pair_address_693) & " wval_725 = "& Convert_SLV_To_Hex_String(wval_725));
          --
        end if; 
        if call_stmt_734_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:setQueueElement:DP:call_stmt_734_call:finished:  outputs: " & " ignore_734= "  & Convert_SLV_To_Hex_String(ignore_734));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_734_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_734_call_req_0;
      call_stmt_734_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_734_call_req_1;
      call_stmt_734_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_727_wire_constant & type_cast_729_wire_constant & bmask_711 & element_pair_address_693 & wval_725;
      ignore_734 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity setQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : in  std_logic_vector(31 downto 0);
    rp : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueuePointers;
architecture setQueuePointers_arch of setQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  -- output port buffer signals
  signal setQueuePointers_CP_470_start: Boolean;
  signal setQueuePointers_CP_470_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_432_call_ack_1 : boolean;
  signal call_stmt_432_call_req_1 : boolean;
  signal call_stmt_432_call_ack_0 : boolean;
  signal call_stmt_432_call_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= wp;
  wp_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= rp;
  rp_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueuePointers_CP_470_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_470_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueuePointers_CP_470_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_470_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,setQueuePointers_CP_470_start,"setQueuePointers cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,setQueuePointers_CP_470_symbol, "setQueuePointers cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueuePointers_CP_470: Block -- control-path 
    signal setQueuePointers_CP_470_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueuePointers_CP_470_elements(0) <= setQueuePointers_CP_470_start;
    setQueuePointers_CP_470_symbol <= setQueuePointers_CP_470_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_432/call_stmt_432_sample_start_
      -- CP-element group 0: 	 call_stmt_432/call_stmt_432_Update/ccr
      -- CP-element group 0: 	 call_stmt_432/call_stmt_432_Update/$entry
      -- CP-element group 0: 	 call_stmt_432/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_432/call_stmt_432_Sample/crr
      -- CP-element group 0: 	 call_stmt_432/call_stmt_432_Sample/$entry
      -- CP-element group 0: 	 call_stmt_432/call_stmt_432_update_start_
      -- 
    -- logger for CP element group setQueuePointers_CP_470_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and setQueuePointers_CP_470_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueuePointers:CP:setQueuePointers_CP_470_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueuePointers:CP:call_stmt_432_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueuePointers:CP:call_stmt_432_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_470_elements(0), ack => call_stmt_432_call_req_0); -- 
    ccr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_470_elements(0), ack => call_stmt_432_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_432/call_stmt_432_sample_completed_
      -- CP-element group 1: 	 call_stmt_432/call_stmt_432_Sample/cra
      -- CP-element group 1: 	 call_stmt_432/call_stmt_432_Sample/$exit
      -- 
    -- logger for CP element group setQueuePointers_CP_470_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and setQueuePointers_CP_470_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueuePointers:CP:setQueuePointers_CP_470_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueuePointers:CP:call_stmt_432_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_432_call_ack_0, ack => setQueuePointers_CP_470_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 call_stmt_432/$exit
      -- CP-element group 2: 	 call_stmt_432/call_stmt_432_Update/cca
      -- CP-element group 2: 	 call_stmt_432/call_stmt_432_Update/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_432/call_stmt_432_update_completed_
      -- 
    -- logger for CP element group setQueuePointers_CP_470_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and setQueuePointers_CP_470_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueuePointers:CP:setQueuePointers_CP_470_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:setQueuePointers:CP:call_stmt_432_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_432_call_ack_1, ack => setQueuePointers_CP_470_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_427_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u32_u64_430_wire : std_logic_vector(63 downto 0);
    signal NOT_u8_u8_424_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_432 : std_logic_vector(63 downto 0);
    signal konst_426_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_419_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_421_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_424_wire_constant <= "11111111";
    konst_426_wire_constant <= "000000000000000000000000000000001000";
    type_cast_419_wire_constant <= "0";
    type_cast_421_wire_constant <= "0";
    -- logger for split-operator ADD_u36_u36_427_inst flow-through 
    process(ADD_u36_u36_427_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueuePointers:DP:ADD_u36_u36_427_inst:flowthrough inputs: " & " q_base_address_buffer = "& Convert_SLV_To_Hex_String(q_base_address_buffer) & " konst_426_wire_constant = "& Convert_SLV_To_Hex_String(konst_426_wire_constant) & " outputs:" & " ADD_u36_u36_427_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_427_wire));
      --
    end process; 
    -- binary operator ADD_u36_u36_427_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_426_wire_constant, tmp_var);
      ADD_u36_u36_427_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u32_u64_430_inst flow-through 
    process(CONCAT_u32_u64_430_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:setQueuePointers:DP:CONCAT_u32_u64_430_inst:flowthrough inputs: " & " wp_buffer = "& Convert_SLV_To_Hex_String(wp_buffer) & " rp_buffer = "& Convert_SLV_To_Hex_String(rp_buffer) & " outputs:" & " CONCAT_u32_u64_430_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u32_u64_430_wire));
      --
    end process; 
    -- binary operator CONCAT_u32_u64_430_inst
    process(wp_buffer, rp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(wp_buffer, rp_buffer, tmp_var);
      CONCAT_u32_u64_430_wire <= tmp_var; --
    end process;
    -- logger for split-operator call_stmt_432_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_432_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:setQueuePointers:DP:call_stmt_432_call:started:  Call to module accessMemory inputs: " & " type_cast_419_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_419_wire_constant) & " type_cast_421_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_421_wire_constant) & " NOT_u8_u8_424_wire_constant = "& Convert_SLV_To_Hex_String(NOT_u8_u8_424_wire_constant) & " ADD_u36_u36_427_wire = "& Convert_SLV_To_Hex_String(ADD_u36_u36_427_wire) & " CONCAT_u32_u64_430_wire = "& Convert_SLV_To_Hex_String(CONCAT_u32_u64_430_wire));
          --
        end if; 
        if call_stmt_432_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:setQueuePointers:DP:call_stmt_432_call:finished:  outputs: " & " ignore_432= "  & Convert_SLV_To_Hex_String(ignore_432));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_432_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_432_call_req_0;
      call_stmt_432_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_432_call_req_1;
      call_stmt_432_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_419_wire_constant & type_cast_421_wire_constant & NOT_u8_u8_424_wire_constant & ADD_u36_u36_427_wire & CONCAT_u32_u64_430_wire;
      ignore_432 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity transmitEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
    getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
    getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
    transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_call_data : out  std_logic_vector(31 downto 0);
    transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
    transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_return_data : in   std_logic_vector(0 downto 0);
    transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitEngineDaemon;
architecture transmitEngineDaemon_arch of transmitEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal transmitEngineDaemon_CP_3152_start: Boolean;
  signal transmitEngineDaemon_CP_3152_symbol: Boolean;
  -- volatile/operator module components. 
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_1 : boolean;
  signal AND_u6_u6_1515_inst_req_0 : boolean;
  signal call_stmt_1524_call_ack_0 : boolean;
  signal AND_u6_u6_1515_inst_ack_0 : boolean;
  signal call_stmt_1536_call_ack_1 : boolean;
  signal call_stmt_1536_call_ack_0 : boolean;
  signal call_stmt_1520_call_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_1 : boolean;
  signal call_stmt_1536_call_req_0 : boolean;
  signal call_stmt_1524_call_req_0 : boolean;
  signal call_stmt_1520_call_req_1 : boolean;
  signal call_stmt_1520_call_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_1 : boolean;
  signal if_stmt_1497_branch_ack_0 : boolean;
  signal do_while_stmt_1504_branch_req_0 : boolean;
  signal call_stmt_1520_call_req_0 : boolean;
  signal call_stmt_1536_call_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_0 : boolean;
  signal if_stmt_1497_branch_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_0 : boolean;
  signal do_while_stmt_1504_branch_ack_0 : boolean;
  signal call_stmt_1524_call_ack_1 : boolean;
  signal call_stmt_1524_call_req_1 : boolean;
  signal do_while_stmt_1504_branch_ack_1 : boolean;
  signal if_stmt_1497_branch_req_0 : boolean;
  signal AND_u6_u6_1515_inst_ack_1 : boolean;
  signal AND_u6_u6_1515_inst_req_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitEngineDaemon_CP_3152_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3152_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3152_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_3152_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,transmitEngineDaemon_CP_3152_start,"transmitEngineDaemon cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,transmitEngineDaemon_CP_3152_symbol, "transmitEngineDaemon cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitEngineDaemon_CP_3152: Block -- control-path 
    signal transmitEngineDaemon_CP_3152_elements: BooleanArray(42 downto 0);
    -- 
  begin -- 
    transmitEngineDaemon_CP_3152_elements(0) <= transmitEngineDaemon_CP_3152_start;
    transmitEngineDaemon_CP_3152_symbol <= transmitEngineDaemon_CP_3152_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_sample_start_
      -- CP-element group 0: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Sample/req
      -- CP-element group 0: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1494/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(0), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Update/req
      -- CP-element group 1: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_update_start_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_0, ack => transmitEngineDaemon_CP_3152_elements(1)); -- 
    req_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(1), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	42 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1495/$entry
      -- CP-element group 2: 	 assign_stmt_1494/WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_Update/ack
      -- CP-element group 2: 	 assign_stmt_1494/$exit
      -- CP-element group 2: 	 branch_block_stmt_1495/merge_stmt_1496_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1495/merge_stmt_1496__entry__
      -- CP-element group 2: 	 branch_block_stmt_1495/branch_block_stmt_1495__entry__
      -- CP-element group 2: 	 branch_block_stmt_1495/merge_stmt_1496__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1495/merge_stmt_1496__entry___PhiReq/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_1, ack => transmitEngineDaemon_CP_3152_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1495/$exit
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_1495/branch_block_stmt_1495__exit__
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	41 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	42 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1495/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_1495/do_while_stmt_1504__exit__
      -- CP-element group 4: 	 branch_block_stmt_1495/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1495/disable_loopback_PhiReq/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(4) <= transmitEngineDaemon_CP_3152_elements(41);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1495/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1495/if_stmt_1497_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1495/if_stmt_1497_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1495/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1495/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(5) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:if_stmt_1497_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    if_choice_transition_3244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1497_branch_ack_1, ack => transmitEngineDaemon_CP_3152_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	42 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_1495/do_while_stmt_1504__entry__
      -- CP-element group 6: 	 branch_block_stmt_1495/if_stmt_1497__exit__
      -- CP-element group 6: 	 branch_block_stmt_1495/if_stmt_1497_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1495/if_stmt_1497_else_link/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(6) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:if_stmt_1497_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    else_choice_transition_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1497_branch_ack_0, ack => transmitEngineDaemon_CP_3152_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504__entry__
      -- CP-element group 7: 	 branch_block_stmt_1495/do_while_stmt_1504/$entry
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(7) <= transmitEngineDaemon_CP_3152_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	41 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504__exit__
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitEngineDaemon_CP_3152_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_back
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitEngineDaemon_CP_3152_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	39 
    -- CP-element group 10: 	40 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1495/do_while_stmt_1504/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_taken/$entry
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(10) <= transmitEngineDaemon_CP_3152_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	38 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_body_done
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(11) <= transmitEngineDaemon_CP_3152_elements(38);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(12) <= transmitEngineDaemon_CP_3152_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(13) <= transmitEngineDaemon_CP_3152_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	37 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/phi_stmt_1506_sample_start_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitEngineDaemon_CP_3152_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	37 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/condition_evaluated
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(15) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:do_while_stmt_1504_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_3264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(15), ack => do_while_stmt_1504_branch_req_0); -- 
    transmitEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(21) & transmitEngineDaemon_CP_3152_elements(37);
      gj_transmitEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	21 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/aggregated_phi_sample_req
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(14) & transmitEngineDaemon_CP_3152_elements(21);
      gj_transmitEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	35 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/phi_stmt_1506_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/aggregated_phi_update_req
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(14) & transmitEngineDaemon_CP_3152_elements(24) & transmitEngineDaemon_CP_3152_elements(35);
      gj_transmitEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_sample_start_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(18) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:AND_u6_u6_1515_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(18), ack => AND_u6_u6_1515_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(16) & transmitEngineDaemon_CP_3152_elements(20);
      gj_transmitEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	21 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Update/cr
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(19) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:AND_u6_u6_1515_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(19), ack => AND_u6_u6_1515_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(17) & transmitEngineDaemon_CP_3152_elements(21);
      gj_transmitEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	38 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/aggregated_phi_sample_ack
      -- CP-element group 20: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/phi_stmt_1506_sample_completed_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:AND_u6_u6_1515_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1515_inst_ack_0, ack => transmitEngineDaemon_CP_3152_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	34 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: 	19 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/phi_stmt_1506_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/AND_u6_u6_1515_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(21) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:AND_u6_u6_1515_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1515_inst_ack_1, ack => transmitEngineDaemon_CP_3152_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: 	33 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Sample/crr
      -- CP-element group 22: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_sample_start_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1520_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(22), ack => call_stmt_1520_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(21) & transmitEngineDaemon_CP_3152_elements(24) & transmitEngineDaemon_CP_3152_elements(33);
      gj_transmitEngineDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	28 
    -- CP-element group 23: 	32 
    -- CP-element group 23: 	33 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Update/ccr
      -- CP-element group 23: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_update_start_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1520_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(23), ack => call_stmt_1520_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(28) & transmitEngineDaemon_CP_3152_elements(32) & transmitEngineDaemon_CP_3152_elements(33);
      gj_transmitEngineDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Sample/cra
      -- CP-element group 24: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_sample_completed_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1520_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1520_call_ack_0, ack => transmitEngineDaemon_CP_3152_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	30 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Update/cca
      -- CP-element group 25: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1520_update_completed_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1520_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1520_call_ack_1, ack => transmitEngineDaemon_CP_3152_elements(25)); -- 
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Sample/crr
      -- CP-element group 26: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_sample_start_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1524_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(26), ack => call_stmt_1524_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(25) & transmitEngineDaemon_CP_3152_elements(28);
      gj_transmitEngineDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	32 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Update/ccr
      -- CP-element group 27: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Update/$entry
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1524_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(27), ack => call_stmt_1524_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3152_elements(32);
      gj_transmitEngineDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Sample/cra
      -- CP-element group 28: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_sample_completed_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1524_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1524_call_ack_0, ack => transmitEngineDaemon_CP_3152_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Update/cca
      -- CP-element group 29: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1524_Update/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1524_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1524_call_ack_1, ack => transmitEngineDaemon_CP_3152_elements(29)); -- 
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	29 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Sample/crr
      -- CP-element group 30: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Sample/$entry
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1536_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(30), ack => call_stmt_1536_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(25) & transmitEngineDaemon_CP_3152_elements(29) & transmitEngineDaemon_CP_3152_elements(32);
      gj_transmitEngineDaemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Update/ccr
      -- CP-element group 31: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Update/$entry
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1536_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(31), ack => call_stmt_1536_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_3152_elements(33);
      gj_transmitEngineDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	27 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Sample/cra
      -- CP-element group 32: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Sample/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1536_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1536_call_ack_0, ack => transmitEngineDaemon_CP_3152_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	38 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	23 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Update/cca
      -- CP-element group 33: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/call_stmt_1536_Update/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:call_stmt_1536_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1536_call_ack_1, ack => transmitEngineDaemon_CP_3152_elements(33)); -- 
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	21 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Sample/req
      -- CP-element group 34: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_sample_start_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(34), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(21) & transmitEngineDaemon_CP_3152_elements(36);
      gj_transmitEngineDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	17 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Update/req
      -- CP-element group 35: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_update_start_
      -- CP-element group 35: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Sample/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_0, ack => transmitEngineDaemon_CP_3152_elements(35)); -- 
    req_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(35), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_1); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_update_completed_
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(36) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_1, ack => transmitEngineDaemon_CP_3152_elements(36)); -- 
    -- CP-element group 37:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	15 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitEngineDaemon_CP_3152_elements(37) is a control-delay.
    cp_element_37_delay: control_delay_element  generic map(name => " 37_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_3152_elements(14), ack => transmitEngineDaemon_CP_3152_elements(37), clk => clk, reset =>reset);
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	20 
    -- CP-element group 38: 	33 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	11 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1495/do_while_stmt_1504/do_while_stmt_1504_loop_body/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_3152_elements(20) & transmitEngineDaemon_CP_3152_elements(33) & transmitEngineDaemon_CP_3152_elements(36);
      gj_transmitEngineDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	10 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_exit/$exit
      -- CP-element group 39: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_exit/ack
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:do_while_stmt_1504_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1504_branch_ack_0, ack => transmitEngineDaemon_CP_3152_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	10 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_taken/$exit
      -- CP-element group 40: 	 branch_block_stmt_1495/do_while_stmt_1504/loop_taken/ack
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:do_while_stmt_1504_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1504_branch_ack_1, ack => transmitEngineDaemon_CP_3152_elements(40)); -- 
    -- CP-element group 41:  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	8 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	4 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1495/do_while_stmt_1504/$exit
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    transmitEngineDaemon_CP_3152_elements(41) <= transmitEngineDaemon_CP_3152_elements(8);
    -- CP-element group 42:  merge  branch  transition  place  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: 	2 
    -- CP-element group 42: 	4 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: 	6 
    -- CP-element group 42:  members (49) 
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Sample/req
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_else_link/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_dead_link/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Update/cr
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_if_link/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/NOT_u1_u1_1501_place
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/branch_req
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Update/cr
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497__entry__
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/SplitProtocol/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Update/ack
      -- CP-element group 42: 	 branch_block_stmt_1495/merge_stmt_1496__exit__
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Update/req
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/SplitProtocol/Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/if_stmt_1497_eval_test/NOT_u1_u1_1501/BITSEL_u32_u1_1500/BITSEL_u32_u1_1500_inputs/RPIPE_CONTROL_REGISTER_1498/Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/merge_stmt_1496_PhiReqMerge
      -- CP-element group 42: 	 branch_block_stmt_1495/merge_stmt_1496_PhiAck/$entry
      -- CP-element group 42: 	 branch_block_stmt_1495/merge_stmt_1496_PhiAck/$exit
      -- CP-element group 42: 	 branch_block_stmt_1495/merge_stmt_1496_PhiAck/dummy
      -- 
    -- logger for CP element group transmitEngineDaemon_CP_3152_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitEngineDaemon_CP_3152_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:transmitEngineDaemon_CP_3152_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitEngineDaemon:CP:if_stmt_1497_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    branch_req_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_3152_elements(42), ack => if_stmt_1497_branch_req_0); -- 
    transmitEngineDaemon_CP_3152_elements(42) <= OrReduce(transmitEngineDaemon_CP_3152_elements(5) & transmitEngineDaemon_CP_3152_elements(2) & transmitEngineDaemon_CP_3152_elements(4));
    transmitEngineDaemon_do_while_stmt_1504_terminator_3353: loop_terminator -- 
      generic map (name => " transmitEngineDaemon_do_while_stmt_1504_terminator_3353", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitEngineDaemon_CP_3152_elements(11),loop_continue => transmitEngineDaemon_CP_3152_elements(40),loop_terminate => transmitEngineDaemon_CP_3152_elements(39),loop_back => transmitEngineDaemon_CP_3152_elements(9),loop_exit => transmitEngineDaemon_CP_3152_elements(8),clk => clk, reset => reset); -- 
    entry_tmerge_3265_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitEngineDaemon_CP_3152_elements(12);
        preds(1)  <= transmitEngineDaemon_CP_3152_elements(13);
        entry_tmerge_3265 : transition_merge -- 
          generic map(name => " entry_tmerge_3265")
          port map (preds => preds, symbol_out => transmitEngineDaemon_CP_3152_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1510_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_1515_wire : std_logic_vector(5 downto 0);
    signal BITSEL_u32_u1_1500_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1543_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1501_wire : std_logic_vector(0 downto 0);
    signal RPIPE_CONTROL_REGISTER_1498_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1541_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1533_wire : std_logic_vector(35 downto 0);
    signal RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1511_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1513_wire : std_logic_vector(31 downto 0);
    signal konst_1493_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1499_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1509_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1512_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1542_wire_constant : std_logic_vector(31 downto 0);
    signal pkt_pointer_1520 : std_logic_vector(31 downto 0);
    signal push_pointer_back_to_free_Q_1529 : std_logic_vector(0 downto 0);
    signal push_status_1536 : std_logic_vector(0 downto 0);
    signal transmitted_flag_1524 : std_logic_vector(0 downto 0);
    signal tx_flag_1520 : std_logic_vector(0 downto 0);
    signal tx_q_index_1506 : std_logic_vector(5 downto 0);
    signal type_cast_1514_wire : std_logic_vector(5 downto 0);
    signal type_cast_1532_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1493_wire_constant <= "000000";
    konst_1499_wire_constant <= "00000000000000000000000000000000";
    konst_1509_wire_constant <= "000001";
    konst_1512_wire_constant <= "00000000000000000000000000000001";
    konst_1542_wire_constant <= "00000000000000000000000000000000";
    type_cast_1532_wire_constant <= "1";
    -- logger for split-operator ssrc_phi_stmt_1506 flow-through 
    process(tx_q_index_1506) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:ssrc_phi_stmt_1506:flowthrough inputs: " & " AND_u6_u6_1515_wire = "& Convert_SLV_To_Hex_String(AND_u6_u6_1515_wire) & " outputs:" & " tx_q_index_1506= "  & Convert_SLV_To_Hex_String(tx_q_index_1506));
      --
    end process; 
    -- interlock ssrc_phi_stmt_1506
    process(AND_u6_u6_1515_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := AND_u6_u6_1515_wire(5 downto 0);
      tx_q_index_1506 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1514_inst flow-through 
    process(type_cast_1514_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:type_cast_1514_inst:flowthrough inputs: " & " SUB_u32_u32_1513_wire = "& Convert_SLV_To_Hex_String(SUB_u32_u32_1513_wire) & " outputs:" & " type_cast_1514_wire= "  & Convert_SLV_To_Hex_String(type_cast_1514_wire));
      --
    end process; 
    -- interlock type_cast_1514_inst
    process(SUB_u32_u32_1513_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1513_wire(5 downto 0);
      type_cast_1514_wire <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1504_branch_req_0," req0 do_while_stmt_1504_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1504_branch_ack_0," ack0 do_while_stmt_1504_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1504_branch_ack_1," ack1 do_while_stmt_1504_branch");
    do_while_stmt_1504_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1543_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1504_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1504_branch_req_0,
          ack0 => do_while_stmt_1504_branch_ack_0,
          ack1 => do_while_stmt_1504_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1497_branch_req_0," req0 if_stmt_1497_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1497_branch_ack_0," ack0 if_stmt_1497_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_1497_branch_ack_1," ack1 if_stmt_1497_branch");
    if_stmt_1497_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1501_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1497_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1497_branch_req_0,
          ack0 => if_stmt_1497_branch_ack_0,
          ack1 => if_stmt_1497_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u6_u6_1510_inst flow-through 
    process(ADD_u6_u6_1510_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:ADD_u6_u6_1510_inst:flowthrough inputs: " & " RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire = "& Convert_SLV_To_Hex_String(RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire) & " konst_1509_wire_constant = "& Convert_SLV_To_Hex_String(konst_1509_wire_constant) & " outputs:" & " ADD_u6_u6_1510_wire= "  & Convert_SLV_To_Hex_String(ADD_u6_u6_1510_wire));
      --
    end process; 
    -- binary operator ADD_u6_u6_1510_inst
    process(RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire, konst_1509_wire_constant, tmp_var);
      ADD_u6_u6_1510_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_1528_inst flow-through 
    process(push_pointer_back_to_free_Q_1529) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:AND_u1_u1_1528_inst:flowthrough inputs: " & " tx_flag_1520 = "& Convert_SLV_To_Hex_String(tx_flag_1520) & " transmitted_flag_1524 = "& Convert_SLV_To_Hex_String(transmitted_flag_1524) & " outputs:" & " push_pointer_back_to_free_Q_1529= "  & Convert_SLV_To_Hex_String(push_pointer_back_to_free_Q_1529));
      --
    end process; 
    -- binary operator AND_u1_u1_1528_inst
    process(tx_flag_1520, transmitted_flag_1524) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tx_flag_1520, transmitted_flag_1524, tmp_var);
      push_pointer_back_to_free_Q_1529 <= tmp_var; --
    end process;
    -- logger for split-operator AND_u6_u6_1515_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if AND_u6_u6_1515_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:AND_u6_u6_1515_inst:started:   inputs: " & " ADD_u6_u6_1510_wire = "& Convert_SLV_To_Hex_String(ADD_u6_u6_1510_wire) & " type_cast_1514_wire = "& Convert_SLV_To_Hex_String(type_cast_1514_wire));
          --
        end if; 
        if AND_u6_u6_1515_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:AND_u6_u6_1515_inst:finished:  outputs: " & " AND_u6_u6_1515_wire= "  & Convert_SLV_To_Hex_String(AND_u6_u6_1515_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (2) : AND_u6_u6_1515_inst 
    ApIntAnd_group_2: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1510_wire & type_cast_1514_wire;
      AND_u6_u6_1515_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1515_inst_req_0;
      AND_u6_u6_1515_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1515_inst_req_1;
      AND_u6_u6_1515_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- logger for split-operator BITSEL_u32_u1_1500_inst flow-through 
    process(BITSEL_u32_u1_1500_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:BITSEL_u32_u1_1500_inst:flowthrough inputs: " & " RPIPE_CONTROL_REGISTER_1498_wire = "& Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_1498_wire) & " konst_1499_wire_constant = "& Convert_SLV_To_Hex_String(konst_1499_wire_constant) & " outputs:" & " BITSEL_u32_u1_1500_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u32_u1_1500_wire));
      --
    end process; 
    -- binary operator BITSEL_u32_u1_1500_inst
    process(RPIPE_CONTROL_REGISTER_1498_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1498_wire, konst_1499_wire_constant, tmp_var);
      BITSEL_u32_u1_1500_wire <= tmp_var; --
    end process;
    -- logger for split-operator BITSEL_u32_u1_1543_inst flow-through 
    process(BITSEL_u32_u1_1543_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:BITSEL_u32_u1_1543_inst:flowthrough inputs: " & " RPIPE_CONTROL_REGISTER_1541_wire = "& Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_1541_wire) & " konst_1542_wire_constant = "& Convert_SLV_To_Hex_String(konst_1542_wire_constant) & " outputs:" & " BITSEL_u32_u1_1543_wire= "  & Convert_SLV_To_Hex_String(BITSEL_u32_u1_1543_wire));
      --
    end process; 
    -- binary operator BITSEL_u32_u1_1543_inst
    process(RPIPE_CONTROL_REGISTER_1541_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1541_wire, konst_1542_wire_constant, tmp_var);
      BITSEL_u32_u1_1543_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_1501_inst flow-through 
    process(NOT_u1_u1_1501_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:NOT_u1_u1_1501_inst:flowthrough inputs: " & " BITSEL_u32_u1_1500_wire = "& Convert_SLV_To_Hex_String(BITSEL_u32_u1_1500_wire) & " outputs:" & " NOT_u1_u1_1501_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_1501_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_1501_inst
    process(BITSEL_u32_u1_1500_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1500_wire, tmp_var);
      NOT_u1_u1_1501_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator SUB_u32_u32_1513_inst flow-through 
    process(SUB_u32_u32_1513_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:SUB_u32_u32_1513_inst:flowthrough inputs: " & " RPIPE_NUMBER_OF_SERVERS_1511_wire = "& Convert_SLV_To_Hex_String(RPIPE_NUMBER_OF_SERVERS_1511_wire) & " konst_1512_wire_constant = "& Convert_SLV_To_Hex_String(konst_1512_wire_constant) & " outputs:" & " SUB_u32_u32_1513_wire= "  & Convert_SLV_To_Hex_String(SUB_u32_u32_1513_wire));
      --
    end process; 
    -- binary operator SUB_u32_u32_1513_inst
    process(RPIPE_NUMBER_OF_SERVERS_1511_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1511_wire, konst_1512_wire_constant, tmp_var);
      SUB_u32_u32_1513_wire <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_CONTROL_REGISTER_1498_inst flow-through 
    process(RPIPE_CONTROL_REGISTER_1498_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:RPIPE_CONTROL_REGISTER_1498_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_CONTROL_REGISTER_1498_wire= "  & Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_1498_wire));
      --
    end process; 
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1498_wire <= CONTROL_REGISTER;
    -- logger for split-operator RPIPE_CONTROL_REGISTER_1541_inst flow-through 
    process(RPIPE_CONTROL_REGISTER_1541_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:RPIPE_CONTROL_REGISTER_1541_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_CONTROL_REGISTER_1541_wire= "  & Convert_SLV_To_Hex_String(RPIPE_CONTROL_REGISTER_1541_wire));
      --
    end process; 
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1541_wire <= CONTROL_REGISTER;
    -- logger for split-operator RPIPE_FREE_Q_1533_inst flow-through 
    process(RPIPE_FREE_Q_1533_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:RPIPE_FREE_Q_1533_inst:flowthrough inputs: " & " push_pointer_back_to_free_Q_1529 (guard)= " & Convert_SLV_To_String(push_pointer_back_to_free_Q_1529) & " outputs:" & " RPIPE_FREE_Q_1533_wire= "  & Convert_SLV_To_Hex_String(RPIPE_FREE_Q_1533_wire));
      --
    end process; 
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1533_wire <= FREE_Q;
    -- logger for split-operator RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_inst flow-through 
    process(RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire= "  & Convert_SLV_To_Hex_String(RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire));
      --
    end process; 
    -- read from input-signal LAST_READ_TX_QUEUE_INDEX
    RPIPE_LAST_READ_TX_QUEUE_INDEX_1508_wire <= LAST_READ_TX_QUEUE_INDEX;
    -- logger for split-operator RPIPE_NUMBER_OF_SERVERS_1511_inst flow-through 
    process(RPIPE_NUMBER_OF_SERVERS_1511_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:RPIPE_NUMBER_OF_SERVERS_1511_inst:flowthrough inputs: " & " no-guard, no-inputs " & " outputs:" & " RPIPE_NUMBER_OF_SERVERS_1511_wire= "  & Convert_SLV_To_Hex_String(RPIPE_NUMBER_OF_SERVERS_1511_wire));
      --
    end process; 
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_1511_wire <= NUMBER_OF_SERVERS;
    -- logger for split-operator WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst:started:   PipeWrite to LAST_READ_TX_QUEUE_INDEX inputs: " & " konst_1493_wire_constant = "& Convert_SLV_To_Hex_String(konst_1493_wire_constant));
          --
        end if; 
        if WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1492_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_1493_wire_constant;
      LAST_READ_TX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 6),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst:started:   PipeWrite to LAST_READ_TX_QUEUE_INDEX inputs: " & " tx_q_index_1506 = "& Convert_SLV_To_Hex_String(tx_q_index_1506));
          --
        end if; 
        if WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (1) : WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_1537_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= tx_q_index_1506;
      LAST_READ_TX_QUEUE_INDEX_write_1_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_1: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logger for split-operator call_stmt_1520_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1520_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:call_stmt_1520_call:started:  Call to module getTxPacketPointerFromServer inputs: " & " tx_q_index_1506 = "& Convert_SLV_To_Hex_String(tx_q_index_1506));
          --
        end if; 
        if call_stmt_1520_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:call_stmt_1520_call:finished:  outputs: " & " pkt_pointer_1520= "  & Convert_SLV_To_Hex_String(pkt_pointer_1520) & " tx_flag_1520= "  & Convert_SLV_To_Hex_String(tx_flag_1520));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1520_call 
    getTxPacketPointerFromServer_call_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1520_call_req_0;
      call_stmt_1520_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1520_call_req_1;
      call_stmt_1520_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTxPacketPointerFromServer_call_group_0_gI: SplitGuardInterface generic map(name => "getTxPacketPointerFromServer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_q_index_1506;
      pkt_pointer_1520 <= data_out(32 downto 1);
      tx_flag_1520 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 6,
        owidth => 6,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTxPacketPointerFromServer_call_reqs(0),
          ackR => getTxPacketPointerFromServer_call_acks(0),
          dataR => getTxPacketPointerFromServer_call_data(5 downto 0),
          tagR => getTxPacketPointerFromServer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTxPacketPointerFromServer_return_acks(0), -- cross-over
          ackL => getTxPacketPointerFromServer_return_reqs(0), -- cross-over
          dataL => getTxPacketPointerFromServer_return_data(32 downto 0),
          tagL => getTxPacketPointerFromServer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_1524_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1524_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:call_stmt_1524_call:started:  Call to module transmitPacket inputs: " & " tx_flag_1520 (guard)= " & Convert_SLV_To_String(tx_flag_1520) & " pkt_pointer_1520 = "& Convert_SLV_To_Hex_String(pkt_pointer_1520));
          --
        end if; 
        if call_stmt_1524_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:call_stmt_1524_call:finished:  outputs: " & " transmitted_flag_1524= "  & Convert_SLV_To_Hex_String(transmitted_flag_1524));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_1524_call 
    transmitPacket_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1524_call_req_0;
      call_stmt_1524_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1524_call_req_1;
      call_stmt_1524_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= tx_flag_1520(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      transmitPacket_call_group_1_gI: SplitGuardInterface generic map(name => "transmitPacket_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pkt_pointer_1520;
      transmitted_flag_1524 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => transmitPacket_call_reqs(0),
          ackR => transmitPacket_call_acks(0),
          dataR => transmitPacket_call_data(31 downto 0),
          tagR => transmitPacket_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => transmitPacket_return_acks(0), -- cross-over
          ackL => transmitPacket_return_reqs(0), -- cross-over
          dataL => transmitPacket_return_data(0 downto 0),
          tagL => transmitPacket_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- logger for split-operator call_stmt_1536_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1536_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:call_stmt_1536_call:started:  Call to module pushIntoQueue inputs: " & " push_pointer_back_to_free_Q_1529 (guard)= " & Convert_SLV_To_String(push_pointer_back_to_free_Q_1529) & " type_cast_1532_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1532_wire_constant) & " RPIPE_FREE_Q_1533_wire = "& Convert_SLV_To_Hex_String(RPIPE_FREE_Q_1533_wire) & " pkt_pointer_1520 = "& Convert_SLV_To_Hex_String(pkt_pointer_1520));
          --
        end if; 
        if call_stmt_1536_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitEngineDaemon:DP:call_stmt_1536_call:finished:  outputs: " & " push_status_1536= "  & Convert_SLV_To_Hex_String(push_status_1536));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (2) : call_stmt_1536_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1536_call_req_0;
      call_stmt_1536_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1536_call_req_1;
      call_stmt_1536_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_1529(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1532_wire_constant & RPIPE_FREE_Q_1533_wire & pkt_pointer_1520;
      push_status_1536 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end transmitEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity transmitPacket is -- 
  generic (tag_length : integer); 
  port ( -- 
    packet_pointer : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_call_acks : in   std_logic_vector(1 downto 0);
    accessMemory_call_data : out  std_logic_vector(219 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_return_acks : in   std_logic_vector(1 downto 0);
    accessMemory_return_data : in   std_logic_vector(127 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitPacket;
architecture transmitPacket_arch of transmitPacket is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal packet_pointer_buffer :  std_logic_vector(31 downto 0);
  signal packet_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal transmitPacket_CP_2898_start: Boolean;
  signal transmitPacket_CP_2898_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1399_call_req_0 : boolean;
  signal call_stmt_1399_call_ack_0 : boolean;
  signal call_stmt_1399_call_req_1 : boolean;
  signal call_stmt_1399_call_ack_1 : boolean;
  signal do_while_stmt_1415_branch_req_0 : boolean;
  signal phi_stmt_1417_req_1 : boolean;
  signal phi_stmt_1417_req_0 : boolean;
  signal phi_stmt_1417_ack_0 : boolean;
  signal packet_size_1409_1419_buf_req_0 : boolean;
  signal packet_size_1409_1419_buf_ack_0 : boolean;
  signal packet_size_1409_1419_buf_req_1 : boolean;
  signal packet_size_1409_1419_buf_ack_1 : boolean;
  signal ncount_down_1450_1420_buf_req_0 : boolean;
  signal ncount_down_1450_1420_buf_ack_0 : boolean;
  signal ncount_down_1450_1420_buf_req_1 : boolean;
  signal ncount_down_1450_1420_buf_ack_1 : boolean;
  signal phi_stmt_1421_req_1 : boolean;
  signal phi_stmt_1421_req_0 : boolean;
  signal phi_stmt_1421_ack_0 : boolean;
  signal ADD_u36_u36_1425_inst_req_0 : boolean;
  signal ADD_u36_u36_1425_inst_ack_0 : boolean;
  signal ADD_u36_u36_1425_inst_req_1 : boolean;
  signal ADD_u36_u36_1425_inst_ack_1 : boolean;
  signal nmem_addr_1455_1426_buf_req_0 : boolean;
  signal nmem_addr_1455_1426_buf_ack_0 : boolean;
  signal nmem_addr_1455_1426_buf_req_1 : boolean;
  signal nmem_addr_1455_1426_buf_ack_1 : boolean;
  signal call_stmt_1437_call_req_0 : boolean;
  signal call_stmt_1437_call_ack_0 : boolean;
  signal call_stmt_1437_call_req_1 : boolean;
  signal call_stmt_1437_call_ack_1 : boolean;
  signal CONCAT_u65_u73_1444_inst_req_0 : boolean;
  signal CONCAT_u65_u73_1444_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_1444_inst_req_1 : boolean;
  signal CONCAT_u65_u73_1444_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_1 : boolean;
  signal do_while_stmt_1415_branch_ack_0 : boolean;
  signal do_while_stmt_1415_branch_ack_1 : boolean;
  signal call_stmt_1472_call_req_0 : boolean;
  signal call_stmt_1472_call_ack_0 : boolean;
  signal call_stmt_1472_call_req_1 : boolean;
  signal call_stmt_1472_call_ack_1 : boolean;
  signal CONCAT_u65_u73_1479_inst_req_0 : boolean;
  signal CONCAT_u65_u73_1479_inst_ack_0 : boolean;
  signal CONCAT_u65_u73_1479_inst_req_1 : boolean;
  signal CONCAT_u65_u73_1479_inst_ack_1 : boolean;
  signal EQ_u12_u1_1487_inst_req_0 : boolean;
  signal EQ_u12_u1_1487_inst_ack_0 : boolean;
  signal EQ_u12_u1_1487_inst_req_1 : boolean;
  signal EQ_u12_u1_1487_inst_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitPacket_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= packet_pointer;
  packet_pointer_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitPacket_CP_2898_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitPacket_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_2898_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitPacket_CP_2898_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_2898_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,transmitPacket_CP_2898_start,"transmitPacket cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,transmitPacket_CP_2898_symbol, "transmitPacket cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitPacket_CP_2898: Block -- control-path 
    signal transmitPacket_CP_2898_elements: BooleanArray(77 downto 0);
    -- 
  begin -- 
    transmitPacket_CP_2898_elements(0) <= transmitPacket_CP_2898_start;
    transmitPacket_CP_2898_symbol <= transmitPacket_CP_2898_elements(77);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1389_to_assign_stmt_1413/$entry
      -- CP-element group 0: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_sample_start_
      -- CP-element group 0: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_update_start_
      -- CP-element group 0: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Update/ccr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1399_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1399_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    ccr_2916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(0), ack => call_stmt_1399_call_req_1); -- 
    crr_2911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(0), ack => call_stmt_1399_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Sample/cra
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1399_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_2912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1399_call_ack_0, ack => transmitPacket_CP_2898_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_1389_to_assign_stmt_1413/$exit
      -- CP-element group 2: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_update_completed_
      -- CP-element group 2: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1389_to_assign_stmt_1413/call_stmt_1399_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1414/$entry
      -- CP-element group 2: 	 branch_block_stmt_1414/branch_block_stmt_1414__entry__
      -- CP-element group 2: 	 branch_block_stmt_1414/do_while_stmt_1415__entry__
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1399_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_2917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1399_call_ack_1, ack => transmitPacket_CP_2898_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	70 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	74 
    -- CP-element group 3: 	75 
    -- CP-element group 3: 	76 
    -- CP-element group 3: 	71 
    -- CP-element group 3: 	72 
    -- CP-element group 3:  members (18) 
      -- CP-element group 3: 	 branch_block_stmt_1414/do_while_stmt_1415__exit__
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488__entry__
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/$entry
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Update/cr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(3) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1472_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1472_call_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1479_inst_req_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:EQ_u12_u1_1487_inst_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:EQ_u12_u1_1487_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_3117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(3), ack => call_stmt_1472_call_req_0); -- 
    ccr_3122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(3), ack => call_stmt_1472_call_req_1); -- 
    cr_3136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(3), ack => CONCAT_u65_u73_1479_inst_req_1); -- 
    rr_3145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(3), ack => EQ_u12_u1_1487_inst_req_0); -- 
    cr_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(3), ack => EQ_u12_u1_1487_inst_req_1); -- 
    transmitPacket_CP_2898_elements(3) <= transmitPacket_CP_2898_elements(70);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_1414/do_while_stmt_1415/$entry
      -- CP-element group 4: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415__entry__
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(4) <= transmitPacket_CP_2898_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	70 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415__exit__
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_back
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	68 
    -- CP-element group 7: 	69 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1414/do_while_stmt_1415/condition_done
      -- CP-element group 7: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_taken/$entry
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(7) <= transmitPacket_CP_2898_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	67 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_body_done
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(8) <= transmitPacket_CP_2898_elements(67);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	21 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(9) <= transmitPacket_CP_2898_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	42 
    -- CP-element group 10: 	23 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(10) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(10) <= transmitPacket_CP_2898_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	66 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/loop_body_start
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	20 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	66 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/condition_evaluated
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(12) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:do_while_stmt_1415_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(12), ack => do_while_stmt_1415_branch_req_0); -- 
    transmitPacket_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(20) & transmitPacket_CP_2898_elements(16) & transmitPacket_CP_2898_elements(66);
      gj_transmitPacket_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	17 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/aggregated_phi_sample_req
      -- CP-element group 13: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_sample_start__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(34) & transmitPacket_CP_2898_elements(17) & transmitPacket_CP_2898_elements(16);
      gj_transmitPacket_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	37 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	67 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	34 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_sample_completed_
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(19) & transmitPacket_CP_2898_elements(37);
      gj_transmitPacket_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	35 
    -- CP-element group 15: 	18 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	38 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/aggregated_phi_update_req
      -- CP-element group 15: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_update_start__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(35) & transmitPacket_CP_2898_elements(18);
      gj_transmitPacket_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	39 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(20) & transmitPacket_CP_2898_elements(39);
      gj_transmitPacket_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_sample_start_
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(11) & transmitPacket_CP_2898_elements(14);
      gj_transmitPacket_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_update_start_
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(11) & transmitPacket_CP_2898_elements(20);
      gj_transmitPacket_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_sample_completed__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	12 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_update_completed__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(20) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_loopback_trigger
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(21) <= transmitPacket_CP_2898_elements(9);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_loopback_sample_req_ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:phi_stmt_1417_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1417_loopback_sample_req_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1417_loopback_sample_req_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(22), ack => phi_stmt_1417_req_1); -- 
    -- Element group transmitPacket_CP_2898_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_entry_trigger
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(23) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(23) <= transmitPacket_CP_2898_elements(10);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_entry_sample_req_ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(24) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:phi_stmt_1417_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1417_entry_sample_req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1417_entry_sample_req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(24), ack => phi_stmt_1417_req_0); -- 
    -- Element group transmitPacket_CP_2898_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1417_phi_mux_ack_ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(25) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:phi_stmt_1417_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1417_phi_mux_ack_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1417_ack_0, ack => transmitPacket_CP_2898_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Sample/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:packet_size_1409_1419_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(26), ack => packet_size_1409_1419_buf_req_0); -- 
    -- Element group transmitPacket_CP_2898_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Update/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:packet_size_1409_1419_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(27), ack => packet_size_1409_1419_buf_req_1); -- 
    -- Element group transmitPacket_CP_2898_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Sample/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:packet_size_1409_1419_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => packet_size_1409_1419_buf_ack_0, ack => transmitPacket_CP_2898_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_packet_size_1419_Update/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:packet_size_1409_1419_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => packet_size_1409_1419_buf_ack_1, ack => transmitPacket_CP_2898_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Sample/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(30) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ncount_down_1450_1420_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_2993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(30), ack => ncount_down_1450_1420_buf_req_0); -- 
    -- Element group transmitPacket_CP_2898_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Update/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(31) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ncount_down_1450_1420_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(31), ack => ncount_down_1450_1420_buf_req_1); -- 
    -- Element group transmitPacket_CP_2898_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Sample/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ncount_down_1450_1420_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_2994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1450_1420_buf_ack_0, ack => transmitPacket_CP_2898_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_ncount_down_1420_Update/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ncount_down_1450_1420_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_1450_1420_buf_ack_1, ack => transmitPacket_CP_2898_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	14 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	13 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_sample_start_
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(34) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(11) & transmitPacket_CP_2898_elements(14);
      gj_transmitPacket_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	57 
    -- CP-element group 35: 	39 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	15 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_update_start_
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(35) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(11) & transmitPacket_CP_2898_elements(57) & transmitPacket_CP_2898_elements(39);
      gj_transmitPacket_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_sample_start__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(36) <= transmitPacket_CP_2898_elements(13);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_sample_completed__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_update_start__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(38) <= transmitPacket_CP_2898_elements(15);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39: 	16 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	35 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_update_completed__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_loopback_trigger
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(40) <= transmitPacket_CP_2898_elements(9);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_loopback_sample_req_ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:phi_stmt_1421_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1421_loopback_sample_req_3010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1421_loopback_sample_req_3010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(41), ack => phi_stmt_1421_req_1); -- 
    -- Element group transmitPacket_CP_2898_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	10 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_entry_trigger
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(42) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(42) <= transmitPacket_CP_2898_elements(10);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_entry_sample_req_ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:phi_stmt_1421_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1421_entry_sample_req_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1421_entry_sample_req_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(43), ack => phi_stmt_1421_req_0); -- 
    -- Element group transmitPacket_CP_2898_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/phi_stmt_1421_phi_mux_ack_ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:phi_stmt_1421_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_1421_phi_mux_ack_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1421_ack_0, ack => transmitPacket_CP_2898_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_sample_start__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_update_start__ps
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Sample/rr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ADD_u36_u36_1425_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(47), ack => ADD_u36_u36_1425_inst_req_0); -- 
    transmitPacket_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(45) & transmitPacket_CP_2898_elements(49);
      gj_transmitPacket_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Update/cr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ADD_u36_u36_1425_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(48), ack => ADD_u36_u36_1425_inst_req_1); -- 
    transmitPacket_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(46) & transmitPacket_CP_2898_elements(50);
      gj_transmitPacket_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Sample/ra
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(49) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ADD_u36_u36_1425_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1425_inst_ack_0, ack => transmitPacket_CP_2898_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/ADD_u36_u36_1425_Update/ca
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(50) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:ADD_u36_u36_1425_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1425_inst_ack_1, ack => transmitPacket_CP_2898_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_sample_start__ps
      -- CP-element group 51: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Sample/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:nmem_addr_1455_1426_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(51), ack => nmem_addr_1455_1426_buf_req_0); -- 
    -- Element group transmitPacket_CP_2898_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_update_start__ps
      -- CP-element group 52: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Update/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:nmem_addr_1455_1426_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(52), ack => nmem_addr_1455_1426_buf_req_1); -- 
    -- Element group transmitPacket_CP_2898_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Sample/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:nmem_addr_1455_1426_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1455_1426_buf_ack_0, ack => transmitPacket_CP_2898_elements(53)); -- 
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/R_nmem_addr_1426_Update/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:nmem_addr_1455_1426_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_1455_1426_buf_ack_1, ack => transmitPacket_CP_2898_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	39 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Sample/crr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(55) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1437_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(55), ack => call_stmt_1437_call_req_0); -- 
    transmitPacket_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(39) & transmitPacket_CP_2898_elements(57);
      gj_transmitPacket_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	61 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Update/ccr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1437_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(56), ack => call_stmt_1437_call_req_1); -- 
    transmitPacket_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(58) & transmitPacket_CP_2898_elements(61);
      gj_transmitPacket_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: 	35 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Sample/cra
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1437_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1437_call_ack_0, ack => transmitPacket_CP_2898_elements(57)); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/call_stmt_1437_Update/cca
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1437_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1437_call_ack_1, ack => transmitPacket_CP_2898_elements(58)); -- 
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Sample/rr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1444_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(59), ack => CONCAT_u65_u73_1444_inst_req_0); -- 
    transmitPacket_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(58) & transmitPacket_CP_2898_elements(61);
      gj_transmitPacket_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: 	64 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Update/cr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1444_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(60), ack => CONCAT_u65_u73_1444_inst_req_1); -- 
    transmitPacket_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(62) & transmitPacket_CP_2898_elements(64);
      gj_transmitPacket_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	56 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Sample/ra
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1444_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1444_inst_ack_0, ack => transmitPacket_CP_2898_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/CONCAT_u65_u73_1444_Update/ca
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1444_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1444_inst_ack_1, ack => transmitPacket_CP_2898_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Sample/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(63), ack => WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_0); -- 
    transmitPacket_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(62) & transmitPacket_CP_2898_elements(65);
      gj_transmitPacket_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	60 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_update_start_
      -- CP-element group 64: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Update/req
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(64) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_0, ack => transmitPacket_CP_2898_elements(64)); -- 
    req_3095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(64), ack => WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/WPIPE_nic_to_mac_transmit_pipe_1438_Update/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(65) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_1, ack => transmitPacket_CP_2898_elements(65)); -- 
    -- CP-element group 66:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	11 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	12 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(66) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group transmitPacket_CP_2898_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => transmitPacket_CP_2898_elements(11), ack => transmitPacket_CP_2898_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  join  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	8 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1414/do_while_stmt_1415/do_while_stmt_1415_loop_body/$exit
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(67) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(14) & transmitPacket_CP_2898_elements(65);
      gj_transmitPacket_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	7 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_exit/$exit
      -- CP-element group 68: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_exit/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(68) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:do_while_stmt_1415_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_3101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1415_branch_ack_0, ack => transmitPacket_CP_2898_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	7 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_taken/$exit
      -- CP-element group 69: 	 branch_block_stmt_1414/do_while_stmt_1415/loop_taken/ack
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(69)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(69)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(69) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:do_while_stmt_1415_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_3105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1415_branch_ack_1, ack => transmitPacket_CP_2898_elements(69)); -- 
    -- CP-element group 70:  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	5 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	3 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1414/do_while_stmt_1415/$exit
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(70)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(70)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(70) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_CP_2898_elements(70) <= transmitPacket_CP_2898_elements(5);
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	3 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Sample/cra
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(71)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(71)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(71) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1472_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_3118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1472_call_ack_0, ack => transmitPacket_CP_2898_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	3 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/call_stmt_1472_Update/cca
      -- CP-element group 72: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Sample/rr
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(72)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(72)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(72) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:call_stmt_1472_call_ack_1 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1479_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    cca_3123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1472_call_ack_1, ack => transmitPacket_CP_2898_elements(72)); -- 
    rr_3131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_2898_elements(72), ack => CONCAT_u65_u73_1479_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Sample/ra
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(73)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(73)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(73) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1479_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1479_inst_ack_0, ack => transmitPacket_CP_2898_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	3 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	77 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/CONCAT_u65_u73_1479_Update/ca
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(74)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(74)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(74) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:CONCAT_u65_u73_1479_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_1479_inst_ack_1, ack => transmitPacket_CP_2898_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	3 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Sample/ra
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(75)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(75)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(75) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:EQ_u12_u1_1487_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_3146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u12_u1_1487_inst_ack_0, ack => transmitPacket_CP_2898_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	3 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/EQ_u12_u1_1487_Update/ca
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(76)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(76)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(76) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:EQ_u12_u1_1487_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u12_u1_1487_inst_ack_1, ack => transmitPacket_CP_2898_elements(76)); -- 
    -- CP-element group 77:  join  transition  place  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 $exit
      -- CP-element group 77: 	 branch_block_stmt_1414/$exit
      -- CP-element group 77: 	 branch_block_stmt_1414/branch_block_stmt_1414__exit__
      -- CP-element group 77: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488__exit__
      -- CP-element group 77: 	 branch_block_stmt_1414/call_stmt_1472_to_assign_stmt_1488/$exit
      -- 
    -- logger for CP element group transmitPacket_CP_2898_elements(77)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and transmitPacket_CP_2898_elements(77)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:transmitPacket:CP:transmitPacket_CP_2898_elements(77) fired."); 
        -- 
      end if; --
    end process; 
    transmitPacket_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_2898_elements(74) & transmitPacket_CP_2898_elements(76);
      gj_transmitPacket_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_2898_elements(77), clk => clk, reset => reset); --
    end block;
    transmitPacket_do_while_stmt_1415_terminator_3106: loop_terminator -- 
      generic map (name => " transmitPacket_do_while_stmt_1415_terminator_3106", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitPacket_CP_2898_elements(8),loop_continue => transmitPacket_CP_2898_elements(69),loop_terminate => transmitPacket_CP_2898_elements(68),loop_back => transmitPacket_CP_2898_elements(6),loop_exit => transmitPacket_CP_2898_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_1417_phi_seq_3000_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_2898_elements(23);
      transmitPacket_CP_2898_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_2898_elements(28);
      transmitPacket_CP_2898_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_2898_elements(29);
      transmitPacket_CP_2898_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_2898_elements(21);
      transmitPacket_CP_2898_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_2898_elements(32);
      transmitPacket_CP_2898_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_2898_elements(33);
      transmitPacket_CP_2898_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1417_phi_seq_3000 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1417_phi_seq_3000") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_2898_elements(13), 
          phi_sample_ack => transmitPacket_CP_2898_elements(19), 
          phi_update_req => transmitPacket_CP_2898_elements(15), 
          phi_update_ack => transmitPacket_CP_2898_elements(20), 
          phi_mux_ack => transmitPacket_CP_2898_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1421_phi_seq_3054_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_2898_elements(42);
      transmitPacket_CP_2898_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_2898_elements(49);
      transmitPacket_CP_2898_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_2898_elements(50);
      transmitPacket_CP_2898_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_2898_elements(40);
      transmitPacket_CP_2898_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_2898_elements(53);
      transmitPacket_CP_2898_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_2898_elements(54);
      transmitPacket_CP_2898_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1421_phi_seq_3054 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1421_phi_seq_3054") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_2898_elements(36), 
          phi_sample_ack => transmitPacket_CP_2898_elements(37), 
          phi_update_req => transmitPacket_CP_2898_elements(38), 
          phi_update_ack => transmitPacket_CP_2898_elements(39), 
          phi_mux_ack => transmitPacket_CP_2898_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2942_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitPacket_CP_2898_elements(9);
        preds(1)  <= transmitPacket_CP_2898_elements(10);
        entry_tmerge_2942 : transition_merge -- 
          generic map(name => " entry_tmerge_2942")
          port map (preds => preds, symbol_out => transmitPacket_CP_2898_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1425_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u1_u65_1442_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u1_u65_1477_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u31_u34_1387_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u65_u73_1444_wire : std_logic_vector(72 downto 0);
    signal R_FULL_BYTE_MASK_1394_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1432_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1443_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_1467_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u36_u36_1485_wire : std_logic_vector(35 downto 0);
    signal control_data_1399 : std_logic_vector(63 downto 0);
    signal control_data_addr_1389 : std_logic_vector(35 downto 0);
    signal count_down_1417 : std_logic_vector(11 downto 0);
    signal data_1437 : std_logic_vector(63 downto 0);
    signal konst_1424_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1448_wire_constant : std_logic_vector(11 downto 0);
    signal konst_1453_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1458_wire_constant : std_logic_vector(11 downto 0);
    signal last_tkeep_1413 : std_logic_vector(7 downto 0);
    signal last_word_1472 : std_logic_vector(63 downto 0);
    signal mem_addr_1421 : std_logic_vector(35 downto 0);
    signal ncount_down_1450 : std_logic_vector(11 downto 0);
    signal ncount_down_1450_1420_buffered : std_logic_vector(11 downto 0);
    signal nic_to_mac_transmit_ppe_1480 : std_logic_vector(72 downto 0);
    signal nmem_addr_1455 : std_logic_vector(35 downto 0);
    signal nmem_addr_1455_1426_buffered : std_logic_vector(35 downto 0);
    signal not_last_word_1460 : std_logic_vector(0 downto 0);
    signal packet_size_1409 : std_logic_vector(11 downto 0);
    signal packet_size_1409_1419_buffered : std_logic_vector(11 downto 0);
    signal slice_1384_wire : std_logic_vector(30 downto 0);
    signal type_cast_1386_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_1391_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1393_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1397_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1429_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1431_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1435_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1440_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1464_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1466_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1470_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1475_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1486_wire : std_logic_vector(11 downto 0);
    signal unused_1404 : std_logic_vector(43 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_1394_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1432_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1443_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_1467_wire_constant <= "11111111";
    konst_1424_wire_constant <= "000000000000000000000000000000010000";
    konst_1448_wire_constant <= "000000001000";
    konst_1453_wire_constant <= "000000000000000000000000000000001000";
    konst_1458_wire_constant <= "000000001000";
    type_cast_1386_wire_constant <= "000";
    type_cast_1391_wire_constant <= "0";
    type_cast_1393_wire_constant <= "1";
    type_cast_1397_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1429_wire_constant <= "0";
    type_cast_1431_wire_constant <= "1";
    type_cast_1435_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1440_wire_constant <= "1";
    type_cast_1464_wire_constant <= "0";
    type_cast_1466_wire_constant <= "1";
    type_cast_1470_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1475_wire_constant <= "1";
    -- logger for phi phi_stmt_1417
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1417_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:transmitPacket:DP:phi_stmt_1417:input-0 packet_size_1409_1419_buffered= " & Convert_SLV_To_Hex_String(packet_size_1409_1419_buffered));
          --
        end if;
        if phi_stmt_1417_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:transmitPacket:DP:phi_stmt_1417:input-1 ncount_down_1450_1420_buffered= " & Convert_SLV_To_Hex_String(ncount_down_1450_1420_buffered));
          --
        end if;
        if phi_stmt_1417_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:transmitPacket:DP:phi_stmt_1417:sample-completed");
          --
        end if;
        if phi_stmt_1417_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:transmitPacket:DP:phi_stmt_1417:output count_down_1417= " & Convert_SLV_To_Hex_String(count_down_1417));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1417: Block -- phi operator 
      signal idata: std_logic_vector(23 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= packet_size_1409_1419_buffered & ncount_down_1450_1420_buffered;
      req <= phi_stmt_1417_req_0 & phi_stmt_1417_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1417",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 12) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1417_ack_0,
          idata => idata,
          odata => count_down_1417,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1417
    -- logger for phi phi_stmt_1421
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_1421_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:transmitPacket:DP:phi_stmt_1421:input-0 ADD_u36_u36_1425_wire= " & Convert_SLV_To_Hex_String(ADD_u36_u36_1425_wire));
          --
        end if;
        if phi_stmt_1421_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:transmitPacket:DP:phi_stmt_1421:input-1 nmem_addr_1455_1426_buffered= " & Convert_SLV_To_Hex_String(nmem_addr_1455_1426_buffered));
          --
        end if;
        if phi_stmt_1421_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:transmitPacket:DP:phi_stmt_1421:sample-completed");
          --
        end if;
        if phi_stmt_1421_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:transmitPacket:DP:phi_stmt_1421:output mem_addr_1421= " & Convert_SLV_To_Hex_String(mem_addr_1421));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_1421: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_1425_wire & nmem_addr_1455_1426_buffered;
      req <= phi_stmt_1421_req_0 & phi_stmt_1421_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1421",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1421_ack_0,
          idata => idata,
          odata => mem_addr_1421,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1421
    -- logger for split-operator slice_1384_inst flow-through 
    process(slice_1384_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:slice_1384_inst:flowthrough inputs: " & " packet_pointer_buffer = "& Convert_SLV_To_Hex_String(packet_pointer_buffer) & " outputs:" & " slice_1384_wire= "  & Convert_SLV_To_Hex_String(slice_1384_wire));
      --
    end process; 
    -- flow-through slice operator slice_1384_inst
    slice_1384_wire <= packet_pointer_buffer(31 downto 1);
    -- logger for split-operator slice_1403_inst flow-through 
    process(unused_1404) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:slice_1403_inst:flowthrough inputs: " & " control_data_1399 = "& Convert_SLV_To_Hex_String(control_data_1399) & " outputs:" & " unused_1404= "  & Convert_SLV_To_Hex_String(unused_1404));
      --
    end process; 
    -- flow-through slice operator slice_1403_inst
    unused_1404 <= control_data_1399(63 downto 20);
    -- logger for split-operator slice_1408_inst flow-through 
    process(packet_size_1409) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:slice_1408_inst:flowthrough inputs: " & " control_data_1399 = "& Convert_SLV_To_Hex_String(control_data_1399) & " outputs:" & " packet_size_1409= "  & Convert_SLV_To_Hex_String(packet_size_1409));
      --
    end process; 
    -- flow-through slice operator slice_1408_inst
    packet_size_1409 <= control_data_1399(19 downto 8);
    -- logger for split-operator slice_1412_inst flow-through 
    process(last_tkeep_1413) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:slice_1412_inst:flowthrough inputs: " & " control_data_1399 = "& Convert_SLV_To_Hex_String(control_data_1399) & " outputs:" & " last_tkeep_1413= "  & Convert_SLV_To_Hex_String(last_tkeep_1413));
      --
    end process; 
    -- flow-through slice operator slice_1412_inst
    last_tkeep_1413 <= control_data_1399(7 downto 0);
    -- logger for split-operator ncount_down_1450_1420_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ncount_down_1450_1420_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:ncount_down_1450_1420_buf:started:   inputs: " & " ncount_down_1450 = "& Convert_SLV_To_Hex_String(ncount_down_1450));
          --
        end if; 
        if ncount_down_1450_1420_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:ncount_down_1450_1420_buf:finished:  outputs: " & " ncount_down_1450_1420_buffered= "  & Convert_SLV_To_Hex_String(ncount_down_1450_1420_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    ncount_down_1450_1420_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_down_1450_1420_buf_req_0;
      ncount_down_1450_1420_buf_ack_0<= wack(0);
      rreq(0) <= ncount_down_1450_1420_buf_req_1;
      ncount_down_1450_1420_buf_ack_1<= rack(0);
      ncount_down_1450_1420_buf : InterlockBuffer generic map ( -- 
        name => "ncount_down_1450_1420_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_down_1450,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_down_1450_1420_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator nmem_addr_1455_1426_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nmem_addr_1455_1426_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:nmem_addr_1455_1426_buf:started:   inputs: " & " nmem_addr_1455 = "& Convert_SLV_To_Hex_String(nmem_addr_1455));
          --
        end if; 
        if nmem_addr_1455_1426_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:nmem_addr_1455_1426_buf:finished:  outputs: " & " nmem_addr_1455_1426_buffered= "  & Convert_SLV_To_Hex_String(nmem_addr_1455_1426_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nmem_addr_1455_1426_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmem_addr_1455_1426_buf_req_0;
      nmem_addr_1455_1426_buf_ack_0<= wack(0);
      rreq(0) <= nmem_addr_1455_1426_buf_req_1;
      nmem_addr_1455_1426_buf_ack_1<= rack(0);
      nmem_addr_1455_1426_buf : InterlockBuffer generic map ( -- 
        name => "nmem_addr_1455_1426_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_1455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmem_addr_1455_1426_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator packet_size_1409_1419_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if packet_size_1409_1419_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:packet_size_1409_1419_buf:started:   inputs: " & " packet_size_1409 = "& Convert_SLV_To_Hex_String(packet_size_1409));
          --
        end if; 
        if packet_size_1409_1419_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:packet_size_1409_1419_buf:finished:  outputs: " & " packet_size_1409_1419_buffered= "  & Convert_SLV_To_Hex_String(packet_size_1409_1419_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    packet_size_1409_1419_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= packet_size_1409_1419_buf_req_0;
      packet_size_1409_1419_buf_ack_0<= wack(0);
      rreq(0) <= packet_size_1409_1419_buf_req_1;
      packet_size_1409_1419_buf_ack_1<= rack(0);
      packet_size_1409_1419_buf : InterlockBuffer generic map ( -- 
        name => "packet_size_1409_1419_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => packet_size_1409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => packet_size_1409_1419_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator type_cast_1388_inst flow-through 
    process(control_data_addr_1389) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:type_cast_1388_inst:flowthrough inputs: " & " CONCAT_u31_u34_1387_wire = "& Convert_SLV_To_Hex_String(CONCAT_u31_u34_1387_wire) & " outputs:" & " control_data_addr_1389= "  & Convert_SLV_To_Hex_String(control_data_addr_1389));
      --
    end process; 
    -- interlock type_cast_1388_inst
    process(CONCAT_u31_u34_1387_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_1387_wire(33 downto 0);
      control_data_addr_1389 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_1486_inst flow-through 
    process(type_cast_1486_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:type_cast_1486_inst:flowthrough inputs: " & " SUB_u36_u36_1485_wire = "& Convert_SLV_To_Hex_String(SUB_u36_u36_1485_wire) & " outputs:" & " type_cast_1486_wire= "  & Convert_SLV_To_Hex_String(type_cast_1486_wire));
      --
    end process; 
    -- interlock type_cast_1486_inst
    process(SUB_u36_u36_1485_wire) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 11 downto 0) := SUB_u36_u36_1485_wire(11 downto 0);
      type_cast_1486_wire <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1415_branch_req_0," req0 do_while_stmt_1415_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1415_branch_ack_0," ack0 do_while_stmt_1415_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_1415_branch_ack_1," ack1 do_while_stmt_1415_branch");
    do_while_stmt_1415_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= not_last_word_1460;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1415_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1415_branch_req_0,
          ack0 => do_while_stmt_1415_branch_ack_0,
          ack1 => do_while_stmt_1415_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u36_u36_1425_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u36_u36_1425_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:ADD_u36_u36_1425_inst:started:   inputs: " & " control_data_addr_1389 = "& Convert_SLV_To_Hex_String(control_data_addr_1389) & " konst_1424_wire_constant = "& Convert_SLV_To_Hex_String(konst_1424_wire_constant));
          --
        end if; 
        if ADD_u36_u36_1425_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:ADD_u36_u36_1425_inst:finished:  outputs: " & " ADD_u36_u36_1425_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_1425_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u36_u36_1425_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= control_data_addr_1389;
      ADD_u36_u36_1425_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1425_inst_req_0;
      ADD_u36_u36_1425_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1425_inst_req_1;
      ADD_u36_u36_1425_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000010000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator ADD_u36_u36_1454_inst flow-through 
    process(nmem_addr_1455) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:ADD_u36_u36_1454_inst:flowthrough inputs: " & " mem_addr_1421 = "& Convert_SLV_To_Hex_String(mem_addr_1421) & " konst_1453_wire_constant = "& Convert_SLV_To_Hex_String(konst_1453_wire_constant) & " outputs:" & " nmem_addr_1455= "  & Convert_SLV_To_Hex_String(nmem_addr_1455));
      --
    end process; 
    -- binary operator ADD_u36_u36_1454_inst
    process(mem_addr_1421) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mem_addr_1421, konst_1453_wire_constant, tmp_var);
      nmem_addr_1455 <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u65_1442_inst flow-through 
    process(CONCAT_u1_u65_1442_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:CONCAT_u1_u65_1442_inst:flowthrough inputs: " & " type_cast_1440_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1440_wire_constant) & " data_1437 = "& Convert_SLV_To_Hex_String(data_1437) & " outputs:" & " CONCAT_u1_u65_1442_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u65_1442_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u65_1442_inst
    process(type_cast_1440_wire_constant, data_1437) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1440_wire_constant, data_1437, tmp_var);
      CONCAT_u1_u65_1442_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u1_u65_1477_inst flow-through 
    process(CONCAT_u1_u65_1477_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:CONCAT_u1_u65_1477_inst:flowthrough inputs: " & " type_cast_1475_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1475_wire_constant) & " last_word_1472 = "& Convert_SLV_To_Hex_String(last_word_1472) & " outputs:" & " CONCAT_u1_u65_1477_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u1_u65_1477_wire));
      --
    end process; 
    -- binary operator CONCAT_u1_u65_1477_inst
    process(type_cast_1475_wire_constant, last_word_1472) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1475_wire_constant, last_word_1472, tmp_var);
      CONCAT_u1_u65_1477_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u31_u34_1387_inst flow-through 
    process(CONCAT_u31_u34_1387_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:CONCAT_u31_u34_1387_inst:flowthrough inputs: " & " slice_1384_wire = "& Convert_SLV_To_Hex_String(slice_1384_wire) & " type_cast_1386_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1386_wire_constant) & " outputs:" & " CONCAT_u31_u34_1387_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u31_u34_1387_wire));
      --
    end process; 
    -- binary operator CONCAT_u31_u34_1387_inst
    process(slice_1384_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1384_wire, type_cast_1386_wire_constant, tmp_var);
      CONCAT_u31_u34_1387_wire <= tmp_var; --
    end process;
    -- logger for split-operator CONCAT_u65_u73_1444_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u65_u73_1444_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:CONCAT_u65_u73_1444_inst:started:   inputs: " & " CONCAT_u1_u65_1442_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u65_1442_wire) & " R_FULL_BYTE_MASK_1443_wire_constant = "& Convert_SLV_To_Hex_String(R_FULL_BYTE_MASK_1443_wire_constant));
          --
        end if; 
        if CONCAT_u65_u73_1444_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:CONCAT_u65_u73_1444_inst:finished:  outputs: " & " CONCAT_u65_u73_1444_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u65_u73_1444_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (5) : CONCAT_u65_u73_1444_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_1442_wire;
      CONCAT_u65_u73_1444_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_1444_inst_req_0;
      CONCAT_u65_u73_1444_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_1444_inst_req_1;
      CONCAT_u65_u73_1444_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- logger for split-operator CONCAT_u65_u73_1479_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if CONCAT_u65_u73_1479_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:CONCAT_u65_u73_1479_inst:started:   inputs: " & " CONCAT_u1_u65_1477_wire = "& Convert_SLV_To_Hex_String(CONCAT_u1_u65_1477_wire) & " last_tkeep_1413 = "& Convert_SLV_To_Hex_String(last_tkeep_1413));
          --
        end if; 
        if CONCAT_u65_u73_1479_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:CONCAT_u65_u73_1479_inst:finished:  outputs: " & " nic_to_mac_transmit_ppe_1480= "  & Convert_SLV_To_Hex_String(nic_to_mac_transmit_ppe_1480));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (6) : CONCAT_u65_u73_1479_inst 
    ApConcat_group_6: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_1477_wire & last_tkeep_1413;
      nic_to_mac_transmit_ppe_1480 <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_1479_inst_req_0;
      CONCAT_u65_u73_1479_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_1479_inst_req_1;
      CONCAT_u65_u73_1479_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_6_gI: SplitGuardInterface generic map(name => "ApConcat_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- logger for split-operator EQ_u12_u1_1487_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if EQ_u12_u1_1487_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:EQ_u12_u1_1487_inst:started:   inputs: " & " packet_size_1409 = "& Convert_SLV_To_Hex_String(packet_size_1409) & " type_cast_1486_wire = "& Convert_SLV_To_Hex_String(type_cast_1486_wire));
          --
        end if; 
        if EQ_u12_u1_1487_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:EQ_u12_u1_1487_inst:finished:  outputs: " & " status_buffer= "  & Convert_SLV_To_Hex_String(status_buffer));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (7) : EQ_u12_u1_1487_inst 
    ApIntEq_group_7: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_1409 & type_cast_1486_wire;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u12_u1_1487_inst_req_0;
      EQ_u12_u1_1487_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u12_u1_1487_inst_req_1;
      EQ_u12_u1_1487_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_7_gI: SplitGuardInterface generic map(name => "ApIntEq_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 12,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 12, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- logger for split-operator SUB_u12_u12_1449_inst flow-through 
    process(ncount_down_1450) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:SUB_u12_u12_1449_inst:flowthrough inputs: " & " count_down_1417 = "& Convert_SLV_To_Hex_String(count_down_1417) & " konst_1448_wire_constant = "& Convert_SLV_To_Hex_String(konst_1448_wire_constant) & " outputs:" & " ncount_down_1450= "  & Convert_SLV_To_Hex_String(ncount_down_1450));
      --
    end process; 
    -- binary operator SUB_u12_u12_1449_inst
    process(count_down_1417) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_1417, konst_1448_wire_constant, tmp_var);
      ncount_down_1450 <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u36_u36_1485_inst flow-through 
    process(SUB_u36_u36_1485_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:SUB_u36_u36_1485_inst:flowthrough inputs: " & " nmem_addr_1455 = "& Convert_SLV_To_Hex_String(nmem_addr_1455) & " control_data_addr_1389 = "& Convert_SLV_To_Hex_String(control_data_addr_1389) & " outputs:" & " SUB_u36_u36_1485_wire= "  & Convert_SLV_To_Hex_String(SUB_u36_u36_1485_wire));
      --
    end process; 
    -- binary operator SUB_u36_u36_1485_inst
    process(nmem_addr_1455, control_data_addr_1389) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(nmem_addr_1455, control_data_addr_1389, tmp_var);
      SUB_u36_u36_1485_wire <= tmp_var; --
    end process;
    -- logger for split-operator UGT_u12_u1_1459_inst flow-through 
    process(not_last_word_1460) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:UGT_u12_u1_1459_inst:flowthrough inputs: " & " ncount_down_1450 = "& Convert_SLV_To_Hex_String(ncount_down_1450) & " konst_1458_wire_constant = "& Convert_SLV_To_Hex_String(konst_1458_wire_constant) & " outputs:" & " not_last_word_1460= "  & Convert_SLV_To_Hex_String(not_last_word_1460));
      --
    end process; 
    -- binary operator UGT_u12_u1_1459_inst
    process(ncount_down_1450) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ncount_down_1450, konst_1458_wire_constant, tmp_var);
      not_last_word_1460 <= tmp_var; --
    end process;
    -- logger for split-operator WPIPE_nic_to_mac_transmit_pipe_1438_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:WPIPE_nic_to_mac_transmit_pipe_1438_inst:started:   PipeWrite to nic_to_mac_transmit_pipe inputs: " & " CONCAT_u65_u73_1444_wire = "& Convert_SLV_To_Hex_String(CONCAT_u65_u73_1444_wire));
          --
        end if; 
        if WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:WPIPE_nic_to_mac_transmit_pipe_1438_inst:finished:  outputs: " & " no-outputs ");
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared outport operator group (0) : WPIPE_nic_to_mac_transmit_pipe_1438_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_1438_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_1438_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_1444_wire;
      nic_to_mac_transmit_pipe_write_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logger for split-operator call_stmt_1472_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1472_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:call_stmt_1472_call:started:  Call to module accessMemory inputs: " & " type_cast_1464_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1464_wire_constant) & " type_cast_1466_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1466_wire_constant) & " R_FULL_BYTE_MASK_1467_wire_constant = "& Convert_SLV_To_Hex_String(R_FULL_BYTE_MASK_1467_wire_constant) & " nmem_addr_1455 = "& Convert_SLV_To_Hex_String(nmem_addr_1455) & " type_cast_1470_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1470_wire_constant));
          --
        end if; 
        if call_stmt_1472_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:call_stmt_1472_call:finished:  outputs: " & " last_word_1472= "  & Convert_SLV_To_Hex_String(last_word_1472));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- logger for split-operator call_stmt_1399_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1399_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:call_stmt_1399_call:started:  Call to module accessMemory inputs: " & " type_cast_1391_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1391_wire_constant) & " type_cast_1393_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1393_wire_constant) & " R_FULL_BYTE_MASK_1394_wire_constant = "& Convert_SLV_To_Hex_String(R_FULL_BYTE_MASK_1394_wire_constant) & " control_data_addr_1389 = "& Convert_SLV_To_Hex_String(control_data_addr_1389) & " type_cast_1397_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1397_wire_constant));
          --
        end if; 
        if call_stmt_1399_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:call_stmt_1399_call:finished:  outputs: " & " control_data_1399= "  & Convert_SLV_To_Hex_String(control_data_1399));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_1472_call call_stmt_1399_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1472_call_req_0;
      reqL_unguarded(0) <= call_stmt_1399_call_req_0;
      call_stmt_1472_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1399_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1472_call_req_1;
      reqR_unguarded(0) <= call_stmt_1399_call_req_1;
      call_stmt_1472_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1399_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1464_wire_constant & type_cast_1466_wire_constant & R_FULL_BYTE_MASK_1467_wire_constant & nmem_addr_1455 & type_cast_1470_wire_constant & type_cast_1391_wire_constant & type_cast_1393_wire_constant & R_FULL_BYTE_MASK_1394_wire_constant & control_data_addr_1389 & type_cast_1397_wire_constant;
      last_word_1472 <= data_out(127 downto 64);
      control_data_1399 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(1),
          ackR => accessMemory_call_acks(1),
          dataR => accessMemory_call_data(219 downto 110),
          tagR => accessMemory_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(1), -- cross-over
          ackL => accessMemory_return_reqs(1), -- cross-over
          dataL => accessMemory_return_data(127 downto 64),
          tagL => accessMemory_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- logger for split-operator call_stmt_1437_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_1437_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:call_stmt_1437_call:started:  Call to module accessMemory inputs: " & " type_cast_1429_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1429_wire_constant) & " type_cast_1431_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1431_wire_constant) & " R_FULL_BYTE_MASK_1432_wire_constant = "& Convert_SLV_To_Hex_String(R_FULL_BYTE_MASK_1432_wire_constant) & " mem_addr_1421 = "& Convert_SLV_To_Hex_String(mem_addr_1421) & " type_cast_1435_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_1435_wire_constant));
          --
        end if; 
        if call_stmt_1437_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:transmitPacket:DP:call_stmt_1437_call:finished:  outputs: " & " data_1437= "  & Convert_SLV_To_Hex_String(data_1437));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (1) : call_stmt_1437_call 
    accessMemory_call_group_1: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1437_call_req_0;
      call_stmt_1437_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1437_call_req_1;
      call_stmt_1437_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1429_wire_constant & type_cast_1431_wire_constant & R_FULL_BYTE_MASK_1432_wire_constant & mem_addr_1421 & type_cast_1435_wire_constant;
      data_1437 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end transmitPacket_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity writeControlInformationToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buffer_pointer : in  std_logic_vector(35 downto 0);
    packet_size : in  std_logic_vector(7 downto 0);
    last_keep : in  std_logic_vector(7 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeControlInformationToMem;
architecture writeControlInformationToMem_arch of writeControlInformationToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 52)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buffer_pointer_update_enable: Boolean;
  signal packet_size_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  -- output port buffer signals
  signal writeControlInformationToMem_CP_905_start: Boolean;
  signal writeControlInformationToMem_CP_905_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_654_call_ack_1 : boolean;
  signal call_stmt_654_call_req_1 : boolean;
  signal call_stmt_654_call_ack_0 : boolean;
  signal call_stmt_654_call_req_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeControlInformationToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 52) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buffer_pointer;
  base_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(43 downto 36) <= packet_size;
  packet_size_buffer <= in_buffer_data_out(43 downto 36);
  in_buffer_data_in(51 downto 44) <= last_keep;
  last_keep_buffer <= in_buffer_data_out(51 downto 44);
  in_buffer_data_in(tag_length + 51 downto 52) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 51 downto 52);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeControlInformationToMem_CP_905_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeControlInformationToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_905_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_905_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_905_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,writeControlInformationToMem_CP_905_start,"writeControlInformationToMem cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,writeControlInformationToMem_CP_905_symbol, "writeControlInformationToMem cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeControlInformationToMem_CP_905: Block -- control-path 
    signal writeControlInformationToMem_CP_905_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeControlInformationToMem_CP_905_elements(0) <= writeControlInformationToMem_CP_905_start;
    writeControlInformationToMem_CP_905_symbol <= writeControlInformationToMem_CP_905_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Update/ccr
      -- CP-element group 0: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Update/$entry
      -- CP-element group 0: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_update_start_
      -- CP-element group 0: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Sample/crr
      -- CP-element group 0: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_sample_start_
      -- CP-element group 0: 	 assign_stmt_645_to_call_stmt_654/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group writeControlInformationToMem_CP_905_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeControlInformationToMem_CP_905_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeControlInformationToMem:CP:writeControlInformationToMem_CP_905_elements(0) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeControlInformationToMem:CP:call_stmt_654_call_req_0 fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeControlInformationToMem:CP:call_stmt_654_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    crr_918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_905_elements(0), ack => call_stmt_654_call_req_0); -- 
    ccr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_905_elements(0), ack => call_stmt_654_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_sample_completed_
      -- CP-element group 1: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Sample/cra
      -- 
    -- logger for CP element group writeControlInformationToMem_CP_905_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeControlInformationToMem_CP_905_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeControlInformationToMem:CP:writeControlInformationToMem_CP_905_elements(1) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeControlInformationToMem:CP:call_stmt_654_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_654_call_ack_0, ack => writeControlInformationToMem_CP_905_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Update/cca
      -- CP-element group 2: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_update_completed_
      -- CP-element group 2: 	 assign_stmt_645_to_call_stmt_654/call_stmt_654_Update/$exit
      -- CP-element group 2: 	 assign_stmt_645_to_call_stmt_654/$exit
      -- CP-element group 2: 	 $exit
      -- 
    -- logger for CP element group writeControlInformationToMem_CP_905_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeControlInformationToMem_CP_905_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeControlInformationToMem:CP:writeControlInformationToMem_CP_905_elements(2) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeControlInformationToMem:CP:call_stmt_654_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_654_call_ack_1, ack => writeControlInformationToMem_CP_905_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_643_wire : std_logic_vector(15 downto 0);
    signal R_FULL_BYTE_MASK_650_wire_constant : std_logic_vector(7 downto 0);
    signal control_data_645 : std_logic_vector(63 downto 0);
    signal ignore_return_654 : std_logic_vector(63 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_649_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_650_wire_constant <= "11111111";
    type_cast_647_wire_constant <= "0";
    type_cast_649_wire_constant <= "0";
    -- logger for split-operator type_cast_644_inst flow-through 
    process(control_data_645) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeControlInformationToMem:DP:type_cast_644_inst:flowthrough inputs: " & " CONCAT_u8_u16_643_wire = "& Convert_SLV_To_Hex_String(CONCAT_u8_u16_643_wire) & " outputs:" & " control_data_645= "  & Convert_SLV_To_Hex_String(control_data_645));
      --
    end process; 
    -- interlock type_cast_644_inst
    process(CONCAT_u8_u16_643_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := CONCAT_u8_u16_643_wire(15 downto 0);
      control_data_645 <= tmp_var; -- 
    end process;
    -- logger for split-operator CONCAT_u8_u16_643_inst flow-through 
    process(CONCAT_u8_u16_643_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeControlInformationToMem:DP:CONCAT_u8_u16_643_inst:flowthrough inputs: " & " packet_size_buffer = "& Convert_SLV_To_Hex_String(packet_size_buffer) & " last_keep_buffer = "& Convert_SLV_To_Hex_String(last_keep_buffer) & " outputs:" & " CONCAT_u8_u16_643_wire= "  & Convert_SLV_To_Hex_String(CONCAT_u8_u16_643_wire));
      --
    end process; 
    -- binary operator CONCAT_u8_u16_643_inst
    process(packet_size_buffer, last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(packet_size_buffer, last_keep_buffer, tmp_var);
      CONCAT_u8_u16_643_wire <= tmp_var; --
    end process;
    -- logger for split-operator call_stmt_654_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_654_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeControlInformationToMem:DP:call_stmt_654_call:started:  Call to module accessMemory inputs: " & " type_cast_647_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_647_wire_constant) & " type_cast_649_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_649_wire_constant) & " R_FULL_BYTE_MASK_650_wire_constant = "& Convert_SLV_To_Hex_String(R_FULL_BYTE_MASK_650_wire_constant) & " base_buffer_pointer_buffer = "& Convert_SLV_To_Hex_String(base_buffer_pointer_buffer) & " control_data_645 = "& Convert_SLV_To_Hex_String(control_data_645));
          --
        end if; 
        if call_stmt_654_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeControlInformationToMem:DP:call_stmt_654_call:finished:  outputs: " & " ignore_return_654= "  & Convert_SLV_To_Hex_String(ignore_return_654));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_654_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_654_call_req_0;
      call_stmt_654_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_654_call_req_1;
      call_stmt_654_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_647_wire_constant & type_cast_649_wire_constant & R_FULL_BYTE_MASK_650_wire_constant & base_buffer_pointer_buffer & control_data_645;
      ignore_return_654 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeControlInformationToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity writeEthernetHeaderToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    buf_pointer : in  std_logic_vector(35 downto 0);
    buf_position : out  std_logic_vector(35 downto 0);
    nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeEthernetHeaderToMem;
architecture writeEthernetHeaderToMem_arch of writeEthernetHeaderToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal buf_position_buffer :  std_logic_vector(35 downto 0);
  signal buf_position_update_enable: Boolean;
  signal writeEthernetHeaderToMem_CP_606_start: Boolean;
  signal writeEthernetHeaderToMem_CP_606_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u36_u36_517_inst_req_0 : boolean;
  signal ADD_u36_u36_517_inst_ack_0 : boolean;
  signal ADD_u36_u36_517_inst_req_1 : boolean;
  signal do_while_stmt_511_branch_req_0 : boolean;
  signal phi_stmt_513_req_1 : boolean;
  signal phi_stmt_513_req_0 : boolean;
  signal phi_stmt_513_ack_0 : boolean;
  signal ADD_u36_u36_517_inst_ack_1 : boolean;
  signal ADD_u36_u36_520_inst_req_0 : boolean;
  signal ADD_u36_u36_520_inst_ack_0 : boolean;
  signal ADD_u36_u36_520_inst_req_1 : boolean;
  signal ADD_u36_u36_520_inst_ack_1 : boolean;
  signal phi_stmt_521_req_1 : boolean;
  signal phi_stmt_521_req_0 : boolean;
  signal phi_stmt_521_ack_0 : boolean;
  signal nI_557_525_buf_req_0 : boolean;
  signal nI_557_525_buf_ack_0 : boolean;
  signal nI_557_525_buf_req_1 : boolean;
  signal nI_557_525_buf_ack_1 : boolean;
  signal RPIPE_nic_rx_to_header_528_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_header_528_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_528_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_header_528_inst_ack_1 : boolean;
  signal call_stmt_552_call_req_0 : boolean;
  signal call_stmt_552_call_ack_0 : boolean;
  signal call_stmt_552_call_req_1 : boolean;
  signal call_stmt_552_call_ack_1 : boolean;
  signal do_while_stmt_511_branch_ack_0 : boolean;
  signal do_while_stmt_511_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeEthernetHeaderToMem_CP_606_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(35 downto 0) <= buf_position_buffer;
  buf_position <= out_buffer_data_out(35 downto 0);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_606_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_606_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_606_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,writeEthernetHeaderToMem_CP_606_start,"writeEthernetHeaderToMem cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,writeEthernetHeaderToMem_CP_606_symbol, "writeEthernetHeaderToMem cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeEthernetHeaderToMem_CP_606: Block -- control-path 
    signal writeEthernetHeaderToMem_CP_606_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    writeEthernetHeaderToMem_CP_606_elements(0) <= writeEthernetHeaderToMem_CP_606_start;
    writeEthernetHeaderToMem_CP_606_symbol <= writeEthernetHeaderToMem_CP_606_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_510/do_while_stmt_511__entry__
      -- CP-element group 0: 	 branch_block_stmt_510/branch_block_stmt_510__entry__
      -- CP-element group 0: 	 branch_block_stmt_510/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	68 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_510/do_while_stmt_511__exit__
      -- CP-element group 1: 	 branch_block_stmt_510/branch_block_stmt_510__exit__
      -- CP-element group 1: 	 branch_block_stmt_510/$exit
      -- CP-element group 1: 	 $exit
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(1) <= writeEthernetHeaderToMem_CP_606_elements(68);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_510/do_while_stmt_511/$entry
      -- CP-element group 2: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511__entry__
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(2) <= writeEthernetHeaderToMem_CP_606_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	68 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511__exit__
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_510/do_while_stmt_511/loop_back
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	66 
    -- CP-element group 5: 	67 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_510/do_while_stmt_511/condition_done
      -- CP-element group 5: 	 branch_block_stmt_510/do_while_stmt_511/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_510/do_while_stmt_511/loop_taken/$entry
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(5) <= writeEthernetHeaderToMem_CP_606_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	65 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_510/do_while_stmt_511/loop_body_done
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(6) <= writeEthernetHeaderToMem_CP_606_elements(65);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	42 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(7) <= writeEthernetHeaderToMem_CP_606_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	44 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(8) <= writeEthernetHeaderToMem_CP_606_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	64 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_526_sample_start_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	64 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/condition_evaluated
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:do_while_stmt_511_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(10), ack => do_while_stmt_511_branch_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(64) & writeEthernetHeaderToMem_CP_606_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	38 
    -- CP-element group 11: 	56 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_sample_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(15) & writeEthernetHeaderToMem_CP_606_elements(36) & writeEthernetHeaderToMem_CP_606_elements(9) & writeEthernetHeaderToMem_CP_606_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	39 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	36 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_526_sample_completed_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(17) & writeEthernetHeaderToMem_CP_606_elements(39) & writeEthernetHeaderToMem_CP_606_elements(58);
      gj_writeEthernetHeaderToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	55 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	40 
    -- CP-element group 13: 	57 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_update_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(16) & writeEthernetHeaderToMem_CP_606_elements(37) & writeEthernetHeaderToMem_CP_606_elements(55);
      gj_writeEthernetHeaderToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	41 
    -- CP-element group 14: 	59 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(18) & writeEthernetHeaderToMem_CP_606_elements(41) & writeEthernetHeaderToMem_CP_606_elements(59);
      gj_writeEthernetHeaderToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_sample_start_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(9) & writeEthernetHeaderToMem_CP_606_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_update_start_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(9) & writeEthernetHeaderToMem_CP_606_elements(18);
      gj_writeEthernetHeaderToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_sample_completed__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_update_completed__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_loopback_trigger
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(19) <= writeEthernetHeaderToMem_CP_606_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_loopback_sample_req_ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:phi_stmt_513_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_513_loopback_sample_req_645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_513_loopback_sample_req_645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(20), ack => phi_stmt_513_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_entry_trigger
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(21) <= writeEthernetHeaderToMem_CP_606_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_entry_sample_req_ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:phi_stmt_513_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_513_entry_sample_req_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_513_entry_sample_req_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(22), ack => phi_stmt_513_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_513_phi_mux_ack_ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:phi_stmt_513_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_513_phi_mux_ack_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_513_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_sample_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_update_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Sample/rr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_517_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(26), ack => ADD_u36_u36_517_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(24) & writeEthernetHeaderToMem_CP_606_elements(28);
      gj_writeEthernetHeaderToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_update_start_
      -- CP-element group 27: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Update/cr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_517_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(27), ack => ADD_u36_u36_517_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(25) & writeEthernetHeaderToMem_CP_606_elements(29);
      gj_writeEthernetHeaderToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Sample/ra
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_517_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_517_inst_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_517_Update/ca
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_517_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_517_inst_ack_1, ack => writeEthernetHeaderToMem_CP_606_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_sample_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_update_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Sample/rr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_520_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(32), ack => ADD_u36_u36_520_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(30) & writeEthernetHeaderToMem_CP_606_elements(34);
      gj_writeEthernetHeaderToMem_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_update_start_
      -- CP-element group 33: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Update/cr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_520_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(33), ack => ADD_u36_u36_520_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(31) & writeEthernetHeaderToMem_CP_606_elements(35);
      gj_writeEthernetHeaderToMem_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Sample/ra
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_520_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_520_inst_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/ADD_u36_u36_520_Update/ca
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:ADD_u36_u36_520_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_520_inst_ack_1, ack => writeEthernetHeaderToMem_CP_606_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_sample_start_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(9) & writeEthernetHeaderToMem_CP_606_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	41 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_update_start_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(37) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(9) & writeEthernetHeaderToMem_CP_606_elements(41);
      gj_writeEthernetHeaderToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_sample_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(38) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(38) <= writeEthernetHeaderToMem_CP_606_elements(11);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	12 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_sample_completed__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(39) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	13 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_update_start__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(40) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(40) <= writeEthernetHeaderToMem_CP_606_elements(13);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	14 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	37 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_update_completed__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(41) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	7 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_loopback_trigger
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(42) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(42) <= writeEthernetHeaderToMem_CP_606_elements(7);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_loopback_sample_req_ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:phi_stmt_521_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_521_loopback_sample_req_699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_521_loopback_sample_req_699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(43), ack => phi_stmt_521_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	8 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_entry_trigger
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(44) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(44) <= writeEthernetHeaderToMem_CP_606_elements(8);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_entry_sample_req
      -- CP-element group 45: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_entry_sample_req_ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(45) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:phi_stmt_521_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_521_entry_sample_req_702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_521_entry_sample_req_702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(45), ack => phi_stmt_521_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_521_phi_mux_ack_ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(46) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:phi_stmt_521_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_521_phi_mux_ack_705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_521_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_sample_completed_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(47) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_update_start_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(48) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_update_completed__ps
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(49) <= writeEthernetHeaderToMem_CP_606_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/type_cast_524_update_completed_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(50)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(50)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(50) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_606_elements(48), ack => writeEthernetHeaderToMem_CP_606_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_sample_start__ps
      -- CP-element group 51: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Sample/req
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(51)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(51)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(51) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:nI_557_525_buf_req_0 fired."); 
        -- 
      end if; --
    end process; 
    req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(51), ack => nI_557_525_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_update_start__ps
      -- CP-element group 52: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_update_start_
      -- CP-element group 52: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Update/req
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(52)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(52)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(52) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:nI_557_525_buf_req_1 fired."); 
        -- 
      end if; --
    end process; 
    req_731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(52), ack => nI_557_525_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Sample/ack
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(53)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(53)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(53) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:nI_557_525_buf_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_557_525_buf_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(53)); -- 
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/R_nI_525_Update/ack
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(54)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(54)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(54) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:nI_557_525_buf_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_557_525_buf_ack_1, ack => writeEthernetHeaderToMem_CP_606_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	62 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	13 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_526_update_start_
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(55)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(55)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(55) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(9) & writeEthernetHeaderToMem_CP_606_elements(62);
      gj_writeEthernetHeaderToMem_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	11 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	59 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Sample/rr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(56)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(56)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(56) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:RPIPE_nic_rx_to_header_528_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(56), ack => RPIPE_nic_rx_to_header_528_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(11) & writeEthernetHeaderToMem_CP_606_elements(59);
      gj_writeEthernetHeaderToMem_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_update_start_
      -- CP-element group 57: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Update/cr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(57)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(57)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(57) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:RPIPE_nic_rx_to_header_528_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(57), ack => RPIPE_nic_rx_to_header_528_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(58) & writeEthernetHeaderToMem_CP_606_elements(13);
      gj_writeEthernetHeaderToMem_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Sample/ra
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(58)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(58)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(58) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:RPIPE_nic_rx_to_header_528_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_528_inst_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	14 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	56 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/phi_stmt_526_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/RPIPE_nic_rx_to_header_528_Update/ca
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(59)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(59)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(59) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:RPIPE_nic_rx_to_header_528_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_528_inst_ack_1, ack => writeEthernetHeaderToMem_CP_606_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Sample/crr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(60)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(60)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(60) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:call_stmt_552_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(60), ack => call_stmt_552_call_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(59) & writeEthernetHeaderToMem_CP_606_elements(62);
      gj_writeEthernetHeaderToMem_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_update_start_
      -- CP-element group 61: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Update/ccr
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(61)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(61)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(61) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:call_stmt_552_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_606_elements(61), ack => call_stmt_552_call_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_606_elements(63);
      gj_writeEthernetHeaderToMem_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	55 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Sample/cra
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(62)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(62)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(62) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:call_stmt_552_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_552_call_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/call_stmt_552_Update/cca
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(63)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(63)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(63) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:call_stmt_552_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_552_call_ack_1, ack => writeEthernetHeaderToMem_CP_606_elements(63)); -- 
    -- CP-element group 64:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	9 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	10 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(64)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(64)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(64) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writeEthernetHeaderToMem_CP_606_elements(64) is a control-delay.
    cp_element_64_delay: control_delay_element  generic map(name => " 64_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_606_elements(9), ack => writeEthernetHeaderToMem_CP_606_elements(64), clk => clk, reset =>reset);
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	12 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	6 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_510/do_while_stmt_511/do_while_stmt_511_loop_body/$exit
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(65)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(65)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(65) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_606_elements(63) & writeEthernetHeaderToMem_CP_606_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	5 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_510/do_while_stmt_511/loop_exit/$exit
      -- CP-element group 66: 	 branch_block_stmt_510/do_while_stmt_511/loop_exit/ack
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(66)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(66)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(66) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:do_while_stmt_511_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_511_branch_ack_0, ack => writeEthernetHeaderToMem_CP_606_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	5 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_510/do_while_stmt_511/loop_taken/$exit
      -- CP-element group 67: 	 branch_block_stmt_510/do_while_stmt_511/loop_taken/ack
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(67)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(67)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(67) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:do_while_stmt_511_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_511_branch_ack_1, ack => writeEthernetHeaderToMem_CP_606_elements(67)); -- 
    -- CP-element group 68:  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	3 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	1 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_510/do_while_stmt_511/$exit
      -- 
    -- logger for CP element group writeEthernetHeaderToMem_CP_606_elements(68)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writeEthernetHeaderToMem_CP_606_elements(68)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writeEthernetHeaderToMem:CP:writeEthernetHeaderToMem_CP_606_elements(68) fired."); 
        -- 
      end if; --
    end process; 
    writeEthernetHeaderToMem_CP_606_elements(68) <= writeEthernetHeaderToMem_CP_606_elements(3);
    writeEthernetHeaderToMem_do_while_stmt_511_terminator_775: loop_terminator -- 
      generic map (name => " writeEthernetHeaderToMem_do_while_stmt_511_terminator_775", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeEthernetHeaderToMem_CP_606_elements(6),loop_continue => writeEthernetHeaderToMem_CP_606_elements(67),loop_terminate => writeEthernetHeaderToMem_CP_606_elements(66),loop_back => writeEthernetHeaderToMem_CP_606_elements(4),loop_exit => writeEthernetHeaderToMem_CP_606_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_513_phi_seq_689_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_606_elements(21);
      writeEthernetHeaderToMem_CP_606_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_606_elements(28);
      writeEthernetHeaderToMem_CP_606_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_606_elements(29);
      writeEthernetHeaderToMem_CP_606_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_606_elements(19);
      writeEthernetHeaderToMem_CP_606_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_606_elements(34);
      writeEthernetHeaderToMem_CP_606_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_606_elements(35);
      writeEthernetHeaderToMem_CP_606_elements(20) <= phi_mux_reqs(1);
      phi_stmt_513_phi_seq_689 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_513_phi_seq_689") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_606_elements(11), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_606_elements(17), 
          phi_update_req => writeEthernetHeaderToMem_CP_606_elements(13), 
          phi_update_ack => writeEthernetHeaderToMem_CP_606_elements(18), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_606_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_521_phi_seq_733_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_606_elements(44);
      writeEthernetHeaderToMem_CP_606_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_606_elements(47);
      writeEthernetHeaderToMem_CP_606_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_606_elements(49);
      writeEthernetHeaderToMem_CP_606_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_606_elements(42);
      writeEthernetHeaderToMem_CP_606_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_606_elements(53);
      writeEthernetHeaderToMem_CP_606_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_606_elements(54);
      writeEthernetHeaderToMem_CP_606_elements(43) <= phi_mux_reqs(1);
      phi_stmt_521_phi_seq_733 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_521_phi_seq_733") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_606_elements(38), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_606_elements(39), 
          phi_update_req => writeEthernetHeaderToMem_CP_606_elements(40), 
          phi_update_ack => writeEthernetHeaderToMem_CP_606_elements(41), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_606_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_631_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeEthernetHeaderToMem_CP_606_elements(7);
        preds(1)  <= writeEthernetHeaderToMem_CP_606_elements(8);
        entry_tmerge_631 : transition_merge -- 
          generic map(name => " entry_tmerge_631")
          port map (preds => preds, symbol_out => writeEthernetHeaderToMem_CP_606_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_517_wire : std_logic_vector(35 downto 0);
    signal ADD_u36_u36_520_wire : std_logic_vector(35 downto 0);
    signal I_521 : std_logic_vector(3 downto 0);
    signal RPIPE_nic_rx_to_header_528_wire : std_logic_vector(72 downto 0);
    signal ULE_u4_u1_561_wire : std_logic_vector(0 downto 0);
    signal ethernet_header_526 : std_logic_vector(72 downto 0);
    signal ignore_return_552 : std_logic_vector(63 downto 0);
    signal konst_516_wire_constant : std_logic_vector(35 downto 0);
    signal konst_519_wire_constant : std_logic_vector(35 downto 0);
    signal konst_555_wire_constant : std_logic_vector(3 downto 0);
    signal konst_560_wire_constant : std_logic_vector(3 downto 0);
    signal last_bit_535 : std_logic_vector(0 downto 0);
    signal nI_557 : std_logic_vector(3 downto 0);
    signal nI_557_525_buffered : std_logic_vector(3 downto 0);
    signal type_cast_524_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_545_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_547_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_539 : std_logic_vector(63 downto 0);
    signal wkeep_543 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_516_wire_constant <= "000000000000000000000000000000001000";
    konst_519_wire_constant <= "000000000000000000000000000000001000";
    konst_555_wire_constant <= "0001";
    konst_560_wire_constant <= "0001";
    type_cast_524_wire_constant <= "0000";
    type_cast_545_wire_constant <= "0";
    type_cast_547_wire_constant <= "0";
    -- logger for phi phi_stmt_513
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_513_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:writeEthernetHeaderToMem:DP:phi_stmt_513:input-0 ADD_u36_u36_517_wire= " & Convert_SLV_To_Hex_String(ADD_u36_u36_517_wire));
          --
        end if;
        if phi_stmt_513_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:writeEthernetHeaderToMem:DP:phi_stmt_513:input-1 ADD_u36_u36_520_wire= " & Convert_SLV_To_Hex_String(ADD_u36_u36_520_wire));
          --
        end if;
        if phi_stmt_513_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:writeEthernetHeaderToMem:DP:phi_stmt_513:sample-completed");
          --
        end if;
        if phi_stmt_513_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:writeEthernetHeaderToMem:DP:phi_stmt_513:output buf_position_buffer= " & Convert_SLV_To_Hex_String(buf_position_buffer));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_513: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_517_wire & ADD_u36_u36_520_wire;
      req <= phi_stmt_513_req_0 & phi_stmt_513_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_513",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_513_ack_0,
          idata => idata,
          odata => buf_position_buffer,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_513
    -- logger for phi phi_stmt_521
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_521_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:writeEthernetHeaderToMem:DP:phi_stmt_521:input-0 type_cast_524_wire_constant= " & Convert_SLV_To_Hex_String(type_cast_524_wire_constant));
          --
        end if;
        if phi_stmt_521_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:writeEthernetHeaderToMem:DP:phi_stmt_521:input-1 nI_557_525_buffered= " & Convert_SLV_To_Hex_String(nI_557_525_buffered));
          --
        end if;
        if phi_stmt_521_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:writeEthernetHeaderToMem:DP:phi_stmt_521:sample-completed");
          --
        end if;
        if phi_stmt_521_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:writeEthernetHeaderToMem:DP:phi_stmt_521:output I_521= " & Convert_SLV_To_Hex_String(I_521));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_521: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_524_wire_constant & nI_557_525_buffered;
      req <= phi_stmt_521_req_0 & phi_stmt_521_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_521",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_521_ack_0,
          idata => idata,
          odata => I_521,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_521
    -- logger for split-operator slice_534_inst flow-through 
    process(last_bit_535) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:slice_534_inst:flowthrough inputs: " & " ethernet_header_526 = "& Convert_SLV_To_Hex_String(ethernet_header_526) & " outputs:" & " last_bit_535= "  & Convert_SLV_To_Hex_String(last_bit_535));
      --
    end process; 
    -- flow-through slice operator slice_534_inst
    last_bit_535 <= ethernet_header_526(72 downto 72);
    -- logger for split-operator slice_538_inst flow-through 
    process(wdata_539) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:slice_538_inst:flowthrough inputs: " & " ethernet_header_526 = "& Convert_SLV_To_Hex_String(ethernet_header_526) & " outputs:" & " wdata_539= "  & Convert_SLV_To_Hex_String(wdata_539));
      --
    end process; 
    -- flow-through slice operator slice_538_inst
    wdata_539 <= ethernet_header_526(71 downto 8);
    -- logger for split-operator slice_542_inst flow-through 
    process(wkeep_543) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:slice_542_inst:flowthrough inputs: " & " ethernet_header_526 = "& Convert_SLV_To_Hex_String(ethernet_header_526) & " outputs:" & " wkeep_543= "  & Convert_SLV_To_Hex_String(wkeep_543));
      --
    end process; 
    -- flow-through slice operator slice_542_inst
    wkeep_543 <= ethernet_header_526(7 downto 0);
    -- logger for split-operator nI_557_525_buf
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if nI_557_525_buf_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:nI_557_525_buf:started:   inputs: " & " nI_557 = "& Convert_SLV_To_Hex_String(nI_557));
          --
        end if; 
        if nI_557_525_buf_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:nI_557_525_buf:finished:  outputs: " & " nI_557_525_buffered= "  & Convert_SLV_To_Hex_String(nI_557_525_buffered));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    nI_557_525_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_557_525_buf_req_0;
      nI_557_525_buf_ack_0<= wack(0);
      rreq(0) <= nI_557_525_buf_req_1;
      nI_557_525_buf_ack_1<= rack(0);
      nI_557_525_buf : InterlockBuffer generic map ( -- 
        name => "nI_557_525_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_557,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_557_525_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- logger for split-operator ssrc_phi_stmt_526 flow-through 
    process(ethernet_header_526) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:ssrc_phi_stmt_526:flowthrough inputs: " & " RPIPE_nic_rx_to_header_528_wire = "& Convert_SLV_To_Hex_String(RPIPE_nic_rx_to_header_528_wire) & " outputs:" & " ethernet_header_526= "  & Convert_SLV_To_Hex_String(ethernet_header_526));
      --
    end process; 
    -- interlock ssrc_phi_stmt_526
    process(RPIPE_nic_rx_to_header_528_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_header_528_wire(72 downto 0);
      ethernet_header_526 <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_511_branch_req_0," req0 do_while_stmt_511_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_511_branch_ack_0," ack0 do_while_stmt_511_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_511_branch_ack_1," ack1 do_while_stmt_511_branch");
    do_while_stmt_511_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULE_u4_u1_561_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_511_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_511_branch_req_0,
          ack0 => do_while_stmt_511_branch_ack_0,
          ack1 => do_while_stmt_511_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u36_u36_517_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u36_u36_517_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:ADD_u36_u36_517_inst:started:   inputs: " & " buf_pointer_buffer = "& Convert_SLV_To_Hex_String(buf_pointer_buffer) & " konst_516_wire_constant = "& Convert_SLV_To_Hex_String(konst_516_wire_constant));
          --
        end if; 
        if ADD_u36_u36_517_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:ADD_u36_u36_517_inst:finished:  outputs: " & " ADD_u36_u36_517_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_517_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u36_u36_517_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_517_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_517_inst_req_0;
      ADD_u36_u36_517_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_517_inst_req_1;
      ADD_u36_u36_517_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator ADD_u36_u36_520_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u36_u36_520_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:ADD_u36_u36_520_inst:started:   inputs: " & " buf_position_buffer = "& Convert_SLV_To_Hex_String(buf_position_buffer) & " konst_519_wire_constant = "& Convert_SLV_To_Hex_String(konst_519_wire_constant));
          --
        end if; 
        if ADD_u36_u36_520_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:ADD_u36_u36_520_inst:finished:  outputs: " & " ADD_u36_u36_520_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_520_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : ADD_u36_u36_520_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_position_buffer;
      ADD_u36_u36_520_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_520_inst_req_0;
      ADD_u36_u36_520_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_520_inst_req_1;
      ADD_u36_u36_520_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator ADD_u4_u4_556_inst flow-through 
    process(nI_557) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:ADD_u4_u4_556_inst:flowthrough inputs: " & " I_521 = "& Convert_SLV_To_Hex_String(I_521) & " konst_555_wire_constant = "& Convert_SLV_To_Hex_String(konst_555_wire_constant) & " outputs:" & " nI_557= "  & Convert_SLV_To_Hex_String(nI_557));
      --
    end process; 
    -- binary operator ADD_u4_u4_556_inst
    process(I_521) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_521, konst_555_wire_constant, tmp_var);
      nI_557 <= tmp_var; --
    end process;
    -- logger for split-operator ULE_u4_u1_561_inst flow-through 
    process(ULE_u4_u1_561_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:ULE_u4_u1_561_inst:flowthrough inputs: " & " nI_557 = "& Convert_SLV_To_Hex_String(nI_557) & " konst_560_wire_constant = "& Convert_SLV_To_Hex_String(konst_560_wire_constant) & " outputs:" & " ULE_u4_u1_561_wire= "  & Convert_SLV_To_Hex_String(ULE_u4_u1_561_wire));
      --
    end process; 
    -- binary operator ULE_u4_u1_561_inst
    process(nI_557) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(nI_557, konst_560_wire_constant, tmp_var);
      ULE_u4_u1_561_wire <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_nic_rx_to_header_528_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_nic_rx_to_header_528_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:RPIPE_nic_rx_to_header_528_inst:started:   PipeRead from nic_rx_to_header inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_nic_rx_to_header_528_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:RPIPE_nic_rx_to_header_528_inst:finished:  outputs: " & " RPIPE_nic_rx_to_header_528_wire= "  & Convert_SLV_To_Hex_String(RPIPE_nic_rx_to_header_528_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_nic_rx_to_header_528_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_header_528_inst_req_0;
      RPIPE_nic_rx_to_header_528_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_header_528_inst_req_1;
      RPIPE_nic_rx_to_header_528_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_header_528_wire <= data_out(72 downto 0);
      nic_rx_to_header_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_header_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_header_pipe_read_req(0),
          oack => nic_rx_to_header_pipe_read_ack(0),
          odata => nic_rx_to_header_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator call_stmt_552_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_552_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:call_stmt_552_call:started:  Call to module accessMemory inputs: " & " type_cast_545_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_545_wire_constant) & " type_cast_547_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_547_wire_constant) & " wkeep_543 = "& Convert_SLV_To_Hex_String(wkeep_543) & " buf_position_buffer = "& Convert_SLV_To_Hex_String(buf_position_buffer) & " wdata_539 = "& Convert_SLV_To_Hex_String(wdata_539));
          --
        end if; 
        if call_stmt_552_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writeEthernetHeaderToMem:DP:call_stmt_552_call:finished:  outputs: " & " ignore_return_552= "  & Convert_SLV_To_Hex_String(ignore_return_552));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_552_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_552_call_req_0;
      call_stmt_552_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_552_call_req_1;
      call_stmt_552_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_545_wire_constant & type_cast_547_wire_constant & wkeep_543 & buf_position_buffer & wdata_539;
      ignore_return_552 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeEthernetHeaderToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity writePayloadToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buf_pointer : in  std_logic_vector(35 downto 0);
    buf_pointer : in  std_logic_vector(35 downto 0);
    packet_size_32 : out  std_logic_vector(7 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    last_keep : out  std_logic_vector(7 downto 0);
    nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writePayloadToMem;
architecture writePayloadToMem_arch of writePayloadToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 17)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buf_pointer_update_enable: Boolean;
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal packet_size_32_buffer :  std_logic_vector(7 downto 0);
  signal packet_size_32_update_enable: Boolean;
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  signal writePayloadToMem_CP_776_start: Boolean;
  signal writePayloadToMem_CP_776_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_571_branch_req_0 : boolean;
  signal phi_stmt_573_req_1 : boolean;
  signal phi_stmt_573_req_0 : boolean;
  signal phi_stmt_573_ack_0 : boolean;
  signal ADD_u36_u36_577_inst_req_0 : boolean;
  signal ADD_u36_u36_577_inst_ack_0 : boolean;
  signal ADD_u36_u36_577_inst_req_1 : boolean;
  signal ADD_u36_u36_577_inst_ack_1 : boolean;
  signal ADD_u36_u36_580_inst_req_0 : boolean;
  signal ADD_u36_u36_580_inst_ack_0 : boolean;
  signal ADD_u36_u36_580_inst_req_1 : boolean;
  signal ADD_u36_u36_580_inst_ack_1 : boolean;
  signal RPIPE_nic_rx_to_packet_583_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_583_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_583_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_packet_583_inst_ack_1 : boolean;
  signal call_stmt_605_call_req_0 : boolean;
  signal call_stmt_605_call_ack_0 : boolean;
  signal call_stmt_605_call_req_1 : boolean;
  signal call_stmt_605_call_ack_1 : boolean;
  signal do_while_stmt_571_branch_ack_0 : boolean;
  signal do_while_stmt_571_branch_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writePayloadToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buf_pointer;
  base_buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(71 downto 36) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(71 downto 36);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writePayloadToMem_CP_776_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writePayloadToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 17) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= packet_size_32_buffer;
  packet_size_32 <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(8 downto 8) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(8 downto 8);
  out_buffer_data_in(16 downto 9) <= last_keep_buffer;
  last_keep <= out_buffer_data_out(16 downto 9);
  out_buffer_data_in(tag_length + 16 downto 17) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 16 downto 17);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_776_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writePayloadToMem_CP_776_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_776_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  --- logging ------------------------------------------------------
  LogCPEvent(clk,reset,global_clock_cycle_count,writePayloadToMem_CP_776_start,"writePayloadToMem cp_entry_symbol ");
  LogCPEvent(clk,reset,global_clock_cycle_count,writePayloadToMem_CP_776_symbol, "writePayloadToMem cp_exit_symbol ");
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writePayloadToMem_CP_776: Block -- control-path 
    signal writePayloadToMem_CP_776_elements: BooleanArray(49 downto 0);
    -- 
  begin -- 
    writePayloadToMem_CP_776_elements(0) <= writePayloadToMem_CP_776_start;
    writePayloadToMem_CP_776_symbol <= writePayloadToMem_CP_776_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_570/$entry
      -- CP-element group 0: 	 branch_block_stmt_570/branch_block_stmt_570__entry__
      -- CP-element group 0: 	 branch_block_stmt_570/do_while_stmt_571__entry__
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(0)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(0)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(0) fired."); 
        -- 
      end if; --
    end process; 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	49 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_570/$exit
      -- CP-element group 1: 	 branch_block_stmt_570/branch_block_stmt_570__exit__
      -- CP-element group 1: 	 branch_block_stmt_570/do_while_stmt_571__exit__
      -- CP-element group 1: 	 assign_stmt_618_to_assign_stmt_634/$entry
      -- CP-element group 1: 	 assign_stmt_618_to_assign_stmt_634/$exit
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(1)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(1)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(1) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(1) <= writePayloadToMem_CP_776_elements(49);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_570/do_while_stmt_571/$entry
      -- CP-element group 2: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571__entry__
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(2)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(2)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(2) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(2) <= writePayloadToMem_CP_776_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	49 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571__exit__
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(3)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(3)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(3) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_570/do_while_stmt_571/loop_back
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(4)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(4)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(4) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	47 
    -- CP-element group 5: 	48 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_570/do_while_stmt_571/condition_done
      -- CP-element group 5: 	 branch_block_stmt_570/do_while_stmt_571/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_570/do_while_stmt_571/loop_taken/$entry
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(5)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(5)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(5) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(5) <= writePayloadToMem_CP_776_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	46 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_570/do_while_stmt_571/loop_body_done
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(6)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(6)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(6) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(6) <= writePayloadToMem_CP_776_elements(46);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/back_edge_to_loop_body
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(7)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(7)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(7) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(7) <= writePayloadToMem_CP_776_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/first_time_through_loop_body
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(8)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(8)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(8) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(8) <= writePayloadToMem_CP_776_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	45 
    -- CP-element group 9: 	36 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_581_sample_start_
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(9)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(9)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(9) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	45 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/condition_evaluated
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(10)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(10)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(10) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:do_while_stmt_571_branch_req_0 fired."); 
        -- 
      end if; --
    end process; 
    condition_evaluated_800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(10), ack => do_while_stmt_571_branch_req_0); -- 
    writePayloadToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(14) & writePayloadToMem_CP_776_elements(45);
      gj_writePayloadToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	37 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_sample_start__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(11)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(11)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(11) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(9) & writePayloadToMem_CP_776_elements(15) & writePayloadToMem_CP_776_elements(14);
      gj_writePayloadToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	39 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	46 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_581_sample_completed_
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(12)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(12)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(12) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(17) & writePayloadToMem_CP_776_elements(39);
      gj_writePayloadToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	36 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_update_start__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(13)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(13)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(13) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(16) & writePayloadToMem_CP_776_elements(36);
      gj_writePayloadToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	40 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/aggregated_phi_update_ack
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(14)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(14)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(14) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(18) & writePayloadToMem_CP_776_elements(40);
      gj_writePayloadToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_sample_start_
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(15)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(15)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(15) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(9) & writePayloadToMem_CP_776_elements(12);
      gj_writePayloadToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	43 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_update_start_
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(16)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(16)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(16) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(9) & writePayloadToMem_CP_776_elements(43);
      gj_writePayloadToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_sample_completed__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(17)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(17)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(17) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_update_completed__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(18)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(18)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(18) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_loopback_trigger
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(19)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(19)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(19) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(19) <= writePayloadToMem_CP_776_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_loopback_sample_req_ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(20)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(20)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(20) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:phi_stmt_573_req_1 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_573_loopback_sample_req_815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_573_loopback_sample_req_815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(20), ack => phi_stmt_573_req_1); -- 
    -- Element group writePayloadToMem_CP_776_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_entry_trigger
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(21)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(21)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(21) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(21) <= writePayloadToMem_CP_776_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_entry_sample_req_ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(22)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(22)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(22) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:phi_stmt_573_req_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_573_entry_sample_req_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_573_entry_sample_req_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(22), ack => phi_stmt_573_req_0); -- 
    -- Element group writePayloadToMem_CP_776_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_573_phi_mux_ack_ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(23)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(23)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(23) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:phi_stmt_573_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    phi_stmt_573_phi_mux_ack_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_573_ack_0, ack => writePayloadToMem_CP_776_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_sample_start__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(24)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(24)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(24) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_update_start__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(25)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(25)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(25) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	28 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Sample/rr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(26)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(26)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(26) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_577_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(26), ack => ADD_u36_u36_577_inst_req_0); -- 
    writePayloadToMem_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(24) & writePayloadToMem_CP_776_elements(28);
      gj_writePayloadToMem_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_update_start_
      -- CP-element group 27: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Update/cr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(27)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(27)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(27) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_577_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(27), ack => ADD_u36_u36_577_inst_req_1); -- 
    writePayloadToMem_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(25) & writePayloadToMem_CP_776_elements(29);
      gj_writePayloadToMem_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	26 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Sample/ra
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(28)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(28)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(28) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_577_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_577_inst_ack_0, ack => writePayloadToMem_CP_776_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_577_Update/ca
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(29)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(29)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(29) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_577_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_577_inst_ack_1, ack => writePayloadToMem_CP_776_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_sample_start__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(30)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(30)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(30) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_update_start__ps
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(31)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(31)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(31) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Sample/rr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(32)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(32)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(32) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_580_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(32), ack => ADD_u36_u36_580_inst_req_0); -- 
    writePayloadToMem_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(30) & writePayloadToMem_CP_776_elements(34);
      gj_writePayloadToMem_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_update_start_
      -- CP-element group 33: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Update/cr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(33)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(33)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(33) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_580_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(33), ack => ADD_u36_u36_580_inst_req_1); -- 
    writePayloadToMem_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(31) & writePayloadToMem_CP_776_elements(35);
      gj_writePayloadToMem_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Sample/ra
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(34)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(34)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(34) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_580_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_580_inst_ack_0, ack => writePayloadToMem_CP_776_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/ADD_u36_u36_580_Update/ca
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(35)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(35)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(35) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:ADD_u36_u36_580_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_580_inst_ack_1, ack => writePayloadToMem_CP_776_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	43 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	13 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_581_update_start_
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(36)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(36)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(36) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(9) & writePayloadToMem_CP_776_elements(43);
      gj_writePayloadToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	40 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Sample/rr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(37)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(37)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(37) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:RPIPE_nic_rx_to_packet_583_inst_req_0 fired."); 
        -- 
      end if; --
    end process; 
    rr_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(37), ack => RPIPE_nic_rx_to_packet_583_inst_req_0); -- 
    writePayloadToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(11) & writePayloadToMem_CP_776_elements(40);
      gj_writePayloadToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_update_start_
      -- CP-element group 38: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Update/cr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(38)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(38)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(38) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:RPIPE_nic_rx_to_packet_583_inst_req_1 fired."); 
        -- 
      end if; --
    end process; 
    cr_876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(38), ack => RPIPE_nic_rx_to_packet_583_inst_req_1); -- 
    writePayloadToMem_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(39) & writePayloadToMem_CP_776_elements(13);
      gj_writePayloadToMem_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	12 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Sample/ra
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(39)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(39)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(39) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:RPIPE_nic_rx_to_packet_583_inst_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ra_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_583_inst_ack_0, ack => writePayloadToMem_CP_776_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	14 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	37 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/phi_stmt_581_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/RPIPE_nic_rx_to_packet_583_Update/ca
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(40)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(40)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(40) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:RPIPE_nic_rx_to_packet_583_inst_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ca_877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_583_inst_ack_1, ack => writePayloadToMem_CP_776_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: 	40 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Sample/crr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(41)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(41)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(41) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:call_stmt_605_call_req_0 fired."); 
        -- 
      end if; --
    end process; 
    crr_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(41), ack => call_stmt_605_call_req_0); -- 
    writePayloadToMem_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(18) & writePayloadToMem_CP_776_elements(40) & writePayloadToMem_CP_776_elements(43);
      gj_writePayloadToMem_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_update_start_
      -- CP-element group 42: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Update/ccr
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(42)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(42)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(42) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:call_stmt_605_call_req_1 fired."); 
        -- 
      end if; --
    end process; 
    ccr_890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_776_elements(42), ack => call_stmt_605_call_req_1); -- 
    writePayloadToMem_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writePayloadToMem_CP_776_elements(44);
      gj_writePayloadToMem_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	16 
    -- CP-element group 43: 	41 
    -- CP-element group 43: 	36 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Sample/cra
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(43)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(43)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(43) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:call_stmt_605_call_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    cra_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_605_call_ack_0, ack => writePayloadToMem_CP_776_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/call_stmt_605_Update/cca
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(44)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(44)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(44) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:call_stmt_605_call_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    cca_891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_605_call_ack_1, ack => writePayloadToMem_CP_776_elements(44)); -- 
    -- CP-element group 45:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	9 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	10 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/loop_body_delay_to_condition_start
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(45)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(45)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(45) fired."); 
        -- 
      end if; --
    end process; 
    -- Element group writePayloadToMem_CP_776_elements(45) is a control-delay.
    cp_element_45_delay: control_delay_element  generic map(name => " 45_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_776_elements(9), ack => writePayloadToMem_CP_776_elements(45), clk => clk, reset =>reset);
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	12 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	6 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_570/do_while_stmt_571/do_while_stmt_571_loop_body/$exit
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(46)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(46)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(46) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_776_elements(12) & writePayloadToMem_CP_776_elements(44);
      gj_writePayloadToMem_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_776_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	5 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_570/do_while_stmt_571/loop_exit/$exit
      -- CP-element group 47: 	 branch_block_stmt_570/do_while_stmt_571/loop_exit/ack
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(47)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(47)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(47) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:do_while_stmt_571_branch_ack_0 fired."); 
        -- 
      end if; --
    end process; 
    ack_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_571_branch_ack_0, ack => writePayloadToMem_CP_776_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	5 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_570/do_while_stmt_571/loop_taken/$exit
      -- CP-element group 48: 	 branch_block_stmt_570/do_while_stmt_571/loop_taken/ack
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(48)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(48)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(48) fired."); 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:do_while_stmt_571_branch_ack_1 fired."); 
        -- 
      end if; --
    end process; 
    ack_900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_571_branch_ack_1, ack => writePayloadToMem_CP_776_elements(48)); -- 
    -- CP-element group 49:  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	3 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	1 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_570/do_while_stmt_571/$exit
      -- 
    -- logger for CP element group writePayloadToMem_CP_776_elements(49)
    process (clk) 
    begin --
      if (clk'event and (clk = '1') and (reset = '0') and writePayloadToMem_CP_776_elements(49)) then -- 
        LogRecordPrint(global_clock_cycle_count,  " logger:writePayloadToMem:CP:writePayloadToMem_CP_776_elements(49) fired."); 
        -- 
      end if; --
    end process; 
    writePayloadToMem_CP_776_elements(49) <= writePayloadToMem_CP_776_elements(3);
    writePayloadToMem_do_while_stmt_571_terminator_901: loop_terminator -- 
      generic map (name => " writePayloadToMem_do_while_stmt_571_terminator_901", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writePayloadToMem_CP_776_elements(6),loop_continue => writePayloadToMem_CP_776_elements(48),loop_terminate => writePayloadToMem_CP_776_elements(47),loop_back => writePayloadToMem_CP_776_elements(4),loop_exit => writePayloadToMem_CP_776_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_573_phi_seq_859_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writePayloadToMem_CP_776_elements(21);
      writePayloadToMem_CP_776_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writePayloadToMem_CP_776_elements(28);
      writePayloadToMem_CP_776_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writePayloadToMem_CP_776_elements(29);
      writePayloadToMem_CP_776_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= writePayloadToMem_CP_776_elements(19);
      writePayloadToMem_CP_776_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writePayloadToMem_CP_776_elements(34);
      writePayloadToMem_CP_776_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= writePayloadToMem_CP_776_elements(35);
      writePayloadToMem_CP_776_elements(20) <= phi_mux_reqs(1);
      phi_stmt_573_phi_seq_859 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_573_phi_seq_859") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writePayloadToMem_CP_776_elements(11), 
          phi_sample_ack => writePayloadToMem_CP_776_elements(17), 
          phi_update_req => writePayloadToMem_CP_776_elements(13), 
          phi_update_ack => writePayloadToMem_CP_776_elements(18), 
          phi_mux_ack => writePayloadToMem_CP_776_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_801_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writePayloadToMem_CP_776_elements(7);
        preds(1)  <= writePayloadToMem_CP_776_elements(8);
        entry_tmerge_801 : transition_merge -- 
          generic map(name => " entry_tmerge_801")
          port map (preds => preds, symbol_out => writePayloadToMem_CP_776_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_577_wire : std_logic_vector(35 downto 0);
    signal ADD_u36_u36_580_wire : std_logic_vector(35 downto 0);
    signal ADD_u36_u36_624_wire : std_logic_vector(35 downto 0);
    signal EQ_u64_u1_613_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_616_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_608_wire : std_logic_vector(0 downto 0);
    signal RPIPE_nic_rx_to_packet_583_wire : std_logic_vector(72 downto 0);
    signal R_BAD_PACKET_DATA_612_wire_constant : std_logic_vector(63 downto 0);
    signal SUB_u36_u36_622_wire : std_logic_vector(35 downto 0);
    signal buf_position_573 : std_logic_vector(35 downto 0);
    signal ignore_return_605 : std_logic_vector(63 downto 0);
    signal konst_576_wire_constant : std_logic_vector(35 downto 0);
    signal konst_579_wire_constant : std_logic_vector(35 downto 0);
    signal konst_615_wire_constant : std_logic_vector(7 downto 0);
    signal konst_623_wire_constant : std_logic_vector(35 downto 0);
    signal konst_629_wire_constant : std_logic_vector(7 downto 0);
    signal last_bit_588 : std_logic_vector(0 downto 0);
    signal packet_size_8_626 : std_logic_vector(7 downto 0);
    signal payload_data_581 : std_logic_vector(72 downto 0);
    signal type_cast_598_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_600_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_592 : std_logic_vector(63 downto 0);
    signal wkeep_596 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_BAD_PACKET_DATA_612_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    konst_576_wire_constant <= "000000000000000000000000000000001000";
    konst_579_wire_constant <= "000000000000000000000000000000001000";
    konst_615_wire_constant <= "00000000";
    konst_623_wire_constant <= "000000000000000000000000000000000001";
    konst_629_wire_constant <= "00000010";
    type_cast_598_wire_constant <= "0";
    type_cast_600_wire_constant <= "0";
    -- logger for phi phi_stmt_573
    process(clk) 
    begin -- 
      if((reset = '0') and (clk'event and clk = '1')) then --
        if phi_stmt_573_req_0 then --
          LogRecordPrint(global_clock_cycle_count, "logger:writePayloadToMem:DP:phi_stmt_573:input-0 ADD_u36_u36_577_wire= " & Convert_SLV_To_Hex_String(ADD_u36_u36_577_wire));
          --
        end if;
        if phi_stmt_573_req_1 then --
          LogRecordPrint(global_clock_cycle_count, "logger:writePayloadToMem:DP:phi_stmt_573:input-1 ADD_u36_u36_580_wire= " & Convert_SLV_To_Hex_String(ADD_u36_u36_580_wire));
          --
        end if;
        if phi_stmt_573_ack_0 then --
          LogRecordPrint(global_clock_cycle_count," logger:writePayloadToMem:DP:phi_stmt_573:sample-completed");
          --
        end if;
        if phi_stmt_573_ack_0 then --
          LogRecordPrint(global_clock_cycle_count,"logger:writePayloadToMem:DP:phi_stmt_573:output buf_position_573= " & Convert_SLV_To_Hex_String(buf_position_573));
          --
        end if;
        --
      end if;
      --
    end process; 
    phi_stmt_573: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_577_wire & ADD_u36_u36_580_wire;
      req <= phi_stmt_573_req_0 & phi_stmt_573_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_573",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_573_ack_0,
          idata => idata,
          odata => buf_position_573,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_573
    -- logger for split-operator slice_587_inst flow-through 
    process(last_bit_588) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:slice_587_inst:flowthrough inputs: " & " payload_data_581 = "& Convert_SLV_To_Hex_String(payload_data_581) & " outputs:" & " last_bit_588= "  & Convert_SLV_To_Hex_String(last_bit_588));
      --
    end process; 
    -- flow-through slice operator slice_587_inst
    last_bit_588 <= payload_data_581(72 downto 72);
    -- logger for split-operator slice_591_inst flow-through 
    process(wdata_592) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:slice_591_inst:flowthrough inputs: " & " payload_data_581 = "& Convert_SLV_To_Hex_String(payload_data_581) & " outputs:" & " wdata_592= "  & Convert_SLV_To_Hex_String(wdata_592));
      --
    end process; 
    -- flow-through slice operator slice_591_inst
    wdata_592 <= payload_data_581(71 downto 8);
    -- logger for split-operator slice_595_inst flow-through 
    process(wkeep_596) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:slice_595_inst:flowthrough inputs: " & " payload_data_581 = "& Convert_SLV_To_Hex_String(payload_data_581) & " outputs:" & " wkeep_596= "  & Convert_SLV_To_Hex_String(wkeep_596));
      --
    end process; 
    -- flow-through slice operator slice_595_inst
    wkeep_596 <= payload_data_581(7 downto 0);
    -- logger for split-operator W_last_keep_632_inst flow-through 
    process(last_keep_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:W_last_keep_632_inst:flowthrough inputs: " & " wkeep_596 = "& Convert_SLV_To_Hex_String(wkeep_596) & " outputs:" & " last_keep_buffer= "  & Convert_SLV_To_Hex_String(last_keep_buffer));
      --
    end process; 
    -- interlock W_last_keep_632_inst
    process(wkeep_596) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := wkeep_596(7 downto 0);
      last_keep_buffer <= tmp_var; -- 
    end process;
    -- logger for split-operator ssrc_phi_stmt_581 flow-through 
    process(payload_data_581) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:ssrc_phi_stmt_581:flowthrough inputs: " & " RPIPE_nic_rx_to_packet_583_wire = "& Convert_SLV_To_Hex_String(RPIPE_nic_rx_to_packet_583_wire) & " outputs:" & " payload_data_581= "  & Convert_SLV_To_Hex_String(payload_data_581));
      --
    end process; 
    -- interlock ssrc_phi_stmt_581
    process(RPIPE_nic_rx_to_packet_583_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_packet_583_wire(72 downto 0);
      payload_data_581 <= tmp_var; -- 
    end process;
    -- logger for split-operator type_cast_625_inst flow-through 
    process(packet_size_8_626) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:type_cast_625_inst:flowthrough inputs: " & " ADD_u36_u36_624_wire = "& Convert_SLV_To_Hex_String(ADD_u36_u36_624_wire) & " outputs:" & " packet_size_8_626= "  & Convert_SLV_To_Hex_String(packet_size_8_626));
      --
    end process; 
    -- interlock type_cast_625_inst
    process(ADD_u36_u36_624_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ADD_u36_u36_624_wire(7 downto 0);
      packet_size_8_626 <= tmp_var; -- 
    end process;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_571_branch_req_0," req0 do_while_stmt_571_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_571_branch_ack_0," ack0 do_while_stmt_571_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_571_branch_ack_1," ack1 do_while_stmt_571_branch");
    do_while_stmt_571_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_608_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_571_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_571_branch_req_0,
          ack0 => do_while_stmt_571_branch_ack_0,
          ack1 => do_while_stmt_571_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- logger for split-operator ADD_u36_u36_577_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u36_u36_577_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:ADD_u36_u36_577_inst:started:   inputs: " & " buf_pointer_buffer = "& Convert_SLV_To_Hex_String(buf_pointer_buffer) & " konst_576_wire_constant = "& Convert_SLV_To_Hex_String(konst_576_wire_constant));
          --
        end if; 
        if ADD_u36_u36_577_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:ADD_u36_u36_577_inst:finished:  outputs: " & " ADD_u36_u36_577_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_577_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (0) : ADD_u36_u36_577_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_577_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_577_inst_req_0;
      ADD_u36_u36_577_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_577_inst_req_1;
      ADD_u36_u36_577_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- logger for split-operator ADD_u36_u36_580_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if ADD_u36_u36_580_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:ADD_u36_u36_580_inst:started:   inputs: " & " buf_position_573 = "& Convert_SLV_To_Hex_String(buf_position_573) & " konst_579_wire_constant = "& Convert_SLV_To_Hex_String(konst_579_wire_constant));
          --
        end if; 
        if ADD_u36_u36_580_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:ADD_u36_u36_580_inst:finished:  outputs: " & " ADD_u36_u36_580_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_580_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared split operator group (1) : ADD_u36_u36_580_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_position_573;
      ADD_u36_u36_580_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_580_inst_req_0;
      ADD_u36_u36_580_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_580_inst_req_1;
      ADD_u36_u36_580_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- logger for split-operator ADD_u36_u36_624_inst flow-through 
    process(ADD_u36_u36_624_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:ADD_u36_u36_624_inst:flowthrough inputs: " & " SUB_u36_u36_622_wire = "& Convert_SLV_To_Hex_String(SUB_u36_u36_622_wire) & " konst_623_wire_constant = "& Convert_SLV_To_Hex_String(konst_623_wire_constant) & " outputs:" & " ADD_u36_u36_624_wire= "  & Convert_SLV_To_Hex_String(ADD_u36_u36_624_wire));
      --
    end process; 
    -- binary operator ADD_u36_u36_624_inst
    process(SUB_u36_u36_622_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(SUB_u36_u36_622_wire, konst_623_wire_constant, tmp_var);
      ADD_u36_u36_624_wire <= tmp_var; --
    end process;
    -- logger for split-operator AND_u1_u1_617_inst flow-through 
    process(bad_packet_identifier_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:AND_u1_u1_617_inst:flowthrough inputs: " & " EQ_u64_u1_613_wire = "& Convert_SLV_To_Hex_String(EQ_u64_u1_613_wire) & " EQ_u8_u1_616_wire = "& Convert_SLV_To_Hex_String(EQ_u8_u1_616_wire) & " outputs:" & " bad_packet_identifier_buffer= "  & Convert_SLV_To_Hex_String(bad_packet_identifier_buffer));
      --
    end process; 
    -- binary operator AND_u1_u1_617_inst
    process(EQ_u64_u1_613_wire, EQ_u8_u1_616_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u64_u1_613_wire, EQ_u8_u1_616_wire, tmp_var);
      bad_packet_identifier_buffer <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u64_u1_613_inst flow-through 
    process(EQ_u64_u1_613_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:EQ_u64_u1_613_inst:flowthrough inputs: " & " wdata_592 = "& Convert_SLV_To_Hex_String(wdata_592) & " R_BAD_PACKET_DATA_612_wire_constant = "& Convert_SLV_To_Hex_String(R_BAD_PACKET_DATA_612_wire_constant) & " outputs:" & " EQ_u64_u1_613_wire= "  & Convert_SLV_To_Hex_String(EQ_u64_u1_613_wire));
      --
    end process; 
    -- binary operator EQ_u64_u1_613_inst
    process(wdata_592) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wdata_592, R_BAD_PACKET_DATA_612_wire_constant, tmp_var);
      EQ_u64_u1_613_wire <= tmp_var; --
    end process;
    -- logger for split-operator EQ_u8_u1_616_inst flow-through 
    process(EQ_u8_u1_616_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:EQ_u8_u1_616_inst:flowthrough inputs: " & " wkeep_596 = "& Convert_SLV_To_Hex_String(wkeep_596) & " konst_615_wire_constant = "& Convert_SLV_To_Hex_String(konst_615_wire_constant) & " outputs:" & " EQ_u8_u1_616_wire= "  & Convert_SLV_To_Hex_String(EQ_u8_u1_616_wire));
      --
    end process; 
    -- binary operator EQ_u8_u1_616_inst
    process(wkeep_596) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wkeep_596, konst_615_wire_constant, tmp_var);
      EQ_u8_u1_616_wire <= tmp_var; --
    end process;
    -- logger for split-operator NOT_u1_u1_608_inst flow-through 
    process(NOT_u1_u1_608_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:NOT_u1_u1_608_inst:flowthrough inputs: " & " last_bit_588 = "& Convert_SLV_To_Hex_String(last_bit_588) & " outputs:" & " NOT_u1_u1_608_wire= "  & Convert_SLV_To_Hex_String(NOT_u1_u1_608_wire));
      --
    end process; 
    -- unary operator NOT_u1_u1_608_inst
    process(last_bit_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_588, tmp_var);
      NOT_u1_u1_608_wire <= tmp_var; -- 
    end process;
    -- logger for split-operator SHL_u8_u8_630_inst flow-through 
    process(packet_size_32_buffer) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:SHL_u8_u8_630_inst:flowthrough inputs: " & " packet_size_8_626 = "& Convert_SLV_To_Hex_String(packet_size_8_626) & " konst_629_wire_constant = "& Convert_SLV_To_Hex_String(konst_629_wire_constant) & " outputs:" & " packet_size_32_buffer= "  & Convert_SLV_To_Hex_String(packet_size_32_buffer));
      --
    end process; 
    -- binary operator SHL_u8_u8_630_inst
    process(packet_size_8_626) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(packet_size_8_626, konst_629_wire_constant, tmp_var);
      packet_size_32_buffer <= tmp_var; --
    end process;
    -- logger for split-operator SUB_u36_u36_622_inst flow-through 
    process(SUB_u36_u36_622_wire) -- 
      --
    begin -- 
      LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:SUB_u36_u36_622_inst:flowthrough inputs: " & " buf_position_573 = "& Convert_SLV_To_Hex_String(buf_position_573) & " base_buf_pointer_buffer = "& Convert_SLV_To_Hex_String(base_buf_pointer_buffer) & " outputs:" & " SUB_u36_u36_622_wire= "  & Convert_SLV_To_Hex_String(SUB_u36_u36_622_wire));
      --
    end process; 
    -- binary operator SUB_u36_u36_622_inst
    process(buf_position_573, base_buf_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(buf_position_573, base_buf_pointer_buffer, tmp_var);
      SUB_u36_u36_622_wire <= tmp_var; --
    end process;
    -- logger for split-operator RPIPE_nic_rx_to_packet_583_inst
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if RPIPE_nic_rx_to_packet_583_inst_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:RPIPE_nic_rx_to_packet_583_inst:started:   PipeRead from nic_rx_to_packet inputs: " & " no-guard, no-inputs ");
          --
        end if; 
        if RPIPE_nic_rx_to_packet_583_inst_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:RPIPE_nic_rx_to_packet_583_inst:finished:  outputs: " & " RPIPE_nic_rx_to_packet_583_wire= "  & Convert_SLV_To_Hex_String(RPIPE_nic_rx_to_packet_583_wire));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared inport operator group (0) : RPIPE_nic_rx_to_packet_583_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_packet_583_inst_req_0;
      RPIPE_nic_rx_to_packet_583_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_packet_583_inst_req_1;
      RPIPE_nic_rx_to_packet_583_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_packet_583_wire <= data_out(72 downto 0);
      nic_rx_to_packet_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_packet_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_packet_pipe_read_req(0),
          oack => nic_rx_to_packet_pipe_read_ack(0),
          odata => nic_rx_to_packet_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logger for split-operator call_stmt_605_call
    process(clk)  
    begin -- 
      if ((reset = '0') and (clk'event and clk = '1')) then -- 
        if call_stmt_605_call_ack_0 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:call_stmt_605_call:started:  Call to module accessMemory inputs: " & " type_cast_598_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_598_wire_constant) & " type_cast_600_wire_constant = "& Convert_SLV_To_Hex_String(type_cast_600_wire_constant) & " wkeep_596 = "& Convert_SLV_To_Hex_String(wkeep_596) & " buf_position_573 = "& Convert_SLV_To_Hex_String(buf_position_573) & " wdata_592 = "& Convert_SLV_To_Hex_String(wdata_592));
          --
        end if; 
        if call_stmt_605_call_ack_1 then -- 
          LogRecordPrint(global_clock_cycle_count,  "logger:writePayloadToMem:DP:call_stmt_605_call:finished:  outputs: " & " ignore_return_605= "  & Convert_SLV_To_Hex_String(ignore_return_605));
          --
        end if; 
        --
      end if; 
      --
    end process; 
    -- shared call operator group (0) : call_stmt_605_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_605_call_req_0;
      call_stmt_605_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_605_call_req_1;
      call_stmt_605_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_598_wire_constant & type_cast_600_wire_constant & wkeep_596 & buf_position_573 & wdata_592;
      ignore_return_605 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writePayloadToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library GhdlLink;
use GhdlLink.LogUtilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data: in std_logic_vector(32 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : in std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : out std_logic_vector(0 downto 0);
    control_word_request_pipe_0_pipe_write_data: in std_logic_vector(31 downto 0);
    control_word_request_pipe_0_pipe_write_req : in std_logic_vector(0 downto 0);
    control_word_request_pipe_0_pipe_write_ack : out std_logic_vector(0 downto 0);
    control_word_request_pipe_1_pipe_write_data: in std_logic_vector(63 downto 0);
    control_word_request_pipe_1_pipe_write_req : in std_logic_vector(0 downto 0);
    control_word_request_pipe_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    control_word_response_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    control_word_response_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    control_word_response_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_0_pipe_write_data: in std_logic_vector(63 downto 0);
    mac_to_nic_data_0_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_0_pipe_write_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_1_pipe_write_data: in std_logic_vector(15 downto 0);
    mac_to_nic_data_1_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_1_pipe_write_ack : out std_logic_vector(0 downto 0);
    mem_req0_pipe0_pipe_read_data: out std_logic_vector(63 downto 0);
    mem_req0_pipe0_pipe_read_req : in std_logic_vector(0 downto 0);
    mem_req0_pipe0_pipe_read_ack : out std_logic_vector(0 downto 0);
    mem_req0_pipe1_pipe_read_data: out std_logic_vector(63 downto 0);
    mem_req0_pipe1_pipe_read_req : in std_logic_vector(0 downto 0);
    mem_req0_pipe1_pipe_read_ack : out std_logic_vector(0 downto 0);
    mem_resp0_pipe0_pipe_write_data: in std_logic_vector(63 downto 0);
    mem_resp0_pipe0_pipe_write_req : in std_logic_vector(0 downto 0);
    mem_resp0_pipe0_pipe_write_ack : out std_logic_vector(0 downto 0);
    mem_resp0_pipe1_pipe_write_data: in std_logic_vector(7 downto 0);
    mem_resp0_pipe1_pipe_write_req : in std_logic_vector(0 downto 0);
    mem_resp0_pipe1_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(11 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(5 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module AccessRegister
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module AccessRegister
  signal AccessRegister_rwbar :  std_logic_vector(0 downto 0);
  signal AccessRegister_bmask :  std_logic_vector(3 downto 0);
  signal AccessRegister_register_index :  std_logic_vector(5 downto 0);
  signal AccessRegister_wdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_rdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_in_args    : std_logic_vector(42 downto 0);
  signal AccessRegister_out_args   : std_logic_vector(31 downto 0);
  signal AccessRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal AccessRegister_tag_out   : std_logic_vector(2 downto 0);
  signal AccessRegister_start_req : std_logic;
  signal AccessRegister_start_ack : std_logic;
  signal AccessRegister_fin_req   : std_logic;
  signal AccessRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module AccessRegister
  signal AccessRegister_call_reqs: std_logic_vector(1 downto 0);
  signal AccessRegister_call_acks: std_logic_vector(1 downto 0);
  signal AccessRegister_return_reqs: std_logic_vector(1 downto 0);
  signal AccessRegister_return_acks: std_logic_vector(1 downto 0);
  signal AccessRegister_call_data: std_logic_vector(85 downto 0);
  signal AccessRegister_call_tag: std_logic_vector(1 downto 0);
  signal AccessRegister_return_data: std_logic_vector(63 downto 0);
  signal AccessRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module NicRegisterAccessDaemon
  component NicRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module NicRegisterAccessDaemon
  signal NicRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal NicRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal NicRegisterAccessDaemon_start_req : std_logic;
  signal NicRegisterAccessDaemon_start_ack : std_logic;
  signal NicRegisterAccessDaemon_fin_req   : std_logic;
  signal NicRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module ReceiveEngineDaemon
  component ReceiveEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_call_data : out  std_logic_vector(35 downto 0);
      loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
      loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_return_data : in   std_logic_vector(0 downto 0);
      loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
      populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ReceiveEngineDaemon
  signal ReceiveEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ReceiveEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal ReceiveEngineDaemon_start_req : std_logic;
  signal ReceiveEngineDaemon_start_ack : std_logic;
  signal ReceiveEngineDaemon_fin_req   : std_logic;
  signal ReceiveEngineDaemon_fin_ack : std_logic;
  -- declarations related to module SoftwareRegisterAccessDaemon
  component SoftwareRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
      CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
      AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
      NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module SoftwareRegisterAccessDaemon
  signal SoftwareRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal SoftwareRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal SoftwareRegisterAccessDaemon_start_req : std_logic;
  signal SoftwareRegisterAccessDaemon_start_ack : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_req   : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module UpdateRegister
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module UpdateRegister
  signal UpdateRegister_bmask :  std_logic_vector(3 downto 0);
  signal UpdateRegister_rval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_wdata :  std_logic_vector(31 downto 0);
  signal UpdateRegister_index :  std_logic_vector(5 downto 0);
  signal UpdateRegister_wval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_in_args    : std_logic_vector(73 downto 0);
  signal UpdateRegister_out_args   : std_logic_vector(31 downto 0);
  signal UpdateRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal UpdateRegister_tag_out   : std_logic_vector(2 downto 0);
  signal UpdateRegister_start_req : std_logic;
  signal UpdateRegister_start_ack : std_logic;
  signal UpdateRegister_fin_req   : std_logic;
  signal UpdateRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module UpdateRegister
  signal UpdateRegister_call_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_data: std_logic_vector(147 downto 0);
  signal UpdateRegister_call_tag: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_data: std_logic_vector(63 downto 0);
  signal UpdateRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMemory
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemory
  signal accessMemory_lock :  std_logic_vector(0 downto 0);
  signal accessMemory_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemory_bmask :  std_logic_vector(7 downto 0);
  signal accessMemory_addr :  std_logic_vector(35 downto 0);
  signal accessMemory_wdata :  std_logic_vector(63 downto 0);
  signal accessMemory_rdata :  std_logic_vector(63 downto 0);
  signal accessMemory_in_args    : std_logic_vector(109 downto 0);
  signal accessMemory_out_args   : std_logic_vector(63 downto 0);
  signal accessMemory_tag_in    : std_logic_vector(5 downto 0) := (others => '0');
  signal accessMemory_tag_out   : std_logic_vector(5 downto 0);
  signal accessMemory_start_req : std_logic;
  signal accessMemory_start_ack : std_logic;
  signal accessMemory_fin_req   : std_logic;
  signal accessMemory_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemory
  signal accessMemory_call_reqs: std_logic_vector(10 downto 0);
  signal accessMemory_call_acks: std_logic_vector(10 downto 0);
  signal accessMemory_return_reqs: std_logic_vector(10 downto 0);
  signal accessMemory_return_acks: std_logic_vector(10 downto 0);
  signal accessMemory_call_data: std_logic_vector(1209 downto 0);
  signal accessMemory_call_tag: std_logic_vector(21 downto 0);
  signal accessMemory_return_data: std_logic_vector(703 downto 0);
  signal accessMemory_return_tag: std_logic_vector(21 downto 0);
  -- declarations related to module acquireMutex
  component acquireMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module acquireMutex
  signal acquireMutex_q_base_address :  std_logic_vector(35 downto 0);
  signal acquireMutex_m_ok :  std_logic_vector(0 downto 0);
  signal acquireMutex_in_args    : std_logic_vector(35 downto 0);
  signal acquireMutex_out_args   : std_logic_vector(0 downto 0);
  signal acquireMutex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal acquireMutex_tag_out   : std_logic_vector(2 downto 0);
  signal acquireMutex_start_req : std_logic;
  signal acquireMutex_start_ack : std_logic;
  signal acquireMutex_fin_req   : std_logic;
  signal acquireMutex_fin_ack : std_logic;
  -- caller side aggregated signals for module acquireMutex
  signal acquireMutex_call_reqs: std_logic_vector(1 downto 0);
  signal acquireMutex_call_acks: std_logic_vector(1 downto 0);
  signal acquireMutex_return_reqs: std_logic_vector(1 downto 0);
  signal acquireMutex_return_acks: std_logic_vector(1 downto 0);
  signal acquireMutex_call_data: std_logic_vector(71 downto 0);
  signal acquireMutex_call_tag: std_logic_vector(1 downto 0);
  signal acquireMutex_return_data: std_logic_vector(1 downto 0);
  signal acquireMutex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module delay_time
  -- declarations related to module getQueueElement
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_pointer : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueElement
  signal getQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueElement_read_pointer :  std_logic_vector(31 downto 0);
  signal getQueueElement_q_r_data :  std_logic_vector(31 downto 0);
  signal getQueueElement_in_args    : std_logic_vector(67 downto 0);
  signal getQueueElement_out_args   : std_logic_vector(31 downto 0);
  signal getQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal getQueueElement_start_req : std_logic;
  signal getQueueElement_start_ack : std_logic;
  signal getQueueElement_fin_req   : std_logic;
  signal getQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueElement
  signal getQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_call_data: std_logic_vector(67 downto 0);
  signal getQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal getQueueElement_return_data: std_logic_vector(31 downto 0);
  signal getQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module getQueuePointers
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointers
  signal getQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_in_args    : std_logic_vector(35 downto 0);
  signal getQueuePointers_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointers_start_req : std_logic;
  signal getQueuePointers_start_ack : std_logic;
  signal getQueuePointers_fin_req   : std_logic;
  signal getQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointers
  signal getQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_data: std_logic_vector(71 downto 0);
  signal getQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTxPacketPointerFromServer
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_queue_index :  std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_pkt_pointer :  std_logic_vector(31 downto 0);
  signal getTxPacketPointerFromServer_status :  std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_in_args    : std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_out_args   : std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getTxPacketPointerFromServer_tag_out   : std_logic_vector(1 downto 0);
  signal getTxPacketPointerFromServer_start_req : std_logic;
  signal getTxPacketPointerFromServer_start_ack : std_logic;
  signal getTxPacketPointerFromServer_fin_req   : std_logic;
  signal getTxPacketPointerFromServer_fin_ack : std_logic;
  -- caller side aggregated signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_call_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_data: std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_call_tag: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_data: std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module loadBuffer
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(51 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(16 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadBuffer
  signal loadBuffer_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal loadBuffer_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal loadBuffer_in_args    : std_logic_vector(35 downto 0);
  signal loadBuffer_out_args   : std_logic_vector(0 downto 0);
  signal loadBuffer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadBuffer_tag_out   : std_logic_vector(1 downto 0);
  signal loadBuffer_start_req : std_logic;
  signal loadBuffer_start_ack : std_logic;
  signal loadBuffer_fin_req   : std_logic;
  signal loadBuffer_fin_ack : std_logic;
  -- caller side aggregated signals for module loadBuffer
  signal loadBuffer_call_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_call_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_return_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_return_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_call_data: std_logic_vector(35 downto 0);
  signal loadBuffer_call_tag: std_logic_vector(0 downto 0);
  signal loadBuffer_return_data: std_logic_vector(0 downto 0);
  signal loadBuffer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module macToNicInterface
  component macToNicInterface is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_0_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_0_pipe_read_data : in   std_logic_vector(63 downto 0);
      mac_to_nic_data_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_1_pipe_read_data : in   std_logic_vector(15 downto 0);
      mac_to_nic_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_write_data : out  std_logic_vector(72 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module macToNicInterface
  signal macToNicInterface_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal macToNicInterface_tag_out   : std_logic_vector(1 downto 0);
  signal macToNicInterface_start_req : std_logic;
  signal macToNicInterface_start_ack : std_logic;
  signal macToNicInterface_fin_req   : std_logic;
  signal macToNicInterface_fin_ack : std_logic;
  -- declarations related to module memoryToNicInterface
  component memoryToNicInterface is -- 
    generic (tag_length : integer); 
    port ( -- 
      mem_resp0_pipe0_pipe_read_req : out  std_logic_vector(0 downto 0);
      mem_resp0_pipe0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mem_resp0_pipe0_pipe_read_data : in   std_logic_vector(63 downto 0);
      mem_resp0_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      mem_resp0_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mem_resp0_pipe1_pipe_read_data : in   std_logic_vector(7 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(64 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module memoryToNicInterface
  signal memoryToNicInterface_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal memoryToNicInterface_tag_out   : std_logic_vector(1 downto 0);
  signal memoryToNicInterface_start_req : std_logic;
  signal memoryToNicInterface_start_ack : std_logic;
  signal memoryToNicInterface_fin_req   : std_logic;
  signal memoryToNicInterface_fin_ack : std_logic;
  -- declarations related to module nextLSTATE
  -- declarations related to module nicRxFromMacDaemon
  component nicRxFromMacDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
      nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
      nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicRxFromMacDaemon
  signal nicRxFromMacDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicRxFromMacDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal nicRxFromMacDaemon_start_req : std_logic;
  signal nicRxFromMacDaemon_start_ack : std_logic;
  signal nicRxFromMacDaemon_fin_req   : std_logic;
  signal nicRxFromMacDaemon_fin_ack : std_logic;
  -- declarations related to module nicToMacInterface
  component nicToMacInterface is -- 
    generic (tag_length : integer); 
    port ( -- 
      nic_to_mac_transmit_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_read_data : in   std_logic_vector(72 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicToMacInterface
  signal nicToMacInterface_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicToMacInterface_tag_out   : std_logic_vector(1 downto 0);
  signal nicToMacInterface_start_req : std_logic;
  signal nicToMacInterface_start_ack : std_logic;
  signal nicToMacInterface_fin_req   : std_logic;
  signal nicToMacInterface_fin_ack : std_logic;
  -- declarations related to module nicToMemoryInterface
  component nicToMemoryInterface is -- 
    generic (tag_length : integer); 
    port ( -- 
      NIC_TO_MEMORY_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_read_data : in   std_logic_vector(109 downto 0);
      mem_req0_pipe0_pipe_write_req : out  std_logic_vector(0 downto 0);
      mem_req0_pipe0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      mem_req0_pipe0_pipe_write_data : out  std_logic_vector(63 downto 0);
      mem_req0_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      mem_req0_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      mem_req0_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicToMemoryInterface
  signal nicToMemoryInterface_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicToMemoryInterface_tag_out   : std_logic_vector(1 downto 0);
  signal nicToMemoryInterface_start_req : std_logic;
  signal nicToMemoryInterface_start_ack : std_logic;
  signal nicToMemoryInterface_fin_req   : std_logic;
  signal nicToMemoryInterface_fin_ack : std_logic;
  -- declarations related to module nicToProcessorInterface
  component nicToProcessorInterface is -- 
    generic (tag_length : integer); 
    port ( -- 
      AFB_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(32 downto 0);
      control_word_response_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      control_word_response_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      control_word_response_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicToProcessorInterface
  signal nicToProcessorInterface_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicToProcessorInterface_tag_out   : std_logic_vector(1 downto 0);
  signal nicToProcessorInterface_start_req : std_logic;
  signal nicToProcessorInterface_start_ack : std_logic;
  signal nicToProcessorInterface_fin_req   : std_logic;
  signal nicToProcessorInterface_fin_ack : std_logic;
  -- declarations related to module popFromQueue
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module popFromQueue
  signal popFromQueue_lock :  std_logic_vector(0 downto 0);
  signal popFromQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal popFromQueue_q_r_data :  std_logic_vector(31 downto 0);
  signal popFromQueue_status :  std_logic_vector(0 downto 0);
  signal popFromQueue_in_args    : std_logic_vector(36 downto 0);
  signal popFromQueue_out_args   : std_logic_vector(32 downto 0);
  signal popFromQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal popFromQueue_tag_out   : std_logic_vector(2 downto 0);
  signal popFromQueue_start_req : std_logic;
  signal popFromQueue_start_ack : std_logic;
  signal popFromQueue_fin_req   : std_logic;
  signal popFromQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module popFromQueue
  signal popFromQueue_call_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_call_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_return_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_return_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_call_data: std_logic_vector(73 downto 0);
  signal popFromQueue_call_tag: std_logic_vector(1 downto 0);
  signal popFromQueue_return_data: std_logic_vector(65 downto 0);
  signal popFromQueue_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module populateRxQueue
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module populateRxQueue
  signal populateRxQueue_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal populateRxQueue_in_args    : std_logic_vector(35 downto 0);
  signal populateRxQueue_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal populateRxQueue_tag_out   : std_logic_vector(1 downto 0);
  signal populateRxQueue_start_req : std_logic;
  signal populateRxQueue_start_ack : std_logic;
  signal populateRxQueue_fin_req   : std_logic;
  signal populateRxQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module populateRxQueue
  signal populateRxQueue_call_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_data: std_logic_vector(35 downto 0);
  signal populateRxQueue_call_tag: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module processorToNicInterface
  component processorToNicInterface is -- 
    generic (tag_length : integer); 
    port ( -- 
      control_word_request_pipe_1_pipe_read_req : out  std_logic_vector(0 downto 0);
      control_word_request_pipe_1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      control_word_request_pipe_1_pipe_read_data : in   std_logic_vector(63 downto 0);
      control_word_request_pipe_0_pipe_read_req : out  std_logic_vector(0 downto 0);
      control_word_request_pipe_0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      control_word_request_pipe_0_pipe_read_data : in   std_logic_vector(31 downto 0);
      AFB_NIC_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_write_data : out  std_logic_vector(73 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module processorToNicInterface
  signal processorToNicInterface_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal processorToNicInterface_tag_out   : std_logic_vector(1 downto 0);
  signal processorToNicInterface_start_req : std_logic;
  signal processorToNicInterface_start_ack : std_logic;
  signal processorToNicInterface_fin_req   : std_logic;
  signal processorToNicInterface_fin_ack : std_logic;
  -- declarations related to module pushIntoQueue
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      releaseMutex_call_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_call_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_call_data : out  std_logic_vector(35 downto 0);
      releaseMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseMutex_return_reqs : out  std_logic_vector(0 downto 0);
      releaseMutex_return_acks : in   std_logic_vector(0 downto 0);
      releaseMutex_return_tag :  in   std_logic_vector(0 downto 0);
      acquireMutex_call_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_call_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_call_data : out  std_logic_vector(35 downto 0);
      acquireMutex_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireMutex_return_reqs : out  std_logic_vector(0 downto 0);
      acquireMutex_return_acks : in   std_logic_vector(0 downto 0);
      acquireMutex_return_data : in   std_logic_vector(0 downto 0);
      acquireMutex_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module pushIntoQueue
  signal pushIntoQueue_lock :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal pushIntoQueue_q_w_data :  std_logic_vector(31 downto 0);
  signal pushIntoQueue_status :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_in_args    : std_logic_vector(68 downto 0);
  signal pushIntoQueue_out_args   : std_logic_vector(0 downto 0);
  signal pushIntoQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal pushIntoQueue_tag_out   : std_logic_vector(2 downto 0);
  signal pushIntoQueue_start_req : std_logic;
  signal pushIntoQueue_start_ack : std_logic;
  signal pushIntoQueue_fin_req   : std_logic;
  signal pushIntoQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module pushIntoQueue
  signal pushIntoQueue_call_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_data: std_logic_vector(206 downto 0);
  signal pushIntoQueue_call_tag: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_data: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module releaseMutex
  component releaseMutex is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module releaseMutex
  signal releaseMutex_q_base_address :  std_logic_vector(35 downto 0);
  signal releaseMutex_in_args    : std_logic_vector(35 downto 0);
  signal releaseMutex_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal releaseMutex_tag_out   : std_logic_vector(2 downto 0);
  signal releaseMutex_start_req : std_logic;
  signal releaseMutex_start_ack : std_logic;
  signal releaseMutex_fin_req   : std_logic;
  signal releaseMutex_fin_ack : std_logic;
  -- caller side aggregated signals for module releaseMutex
  signal releaseMutex_call_reqs: std_logic_vector(1 downto 0);
  signal releaseMutex_call_acks: std_logic_vector(1 downto 0);
  signal releaseMutex_return_reqs: std_logic_vector(1 downto 0);
  signal releaseMutex_return_acks: std_logic_vector(1 downto 0);
  signal releaseMutex_call_data: std_logic_vector(71 downto 0);
  signal releaseMutex_call_tag: std_logic_vector(1 downto 0);
  signal releaseMutex_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setQueueElement
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_pointer : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueueElement
  signal setQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueueElement_write_pointer :  std_logic_vector(31 downto 0);
  signal setQueueElement_q_w_data :  std_logic_vector(31 downto 0);
  signal setQueueElement_in_args    : std_logic_vector(99 downto 0);
  signal setQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal setQueueElement_start_req : std_logic;
  signal setQueueElement_start_ack : std_logic;
  signal setQueueElement_fin_req   : std_logic;
  signal setQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueueElement
  signal setQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_call_data: std_logic_vector(99 downto 0);
  signal setQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal setQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueuePointers
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueuePointers
  signal setQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_in_args    : std_logic_vector(99 downto 0);
  signal setQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal setQueuePointers_start_req : std_logic;
  signal setQueuePointers_start_ack : std_logic;
  signal setQueuePointers_fin_req   : std_logic;
  signal setQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueuePointers
  signal setQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_data: std_logic_vector(199 downto 0);
  signal setQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module transmitEngineDaemon
  component transmitEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
      getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
      getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
      transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_call_data : out  std_logic_vector(31 downto 0);
      transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
      transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_return_data : in   std_logic_vector(0 downto 0);
      transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitEngineDaemon
  signal transmitEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal transmitEngineDaemon_start_req : std_logic;
  signal transmitEngineDaemon_start_ack : std_logic;
  signal transmitEngineDaemon_fin_req   : std_logic;
  signal transmitEngineDaemon_fin_ack : std_logic;
  -- declarations related to module transmitPacket
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(3 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitPacket
  signal transmitPacket_packet_pointer :  std_logic_vector(31 downto 0);
  signal transmitPacket_status :  std_logic_vector(0 downto 0);
  signal transmitPacket_in_args    : std_logic_vector(31 downto 0);
  signal transmitPacket_out_args   : std_logic_vector(0 downto 0);
  signal transmitPacket_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitPacket_tag_out   : std_logic_vector(1 downto 0);
  signal transmitPacket_start_req : std_logic;
  signal transmitPacket_start_ack : std_logic;
  signal transmitPacket_fin_req   : std_logic;
  signal transmitPacket_fin_ack : std_logic;
  -- caller side aggregated signals for module transmitPacket
  signal transmitPacket_call_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_call_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_return_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_return_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_call_data: std_logic_vector(31 downto 0);
  signal transmitPacket_call_tag: std_logic_vector(0 downto 0);
  signal transmitPacket_return_data: std_logic_vector(0 downto 0);
  signal transmitPacket_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeControlInformationToMem
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(7 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeControlInformationToMem
  signal writeControlInformationToMem_base_buffer_pointer :  std_logic_vector(35 downto 0);
  signal writeControlInformationToMem_packet_size :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_in_args    : std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeControlInformationToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeControlInformationToMem_start_req : std_logic;
  signal writeControlInformationToMem_start_ack : std_logic;
  signal writeControlInformationToMem_fin_req   : std_logic;
  signal writeControlInformationToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeControlInformationToMem
  signal writeControlInformationToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_data: std_logic_vector(51 downto 0);
  signal writeControlInformationToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeEthernetHeaderToMem
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_buf_position :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_in_args    : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_out_args   : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeEthernetHeaderToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeEthernetHeaderToMem_start_req : std_logic;
  signal writeEthernetHeaderToMem_start_ack : std_logic;
  signal writeEthernetHeaderToMem_fin_req   : std_logic;
  signal writeEthernetHeaderToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writePayloadToMem
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(7 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(1 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writePayloadToMem
  signal writePayloadToMem_base_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_packet_size_32 :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal writePayloadToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_in_args    : std_logic_vector(71 downto 0);
  signal writePayloadToMem_out_args   : std_logic_vector(16 downto 0);
  signal writePayloadToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writePayloadToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writePayloadToMem_start_req : std_logic;
  signal writePayloadToMem_start_ack : std_logic;
  signal writePayloadToMem_fin_req   : std_logic;
  signal writePayloadToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writePayloadToMem
  signal writePayloadToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_data: std_logic_vector(71 downto 0);
  signal writePayloadToMem_call_tag: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_data: std_logic_vector(16 downto 0);
  signal writePayloadToMem_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_write_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_read_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_write_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_read_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe CONTROL_REGISTER
  signal CONTROL_REGISTER_pipe_write_data: std_logic_vector(31 downto 0);
  signal CONTROL_REGISTER_pipe_write_req: std_logic_vector(0 downto 0);
  signal CONTROL_REGISTER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe CONTROL_REGISTER
  signal CONTROL_REGISTER: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe FREE_Q
  signal FREE_Q_pipe_write_data: std_logic_vector(35 downto 0);
  signal FREE_Q_pipe_write_req: std_logic_vector(0 downto 0);
  signal FREE_Q_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe FREE_Q
  signal FREE_Q: std_logic_vector(35 downto 0);
  -- aggregate signals for write to pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_write_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_read_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS_pipe_write_data: std_logic_vector(31 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_req: std_logic_vector(0 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS: std_logic_vector(31 downto 0);
  -- aggregate signals for read from pipe control_word_request_pipe_0
  signal control_word_request_pipe_0_pipe_read_data: std_logic_vector(31 downto 0);
  signal control_word_request_pipe_0_pipe_read_req: std_logic_vector(0 downto 0);
  signal control_word_request_pipe_0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe control_word_request_pipe_1
  signal control_word_request_pipe_1_pipe_read_data: std_logic_vector(63 downto 0);
  signal control_word_request_pipe_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal control_word_request_pipe_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe control_word_response_pipe
  signal control_word_response_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal control_word_response_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal control_word_response_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_write_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_read_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data_0
  signal mac_to_nic_data_0_pipe_read_data: std_logic_vector(63 downto 0);
  signal mac_to_nic_data_0_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data_1
  signal mac_to_nic_data_1_pipe_read_data: std_logic_vector(15 downto 0);
  signal mac_to_nic_data_1_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe mem_req0_pipe0
  signal mem_req0_pipe0_pipe_write_data: std_logic_vector(63 downto 0);
  signal mem_req0_pipe0_pipe_write_req: std_logic_vector(0 downto 0);
  signal mem_req0_pipe0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe mem_req0_pipe1
  signal mem_req0_pipe1_pipe_write_data: std_logic_vector(63 downto 0);
  signal mem_req0_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal mem_req0_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mem_resp0_pipe0
  signal mem_resp0_pipe0_pipe_read_data: std_logic_vector(63 downto 0);
  signal mem_resp0_pipe0_pipe_read_req: std_logic_vector(0 downto 0);
  signal mem_resp0_pipe0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mem_resp0_pipe1
  signal mem_resp0_pipe1_pipe_read_data: std_logic_vector(7 downto 0);
  signal mem_resp0_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal mem_resp0_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module AccessRegister
  AccessRegister_rwbar <= AccessRegister_in_args(42 downto 42);
  AccessRegister_bmask <= AccessRegister_in_args(41 downto 38);
  AccessRegister_register_index <= AccessRegister_in_args(37 downto 32);
  AccessRegister_wdata <= AccessRegister_in_args(31 downto 0);
  AccessRegister_out_args <= AccessRegister_rdata ;
  -- call arbiter for module AccessRegister
  AccessRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 43,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => AccessRegister_call_reqs,
      call_acks => AccessRegister_call_acks,
      return_reqs => AccessRegister_return_reqs,
      return_acks => AccessRegister_return_acks,
      call_data  => AccessRegister_call_data,
      call_tag  => AccessRegister_call_tag,
      return_tag  => AccessRegister_return_tag,
      call_mtag => AccessRegister_tag_in,
      return_mtag => AccessRegister_tag_out,
      return_data =>AccessRegister_return_data,
      call_mreq => AccessRegister_start_req,
      call_mack => AccessRegister_start_ack,
      return_mreq => AccessRegister_fin_req,
      return_mack => AccessRegister_fin_ack,
      call_mdata => AccessRegister_in_args,
      return_mdata => AccessRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  AccessRegister_instance:AccessRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      rwbar => AccessRegister_rwbar,
      bmask => AccessRegister_bmask,
      register_index => AccessRegister_register_index,
      wdata => AccessRegister_wdata,
      rdata => AccessRegister_rdata,
      start_req => AccessRegister_start_req,
      start_ack => AccessRegister_start_ack,
      fin_req => AccessRegister_fin_req,
      fin_ack => AccessRegister_fin_ack,
      clk => clk,
      reset => reset,
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
      tag_in => AccessRegister_tag_in,
      tag_out => AccessRegister_tag_out-- 
    ); -- 
  -- module NicRegisterAccessDaemon
  NicRegisterAccessDaemon_instance:NicRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => NicRegisterAccessDaemon_start_req,
      start_ack => NicRegisterAccessDaemon_start_ack,
      fin_req => NicRegisterAccessDaemon_fin_req,
      fin_ack => NicRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(11 downto 6),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(1 downto 1),
      UpdateRegister_call_acks => UpdateRegister_call_acks(1 downto 1),
      UpdateRegister_call_data => UpdateRegister_call_data(147 downto 74),
      UpdateRegister_call_tag => UpdateRegister_call_tag(1 downto 1),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(1 downto 1),
      UpdateRegister_return_acks => UpdateRegister_return_acks(1 downto 1),
      UpdateRegister_return_data => UpdateRegister_return_data(63 downto 32),
      UpdateRegister_return_tag => UpdateRegister_return_tag(1 downto 1),
      tag_in => NicRegisterAccessDaemon_tag_in,
      tag_out => NicRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  NicRegisterAccessDaemon_tag_in <= (others => '0');
  NicRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => NicRegisterAccessDaemon_start_req, start_ack => NicRegisterAccessDaemon_start_ack,  fin_req => NicRegisterAccessDaemon_fin_req,  fin_ack => NicRegisterAccessDaemon_fin_ack);
  -- module ReceiveEngineDaemon
  ReceiveEngineDaemon_instance:ReceiveEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ReceiveEngineDaemon_start_req,
      start_ack => ReceiveEngineDaemon_start_ack,
      fin_req => ReceiveEngineDaemon_fin_req,
      fin_ack => ReceiveEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      FREE_Q => FREE_Q,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(11 downto 6),
      popFromQueue_call_reqs => popFromQueue_call_reqs(1 downto 1),
      popFromQueue_call_acks => popFromQueue_call_acks(1 downto 1),
      popFromQueue_call_data => popFromQueue_call_data(73 downto 37),
      popFromQueue_call_tag => popFromQueue_call_tag(1 downto 1),
      popFromQueue_return_reqs => popFromQueue_return_reqs(1 downto 1),
      popFromQueue_return_acks => popFromQueue_return_acks(1 downto 1),
      popFromQueue_return_data => popFromQueue_return_data(65 downto 33),
      popFromQueue_return_tag => popFromQueue_return_tag(1 downto 1),
      loadBuffer_call_reqs => loadBuffer_call_reqs(0 downto 0),
      loadBuffer_call_acks => loadBuffer_call_acks(0 downto 0),
      loadBuffer_call_data => loadBuffer_call_data(35 downto 0),
      loadBuffer_call_tag => loadBuffer_call_tag(0 downto 0),
      loadBuffer_return_reqs => loadBuffer_return_reqs(0 downto 0),
      loadBuffer_return_acks => loadBuffer_return_acks(0 downto 0),
      loadBuffer_return_data => loadBuffer_return_data(0 downto 0),
      loadBuffer_return_tag => loadBuffer_return_tag(0 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(2 downto 2),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(2 downto 2),
      pushIntoQueue_call_data => pushIntoQueue_call_data(206 downto 138),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(2 downto 2),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(2 downto 2),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(2 downto 2),
      pushIntoQueue_return_data => pushIntoQueue_return_data(2 downto 2),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(2 downto 2),
      populateRxQueue_call_reqs => populateRxQueue_call_reqs(0 downto 0),
      populateRxQueue_call_acks => populateRxQueue_call_acks(0 downto 0),
      populateRxQueue_call_data => populateRxQueue_call_data(35 downto 0),
      populateRxQueue_call_tag => populateRxQueue_call_tag(0 downto 0),
      populateRxQueue_return_reqs => populateRxQueue_return_reqs(0 downto 0),
      populateRxQueue_return_acks => populateRxQueue_return_acks(0 downto 0),
      populateRxQueue_return_tag => populateRxQueue_return_tag(0 downto 0),
      tag_in => ReceiveEngineDaemon_tag_in,
      tag_out => ReceiveEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  ReceiveEngineDaemon_tag_in <= (others => '0');
  ReceiveEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ReceiveEngineDaemon_start_req, start_ack => ReceiveEngineDaemon_start_ack,  fin_req => ReceiveEngineDaemon_fin_req,  fin_ack => ReceiveEngineDaemon_fin_ack);
  -- module SoftwareRegisterAccessDaemon
  SoftwareRegisterAccessDaemon_instance:SoftwareRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => SoftwareRegisterAccessDaemon_start_req,
      start_ack => SoftwareRegisterAccessDaemon_start_ack,
      fin_req => SoftwareRegisterAccessDaemon_fin_req,
      fin_ack => SoftwareRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(5 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      AFB_NIC_REQUEST_pipe_read_req => AFB_NIC_REQUEST_pipe_read_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_ack => AFB_NIC_REQUEST_pipe_read_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_data => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
      CONTROL_REGISTER_pipe_write_req => CONTROL_REGISTER_pipe_write_req(0 downto 0),
      CONTROL_REGISTER_pipe_write_ack => CONTROL_REGISTER_pipe_write_ack(0 downto 0),
      CONTROL_REGISTER_pipe_write_data => CONTROL_REGISTER_pipe_write_data(31 downto 0),
      FREE_Q_pipe_write_req => FREE_Q_pipe_write_req(0 downto 0),
      FREE_Q_pipe_write_ack => FREE_Q_pipe_write_ack(0 downto 0),
      FREE_Q_pipe_write_data => FREE_Q_pipe_write_data(35 downto 0),
      AFB_NIC_RESPONSE_pipe_write_req => AFB_NIC_RESPONSE_pipe_write_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_ack => AFB_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_data => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
      NUMBER_OF_SERVERS_pipe_write_req => NUMBER_OF_SERVERS_pipe_write_req(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_ack => NUMBER_OF_SERVERS_pipe_write_ack(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_data => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(0 downto 0),
      UpdateRegister_call_acks => UpdateRegister_call_acks(0 downto 0),
      UpdateRegister_call_data => UpdateRegister_call_data(73 downto 0),
      UpdateRegister_call_tag => UpdateRegister_call_tag(0 downto 0),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(0 downto 0),
      UpdateRegister_return_acks => UpdateRegister_return_acks(0 downto 0),
      UpdateRegister_return_data => UpdateRegister_return_data(31 downto 0),
      UpdateRegister_return_tag => UpdateRegister_return_tag(0 downto 0),
      tag_in => SoftwareRegisterAccessDaemon_tag_in,
      tag_out => SoftwareRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  SoftwareRegisterAccessDaemon_tag_in <= (others => '0');
  SoftwareRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => SoftwareRegisterAccessDaemon_start_req, start_ack => SoftwareRegisterAccessDaemon_start_ack,  fin_req => SoftwareRegisterAccessDaemon_fin_req,  fin_ack => SoftwareRegisterAccessDaemon_fin_ack);
  -- module UpdateRegister
  UpdateRegister_bmask <= UpdateRegister_in_args(73 downto 70);
  UpdateRegister_rval <= UpdateRegister_in_args(69 downto 38);
  UpdateRegister_wdata <= UpdateRegister_in_args(37 downto 6);
  UpdateRegister_index <= UpdateRegister_in_args(5 downto 0);
  UpdateRegister_out_args <= UpdateRegister_wval ;
  -- call arbiter for module UpdateRegister
  UpdateRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 74,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => UpdateRegister_call_reqs,
      call_acks => UpdateRegister_call_acks,
      return_reqs => UpdateRegister_return_reqs,
      return_acks => UpdateRegister_return_acks,
      call_data  => UpdateRegister_call_data,
      call_tag  => UpdateRegister_call_tag,
      return_tag  => UpdateRegister_return_tag,
      call_mtag => UpdateRegister_tag_in,
      return_mtag => UpdateRegister_tag_out,
      return_data =>UpdateRegister_return_data,
      call_mreq => UpdateRegister_start_req,
      call_mack => UpdateRegister_start_ack,
      return_mreq => UpdateRegister_fin_req,
      return_mack => UpdateRegister_fin_ack,
      call_mdata => UpdateRegister_in_args,
      return_mdata => UpdateRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  UpdateRegister_instance:UpdateRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      bmask => UpdateRegister_bmask,
      rval => UpdateRegister_rval,
      wdata => UpdateRegister_wdata,
      index => UpdateRegister_index,
      wval => UpdateRegister_wval,
      start_req => UpdateRegister_start_req,
      start_ack => UpdateRegister_start_ack,
      fin_req => UpdateRegister_fin_req,
      fin_ack => UpdateRegister_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(5 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => UpdateRegister_tag_in,
      tag_out => UpdateRegister_tag_out-- 
    ); -- 
  -- module accessMemory
  accessMemory_lock <= accessMemory_in_args(109 downto 109);
  accessMemory_rwbar <= accessMemory_in_args(108 downto 108);
  accessMemory_bmask <= accessMemory_in_args(107 downto 100);
  accessMemory_addr <= accessMemory_in_args(99 downto 64);
  accessMemory_wdata <= accessMemory_in_args(63 downto 0);
  accessMemory_out_args <= accessMemory_rdata ;
  -- call arbiter for module accessMemory
  accessMemory_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 11,
      call_data_width => 110,
      return_data_width => 64,
      callee_tag_length => 4,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => accessMemory_call_reqs,
      call_acks => accessMemory_call_acks,
      return_reqs => accessMemory_return_reqs,
      return_acks => accessMemory_return_acks,
      call_data  => accessMemory_call_data,
      call_tag  => accessMemory_call_tag,
      return_tag  => accessMemory_return_tag,
      call_mtag => accessMemory_tag_in,
      return_mtag => accessMemory_tag_out,
      return_data =>accessMemory_return_data,
      call_mreq => accessMemory_start_req,
      call_mack => accessMemory_start_ack,
      return_mreq => accessMemory_fin_req,
      return_mack => accessMemory_fin_ack,
      call_mdata => accessMemory_in_args,
      return_mdata => accessMemory_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemory_instance:accessMemory-- 
    generic map(tag_length => 6)
    port map(-- 
      lock => accessMemory_lock,
      rwbar => accessMemory_rwbar,
      bmask => accessMemory_bmask,
      addr => accessMemory_addr,
      wdata => accessMemory_wdata,
      rdata => accessMemory_rdata,
      start_req => accessMemory_start_req,
      start_ack => accessMemory_start_ack,
      fin_req => accessMemory_fin_req,
      fin_ack => accessMemory_fin_ack,
      clk => clk,
      reset => reset,
      MEMORY_TO_NIC_RESPONSE_pipe_read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessMemory_tag_in,
      tag_out => accessMemory_tag_out-- 
    ); -- 
  -- module acquireMutex
  acquireMutex_q_base_address <= acquireMutex_in_args(35 downto 0);
  acquireMutex_out_args <= acquireMutex_m_ok ;
  -- call arbiter for module acquireMutex
  acquireMutex_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => acquireMutex_call_reqs,
      call_acks => acquireMutex_call_acks,
      return_reqs => acquireMutex_return_reqs,
      return_acks => acquireMutex_return_acks,
      call_data  => acquireMutex_call_data,
      call_tag  => acquireMutex_call_tag,
      return_tag  => acquireMutex_return_tag,
      call_mtag => acquireMutex_tag_in,
      return_mtag => acquireMutex_tag_out,
      return_data =>acquireMutex_return_data,
      call_mreq => acquireMutex_start_req,
      call_mack => acquireMutex_start_ack,
      return_mreq => acquireMutex_fin_req,
      return_mack => acquireMutex_fin_ack,
      call_mdata => acquireMutex_in_args,
      return_mdata => acquireMutex_out_args,
      clk => clk, 
      reset => reset --
    ); --
  acquireMutex_instance:acquireMutex-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => acquireMutex_q_base_address,
      m_ok => acquireMutex_m_ok,
      start_req => acquireMutex_start_req,
      start_ack => acquireMutex_start_ack,
      fin_req => acquireMutex_fin_req,
      fin_ack => acquireMutex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(5 downto 5),
      accessMemory_call_acks => accessMemory_call_acks(5 downto 5),
      accessMemory_call_data => accessMemory_call_data(659 downto 550),
      accessMemory_call_tag => accessMemory_call_tag(11 downto 10),
      accessMemory_return_reqs => accessMemory_return_reqs(5 downto 5),
      accessMemory_return_acks => accessMemory_return_acks(5 downto 5),
      accessMemory_return_data => accessMemory_return_data(383 downto 320),
      accessMemory_return_tag => accessMemory_return_tag(11 downto 10),
      tag_in => acquireMutex_tag_in,
      tag_out => acquireMutex_tag_out-- 
    ); -- 
  -- module getQueueElement
  getQueueElement_q_base_address <= getQueueElement_in_args(67 downto 32);
  getQueueElement_read_pointer <= getQueueElement_in_args(31 downto 0);
  getQueueElement_out_args <= getQueueElement_q_r_data ;
  -- call arbiter for module getQueueElement
  getQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 68,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueElement_call_reqs,
      call_acks => getQueueElement_call_acks,
      return_reqs => getQueueElement_return_reqs,
      return_acks => getQueueElement_return_acks,
      call_data  => getQueueElement_call_data,
      call_tag  => getQueueElement_call_tag,
      return_tag  => getQueueElement_return_tag,
      call_mtag => getQueueElement_tag_in,
      return_mtag => getQueueElement_tag_out,
      return_data =>getQueueElement_return_data,
      call_mreq => getQueueElement_start_req,
      call_mack => getQueueElement_start_ack,
      return_mreq => getQueueElement_fin_req,
      return_mack => getQueueElement_fin_ack,
      call_mdata => getQueueElement_in_args,
      return_mdata => getQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueElement_instance:getQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => getQueueElement_q_base_address,
      read_pointer => getQueueElement_read_pointer,
      q_r_data => getQueueElement_q_r_data,
      start_req => getQueueElement_start_req,
      start_ack => getQueueElement_start_ack,
      fin_req => getQueueElement_fin_req,
      fin_ack => getQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(7 downto 7),
      accessMemory_call_acks => accessMemory_call_acks(7 downto 7),
      accessMemory_call_data => accessMemory_call_data(879 downto 770),
      accessMemory_call_tag => accessMemory_call_tag(15 downto 14),
      accessMemory_return_reqs => accessMemory_return_reqs(7 downto 7),
      accessMemory_return_acks => accessMemory_return_acks(7 downto 7),
      accessMemory_return_data => accessMemory_return_data(511 downto 448),
      accessMemory_return_tag => accessMemory_return_tag(15 downto 14),
      tag_in => getQueueElement_tag_in,
      tag_out => getQueueElement_tag_out-- 
    ); -- 
  -- module getQueuePointers
  getQueuePointers_q_base_address <= getQueuePointers_in_args(35 downto 0);
  getQueuePointers_out_args <= getQueuePointers_wp & getQueuePointers_rp ;
  -- call arbiter for module getQueuePointers
  getQueuePointers_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointers_call_reqs,
      call_acks => getQueuePointers_call_acks,
      return_reqs => getQueuePointers_return_reqs,
      return_acks => getQueuePointers_return_acks,
      call_data  => getQueuePointers_call_data,
      call_tag  => getQueuePointers_call_tag,
      return_tag  => getQueuePointers_return_tag,
      call_mtag => getQueuePointers_tag_in,
      return_mtag => getQueuePointers_tag_out,
      return_data =>getQueuePointers_return_data,
      call_mreq => getQueuePointers_start_req,
      call_mack => getQueuePointers_start_ack,
      return_mreq => getQueuePointers_fin_req,
      return_mack => getQueuePointers_fin_ack,
      call_mdata => getQueuePointers_in_args,
      return_mdata => getQueuePointers_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointers_instance:getQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueuePointers_q_base_address,
      wp => getQueuePointers_wp,
      rp => getQueuePointers_rp,
      start_req => getQueuePointers_start_req,
      start_ack => getQueuePointers_start_ack,
      fin_req => getQueuePointers_fin_req,
      fin_ack => getQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(4 downto 4),
      accessMemory_call_acks => accessMemory_call_acks(4 downto 4),
      accessMemory_call_data => accessMemory_call_data(549 downto 440),
      accessMemory_call_tag => accessMemory_call_tag(9 downto 8),
      accessMemory_return_reqs => accessMemory_return_reqs(4 downto 4),
      accessMemory_return_acks => accessMemory_return_acks(4 downto 4),
      accessMemory_return_data => accessMemory_return_data(319 downto 256),
      accessMemory_return_tag => accessMemory_return_tag(9 downto 8),
      tag_in => getQueuePointers_tag_in,
      tag_out => getQueuePointers_tag_out-- 
    ); -- 
  -- module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_queue_index <= getTxPacketPointerFromServer_in_args(5 downto 0);
  getTxPacketPointerFromServer_out_args <= getTxPacketPointerFromServer_pkt_pointer & getTxPacketPointerFromServer_status ;
  -- call arbiter for module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 6,
      return_data_width => 33,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTxPacketPointerFromServer_call_reqs,
      call_acks => getTxPacketPointerFromServer_call_acks,
      return_reqs => getTxPacketPointerFromServer_return_reqs,
      return_acks => getTxPacketPointerFromServer_return_acks,
      call_data  => getTxPacketPointerFromServer_call_data,
      call_tag  => getTxPacketPointerFromServer_call_tag,
      return_tag  => getTxPacketPointerFromServer_return_tag,
      call_mtag => getTxPacketPointerFromServer_tag_in,
      return_mtag => getTxPacketPointerFromServer_tag_out,
      return_data =>getTxPacketPointerFromServer_return_data,
      call_mreq => getTxPacketPointerFromServer_start_req,
      call_mack => getTxPacketPointerFromServer_start_ack,
      return_mreq => getTxPacketPointerFromServer_fin_req,
      return_mack => getTxPacketPointerFromServer_fin_ack,
      call_mdata => getTxPacketPointerFromServer_in_args,
      return_mdata => getTxPacketPointerFromServer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTxPacketPointerFromServer_instance:getTxPacketPointerFromServer-- 
    generic map(tag_length => 2)
    port map(-- 
      queue_index => getTxPacketPointerFromServer_queue_index,
      pkt_pointer => getTxPacketPointerFromServer_pkt_pointer,
      status => getTxPacketPointerFromServer_status,
      start_req => getTxPacketPointerFromServer_start_req,
      start_ack => getTxPacketPointerFromServer_start_ack,
      fin_req => getTxPacketPointerFromServer_fin_req,
      fin_ack => getTxPacketPointerFromServer_fin_ack,
      clk => clk,
      reset => reset,
      AccessRegister_call_reqs => AccessRegister_call_reqs(0 downto 0),
      AccessRegister_call_acks => AccessRegister_call_acks(0 downto 0),
      AccessRegister_call_data => AccessRegister_call_data(42 downto 0),
      AccessRegister_call_tag => AccessRegister_call_tag(0 downto 0),
      AccessRegister_return_reqs => AccessRegister_return_reqs(0 downto 0),
      AccessRegister_return_acks => AccessRegister_return_acks(0 downto 0),
      AccessRegister_return_data => AccessRegister_return_data(31 downto 0),
      AccessRegister_return_tag => AccessRegister_return_tag(0 downto 0),
      popFromQueue_call_reqs => popFromQueue_call_reqs(0 downto 0),
      popFromQueue_call_acks => popFromQueue_call_acks(0 downto 0),
      popFromQueue_call_data => popFromQueue_call_data(36 downto 0),
      popFromQueue_call_tag => popFromQueue_call_tag(0 downto 0),
      popFromQueue_return_reqs => popFromQueue_return_reqs(0 downto 0),
      popFromQueue_return_acks => popFromQueue_return_acks(0 downto 0),
      popFromQueue_return_data => popFromQueue_return_data(32 downto 0),
      popFromQueue_return_tag => popFromQueue_return_tag(0 downto 0),
      tag_in => getTxPacketPointerFromServer_tag_in,
      tag_out => getTxPacketPointerFromServer_tag_out-- 
    ); -- 
  -- module loadBuffer
  loadBuffer_rx_buffer_pointer <= loadBuffer_in_args(35 downto 0);
  loadBuffer_out_args <= loadBuffer_bad_packet_identifier ;
  -- call arbiter for module loadBuffer
  loadBuffer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadBuffer_call_reqs,
      call_acks => loadBuffer_call_acks,
      return_reqs => loadBuffer_return_reqs,
      return_acks => loadBuffer_return_acks,
      call_data  => loadBuffer_call_data,
      call_tag  => loadBuffer_call_tag,
      return_tag  => loadBuffer_return_tag,
      call_mtag => loadBuffer_tag_in,
      return_mtag => loadBuffer_tag_out,
      return_data =>loadBuffer_return_data,
      call_mreq => loadBuffer_start_req,
      call_mack => loadBuffer_start_ack,
      return_mreq => loadBuffer_fin_req,
      return_mack => loadBuffer_fin_ack,
      call_mdata => loadBuffer_in_args,
      return_mdata => loadBuffer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  loadBuffer_instance:loadBuffer-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => loadBuffer_rx_buffer_pointer,
      bad_packet_identifier => loadBuffer_bad_packet_identifier,
      start_req => loadBuffer_start_req,
      start_ack => loadBuffer_start_ack,
      fin_req => loadBuffer_fin_req,
      fin_ack => loadBuffer_fin_ack,
      clk => clk,
      reset => reset,
      writeEthernetHeaderToMem_call_reqs => writeEthernetHeaderToMem_call_reqs(0 downto 0),
      writeEthernetHeaderToMem_call_acks => writeEthernetHeaderToMem_call_acks(0 downto 0),
      writeEthernetHeaderToMem_call_data => writeEthernetHeaderToMem_call_data(35 downto 0),
      writeEthernetHeaderToMem_call_tag => writeEthernetHeaderToMem_call_tag(0 downto 0),
      writeEthernetHeaderToMem_return_reqs => writeEthernetHeaderToMem_return_reqs(0 downto 0),
      writeEthernetHeaderToMem_return_acks => writeEthernetHeaderToMem_return_acks(0 downto 0),
      writeEthernetHeaderToMem_return_data => writeEthernetHeaderToMem_return_data(35 downto 0),
      writeEthernetHeaderToMem_return_tag => writeEthernetHeaderToMem_return_tag(0 downto 0),
      writePayloadToMem_call_reqs => writePayloadToMem_call_reqs(0 downto 0),
      writePayloadToMem_call_acks => writePayloadToMem_call_acks(0 downto 0),
      writePayloadToMem_call_data => writePayloadToMem_call_data(71 downto 0),
      writePayloadToMem_call_tag => writePayloadToMem_call_tag(0 downto 0),
      writePayloadToMem_return_reqs => writePayloadToMem_return_reqs(0 downto 0),
      writePayloadToMem_return_acks => writePayloadToMem_return_acks(0 downto 0),
      writePayloadToMem_return_data => writePayloadToMem_return_data(16 downto 0),
      writePayloadToMem_return_tag => writePayloadToMem_return_tag(0 downto 0),
      writeControlInformationToMem_call_reqs => writeControlInformationToMem_call_reqs(0 downto 0),
      writeControlInformationToMem_call_acks => writeControlInformationToMem_call_acks(0 downto 0),
      writeControlInformationToMem_call_data => writeControlInformationToMem_call_data(51 downto 0),
      writeControlInformationToMem_call_tag => writeControlInformationToMem_call_tag(0 downto 0),
      writeControlInformationToMem_return_reqs => writeControlInformationToMem_return_reqs(0 downto 0),
      writeControlInformationToMem_return_acks => writeControlInformationToMem_return_acks(0 downto 0),
      writeControlInformationToMem_return_tag => writeControlInformationToMem_return_tag(0 downto 0),
      tag_in => loadBuffer_tag_in,
      tag_out => loadBuffer_tag_out-- 
    ); -- 
  -- module macToNicInterface
  macToNicInterface_instance:macToNicInterface-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => macToNicInterface_start_req,
      start_ack => macToNicInterface_start_ack,
      fin_req => macToNicInterface_fin_req,
      fin_ack => macToNicInterface_fin_ack,
      clk => clk,
      reset => reset,
      mac_to_nic_data_0_pipe_read_req => mac_to_nic_data_0_pipe_read_req(0 downto 0),
      mac_to_nic_data_0_pipe_read_ack => mac_to_nic_data_0_pipe_read_ack(0 downto 0),
      mac_to_nic_data_0_pipe_read_data => mac_to_nic_data_0_pipe_read_data(63 downto 0),
      mac_to_nic_data_1_pipe_read_req => mac_to_nic_data_1_pipe_read_req(0 downto 0),
      mac_to_nic_data_1_pipe_read_ack => mac_to_nic_data_1_pipe_read_ack(0 downto 0),
      mac_to_nic_data_1_pipe_read_data => mac_to_nic_data_1_pipe_read_data(15 downto 0),
      mac_to_nic_data_pipe_write_req => mac_to_nic_data_pipe_write_req(0 downto 0),
      mac_to_nic_data_pipe_write_ack => mac_to_nic_data_pipe_write_ack(0 downto 0),
      mac_to_nic_data_pipe_write_data => mac_to_nic_data_pipe_write_data(72 downto 0),
      tag_in => macToNicInterface_tag_in,
      tag_out => macToNicInterface_tag_out-- 
    ); -- 
  -- module will be run forever 
  macToNicInterface_tag_in <= (others => '0');
  macToNicInterface_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => macToNicInterface_start_req, start_ack => macToNicInterface_start_ack,  fin_req => macToNicInterface_fin_req,  fin_ack => macToNicInterface_fin_ack);
  -- module memoryToNicInterface
  memoryToNicInterface_instance:memoryToNicInterface-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => memoryToNicInterface_start_req,
      start_ack => memoryToNicInterface_start_ack,
      fin_req => memoryToNicInterface_fin_req,
      fin_ack => memoryToNicInterface_fin_ack,
      clk => clk,
      reset => reset,
      mem_resp0_pipe0_pipe_read_req => mem_resp0_pipe0_pipe_read_req(0 downto 0),
      mem_resp0_pipe0_pipe_read_ack => mem_resp0_pipe0_pipe_read_ack(0 downto 0),
      mem_resp0_pipe0_pipe_read_data => mem_resp0_pipe0_pipe_read_data(63 downto 0),
      mem_resp0_pipe1_pipe_read_req => mem_resp0_pipe1_pipe_read_req(0 downto 0),
      mem_resp0_pipe1_pipe_read_ack => mem_resp0_pipe1_pipe_read_ack(0 downto 0),
      mem_resp0_pipe1_pipe_read_data => mem_resp0_pipe1_pipe_read_data(7 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data(64 downto 0),
      tag_in => memoryToNicInterface_tag_in,
      tag_out => memoryToNicInterface_tag_out-- 
    ); -- 
  -- module will be run forever 
  memoryToNicInterface_tag_in <= (others => '0');
  memoryToNicInterface_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => memoryToNicInterface_start_req, start_ack => memoryToNicInterface_start_ack,  fin_req => memoryToNicInterface_fin_req,  fin_ack => memoryToNicInterface_fin_ack);
  -- module nicRxFromMacDaemon
  nicRxFromMacDaemon_instance:nicRxFromMacDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicRxFromMacDaemon_start_req,
      start_ack => nicRxFromMacDaemon_start_ack,
      fin_req => nicRxFromMacDaemon_fin_req,
      fin_ack => nicRxFromMacDaemon_fin_ack,
      clk => clk,
      reset => reset,
      mac_to_nic_data_pipe_read_req => mac_to_nic_data_pipe_read_req(0 downto 0),
      mac_to_nic_data_pipe_read_ack => mac_to_nic_data_pipe_read_ack(0 downto 0),
      mac_to_nic_data_pipe_read_data => mac_to_nic_data_pipe_read_data(72 downto 0),
      nic_rx_to_header_pipe_write_req => nic_rx_to_header_pipe_write_req(0 downto 0),
      nic_rx_to_header_pipe_write_ack => nic_rx_to_header_pipe_write_ack(0 downto 0),
      nic_rx_to_header_pipe_write_data => nic_rx_to_header_pipe_write_data(72 downto 0),
      nic_rx_to_packet_pipe_write_req => nic_rx_to_packet_pipe_write_req(0 downto 0),
      nic_rx_to_packet_pipe_write_ack => nic_rx_to_packet_pipe_write_ack(0 downto 0),
      nic_rx_to_packet_pipe_write_data => nic_rx_to_packet_pipe_write_data(72 downto 0),
      tag_in => nicRxFromMacDaemon_tag_in,
      tag_out => nicRxFromMacDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicRxFromMacDaemon_tag_in <= (others => '0');
  nicRxFromMacDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicRxFromMacDaemon_start_req, start_ack => nicRxFromMacDaemon_start_ack,  fin_req => nicRxFromMacDaemon_fin_req,  fin_ack => nicRxFromMacDaemon_fin_ack);
  -- module nicToMacInterface
  nicToMacInterface_instance:nicToMacInterface-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicToMacInterface_start_req,
      start_ack => nicToMacInterface_start_ack,
      fin_req => nicToMacInterface_fin_req,
      fin_ack => nicToMacInterface_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_read_req => nic_to_mac_transmit_pipe_pipe_read_req(0 downto 0),
      nic_to_mac_transmit_pipe_pipe_read_ack => nic_to_mac_transmit_pipe_pipe_read_ack(0 downto 0),
      nic_to_mac_transmit_pipe_pipe_read_data => nic_to_mac_transmit_pipe_pipe_read_data(72 downto 0),
      tag_in => nicToMacInterface_tag_in,
      tag_out => nicToMacInterface_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicToMacInterface_tag_in <= (others => '0');
  nicToMacInterface_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicToMacInterface_start_req, start_ack => nicToMacInterface_start_ack,  fin_req => nicToMacInterface_fin_req,  fin_ack => nicToMacInterface_fin_ack);
  -- module nicToMemoryInterface
  nicToMemoryInterface_instance:nicToMemoryInterface-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicToMemoryInterface_start_req,
      start_ack => nicToMemoryInterface_start_ack,
      fin_req => nicToMemoryInterface_fin_req,
      fin_ack => nicToMemoryInterface_fin_ack,
      clk => clk,
      reset => reset,
      NIC_TO_MEMORY_REQUEST_pipe_read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data(109 downto 0),
      mem_req0_pipe0_pipe_write_req => mem_req0_pipe0_pipe_write_req(0 downto 0),
      mem_req0_pipe0_pipe_write_ack => mem_req0_pipe0_pipe_write_ack(0 downto 0),
      mem_req0_pipe0_pipe_write_data => mem_req0_pipe0_pipe_write_data(63 downto 0),
      mem_req0_pipe1_pipe_write_req => mem_req0_pipe1_pipe_write_req(0 downto 0),
      mem_req0_pipe1_pipe_write_ack => mem_req0_pipe1_pipe_write_ack(0 downto 0),
      mem_req0_pipe1_pipe_write_data => mem_req0_pipe1_pipe_write_data(63 downto 0),
      tag_in => nicToMemoryInterface_tag_in,
      tag_out => nicToMemoryInterface_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicToMemoryInterface_tag_in <= (others => '0');
  nicToMemoryInterface_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicToMemoryInterface_start_req, start_ack => nicToMemoryInterface_start_ack,  fin_req => nicToMemoryInterface_fin_req,  fin_ack => nicToMemoryInterface_fin_ack);
  -- module nicToProcessorInterface
  nicToProcessorInterface_instance:nicToProcessorInterface-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicToProcessorInterface_start_req,
      start_ack => nicToProcessorInterface_start_ack,
      fin_req => nicToProcessorInterface_fin_req,
      fin_ack => nicToProcessorInterface_fin_ack,
      clk => clk,
      reset => reset,
      AFB_NIC_RESPONSE_pipe_read_req => AFB_NIC_RESPONSE_pipe_read_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_read_ack => AFB_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_read_data => AFB_NIC_RESPONSE_pipe_read_data(32 downto 0),
      control_word_response_pipe_pipe_write_req => control_word_response_pipe_pipe_write_req(0 downto 0),
      control_word_response_pipe_pipe_write_ack => control_word_response_pipe_pipe_write_ack(0 downto 0),
      control_word_response_pipe_pipe_write_data => control_word_response_pipe_pipe_write_data(63 downto 0),
      tag_in => nicToProcessorInterface_tag_in,
      tag_out => nicToProcessorInterface_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicToProcessorInterface_tag_in <= (others => '0');
  nicToProcessorInterface_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicToProcessorInterface_start_req, start_ack => nicToProcessorInterface_start_ack,  fin_req => nicToProcessorInterface_fin_req,  fin_ack => nicToProcessorInterface_fin_ack);
  -- module popFromQueue
  popFromQueue_lock <= popFromQueue_in_args(36 downto 36);
  popFromQueue_q_base_address <= popFromQueue_in_args(35 downto 0);
  popFromQueue_out_args <= popFromQueue_q_r_data & popFromQueue_status ;
  -- call arbiter for module popFromQueue
  popFromQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 37,
      return_data_width => 33,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => popFromQueue_call_reqs,
      call_acks => popFromQueue_call_acks,
      return_reqs => popFromQueue_return_reqs,
      return_acks => popFromQueue_return_acks,
      call_data  => popFromQueue_call_data,
      call_tag  => popFromQueue_call_tag,
      return_tag  => popFromQueue_return_tag,
      call_mtag => popFromQueue_tag_in,
      return_mtag => popFromQueue_tag_out,
      return_data =>popFromQueue_return_data,
      call_mreq => popFromQueue_start_req,
      call_mack => popFromQueue_start_ack,
      return_mreq => popFromQueue_fin_req,
      return_mack => popFromQueue_fin_ack,
      call_mdata => popFromQueue_in_args,
      return_mdata => popFromQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  popFromQueue_instance:popFromQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => popFromQueue_lock,
      q_base_address => popFromQueue_q_base_address,
      q_r_data => popFromQueue_q_r_data,
      status => popFromQueue_status,
      start_req => popFromQueue_start_req,
      start_ack => popFromQueue_start_ack,
      fin_req => popFromQueue_fin_req,
      fin_ack => popFromQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireMutex_call_reqs => acquireMutex_call_reqs(0 downto 0),
      acquireMutex_call_acks => acquireMutex_call_acks(0 downto 0),
      acquireMutex_call_data => acquireMutex_call_data(35 downto 0),
      acquireMutex_call_tag => acquireMutex_call_tag(0 downto 0),
      acquireMutex_return_reqs => acquireMutex_return_reqs(0 downto 0),
      acquireMutex_return_acks => acquireMutex_return_acks(0 downto 0),
      acquireMutex_return_data => acquireMutex_return_data(0 downto 0),
      acquireMutex_return_tag => acquireMutex_return_tag(0 downto 0),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(0 downto 0),
      getQueuePointers_call_acks => getQueuePointers_call_acks(0 downto 0),
      getQueuePointers_call_data => getQueuePointers_call_data(35 downto 0),
      getQueuePointers_call_tag => getQueuePointers_call_tag(0 downto 0),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(0 downto 0),
      getQueuePointers_return_acks => getQueuePointers_return_acks(0 downto 0),
      getQueuePointers_return_data => getQueuePointers_return_data(63 downto 0),
      getQueuePointers_return_tag => getQueuePointers_return_tag(0 downto 0),
      getQueueElement_call_reqs => getQueueElement_call_reqs(0 downto 0),
      getQueueElement_call_acks => getQueueElement_call_acks(0 downto 0),
      getQueueElement_call_data => getQueueElement_call_data(67 downto 0),
      getQueueElement_call_tag => getQueueElement_call_tag(0 downto 0),
      getQueueElement_return_reqs => getQueueElement_return_reqs(0 downto 0),
      getQueueElement_return_acks => getQueueElement_return_acks(0 downto 0),
      getQueueElement_return_data => getQueueElement_return_data(31 downto 0),
      getQueueElement_return_tag => getQueueElement_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(0 downto 0),
      setQueuePointers_call_acks => setQueuePointers_call_acks(0 downto 0),
      setQueuePointers_call_data => setQueuePointers_call_data(99 downto 0),
      setQueuePointers_call_tag => setQueuePointers_call_tag(0 downto 0),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(0 downto 0),
      setQueuePointers_return_acks => setQueuePointers_return_acks(0 downto 0),
      setQueuePointers_return_tag => setQueuePointers_return_tag(0 downto 0),
      releaseMutex_call_reqs => releaseMutex_call_reqs(0 downto 0),
      releaseMutex_call_acks => releaseMutex_call_acks(0 downto 0),
      releaseMutex_call_data => releaseMutex_call_data(35 downto 0),
      releaseMutex_call_tag => releaseMutex_call_tag(0 downto 0),
      releaseMutex_return_reqs => releaseMutex_return_reqs(0 downto 0),
      releaseMutex_return_acks => releaseMutex_return_acks(0 downto 0),
      releaseMutex_return_tag => releaseMutex_return_tag(0 downto 0),
      tag_in => popFromQueue_tag_in,
      tag_out => popFromQueue_tag_out-- 
    ); -- 
  -- module populateRxQueue
  populateRxQueue_rx_buffer_pointer <= populateRxQueue_in_args(35 downto 0);
  -- call arbiter for module populateRxQueue
  populateRxQueue_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => populateRxQueue_call_reqs,
      call_acks => populateRxQueue_call_acks,
      return_reqs => populateRxQueue_return_reqs,
      return_acks => populateRxQueue_return_acks,
      call_data  => populateRxQueue_call_data,
      call_tag  => populateRxQueue_call_tag,
      return_tag  => populateRxQueue_return_tag,
      call_mtag => populateRxQueue_tag_in,
      return_mtag => populateRxQueue_tag_out,
      call_mreq => populateRxQueue_start_req,
      call_mack => populateRxQueue_start_ack,
      return_mreq => populateRxQueue_fin_req,
      return_mack => populateRxQueue_fin_ack,
      call_mdata => populateRxQueue_in_args,
      clk => clk, 
      reset => reset --
    ); --
  populateRxQueue_instance:populateRxQueue-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => populateRxQueue_rx_buffer_pointer,
      start_req => populateRxQueue_start_req,
      start_ack => populateRxQueue_start_ack,
      fin_req => populateRxQueue_fin_req,
      fin_ack => populateRxQueue_fin_ack,
      clk => clk,
      reset => reset,
      LAST_WRITTEN_RX_QUEUE_INDEX => LAST_WRITTEN_RX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(1 downto 1),
      AccessRegister_call_acks => AccessRegister_call_acks(1 downto 1),
      AccessRegister_call_data => AccessRegister_call_data(85 downto 43),
      AccessRegister_call_tag => AccessRegister_call_tag(1 downto 1),
      AccessRegister_return_reqs => AccessRegister_return_reqs(1 downto 1),
      AccessRegister_return_acks => AccessRegister_return_acks(1 downto 1),
      AccessRegister_return_data => AccessRegister_return_data(63 downto 32),
      AccessRegister_return_tag => AccessRegister_return_tag(1 downto 1),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(1 downto 1),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(1 downto 1),
      pushIntoQueue_call_data => pushIntoQueue_call_data(137 downto 69),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(1 downto 1),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(1 downto 1),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(1 downto 1),
      pushIntoQueue_return_data => pushIntoQueue_return_data(1 downto 1),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(1 downto 1),
      tag_in => populateRxQueue_tag_in,
      tag_out => populateRxQueue_tag_out-- 
    ); -- 
  -- module processorToNicInterface
  processorToNicInterface_instance:processorToNicInterface-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => processorToNicInterface_start_req,
      start_ack => processorToNicInterface_start_ack,
      fin_req => processorToNicInterface_fin_req,
      fin_ack => processorToNicInterface_fin_ack,
      clk => clk,
      reset => reset,
      control_word_request_pipe_1_pipe_read_req => control_word_request_pipe_1_pipe_read_req(0 downto 0),
      control_word_request_pipe_1_pipe_read_ack => control_word_request_pipe_1_pipe_read_ack(0 downto 0),
      control_word_request_pipe_1_pipe_read_data => control_word_request_pipe_1_pipe_read_data(63 downto 0),
      control_word_request_pipe_0_pipe_read_req => control_word_request_pipe_0_pipe_read_req(0 downto 0),
      control_word_request_pipe_0_pipe_read_ack => control_word_request_pipe_0_pipe_read_ack(0 downto 0),
      control_word_request_pipe_0_pipe_read_data => control_word_request_pipe_0_pipe_read_data(31 downto 0),
      AFB_NIC_REQUEST_pipe_write_req => AFB_NIC_REQUEST_pipe_write_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_write_ack => AFB_NIC_REQUEST_pipe_write_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_write_data => AFB_NIC_REQUEST_pipe_write_data(73 downto 0),
      tag_in => processorToNicInterface_tag_in,
      tag_out => processorToNicInterface_tag_out-- 
    ); -- 
  -- module will be run forever 
  processorToNicInterface_tag_in <= (others => '0');
  processorToNicInterface_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => processorToNicInterface_start_req, start_ack => processorToNicInterface_start_ack,  fin_req => processorToNicInterface_fin_req,  fin_ack => processorToNicInterface_fin_ack);
  -- module pushIntoQueue
  pushIntoQueue_lock <= pushIntoQueue_in_args(68 downto 68);
  pushIntoQueue_q_base_address <= pushIntoQueue_in_args(67 downto 32);
  pushIntoQueue_q_w_data <= pushIntoQueue_in_args(31 downto 0);
  pushIntoQueue_out_args <= pushIntoQueue_status ;
  -- call arbiter for module pushIntoQueue
  pushIntoQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 69,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => pushIntoQueue_call_reqs,
      call_acks => pushIntoQueue_call_acks,
      return_reqs => pushIntoQueue_return_reqs,
      return_acks => pushIntoQueue_return_acks,
      call_data  => pushIntoQueue_call_data,
      call_tag  => pushIntoQueue_call_tag,
      return_tag  => pushIntoQueue_return_tag,
      call_mtag => pushIntoQueue_tag_in,
      return_mtag => pushIntoQueue_tag_out,
      return_data =>pushIntoQueue_return_data,
      call_mreq => pushIntoQueue_start_req,
      call_mack => pushIntoQueue_start_ack,
      return_mreq => pushIntoQueue_fin_req,
      return_mack => pushIntoQueue_fin_ack,
      call_mdata => pushIntoQueue_in_args,
      return_mdata => pushIntoQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  pushIntoQueue_instance:pushIntoQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => pushIntoQueue_lock,
      q_base_address => pushIntoQueue_q_base_address,
      q_w_data => pushIntoQueue_q_w_data,
      status => pushIntoQueue_status,
      start_req => pushIntoQueue_start_req,
      start_ack => pushIntoQueue_start_ack,
      fin_req => pushIntoQueue_fin_req,
      fin_ack => pushIntoQueue_fin_ack,
      clk => clk,
      reset => reset,
      acquireMutex_call_reqs => acquireMutex_call_reqs(1 downto 1),
      acquireMutex_call_acks => acquireMutex_call_acks(1 downto 1),
      acquireMutex_call_data => acquireMutex_call_data(71 downto 36),
      acquireMutex_call_tag => acquireMutex_call_tag(1 downto 1),
      acquireMutex_return_reqs => acquireMutex_return_reqs(1 downto 1),
      acquireMutex_return_acks => acquireMutex_return_acks(1 downto 1),
      acquireMutex_return_data => acquireMutex_return_data(1 downto 1),
      acquireMutex_return_tag => acquireMutex_return_tag(1 downto 1),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(1 downto 1),
      getQueuePointers_call_acks => getQueuePointers_call_acks(1 downto 1),
      getQueuePointers_call_data => getQueuePointers_call_data(71 downto 36),
      getQueuePointers_call_tag => getQueuePointers_call_tag(1 downto 1),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(1 downto 1),
      getQueuePointers_return_acks => getQueuePointers_return_acks(1 downto 1),
      getQueuePointers_return_data => getQueuePointers_return_data(127 downto 64),
      getQueuePointers_return_tag => getQueuePointers_return_tag(1 downto 1),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(1 downto 1),
      setQueuePointers_call_acks => setQueuePointers_call_acks(1 downto 1),
      setQueuePointers_call_data => setQueuePointers_call_data(199 downto 100),
      setQueuePointers_call_tag => setQueuePointers_call_tag(1 downto 1),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(1 downto 1),
      setQueuePointers_return_acks => setQueuePointers_return_acks(1 downto 1),
      setQueuePointers_return_tag => setQueuePointers_return_tag(1 downto 1),
      releaseMutex_call_reqs => releaseMutex_call_reqs(1 downto 1),
      releaseMutex_call_acks => releaseMutex_call_acks(1 downto 1),
      releaseMutex_call_data => releaseMutex_call_data(71 downto 36),
      releaseMutex_call_tag => releaseMutex_call_tag(1 downto 1),
      releaseMutex_return_reqs => releaseMutex_return_reqs(1 downto 1),
      releaseMutex_return_acks => releaseMutex_return_acks(1 downto 1),
      releaseMutex_return_tag => releaseMutex_return_tag(1 downto 1),
      setQueueElement_call_reqs => setQueueElement_call_reqs(0 downto 0),
      setQueueElement_call_acks => setQueueElement_call_acks(0 downto 0),
      setQueueElement_call_data => setQueueElement_call_data(99 downto 0),
      setQueueElement_call_tag => setQueueElement_call_tag(0 downto 0),
      setQueueElement_return_reqs => setQueueElement_return_reqs(0 downto 0),
      setQueueElement_return_acks => setQueueElement_return_acks(0 downto 0),
      setQueueElement_return_tag => setQueueElement_return_tag(0 downto 0),
      tag_in => pushIntoQueue_tag_in,
      tag_out => pushIntoQueue_tag_out-- 
    ); -- 
  -- module releaseMutex
  releaseMutex_q_base_address <= releaseMutex_in_args(35 downto 0);
  -- call arbiter for module releaseMutex
  releaseMutex_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 36,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => releaseMutex_call_reqs,
      call_acks => releaseMutex_call_acks,
      return_reqs => releaseMutex_return_reqs,
      return_acks => releaseMutex_return_acks,
      call_data  => releaseMutex_call_data,
      call_tag  => releaseMutex_call_tag,
      return_tag  => releaseMutex_return_tag,
      call_mtag => releaseMutex_tag_in,
      return_mtag => releaseMutex_tag_out,
      call_mreq => releaseMutex_start_req,
      call_mack => releaseMutex_start_ack,
      return_mreq => releaseMutex_fin_req,
      return_mack => releaseMutex_fin_ack,
      call_mdata => releaseMutex_in_args,
      clk => clk, 
      reset => reset --
    ); --
  releaseMutex_instance:releaseMutex-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => releaseMutex_q_base_address,
      start_req => releaseMutex_start_req,
      start_ack => releaseMutex_start_ack,
      fin_req => releaseMutex_fin_req,
      fin_ack => releaseMutex_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(6 downto 6),
      accessMemory_call_acks => accessMemory_call_acks(6 downto 6),
      accessMemory_call_data => accessMemory_call_data(769 downto 660),
      accessMemory_call_tag => accessMemory_call_tag(13 downto 12),
      accessMemory_return_reqs => accessMemory_return_reqs(6 downto 6),
      accessMemory_return_acks => accessMemory_return_acks(6 downto 6),
      accessMemory_return_data => accessMemory_return_data(447 downto 384),
      accessMemory_return_tag => accessMemory_return_tag(13 downto 12),
      tag_in => releaseMutex_tag_in,
      tag_out => releaseMutex_tag_out-- 
    ); -- 
  -- module setQueueElement
  setQueueElement_q_base_address <= setQueueElement_in_args(99 downto 64);
  setQueueElement_write_pointer <= setQueueElement_in_args(63 downto 32);
  setQueueElement_q_w_data <= setQueueElement_in_args(31 downto 0);
  -- call arbiter for module setQueueElement
  setQueueElement_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 100,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueueElement_call_reqs,
      call_acks => setQueueElement_call_acks,
      return_reqs => setQueueElement_return_reqs,
      return_acks => setQueueElement_return_acks,
      call_data  => setQueueElement_call_data,
      call_tag  => setQueueElement_call_tag,
      return_tag  => setQueueElement_return_tag,
      call_mtag => setQueueElement_tag_in,
      return_mtag => setQueueElement_tag_out,
      call_mreq => setQueueElement_start_req,
      call_mack => setQueueElement_start_ack,
      return_mreq => setQueueElement_fin_req,
      return_mack => setQueueElement_fin_ack,
      call_mdata => setQueueElement_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueueElement_instance:setQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => setQueueElement_q_base_address,
      write_pointer => setQueueElement_write_pointer,
      q_w_data => setQueueElement_q_w_data,
      start_req => setQueueElement_start_req,
      start_ack => setQueueElement_start_ack,
      fin_req => setQueueElement_fin_req,
      fin_ack => setQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(9 downto 9),
      accessMemory_call_acks => accessMemory_call_acks(9 downto 9),
      accessMemory_call_data => accessMemory_call_data(1099 downto 990),
      accessMemory_call_tag => accessMemory_call_tag(19 downto 18),
      accessMemory_return_reqs => accessMemory_return_reqs(9 downto 9),
      accessMemory_return_acks => accessMemory_return_acks(9 downto 9),
      accessMemory_return_data => accessMemory_return_data(639 downto 576),
      accessMemory_return_tag => accessMemory_return_tag(19 downto 18),
      tag_in => setQueueElement_tag_in,
      tag_out => setQueueElement_tag_out-- 
    ); -- 
  -- module setQueuePointers
  setQueuePointers_q_base_address <= setQueuePointers_in_args(99 downto 64);
  setQueuePointers_wp <= setQueuePointers_in_args(63 downto 32);
  setQueuePointers_rp <= setQueuePointers_in_args(31 downto 0);
  -- call arbiter for module setQueuePointers
  setQueuePointers_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 100,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueuePointers_call_reqs,
      call_acks => setQueuePointers_call_acks,
      return_reqs => setQueuePointers_return_reqs,
      return_acks => setQueuePointers_return_acks,
      call_data  => setQueuePointers_call_data,
      call_tag  => setQueuePointers_call_tag,
      return_tag  => setQueuePointers_return_tag,
      call_mtag => setQueuePointers_tag_in,
      return_mtag => setQueuePointers_tag_out,
      call_mreq => setQueuePointers_start_req,
      call_mack => setQueuePointers_start_ack,
      return_mreq => setQueuePointers_fin_req,
      return_mack => setQueuePointers_fin_ack,
      call_mdata => setQueuePointers_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueuePointers_instance:setQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => setQueuePointers_q_base_address,
      wp => setQueuePointers_wp,
      rp => setQueuePointers_rp,
      start_req => setQueuePointers_start_req,
      start_ack => setQueuePointers_start_ack,
      fin_req => setQueuePointers_fin_req,
      fin_ack => setQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(8 downto 8),
      accessMemory_call_acks => accessMemory_call_acks(8 downto 8),
      accessMemory_call_data => accessMemory_call_data(989 downto 880),
      accessMemory_call_tag => accessMemory_call_tag(17 downto 16),
      accessMemory_return_reqs => accessMemory_return_reqs(8 downto 8),
      accessMemory_return_acks => accessMemory_return_acks(8 downto 8),
      accessMemory_return_data => accessMemory_return_data(575 downto 512),
      accessMemory_return_tag => accessMemory_return_tag(17 downto 16),
      tag_in => setQueuePointers_tag_in,
      tag_out => setQueuePointers_tag_out-- 
    ); -- 
  -- module transmitEngineDaemon
  transmitEngineDaemon_instance:transmitEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => transmitEngineDaemon_start_req,
      start_ack => transmitEngineDaemon_start_ack,
      fin_req => transmitEngineDaemon_fin_req,
      fin_ack => transmitEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      FREE_Q => FREE_Q,
      LAST_READ_TX_QUEUE_INDEX => LAST_READ_TX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(0 downto 0),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(0 downto 0),
      pushIntoQueue_call_data => pushIntoQueue_call_data(68 downto 0),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(0 downto 0),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(0 downto 0),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(0 downto 0),
      pushIntoQueue_return_data => pushIntoQueue_return_data(0 downto 0),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(0 downto 0),
      getTxPacketPointerFromServer_call_reqs => getTxPacketPointerFromServer_call_reqs(0 downto 0),
      getTxPacketPointerFromServer_call_acks => getTxPacketPointerFromServer_call_acks(0 downto 0),
      getTxPacketPointerFromServer_call_data => getTxPacketPointerFromServer_call_data(5 downto 0),
      getTxPacketPointerFromServer_call_tag => getTxPacketPointerFromServer_call_tag(0 downto 0),
      getTxPacketPointerFromServer_return_reqs => getTxPacketPointerFromServer_return_reqs(0 downto 0),
      getTxPacketPointerFromServer_return_acks => getTxPacketPointerFromServer_return_acks(0 downto 0),
      getTxPacketPointerFromServer_return_data => getTxPacketPointerFromServer_return_data(32 downto 0),
      getTxPacketPointerFromServer_return_tag => getTxPacketPointerFromServer_return_tag(0 downto 0),
      transmitPacket_call_reqs => transmitPacket_call_reqs(0 downto 0),
      transmitPacket_call_acks => transmitPacket_call_acks(0 downto 0),
      transmitPacket_call_data => transmitPacket_call_data(31 downto 0),
      transmitPacket_call_tag => transmitPacket_call_tag(0 downto 0),
      transmitPacket_return_reqs => transmitPacket_return_reqs(0 downto 0),
      transmitPacket_return_acks => transmitPacket_return_acks(0 downto 0),
      transmitPacket_return_data => transmitPacket_return_data(0 downto 0),
      transmitPacket_return_tag => transmitPacket_return_tag(0 downto 0),
      tag_in => transmitEngineDaemon_tag_in,
      tag_out => transmitEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  transmitEngineDaemon_tag_in <= (others => '0');
  transmitEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => transmitEngineDaemon_start_req, start_ack => transmitEngineDaemon_start_ack,  fin_req => transmitEngineDaemon_fin_req,  fin_ack => transmitEngineDaemon_fin_ack);
  -- module transmitPacket
  transmitPacket_packet_pointer <= transmitPacket_in_args(31 downto 0);
  transmitPacket_out_args <= transmitPacket_status ;
  -- call arbiter for module transmitPacket
  transmitPacket_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => transmitPacket_call_reqs,
      call_acks => transmitPacket_call_acks,
      return_reqs => transmitPacket_return_reqs,
      return_acks => transmitPacket_return_acks,
      call_data  => transmitPacket_call_data,
      call_tag  => transmitPacket_call_tag,
      return_tag  => transmitPacket_return_tag,
      call_mtag => transmitPacket_tag_in,
      return_mtag => transmitPacket_tag_out,
      return_data =>transmitPacket_return_data,
      call_mreq => transmitPacket_start_req,
      call_mack => transmitPacket_start_ack,
      return_mreq => transmitPacket_fin_req,
      return_mack => transmitPacket_fin_ack,
      call_mdata => transmitPacket_in_args,
      return_mdata => transmitPacket_out_args,
      clk => clk, 
      reset => reset --
    ); --
  transmitPacket_instance:transmitPacket-- 
    generic map(tag_length => 2)
    port map(-- 
      packet_pointer => transmitPacket_packet_pointer,
      status => transmitPacket_status,
      start_req => transmitPacket_start_req,
      start_ack => transmitPacket_start_ack,
      fin_req => transmitPacket_fin_req,
      fin_ack => transmitPacket_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_write_req => nic_to_mac_transmit_pipe_pipe_write_req(0 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_ack => nic_to_mac_transmit_pipe_pipe_write_ack(0 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_data => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(1 downto 0),
      accessMemory_call_acks => accessMemory_call_acks(1 downto 0),
      accessMemory_call_data => accessMemory_call_data(219 downto 0),
      accessMemory_call_tag => accessMemory_call_tag(3 downto 0),
      accessMemory_return_reqs => accessMemory_return_reqs(1 downto 0),
      accessMemory_return_acks => accessMemory_return_acks(1 downto 0),
      accessMemory_return_data => accessMemory_return_data(127 downto 0),
      accessMemory_return_tag => accessMemory_return_tag(3 downto 0),
      tag_in => transmitPacket_tag_in,
      tag_out => transmitPacket_tag_out-- 
    ); -- 
  -- module writeControlInformationToMem
  writeControlInformationToMem_base_buffer_pointer <= writeControlInformationToMem_in_args(51 downto 16);
  writeControlInformationToMem_packet_size <= writeControlInformationToMem_in_args(15 downto 8);
  writeControlInformationToMem_last_keep <= writeControlInformationToMem_in_args(7 downto 0);
  -- call arbiter for module writeControlInformationToMem
  writeControlInformationToMem_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 52,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeControlInformationToMem_call_reqs,
      call_acks => writeControlInformationToMem_call_acks,
      return_reqs => writeControlInformationToMem_return_reqs,
      return_acks => writeControlInformationToMem_return_acks,
      call_data  => writeControlInformationToMem_call_data,
      call_tag  => writeControlInformationToMem_call_tag,
      return_tag  => writeControlInformationToMem_return_tag,
      call_mtag => writeControlInformationToMem_tag_in,
      return_mtag => writeControlInformationToMem_tag_out,
      call_mreq => writeControlInformationToMem_start_req,
      call_mack => writeControlInformationToMem_start_ack,
      return_mreq => writeControlInformationToMem_fin_req,
      return_mack => writeControlInformationToMem_fin_ack,
      call_mdata => writeControlInformationToMem_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeControlInformationToMem_instance:writeControlInformationToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buffer_pointer => writeControlInformationToMem_base_buffer_pointer,
      packet_size => writeControlInformationToMem_packet_size,
      last_keep => writeControlInformationToMem_last_keep,
      start_req => writeControlInformationToMem_start_req,
      start_ack => writeControlInformationToMem_start_ack,
      fin_req => writeControlInformationToMem_fin_req,
      fin_ack => writeControlInformationToMem_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(3 downto 3),
      accessMemory_call_acks => accessMemory_call_acks(3 downto 3),
      accessMemory_call_data => accessMemory_call_data(439 downto 330),
      accessMemory_call_tag => accessMemory_call_tag(7 downto 6),
      accessMemory_return_reqs => accessMemory_return_reqs(3 downto 3),
      accessMemory_return_acks => accessMemory_return_acks(3 downto 3),
      accessMemory_return_data => accessMemory_return_data(255 downto 192),
      accessMemory_return_tag => accessMemory_return_tag(7 downto 6),
      tag_in => writeControlInformationToMem_tag_in,
      tag_out => writeControlInformationToMem_tag_out-- 
    ); -- 
  -- module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_buf_pointer <= writeEthernetHeaderToMem_in_args(35 downto 0);
  writeEthernetHeaderToMem_out_args <= writeEthernetHeaderToMem_buf_position ;
  -- call arbiter for module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeEthernetHeaderToMem_call_reqs,
      call_acks => writeEthernetHeaderToMem_call_acks,
      return_reqs => writeEthernetHeaderToMem_return_reqs,
      return_acks => writeEthernetHeaderToMem_return_acks,
      call_data  => writeEthernetHeaderToMem_call_data,
      call_tag  => writeEthernetHeaderToMem_call_tag,
      return_tag  => writeEthernetHeaderToMem_return_tag,
      call_mtag => writeEthernetHeaderToMem_tag_in,
      return_mtag => writeEthernetHeaderToMem_tag_out,
      return_data =>writeEthernetHeaderToMem_return_data,
      call_mreq => writeEthernetHeaderToMem_start_req,
      call_mack => writeEthernetHeaderToMem_start_ack,
      return_mreq => writeEthernetHeaderToMem_fin_req,
      return_mack => writeEthernetHeaderToMem_fin_ack,
      call_mdata => writeEthernetHeaderToMem_in_args,
      return_mdata => writeEthernetHeaderToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeEthernetHeaderToMem_instance:writeEthernetHeaderToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      buf_pointer => writeEthernetHeaderToMem_buf_pointer,
      buf_position => writeEthernetHeaderToMem_buf_position,
      start_req => writeEthernetHeaderToMem_start_req,
      start_ack => writeEthernetHeaderToMem_start_ack,
      fin_req => writeEthernetHeaderToMem_fin_req,
      fin_ack => writeEthernetHeaderToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_header_pipe_read_req => nic_rx_to_header_pipe_read_req(0 downto 0),
      nic_rx_to_header_pipe_read_ack => nic_rx_to_header_pipe_read_ack(0 downto 0),
      nic_rx_to_header_pipe_read_data => nic_rx_to_header_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(10 downto 10),
      accessMemory_call_acks => accessMemory_call_acks(10 downto 10),
      accessMemory_call_data => accessMemory_call_data(1209 downto 1100),
      accessMemory_call_tag => accessMemory_call_tag(21 downto 20),
      accessMemory_return_reqs => accessMemory_return_reqs(10 downto 10),
      accessMemory_return_acks => accessMemory_return_acks(10 downto 10),
      accessMemory_return_data => accessMemory_return_data(703 downto 640),
      accessMemory_return_tag => accessMemory_return_tag(21 downto 20),
      tag_in => writeEthernetHeaderToMem_tag_in,
      tag_out => writeEthernetHeaderToMem_tag_out-- 
    ); -- 
  -- module writePayloadToMem
  writePayloadToMem_base_buf_pointer <= writePayloadToMem_in_args(71 downto 36);
  writePayloadToMem_buf_pointer <= writePayloadToMem_in_args(35 downto 0);
  writePayloadToMem_out_args <= writePayloadToMem_packet_size_32 & writePayloadToMem_bad_packet_identifier & writePayloadToMem_last_keep ;
  -- call arbiter for module writePayloadToMem
  writePayloadToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 17,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writePayloadToMem_call_reqs,
      call_acks => writePayloadToMem_call_acks,
      return_reqs => writePayloadToMem_return_reqs,
      return_acks => writePayloadToMem_return_acks,
      call_data  => writePayloadToMem_call_data,
      call_tag  => writePayloadToMem_call_tag,
      return_tag  => writePayloadToMem_return_tag,
      call_mtag => writePayloadToMem_tag_in,
      return_mtag => writePayloadToMem_tag_out,
      return_data =>writePayloadToMem_return_data,
      call_mreq => writePayloadToMem_start_req,
      call_mack => writePayloadToMem_start_ack,
      return_mreq => writePayloadToMem_fin_req,
      return_mack => writePayloadToMem_fin_ack,
      call_mdata => writePayloadToMem_in_args,
      return_mdata => writePayloadToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writePayloadToMem_instance:writePayloadToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buf_pointer => writePayloadToMem_base_buf_pointer,
      buf_pointer => writePayloadToMem_buf_pointer,
      packet_size_32 => writePayloadToMem_packet_size_32,
      bad_packet_identifier => writePayloadToMem_bad_packet_identifier,
      last_keep => writePayloadToMem_last_keep,
      start_req => writePayloadToMem_start_req,
      start_ack => writePayloadToMem_start_ack,
      fin_req => writePayloadToMem_fin_req,
      fin_ack => writePayloadToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_packet_pipe_read_req => nic_rx_to_packet_pipe_read_req(0 downto 0),
      nic_rx_to_packet_pipe_read_ack => nic_rx_to_packet_pipe_read_ack(0 downto 0),
      nic_rx_to_packet_pipe_read_data => nic_rx_to_packet_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(2 downto 2),
      accessMemory_call_acks => accessMemory_call_acks(2 downto 2),
      accessMemory_call_data => accessMemory_call_data(329 downto 220),
      accessMemory_call_tag => accessMemory_call_tag(5 downto 4),
      accessMemory_return_reqs => accessMemory_return_reqs(2 downto 2),
      accessMemory_return_acks => accessMemory_return_acks(2 downto 2),
      accessMemory_return_data => accessMemory_return_data(191 downto 128),
      accessMemory_return_tag => accessMemory_return_tag(5 downto 4),
      tag_in => writePayloadToMem_tag_in,
      tag_out => writePayloadToMem_tag_out-- 
    ); -- 
  AFB_NIC_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 74,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => AFB_NIC_REQUEST_pipe_read_req,
      read_ack => AFB_NIC_REQUEST_pipe_read_ack,
      read_data => AFB_NIC_REQUEST_pipe_read_data,
      write_req => AFB_NIC_REQUEST_pipe_write_req,
      write_ack => AFB_NIC_REQUEST_pipe_write_ack,
      write_data => AFB_NIC_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  AFB_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => AFB_NIC_RESPONSE_pipe_read_req,
      read_ack => AFB_NIC_RESPONSE_pipe_read_ack,
      read_data => AFB_NIC_RESPONSE_pipe_read_data,
      write_req => AFB_NIC_RESPONSE_pipe_write_req,
      write_ack => AFB_NIC_RESPONSE_pipe_write_ack,
      write_data => AFB_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  CONTROL_REGISTER_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe CONTROL_REGISTER",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => CONTROL_REGISTER,
      write_req => CONTROL_REGISTER_pipe_write_req,
      write_ack => CONTROL_REGISTER_pipe_write_ack,
      write_data => CONTROL_REGISTER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  FREE_Q_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe FREE_Q",
      volatile_flag => false,
      num_writes => 1,
      data_width => 36 --
    ) 
    port map( -- 
      read_data => FREE_Q,
      write_req => FREE_Q_pipe_write_req,
      write_ack => FREE_Q_pipe_write_ack,
      write_data => FREE_Q_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_READ_TX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_READ_TX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_READ_TX_QUEUE_INDEX,
      write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_WRITTEN_RX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_WRITTEN_RX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_WRITTEN_RX_QUEUE_INDEX,
      write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEMORY_TO_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEMORY_TO_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req,
      read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack,
      read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data,
      write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req,
      write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack,
      write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_REQUEST_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_REQUEST_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 43,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_RESPONSE_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_TO_MEMORY_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_TO_MEMORY_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req,
      read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack,
      read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data,
      write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req,
      write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack,
      write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NUMBER_OF_SERVERS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NUMBER_OF_SERVERS",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => NUMBER_OF_SERVERS,
      write_req => NUMBER_OF_SERVERS_pipe_write_req,
      write_ack => NUMBER_OF_SERVERS_pipe_write_ack,
      write_data => NUMBER_OF_SERVERS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  control_word_request_pipe_0_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe control_word_request_pipe_0",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => control_word_request_pipe_0_pipe_read_req,
      read_ack => control_word_request_pipe_0_pipe_read_ack,
      read_data => control_word_request_pipe_0_pipe_read_data,
      write_req => control_word_request_pipe_0_pipe_write_req,
      write_ack => control_word_request_pipe_0_pipe_write_ack,
      write_data => control_word_request_pipe_0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  control_word_request_pipe_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe control_word_request_pipe_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => control_word_request_pipe_1_pipe_read_req,
      read_ack => control_word_request_pipe_1_pipe_read_ack,
      read_data => control_word_request_pipe_1_pipe_read_data,
      write_req => control_word_request_pipe_1_pipe_write_req,
      write_ack => control_word_request_pipe_1_pipe_write_ack,
      write_data => control_word_request_pipe_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  control_word_response_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe control_word_response_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => control_word_response_pipe_pipe_read_req,
      read_ack => control_word_response_pipe_pipe_read_ack,
      read_data => control_word_response_pipe_pipe_read_data,
      write_req => control_word_response_pipe_pipe_write_req,
      write_ack => control_word_response_pipe_pipe_write_ack,
      write_data => control_word_response_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mac_to_nic_data_pipe_read_req,
      read_ack => mac_to_nic_data_pipe_read_ack,
      read_data => mac_to_nic_data_pipe_read_data,
      write_req => mac_to_nic_data_pipe_write_req,
      write_ack => mac_to_nic_data_pipe_write_ack,
      write_data => mac_to_nic_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_0_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data_0",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mac_to_nic_data_0_pipe_read_req,
      read_ack => mac_to_nic_data_0_pipe_read_ack,
      read_data => mac_to_nic_data_0_pipe_read_data,
      write_req => mac_to_nic_data_0_pipe_write_req,
      write_ack => mac_to_nic_data_0_pipe_write_ack,
      write_data => mac_to_nic_data_0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data_1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mac_to_nic_data_1_pipe_read_req,
      read_ack => mac_to_nic_data_1_pipe_read_ack,
      read_data => mac_to_nic_data_1_pipe_read_data,
      write_req => mac_to_nic_data_1_pipe_write_req,
      write_ack => mac_to_nic_data_1_pipe_write_ack,
      write_data => mac_to_nic_data_1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mem_req0_pipe0_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mem_req0_pipe0",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mem_req0_pipe0_pipe_read_req,
      read_ack => mem_req0_pipe0_pipe_read_ack,
      read_data => mem_req0_pipe0_pipe_read_data,
      write_req => mem_req0_pipe0_pipe_write_req,
      write_ack => mem_req0_pipe0_pipe_write_ack,
      write_data => mem_req0_pipe0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mem_req0_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mem_req0_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mem_req0_pipe1_pipe_read_req,
      read_ack => mem_req0_pipe1_pipe_read_ack,
      read_data => mem_req0_pipe1_pipe_read_data,
      write_req => mem_req0_pipe1_pipe_write_req,
      write_ack => mem_req0_pipe1_pipe_write_ack,
      write_data => mem_req0_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mem_resp0_pipe0_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mem_resp0_pipe0",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mem_resp0_pipe0_pipe_read_req,
      read_ack => mem_resp0_pipe0_pipe_read_ack,
      read_data => mem_resp0_pipe0_pipe_read_data,
      write_req => mem_resp0_pipe0_pipe_write_req,
      write_ack => mem_resp0_pipe0_pipe_write_ack,
      write_data => mem_resp0_pipe0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mem_resp0_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mem_resp0_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mem_resp0_pipe1_pipe_read_req,
      read_ack => mem_resp0_pipe1_pipe_read_ack,
      read_data => mem_resp0_pipe1_pipe_read_data,
      write_req => mem_resp0_pipe1_pipe_write_req,
      write_ack => mem_resp0_pipe1_pipe_write_ack,
      write_data => mem_resp0_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_header_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_header",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_header_pipe_read_req,
      read_ack => nic_rx_to_header_pipe_read_ack,
      read_data => nic_rx_to_header_pipe_read_data,
      write_req => nic_rx_to_header_pipe_write_req,
      write_ack => nic_rx_to_header_pipe_write_ack,
      write_data => nic_rx_to_header_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_packet_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_packet",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_packet_pipe_read_req,
      read_ack => nic_rx_to_packet_pipe_read_ack,
      read_data => nic_rx_to_packet_pipe_read_data,
      write_req => nic_rx_to_packet_pipe_write_req,
      write_ack => nic_rx_to_packet_pipe_write_ack,
      write_data => nic_rx_to_packet_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_to_mac_transmit_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_to_mac_transmit_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_to_mac_transmit_pipe_pipe_read_req,
      read_ack => nic_to_mac_transmit_pipe_pipe_read_ack,
      read_data => nic_to_mac_transmit_pipe_pipe_read_data,
      write_req => nic_to_mac_transmit_pipe_pipe_write_req,
      write_ack => nic_to_mac_transmit_pipe_pipe_write_ack,
      write_data => nic_to_mac_transmit_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 6,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 6,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
